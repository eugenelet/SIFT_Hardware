module detect_keypoint(
  top_0,
  top_1,
  top_2,
  mid_0,
  mid_1,
  mid_2,
  btm_0,
  btm_1,
  btm_2,
  is_keypoint
);

input       [5119:0]	top_0,
						top_1,
						top_2,
						mid_0,
						mid_1,
						mid_2,
						btm_0,
						btm_1,
						btm_2;
output reg 	 [637:0]	is_keypoint;

wire	[25:0]		detect_max[0:637];
assign detect_max[0][0] = (mid_1[15:8] > top_0[7:0]) ? 1 : 0;
assign detect_max[0][1] = (mid_1[15:8] > top_0[15:8]) ? 1 : 0;
assign detect_max[0][2] = (mid_1[15:8] > top_0[23:16]) ? 1 : 0;
assign detect_max[0][3] = (mid_1[15:8] > top_1[7:0]) ? 1 : 0;
assign detect_max[0][4] = (mid_1[15:8] > top_1[15:8]) ? 1 : 0;
assign detect_max[0][5] = (mid_1[15:8] > top_1[23:16]) ? 1 : 0;
assign detect_max[0][6] = (mid_1[15:8] > top_2[7:0]) ? 1 : 0;
assign detect_max[0][7] = (mid_1[15:8] > top_2[15:8]) ? 1 : 0;
assign detect_max[0][8] = (mid_1[15:8] > top_2[23:16]) ? 1 : 0;
assign detect_max[0][9] = (mid_1[15:8] > mid_0[7:0]) ? 1 : 0;
assign detect_max[0][10] = (mid_1[15:8] > mid_0[15:8]) ? 1 : 0;
assign detect_max[0][11] = (mid_1[15:8] > mid_0[23:16]) ? 1 : 0;
assign detect_max[0][12] = (mid_1[15:8] > mid_1[7:0]) ? 1 : 0;
assign detect_max[0][13] = (mid_1[15:8] > mid_1[23:16]) ? 1 : 0;
assign detect_max[0][14] = (mid_1[15:8] > mid_2[7:0]) ? 1 : 0;
assign detect_max[0][15] = (mid_1[15:8] > mid_2[15:8]) ? 1 : 0;
assign detect_max[0][16] = (mid_1[15:8] > mid_2[23:16]) ? 1 : 0;
assign detect_max[0][17] = (mid_1[15:8] > btm_0[7:0]) ? 1 : 0;
assign detect_max[0][18] = (mid_1[15:8] > btm_0[15:8]) ? 1 : 0;
assign detect_max[0][19] = (mid_1[15:8] > btm_0[23:16]) ? 1 : 0;
assign detect_max[0][20] = (mid_1[15:8] > btm_1[7:0]) ? 1 : 0;
assign detect_max[0][21] = (mid_1[15:8] > btm_1[15:8]) ? 1 : 0;
assign detect_max[0][22] = (mid_1[15:8] > btm_1[23:16]) ? 1 : 0;
assign detect_max[0][23] = (mid_1[15:8] > btm_2[7:0]) ? 1 : 0;
assign detect_max[0][24] = (mid_1[15:8] > btm_2[15:8]) ? 1 : 0;
assign detect_max[0][25] = (mid_1[15:8] > btm_2[23:16]) ? 1 : 0;

assign detect_max[1][0] = (mid_1[23:16] > top_0[15:8]) ? 1 : 0;
assign detect_max[1][1] = (mid_1[23:16] > top_0[23:16]) ? 1 : 0;
assign detect_max[1][2] = (mid_1[23:16] > top_0[31:24]) ? 1 : 0;
assign detect_max[1][3] = (mid_1[23:16] > top_1[15:8]) ? 1 : 0;
assign detect_max[1][4] = (mid_1[23:16] > top_1[23:16]) ? 1 : 0;
assign detect_max[1][5] = (mid_1[23:16] > top_1[31:24]) ? 1 : 0;
assign detect_max[1][6] = (mid_1[23:16] > top_2[15:8]) ? 1 : 0;
assign detect_max[1][7] = (mid_1[23:16] > top_2[23:16]) ? 1 : 0;
assign detect_max[1][8] = (mid_1[23:16] > top_2[31:24]) ? 1 : 0;
assign detect_max[1][9] = (mid_1[23:16] > mid_0[15:8]) ? 1 : 0;
assign detect_max[1][10] = (mid_1[23:16] > mid_0[23:16]) ? 1 : 0;
assign detect_max[1][11] = (mid_1[23:16] > mid_0[31:24]) ? 1 : 0;
assign detect_max[1][12] = (mid_1[23:16] > mid_1[15:8]) ? 1 : 0;
assign detect_max[1][13] = (mid_1[23:16] > mid_1[31:24]) ? 1 : 0;
assign detect_max[1][14] = (mid_1[23:16] > mid_2[15:8]) ? 1 : 0;
assign detect_max[1][15] = (mid_1[23:16] > mid_2[23:16]) ? 1 : 0;
assign detect_max[1][16] = (mid_1[23:16] > mid_2[31:24]) ? 1 : 0;
assign detect_max[1][17] = (mid_1[23:16] > btm_0[15:8]) ? 1 : 0;
assign detect_max[1][18] = (mid_1[23:16] > btm_0[23:16]) ? 1 : 0;
assign detect_max[1][19] = (mid_1[23:16] > btm_0[31:24]) ? 1 : 0;
assign detect_max[1][20] = (mid_1[23:16] > btm_1[15:8]) ? 1 : 0;
assign detect_max[1][21] = (mid_1[23:16] > btm_1[23:16]) ? 1 : 0;
assign detect_max[1][22] = (mid_1[23:16] > btm_1[31:24]) ? 1 : 0;
assign detect_max[1][23] = (mid_1[23:16] > btm_2[15:8]) ? 1 : 0;
assign detect_max[1][24] = (mid_1[23:16] > btm_2[23:16]) ? 1 : 0;
assign detect_max[1][25] = (mid_1[23:16] > btm_2[31:24]) ? 1 : 0;

assign detect_max[2][0] = (mid_1[31:24] > top_0[23:16]) ? 1 : 0;
assign detect_max[2][1] = (mid_1[31:24] > top_0[31:24]) ? 1 : 0;
assign detect_max[2][2] = (mid_1[31:24] > top_0[39:32]) ? 1 : 0;
assign detect_max[2][3] = (mid_1[31:24] > top_1[23:16]) ? 1 : 0;
assign detect_max[2][4] = (mid_1[31:24] > top_1[31:24]) ? 1 : 0;
assign detect_max[2][5] = (mid_1[31:24] > top_1[39:32]) ? 1 : 0;
assign detect_max[2][6] = (mid_1[31:24] > top_2[23:16]) ? 1 : 0;
assign detect_max[2][7] = (mid_1[31:24] > top_2[31:24]) ? 1 : 0;
assign detect_max[2][8] = (mid_1[31:24] > top_2[39:32]) ? 1 : 0;
assign detect_max[2][9] = (mid_1[31:24] > mid_0[23:16]) ? 1 : 0;
assign detect_max[2][10] = (mid_1[31:24] > mid_0[31:24]) ? 1 : 0;
assign detect_max[2][11] = (mid_1[31:24] > mid_0[39:32]) ? 1 : 0;
assign detect_max[2][12] = (mid_1[31:24] > mid_1[23:16]) ? 1 : 0;
assign detect_max[2][13] = (mid_1[31:24] > mid_1[39:32]) ? 1 : 0;
assign detect_max[2][14] = (mid_1[31:24] > mid_2[23:16]) ? 1 : 0;
assign detect_max[2][15] = (mid_1[31:24] > mid_2[31:24]) ? 1 : 0;
assign detect_max[2][16] = (mid_1[31:24] > mid_2[39:32]) ? 1 : 0;
assign detect_max[2][17] = (mid_1[31:24] > btm_0[23:16]) ? 1 : 0;
assign detect_max[2][18] = (mid_1[31:24] > btm_0[31:24]) ? 1 : 0;
assign detect_max[2][19] = (mid_1[31:24] > btm_0[39:32]) ? 1 : 0;
assign detect_max[2][20] = (mid_1[31:24] > btm_1[23:16]) ? 1 : 0;
assign detect_max[2][21] = (mid_1[31:24] > btm_1[31:24]) ? 1 : 0;
assign detect_max[2][22] = (mid_1[31:24] > btm_1[39:32]) ? 1 : 0;
assign detect_max[2][23] = (mid_1[31:24] > btm_2[23:16]) ? 1 : 0;
assign detect_max[2][24] = (mid_1[31:24] > btm_2[31:24]) ? 1 : 0;
assign detect_max[2][25] = (mid_1[31:24] > btm_2[39:32]) ? 1 : 0;

assign detect_max[3][0] = (mid_1[39:32] > top_0[31:24]) ? 1 : 0;
assign detect_max[3][1] = (mid_1[39:32] > top_0[39:32]) ? 1 : 0;
assign detect_max[3][2] = (mid_1[39:32] > top_0[47:40]) ? 1 : 0;
assign detect_max[3][3] = (mid_1[39:32] > top_1[31:24]) ? 1 : 0;
assign detect_max[3][4] = (mid_1[39:32] > top_1[39:32]) ? 1 : 0;
assign detect_max[3][5] = (mid_1[39:32] > top_1[47:40]) ? 1 : 0;
assign detect_max[3][6] = (mid_1[39:32] > top_2[31:24]) ? 1 : 0;
assign detect_max[3][7] = (mid_1[39:32] > top_2[39:32]) ? 1 : 0;
assign detect_max[3][8] = (mid_1[39:32] > top_2[47:40]) ? 1 : 0;
assign detect_max[3][9] = (mid_1[39:32] > mid_0[31:24]) ? 1 : 0;
assign detect_max[3][10] = (mid_1[39:32] > mid_0[39:32]) ? 1 : 0;
assign detect_max[3][11] = (mid_1[39:32] > mid_0[47:40]) ? 1 : 0;
assign detect_max[3][12] = (mid_1[39:32] > mid_1[31:24]) ? 1 : 0;
assign detect_max[3][13] = (mid_1[39:32] > mid_1[47:40]) ? 1 : 0;
assign detect_max[3][14] = (mid_1[39:32] > mid_2[31:24]) ? 1 : 0;
assign detect_max[3][15] = (mid_1[39:32] > mid_2[39:32]) ? 1 : 0;
assign detect_max[3][16] = (mid_1[39:32] > mid_2[47:40]) ? 1 : 0;
assign detect_max[3][17] = (mid_1[39:32] > btm_0[31:24]) ? 1 : 0;
assign detect_max[3][18] = (mid_1[39:32] > btm_0[39:32]) ? 1 : 0;
assign detect_max[3][19] = (mid_1[39:32] > btm_0[47:40]) ? 1 : 0;
assign detect_max[3][20] = (mid_1[39:32] > btm_1[31:24]) ? 1 : 0;
assign detect_max[3][21] = (mid_1[39:32] > btm_1[39:32]) ? 1 : 0;
assign detect_max[3][22] = (mid_1[39:32] > btm_1[47:40]) ? 1 : 0;
assign detect_max[3][23] = (mid_1[39:32] > btm_2[31:24]) ? 1 : 0;
assign detect_max[3][24] = (mid_1[39:32] > btm_2[39:32]) ? 1 : 0;
assign detect_max[3][25] = (mid_1[39:32] > btm_2[47:40]) ? 1 : 0;

assign detect_max[4][0] = (mid_1[47:40] > top_0[39:32]) ? 1 : 0;
assign detect_max[4][1] = (mid_1[47:40] > top_0[47:40]) ? 1 : 0;
assign detect_max[4][2] = (mid_1[47:40] > top_0[55:48]) ? 1 : 0;
assign detect_max[4][3] = (mid_1[47:40] > top_1[39:32]) ? 1 : 0;
assign detect_max[4][4] = (mid_1[47:40] > top_1[47:40]) ? 1 : 0;
assign detect_max[4][5] = (mid_1[47:40] > top_1[55:48]) ? 1 : 0;
assign detect_max[4][6] = (mid_1[47:40] > top_2[39:32]) ? 1 : 0;
assign detect_max[4][7] = (mid_1[47:40] > top_2[47:40]) ? 1 : 0;
assign detect_max[4][8] = (mid_1[47:40] > top_2[55:48]) ? 1 : 0;
assign detect_max[4][9] = (mid_1[47:40] > mid_0[39:32]) ? 1 : 0;
assign detect_max[4][10] = (mid_1[47:40] > mid_0[47:40]) ? 1 : 0;
assign detect_max[4][11] = (mid_1[47:40] > mid_0[55:48]) ? 1 : 0;
assign detect_max[4][12] = (mid_1[47:40] > mid_1[39:32]) ? 1 : 0;
assign detect_max[4][13] = (mid_1[47:40] > mid_1[55:48]) ? 1 : 0;
assign detect_max[4][14] = (mid_1[47:40] > mid_2[39:32]) ? 1 : 0;
assign detect_max[4][15] = (mid_1[47:40] > mid_2[47:40]) ? 1 : 0;
assign detect_max[4][16] = (mid_1[47:40] > mid_2[55:48]) ? 1 : 0;
assign detect_max[4][17] = (mid_1[47:40] > btm_0[39:32]) ? 1 : 0;
assign detect_max[4][18] = (mid_1[47:40] > btm_0[47:40]) ? 1 : 0;
assign detect_max[4][19] = (mid_1[47:40] > btm_0[55:48]) ? 1 : 0;
assign detect_max[4][20] = (mid_1[47:40] > btm_1[39:32]) ? 1 : 0;
assign detect_max[4][21] = (mid_1[47:40] > btm_1[47:40]) ? 1 : 0;
assign detect_max[4][22] = (mid_1[47:40] > btm_1[55:48]) ? 1 : 0;
assign detect_max[4][23] = (mid_1[47:40] > btm_2[39:32]) ? 1 : 0;
assign detect_max[4][24] = (mid_1[47:40] > btm_2[47:40]) ? 1 : 0;
assign detect_max[4][25] = (mid_1[47:40] > btm_2[55:48]) ? 1 : 0;

assign detect_max[5][0] = (mid_1[55:48] > top_0[47:40]) ? 1 : 0;
assign detect_max[5][1] = (mid_1[55:48] > top_0[55:48]) ? 1 : 0;
assign detect_max[5][2] = (mid_1[55:48] > top_0[63:56]) ? 1 : 0;
assign detect_max[5][3] = (mid_1[55:48] > top_1[47:40]) ? 1 : 0;
assign detect_max[5][4] = (mid_1[55:48] > top_1[55:48]) ? 1 : 0;
assign detect_max[5][5] = (mid_1[55:48] > top_1[63:56]) ? 1 : 0;
assign detect_max[5][6] = (mid_1[55:48] > top_2[47:40]) ? 1 : 0;
assign detect_max[5][7] = (mid_1[55:48] > top_2[55:48]) ? 1 : 0;
assign detect_max[5][8] = (mid_1[55:48] > top_2[63:56]) ? 1 : 0;
assign detect_max[5][9] = (mid_1[55:48] > mid_0[47:40]) ? 1 : 0;
assign detect_max[5][10] = (mid_1[55:48] > mid_0[55:48]) ? 1 : 0;
assign detect_max[5][11] = (mid_1[55:48] > mid_0[63:56]) ? 1 : 0;
assign detect_max[5][12] = (mid_1[55:48] > mid_1[47:40]) ? 1 : 0;
assign detect_max[5][13] = (mid_1[55:48] > mid_1[63:56]) ? 1 : 0;
assign detect_max[5][14] = (mid_1[55:48] > mid_2[47:40]) ? 1 : 0;
assign detect_max[5][15] = (mid_1[55:48] > mid_2[55:48]) ? 1 : 0;
assign detect_max[5][16] = (mid_1[55:48] > mid_2[63:56]) ? 1 : 0;
assign detect_max[5][17] = (mid_1[55:48] > btm_0[47:40]) ? 1 : 0;
assign detect_max[5][18] = (mid_1[55:48] > btm_0[55:48]) ? 1 : 0;
assign detect_max[5][19] = (mid_1[55:48] > btm_0[63:56]) ? 1 : 0;
assign detect_max[5][20] = (mid_1[55:48] > btm_1[47:40]) ? 1 : 0;
assign detect_max[5][21] = (mid_1[55:48] > btm_1[55:48]) ? 1 : 0;
assign detect_max[5][22] = (mid_1[55:48] > btm_1[63:56]) ? 1 : 0;
assign detect_max[5][23] = (mid_1[55:48] > btm_2[47:40]) ? 1 : 0;
assign detect_max[5][24] = (mid_1[55:48] > btm_2[55:48]) ? 1 : 0;
assign detect_max[5][25] = (mid_1[55:48] > btm_2[63:56]) ? 1 : 0;

assign detect_max[6][0] = (mid_1[63:56] > top_0[55:48]) ? 1 : 0;
assign detect_max[6][1] = (mid_1[63:56] > top_0[63:56]) ? 1 : 0;
assign detect_max[6][2] = (mid_1[63:56] > top_0[71:64]) ? 1 : 0;
assign detect_max[6][3] = (mid_1[63:56] > top_1[55:48]) ? 1 : 0;
assign detect_max[6][4] = (mid_1[63:56] > top_1[63:56]) ? 1 : 0;
assign detect_max[6][5] = (mid_1[63:56] > top_1[71:64]) ? 1 : 0;
assign detect_max[6][6] = (mid_1[63:56] > top_2[55:48]) ? 1 : 0;
assign detect_max[6][7] = (mid_1[63:56] > top_2[63:56]) ? 1 : 0;
assign detect_max[6][8] = (mid_1[63:56] > top_2[71:64]) ? 1 : 0;
assign detect_max[6][9] = (mid_1[63:56] > mid_0[55:48]) ? 1 : 0;
assign detect_max[6][10] = (mid_1[63:56] > mid_0[63:56]) ? 1 : 0;
assign detect_max[6][11] = (mid_1[63:56] > mid_0[71:64]) ? 1 : 0;
assign detect_max[6][12] = (mid_1[63:56] > mid_1[55:48]) ? 1 : 0;
assign detect_max[6][13] = (mid_1[63:56] > mid_1[71:64]) ? 1 : 0;
assign detect_max[6][14] = (mid_1[63:56] > mid_2[55:48]) ? 1 : 0;
assign detect_max[6][15] = (mid_1[63:56] > mid_2[63:56]) ? 1 : 0;
assign detect_max[6][16] = (mid_1[63:56] > mid_2[71:64]) ? 1 : 0;
assign detect_max[6][17] = (mid_1[63:56] > btm_0[55:48]) ? 1 : 0;
assign detect_max[6][18] = (mid_1[63:56] > btm_0[63:56]) ? 1 : 0;
assign detect_max[6][19] = (mid_1[63:56] > btm_0[71:64]) ? 1 : 0;
assign detect_max[6][20] = (mid_1[63:56] > btm_1[55:48]) ? 1 : 0;
assign detect_max[6][21] = (mid_1[63:56] > btm_1[63:56]) ? 1 : 0;
assign detect_max[6][22] = (mid_1[63:56] > btm_1[71:64]) ? 1 : 0;
assign detect_max[6][23] = (mid_1[63:56] > btm_2[55:48]) ? 1 : 0;
assign detect_max[6][24] = (mid_1[63:56] > btm_2[63:56]) ? 1 : 0;
assign detect_max[6][25] = (mid_1[63:56] > btm_2[71:64]) ? 1 : 0;

assign detect_max[7][0] = (mid_1[71:64] > top_0[63:56]) ? 1 : 0;
assign detect_max[7][1] = (mid_1[71:64] > top_0[71:64]) ? 1 : 0;
assign detect_max[7][2] = (mid_1[71:64] > top_0[79:72]) ? 1 : 0;
assign detect_max[7][3] = (mid_1[71:64] > top_1[63:56]) ? 1 : 0;
assign detect_max[7][4] = (mid_1[71:64] > top_1[71:64]) ? 1 : 0;
assign detect_max[7][5] = (mid_1[71:64] > top_1[79:72]) ? 1 : 0;
assign detect_max[7][6] = (mid_1[71:64] > top_2[63:56]) ? 1 : 0;
assign detect_max[7][7] = (mid_1[71:64] > top_2[71:64]) ? 1 : 0;
assign detect_max[7][8] = (mid_1[71:64] > top_2[79:72]) ? 1 : 0;
assign detect_max[7][9] = (mid_1[71:64] > mid_0[63:56]) ? 1 : 0;
assign detect_max[7][10] = (mid_1[71:64] > mid_0[71:64]) ? 1 : 0;
assign detect_max[7][11] = (mid_1[71:64] > mid_0[79:72]) ? 1 : 0;
assign detect_max[7][12] = (mid_1[71:64] > mid_1[63:56]) ? 1 : 0;
assign detect_max[7][13] = (mid_1[71:64] > mid_1[79:72]) ? 1 : 0;
assign detect_max[7][14] = (mid_1[71:64] > mid_2[63:56]) ? 1 : 0;
assign detect_max[7][15] = (mid_1[71:64] > mid_2[71:64]) ? 1 : 0;
assign detect_max[7][16] = (mid_1[71:64] > mid_2[79:72]) ? 1 : 0;
assign detect_max[7][17] = (mid_1[71:64] > btm_0[63:56]) ? 1 : 0;
assign detect_max[7][18] = (mid_1[71:64] > btm_0[71:64]) ? 1 : 0;
assign detect_max[7][19] = (mid_1[71:64] > btm_0[79:72]) ? 1 : 0;
assign detect_max[7][20] = (mid_1[71:64] > btm_1[63:56]) ? 1 : 0;
assign detect_max[7][21] = (mid_1[71:64] > btm_1[71:64]) ? 1 : 0;
assign detect_max[7][22] = (mid_1[71:64] > btm_1[79:72]) ? 1 : 0;
assign detect_max[7][23] = (mid_1[71:64] > btm_2[63:56]) ? 1 : 0;
assign detect_max[7][24] = (mid_1[71:64] > btm_2[71:64]) ? 1 : 0;
assign detect_max[7][25] = (mid_1[71:64] > btm_2[79:72]) ? 1 : 0;

assign detect_max[8][0] = (mid_1[79:72] > top_0[71:64]) ? 1 : 0;
assign detect_max[8][1] = (mid_1[79:72] > top_0[79:72]) ? 1 : 0;
assign detect_max[8][2] = (mid_1[79:72] > top_0[87:80]) ? 1 : 0;
assign detect_max[8][3] = (mid_1[79:72] > top_1[71:64]) ? 1 : 0;
assign detect_max[8][4] = (mid_1[79:72] > top_1[79:72]) ? 1 : 0;
assign detect_max[8][5] = (mid_1[79:72] > top_1[87:80]) ? 1 : 0;
assign detect_max[8][6] = (mid_1[79:72] > top_2[71:64]) ? 1 : 0;
assign detect_max[8][7] = (mid_1[79:72] > top_2[79:72]) ? 1 : 0;
assign detect_max[8][8] = (mid_1[79:72] > top_2[87:80]) ? 1 : 0;
assign detect_max[8][9] = (mid_1[79:72] > mid_0[71:64]) ? 1 : 0;
assign detect_max[8][10] = (mid_1[79:72] > mid_0[79:72]) ? 1 : 0;
assign detect_max[8][11] = (mid_1[79:72] > mid_0[87:80]) ? 1 : 0;
assign detect_max[8][12] = (mid_1[79:72] > mid_1[71:64]) ? 1 : 0;
assign detect_max[8][13] = (mid_1[79:72] > mid_1[87:80]) ? 1 : 0;
assign detect_max[8][14] = (mid_1[79:72] > mid_2[71:64]) ? 1 : 0;
assign detect_max[8][15] = (mid_1[79:72] > mid_2[79:72]) ? 1 : 0;
assign detect_max[8][16] = (mid_1[79:72] > mid_2[87:80]) ? 1 : 0;
assign detect_max[8][17] = (mid_1[79:72] > btm_0[71:64]) ? 1 : 0;
assign detect_max[8][18] = (mid_1[79:72] > btm_0[79:72]) ? 1 : 0;
assign detect_max[8][19] = (mid_1[79:72] > btm_0[87:80]) ? 1 : 0;
assign detect_max[8][20] = (mid_1[79:72] > btm_1[71:64]) ? 1 : 0;
assign detect_max[8][21] = (mid_1[79:72] > btm_1[79:72]) ? 1 : 0;
assign detect_max[8][22] = (mid_1[79:72] > btm_1[87:80]) ? 1 : 0;
assign detect_max[8][23] = (mid_1[79:72] > btm_2[71:64]) ? 1 : 0;
assign detect_max[8][24] = (mid_1[79:72] > btm_2[79:72]) ? 1 : 0;
assign detect_max[8][25] = (mid_1[79:72] > btm_2[87:80]) ? 1 : 0;

assign detect_max[9][0] = (mid_1[87:80] > top_0[79:72]) ? 1 : 0;
assign detect_max[9][1] = (mid_1[87:80] > top_0[87:80]) ? 1 : 0;
assign detect_max[9][2] = (mid_1[87:80] > top_0[95:88]) ? 1 : 0;
assign detect_max[9][3] = (mid_1[87:80] > top_1[79:72]) ? 1 : 0;
assign detect_max[9][4] = (mid_1[87:80] > top_1[87:80]) ? 1 : 0;
assign detect_max[9][5] = (mid_1[87:80] > top_1[95:88]) ? 1 : 0;
assign detect_max[9][6] = (mid_1[87:80] > top_2[79:72]) ? 1 : 0;
assign detect_max[9][7] = (mid_1[87:80] > top_2[87:80]) ? 1 : 0;
assign detect_max[9][8] = (mid_1[87:80] > top_2[95:88]) ? 1 : 0;
assign detect_max[9][9] = (mid_1[87:80] > mid_0[79:72]) ? 1 : 0;
assign detect_max[9][10] = (mid_1[87:80] > mid_0[87:80]) ? 1 : 0;
assign detect_max[9][11] = (mid_1[87:80] > mid_0[95:88]) ? 1 : 0;
assign detect_max[9][12] = (mid_1[87:80] > mid_1[79:72]) ? 1 : 0;
assign detect_max[9][13] = (mid_1[87:80] > mid_1[95:88]) ? 1 : 0;
assign detect_max[9][14] = (mid_1[87:80] > mid_2[79:72]) ? 1 : 0;
assign detect_max[9][15] = (mid_1[87:80] > mid_2[87:80]) ? 1 : 0;
assign detect_max[9][16] = (mid_1[87:80] > mid_2[95:88]) ? 1 : 0;
assign detect_max[9][17] = (mid_1[87:80] > btm_0[79:72]) ? 1 : 0;
assign detect_max[9][18] = (mid_1[87:80] > btm_0[87:80]) ? 1 : 0;
assign detect_max[9][19] = (mid_1[87:80] > btm_0[95:88]) ? 1 : 0;
assign detect_max[9][20] = (mid_1[87:80] > btm_1[79:72]) ? 1 : 0;
assign detect_max[9][21] = (mid_1[87:80] > btm_1[87:80]) ? 1 : 0;
assign detect_max[9][22] = (mid_1[87:80] > btm_1[95:88]) ? 1 : 0;
assign detect_max[9][23] = (mid_1[87:80] > btm_2[79:72]) ? 1 : 0;
assign detect_max[9][24] = (mid_1[87:80] > btm_2[87:80]) ? 1 : 0;
assign detect_max[9][25] = (mid_1[87:80] > btm_2[95:88]) ? 1 : 0;

assign detect_max[10][0] = (mid_1[95:88] > top_0[87:80]) ? 1 : 0;
assign detect_max[10][1] = (mid_1[95:88] > top_0[95:88]) ? 1 : 0;
assign detect_max[10][2] = (mid_1[95:88] > top_0[103:96]) ? 1 : 0;
assign detect_max[10][3] = (mid_1[95:88] > top_1[87:80]) ? 1 : 0;
assign detect_max[10][4] = (mid_1[95:88] > top_1[95:88]) ? 1 : 0;
assign detect_max[10][5] = (mid_1[95:88] > top_1[103:96]) ? 1 : 0;
assign detect_max[10][6] = (mid_1[95:88] > top_2[87:80]) ? 1 : 0;
assign detect_max[10][7] = (mid_1[95:88] > top_2[95:88]) ? 1 : 0;
assign detect_max[10][8] = (mid_1[95:88] > top_2[103:96]) ? 1 : 0;
assign detect_max[10][9] = (mid_1[95:88] > mid_0[87:80]) ? 1 : 0;
assign detect_max[10][10] = (mid_1[95:88] > mid_0[95:88]) ? 1 : 0;
assign detect_max[10][11] = (mid_1[95:88] > mid_0[103:96]) ? 1 : 0;
assign detect_max[10][12] = (mid_1[95:88] > mid_1[87:80]) ? 1 : 0;
assign detect_max[10][13] = (mid_1[95:88] > mid_1[103:96]) ? 1 : 0;
assign detect_max[10][14] = (mid_1[95:88] > mid_2[87:80]) ? 1 : 0;
assign detect_max[10][15] = (mid_1[95:88] > mid_2[95:88]) ? 1 : 0;
assign detect_max[10][16] = (mid_1[95:88] > mid_2[103:96]) ? 1 : 0;
assign detect_max[10][17] = (mid_1[95:88] > btm_0[87:80]) ? 1 : 0;
assign detect_max[10][18] = (mid_1[95:88] > btm_0[95:88]) ? 1 : 0;
assign detect_max[10][19] = (mid_1[95:88] > btm_0[103:96]) ? 1 : 0;
assign detect_max[10][20] = (mid_1[95:88] > btm_1[87:80]) ? 1 : 0;
assign detect_max[10][21] = (mid_1[95:88] > btm_1[95:88]) ? 1 : 0;
assign detect_max[10][22] = (mid_1[95:88] > btm_1[103:96]) ? 1 : 0;
assign detect_max[10][23] = (mid_1[95:88] > btm_2[87:80]) ? 1 : 0;
assign detect_max[10][24] = (mid_1[95:88] > btm_2[95:88]) ? 1 : 0;
assign detect_max[10][25] = (mid_1[95:88] > btm_2[103:96]) ? 1 : 0;

assign detect_max[11][0] = (mid_1[103:96] > top_0[95:88]) ? 1 : 0;
assign detect_max[11][1] = (mid_1[103:96] > top_0[103:96]) ? 1 : 0;
assign detect_max[11][2] = (mid_1[103:96] > top_0[111:104]) ? 1 : 0;
assign detect_max[11][3] = (mid_1[103:96] > top_1[95:88]) ? 1 : 0;
assign detect_max[11][4] = (mid_1[103:96] > top_1[103:96]) ? 1 : 0;
assign detect_max[11][5] = (mid_1[103:96] > top_1[111:104]) ? 1 : 0;
assign detect_max[11][6] = (mid_1[103:96] > top_2[95:88]) ? 1 : 0;
assign detect_max[11][7] = (mid_1[103:96] > top_2[103:96]) ? 1 : 0;
assign detect_max[11][8] = (mid_1[103:96] > top_2[111:104]) ? 1 : 0;
assign detect_max[11][9] = (mid_1[103:96] > mid_0[95:88]) ? 1 : 0;
assign detect_max[11][10] = (mid_1[103:96] > mid_0[103:96]) ? 1 : 0;
assign detect_max[11][11] = (mid_1[103:96] > mid_0[111:104]) ? 1 : 0;
assign detect_max[11][12] = (mid_1[103:96] > mid_1[95:88]) ? 1 : 0;
assign detect_max[11][13] = (mid_1[103:96] > mid_1[111:104]) ? 1 : 0;
assign detect_max[11][14] = (mid_1[103:96] > mid_2[95:88]) ? 1 : 0;
assign detect_max[11][15] = (mid_1[103:96] > mid_2[103:96]) ? 1 : 0;
assign detect_max[11][16] = (mid_1[103:96] > mid_2[111:104]) ? 1 : 0;
assign detect_max[11][17] = (mid_1[103:96] > btm_0[95:88]) ? 1 : 0;
assign detect_max[11][18] = (mid_1[103:96] > btm_0[103:96]) ? 1 : 0;
assign detect_max[11][19] = (mid_1[103:96] > btm_0[111:104]) ? 1 : 0;
assign detect_max[11][20] = (mid_1[103:96] > btm_1[95:88]) ? 1 : 0;
assign detect_max[11][21] = (mid_1[103:96] > btm_1[103:96]) ? 1 : 0;
assign detect_max[11][22] = (mid_1[103:96] > btm_1[111:104]) ? 1 : 0;
assign detect_max[11][23] = (mid_1[103:96] > btm_2[95:88]) ? 1 : 0;
assign detect_max[11][24] = (mid_1[103:96] > btm_2[103:96]) ? 1 : 0;
assign detect_max[11][25] = (mid_1[103:96] > btm_2[111:104]) ? 1 : 0;

assign detect_max[12][0] = (mid_1[111:104] > top_0[103:96]) ? 1 : 0;
assign detect_max[12][1] = (mid_1[111:104] > top_0[111:104]) ? 1 : 0;
assign detect_max[12][2] = (mid_1[111:104] > top_0[119:112]) ? 1 : 0;
assign detect_max[12][3] = (mid_1[111:104] > top_1[103:96]) ? 1 : 0;
assign detect_max[12][4] = (mid_1[111:104] > top_1[111:104]) ? 1 : 0;
assign detect_max[12][5] = (mid_1[111:104] > top_1[119:112]) ? 1 : 0;
assign detect_max[12][6] = (mid_1[111:104] > top_2[103:96]) ? 1 : 0;
assign detect_max[12][7] = (mid_1[111:104] > top_2[111:104]) ? 1 : 0;
assign detect_max[12][8] = (mid_1[111:104] > top_2[119:112]) ? 1 : 0;
assign detect_max[12][9] = (mid_1[111:104] > mid_0[103:96]) ? 1 : 0;
assign detect_max[12][10] = (mid_1[111:104] > mid_0[111:104]) ? 1 : 0;
assign detect_max[12][11] = (mid_1[111:104] > mid_0[119:112]) ? 1 : 0;
assign detect_max[12][12] = (mid_1[111:104] > mid_1[103:96]) ? 1 : 0;
assign detect_max[12][13] = (mid_1[111:104] > mid_1[119:112]) ? 1 : 0;
assign detect_max[12][14] = (mid_1[111:104] > mid_2[103:96]) ? 1 : 0;
assign detect_max[12][15] = (mid_1[111:104] > mid_2[111:104]) ? 1 : 0;
assign detect_max[12][16] = (mid_1[111:104] > mid_2[119:112]) ? 1 : 0;
assign detect_max[12][17] = (mid_1[111:104] > btm_0[103:96]) ? 1 : 0;
assign detect_max[12][18] = (mid_1[111:104] > btm_0[111:104]) ? 1 : 0;
assign detect_max[12][19] = (mid_1[111:104] > btm_0[119:112]) ? 1 : 0;
assign detect_max[12][20] = (mid_1[111:104] > btm_1[103:96]) ? 1 : 0;
assign detect_max[12][21] = (mid_1[111:104] > btm_1[111:104]) ? 1 : 0;
assign detect_max[12][22] = (mid_1[111:104] > btm_1[119:112]) ? 1 : 0;
assign detect_max[12][23] = (mid_1[111:104] > btm_2[103:96]) ? 1 : 0;
assign detect_max[12][24] = (mid_1[111:104] > btm_2[111:104]) ? 1 : 0;
assign detect_max[12][25] = (mid_1[111:104] > btm_2[119:112]) ? 1 : 0;

assign detect_max[13][0] = (mid_1[119:112] > top_0[111:104]) ? 1 : 0;
assign detect_max[13][1] = (mid_1[119:112] > top_0[119:112]) ? 1 : 0;
assign detect_max[13][2] = (mid_1[119:112] > top_0[127:120]) ? 1 : 0;
assign detect_max[13][3] = (mid_1[119:112] > top_1[111:104]) ? 1 : 0;
assign detect_max[13][4] = (mid_1[119:112] > top_1[119:112]) ? 1 : 0;
assign detect_max[13][5] = (mid_1[119:112] > top_1[127:120]) ? 1 : 0;
assign detect_max[13][6] = (mid_1[119:112] > top_2[111:104]) ? 1 : 0;
assign detect_max[13][7] = (mid_1[119:112] > top_2[119:112]) ? 1 : 0;
assign detect_max[13][8] = (mid_1[119:112] > top_2[127:120]) ? 1 : 0;
assign detect_max[13][9] = (mid_1[119:112] > mid_0[111:104]) ? 1 : 0;
assign detect_max[13][10] = (mid_1[119:112] > mid_0[119:112]) ? 1 : 0;
assign detect_max[13][11] = (mid_1[119:112] > mid_0[127:120]) ? 1 : 0;
assign detect_max[13][12] = (mid_1[119:112] > mid_1[111:104]) ? 1 : 0;
assign detect_max[13][13] = (mid_1[119:112] > mid_1[127:120]) ? 1 : 0;
assign detect_max[13][14] = (mid_1[119:112] > mid_2[111:104]) ? 1 : 0;
assign detect_max[13][15] = (mid_1[119:112] > mid_2[119:112]) ? 1 : 0;
assign detect_max[13][16] = (mid_1[119:112] > mid_2[127:120]) ? 1 : 0;
assign detect_max[13][17] = (mid_1[119:112] > btm_0[111:104]) ? 1 : 0;
assign detect_max[13][18] = (mid_1[119:112] > btm_0[119:112]) ? 1 : 0;
assign detect_max[13][19] = (mid_1[119:112] > btm_0[127:120]) ? 1 : 0;
assign detect_max[13][20] = (mid_1[119:112] > btm_1[111:104]) ? 1 : 0;
assign detect_max[13][21] = (mid_1[119:112] > btm_1[119:112]) ? 1 : 0;
assign detect_max[13][22] = (mid_1[119:112] > btm_1[127:120]) ? 1 : 0;
assign detect_max[13][23] = (mid_1[119:112] > btm_2[111:104]) ? 1 : 0;
assign detect_max[13][24] = (mid_1[119:112] > btm_2[119:112]) ? 1 : 0;
assign detect_max[13][25] = (mid_1[119:112] > btm_2[127:120]) ? 1 : 0;

assign detect_max[14][0] = (mid_1[127:120] > top_0[119:112]) ? 1 : 0;
assign detect_max[14][1] = (mid_1[127:120] > top_0[127:120]) ? 1 : 0;
assign detect_max[14][2] = (mid_1[127:120] > top_0[135:128]) ? 1 : 0;
assign detect_max[14][3] = (mid_1[127:120] > top_1[119:112]) ? 1 : 0;
assign detect_max[14][4] = (mid_1[127:120] > top_1[127:120]) ? 1 : 0;
assign detect_max[14][5] = (mid_1[127:120] > top_1[135:128]) ? 1 : 0;
assign detect_max[14][6] = (mid_1[127:120] > top_2[119:112]) ? 1 : 0;
assign detect_max[14][7] = (mid_1[127:120] > top_2[127:120]) ? 1 : 0;
assign detect_max[14][8] = (mid_1[127:120] > top_2[135:128]) ? 1 : 0;
assign detect_max[14][9] = (mid_1[127:120] > mid_0[119:112]) ? 1 : 0;
assign detect_max[14][10] = (mid_1[127:120] > mid_0[127:120]) ? 1 : 0;
assign detect_max[14][11] = (mid_1[127:120] > mid_0[135:128]) ? 1 : 0;
assign detect_max[14][12] = (mid_1[127:120] > mid_1[119:112]) ? 1 : 0;
assign detect_max[14][13] = (mid_1[127:120] > mid_1[135:128]) ? 1 : 0;
assign detect_max[14][14] = (mid_1[127:120] > mid_2[119:112]) ? 1 : 0;
assign detect_max[14][15] = (mid_1[127:120] > mid_2[127:120]) ? 1 : 0;
assign detect_max[14][16] = (mid_1[127:120] > mid_2[135:128]) ? 1 : 0;
assign detect_max[14][17] = (mid_1[127:120] > btm_0[119:112]) ? 1 : 0;
assign detect_max[14][18] = (mid_1[127:120] > btm_0[127:120]) ? 1 : 0;
assign detect_max[14][19] = (mid_1[127:120] > btm_0[135:128]) ? 1 : 0;
assign detect_max[14][20] = (mid_1[127:120] > btm_1[119:112]) ? 1 : 0;
assign detect_max[14][21] = (mid_1[127:120] > btm_1[127:120]) ? 1 : 0;
assign detect_max[14][22] = (mid_1[127:120] > btm_1[135:128]) ? 1 : 0;
assign detect_max[14][23] = (mid_1[127:120] > btm_2[119:112]) ? 1 : 0;
assign detect_max[14][24] = (mid_1[127:120] > btm_2[127:120]) ? 1 : 0;
assign detect_max[14][25] = (mid_1[127:120] > btm_2[135:128]) ? 1 : 0;

assign detect_max[15][0] = (mid_1[135:128] > top_0[127:120]) ? 1 : 0;
assign detect_max[15][1] = (mid_1[135:128] > top_0[135:128]) ? 1 : 0;
assign detect_max[15][2] = (mid_1[135:128] > top_0[143:136]) ? 1 : 0;
assign detect_max[15][3] = (mid_1[135:128] > top_1[127:120]) ? 1 : 0;
assign detect_max[15][4] = (mid_1[135:128] > top_1[135:128]) ? 1 : 0;
assign detect_max[15][5] = (mid_1[135:128] > top_1[143:136]) ? 1 : 0;
assign detect_max[15][6] = (mid_1[135:128] > top_2[127:120]) ? 1 : 0;
assign detect_max[15][7] = (mid_1[135:128] > top_2[135:128]) ? 1 : 0;
assign detect_max[15][8] = (mid_1[135:128] > top_2[143:136]) ? 1 : 0;
assign detect_max[15][9] = (mid_1[135:128] > mid_0[127:120]) ? 1 : 0;
assign detect_max[15][10] = (mid_1[135:128] > mid_0[135:128]) ? 1 : 0;
assign detect_max[15][11] = (mid_1[135:128] > mid_0[143:136]) ? 1 : 0;
assign detect_max[15][12] = (mid_1[135:128] > mid_1[127:120]) ? 1 : 0;
assign detect_max[15][13] = (mid_1[135:128] > mid_1[143:136]) ? 1 : 0;
assign detect_max[15][14] = (mid_1[135:128] > mid_2[127:120]) ? 1 : 0;
assign detect_max[15][15] = (mid_1[135:128] > mid_2[135:128]) ? 1 : 0;
assign detect_max[15][16] = (mid_1[135:128] > mid_2[143:136]) ? 1 : 0;
assign detect_max[15][17] = (mid_1[135:128] > btm_0[127:120]) ? 1 : 0;
assign detect_max[15][18] = (mid_1[135:128] > btm_0[135:128]) ? 1 : 0;
assign detect_max[15][19] = (mid_1[135:128] > btm_0[143:136]) ? 1 : 0;
assign detect_max[15][20] = (mid_1[135:128] > btm_1[127:120]) ? 1 : 0;
assign detect_max[15][21] = (mid_1[135:128] > btm_1[135:128]) ? 1 : 0;
assign detect_max[15][22] = (mid_1[135:128] > btm_1[143:136]) ? 1 : 0;
assign detect_max[15][23] = (mid_1[135:128] > btm_2[127:120]) ? 1 : 0;
assign detect_max[15][24] = (mid_1[135:128] > btm_2[135:128]) ? 1 : 0;
assign detect_max[15][25] = (mid_1[135:128] > btm_2[143:136]) ? 1 : 0;

assign detect_max[16][0] = (mid_1[143:136] > top_0[135:128]) ? 1 : 0;
assign detect_max[16][1] = (mid_1[143:136] > top_0[143:136]) ? 1 : 0;
assign detect_max[16][2] = (mid_1[143:136] > top_0[151:144]) ? 1 : 0;
assign detect_max[16][3] = (mid_1[143:136] > top_1[135:128]) ? 1 : 0;
assign detect_max[16][4] = (mid_1[143:136] > top_1[143:136]) ? 1 : 0;
assign detect_max[16][5] = (mid_1[143:136] > top_1[151:144]) ? 1 : 0;
assign detect_max[16][6] = (mid_1[143:136] > top_2[135:128]) ? 1 : 0;
assign detect_max[16][7] = (mid_1[143:136] > top_2[143:136]) ? 1 : 0;
assign detect_max[16][8] = (mid_1[143:136] > top_2[151:144]) ? 1 : 0;
assign detect_max[16][9] = (mid_1[143:136] > mid_0[135:128]) ? 1 : 0;
assign detect_max[16][10] = (mid_1[143:136] > mid_0[143:136]) ? 1 : 0;
assign detect_max[16][11] = (mid_1[143:136] > mid_0[151:144]) ? 1 : 0;
assign detect_max[16][12] = (mid_1[143:136] > mid_1[135:128]) ? 1 : 0;
assign detect_max[16][13] = (mid_1[143:136] > mid_1[151:144]) ? 1 : 0;
assign detect_max[16][14] = (mid_1[143:136] > mid_2[135:128]) ? 1 : 0;
assign detect_max[16][15] = (mid_1[143:136] > mid_2[143:136]) ? 1 : 0;
assign detect_max[16][16] = (mid_1[143:136] > mid_2[151:144]) ? 1 : 0;
assign detect_max[16][17] = (mid_1[143:136] > btm_0[135:128]) ? 1 : 0;
assign detect_max[16][18] = (mid_1[143:136] > btm_0[143:136]) ? 1 : 0;
assign detect_max[16][19] = (mid_1[143:136] > btm_0[151:144]) ? 1 : 0;
assign detect_max[16][20] = (mid_1[143:136] > btm_1[135:128]) ? 1 : 0;
assign detect_max[16][21] = (mid_1[143:136] > btm_1[143:136]) ? 1 : 0;
assign detect_max[16][22] = (mid_1[143:136] > btm_1[151:144]) ? 1 : 0;
assign detect_max[16][23] = (mid_1[143:136] > btm_2[135:128]) ? 1 : 0;
assign detect_max[16][24] = (mid_1[143:136] > btm_2[143:136]) ? 1 : 0;
assign detect_max[16][25] = (mid_1[143:136] > btm_2[151:144]) ? 1 : 0;

assign detect_max[17][0] = (mid_1[151:144] > top_0[143:136]) ? 1 : 0;
assign detect_max[17][1] = (mid_1[151:144] > top_0[151:144]) ? 1 : 0;
assign detect_max[17][2] = (mid_1[151:144] > top_0[159:152]) ? 1 : 0;
assign detect_max[17][3] = (mid_1[151:144] > top_1[143:136]) ? 1 : 0;
assign detect_max[17][4] = (mid_1[151:144] > top_1[151:144]) ? 1 : 0;
assign detect_max[17][5] = (mid_1[151:144] > top_1[159:152]) ? 1 : 0;
assign detect_max[17][6] = (mid_1[151:144] > top_2[143:136]) ? 1 : 0;
assign detect_max[17][7] = (mid_1[151:144] > top_2[151:144]) ? 1 : 0;
assign detect_max[17][8] = (mid_1[151:144] > top_2[159:152]) ? 1 : 0;
assign detect_max[17][9] = (mid_1[151:144] > mid_0[143:136]) ? 1 : 0;
assign detect_max[17][10] = (mid_1[151:144] > mid_0[151:144]) ? 1 : 0;
assign detect_max[17][11] = (mid_1[151:144] > mid_0[159:152]) ? 1 : 0;
assign detect_max[17][12] = (mid_1[151:144] > mid_1[143:136]) ? 1 : 0;
assign detect_max[17][13] = (mid_1[151:144] > mid_1[159:152]) ? 1 : 0;
assign detect_max[17][14] = (mid_1[151:144] > mid_2[143:136]) ? 1 : 0;
assign detect_max[17][15] = (mid_1[151:144] > mid_2[151:144]) ? 1 : 0;
assign detect_max[17][16] = (mid_1[151:144] > mid_2[159:152]) ? 1 : 0;
assign detect_max[17][17] = (mid_1[151:144] > btm_0[143:136]) ? 1 : 0;
assign detect_max[17][18] = (mid_1[151:144] > btm_0[151:144]) ? 1 : 0;
assign detect_max[17][19] = (mid_1[151:144] > btm_0[159:152]) ? 1 : 0;
assign detect_max[17][20] = (mid_1[151:144] > btm_1[143:136]) ? 1 : 0;
assign detect_max[17][21] = (mid_1[151:144] > btm_1[151:144]) ? 1 : 0;
assign detect_max[17][22] = (mid_1[151:144] > btm_1[159:152]) ? 1 : 0;
assign detect_max[17][23] = (mid_1[151:144] > btm_2[143:136]) ? 1 : 0;
assign detect_max[17][24] = (mid_1[151:144] > btm_2[151:144]) ? 1 : 0;
assign detect_max[17][25] = (mid_1[151:144] > btm_2[159:152]) ? 1 : 0;

assign detect_max[18][0] = (mid_1[159:152] > top_0[151:144]) ? 1 : 0;
assign detect_max[18][1] = (mid_1[159:152] > top_0[159:152]) ? 1 : 0;
assign detect_max[18][2] = (mid_1[159:152] > top_0[167:160]) ? 1 : 0;
assign detect_max[18][3] = (mid_1[159:152] > top_1[151:144]) ? 1 : 0;
assign detect_max[18][4] = (mid_1[159:152] > top_1[159:152]) ? 1 : 0;
assign detect_max[18][5] = (mid_1[159:152] > top_1[167:160]) ? 1 : 0;
assign detect_max[18][6] = (mid_1[159:152] > top_2[151:144]) ? 1 : 0;
assign detect_max[18][7] = (mid_1[159:152] > top_2[159:152]) ? 1 : 0;
assign detect_max[18][8] = (mid_1[159:152] > top_2[167:160]) ? 1 : 0;
assign detect_max[18][9] = (mid_1[159:152] > mid_0[151:144]) ? 1 : 0;
assign detect_max[18][10] = (mid_1[159:152] > mid_0[159:152]) ? 1 : 0;
assign detect_max[18][11] = (mid_1[159:152] > mid_0[167:160]) ? 1 : 0;
assign detect_max[18][12] = (mid_1[159:152] > mid_1[151:144]) ? 1 : 0;
assign detect_max[18][13] = (mid_1[159:152] > mid_1[167:160]) ? 1 : 0;
assign detect_max[18][14] = (mid_1[159:152] > mid_2[151:144]) ? 1 : 0;
assign detect_max[18][15] = (mid_1[159:152] > mid_2[159:152]) ? 1 : 0;
assign detect_max[18][16] = (mid_1[159:152] > mid_2[167:160]) ? 1 : 0;
assign detect_max[18][17] = (mid_1[159:152] > btm_0[151:144]) ? 1 : 0;
assign detect_max[18][18] = (mid_1[159:152] > btm_0[159:152]) ? 1 : 0;
assign detect_max[18][19] = (mid_1[159:152] > btm_0[167:160]) ? 1 : 0;
assign detect_max[18][20] = (mid_1[159:152] > btm_1[151:144]) ? 1 : 0;
assign detect_max[18][21] = (mid_1[159:152] > btm_1[159:152]) ? 1 : 0;
assign detect_max[18][22] = (mid_1[159:152] > btm_1[167:160]) ? 1 : 0;
assign detect_max[18][23] = (mid_1[159:152] > btm_2[151:144]) ? 1 : 0;
assign detect_max[18][24] = (mid_1[159:152] > btm_2[159:152]) ? 1 : 0;
assign detect_max[18][25] = (mid_1[159:152] > btm_2[167:160]) ? 1 : 0;

assign detect_max[19][0] = (mid_1[167:160] > top_0[159:152]) ? 1 : 0;
assign detect_max[19][1] = (mid_1[167:160] > top_0[167:160]) ? 1 : 0;
assign detect_max[19][2] = (mid_1[167:160] > top_0[175:168]) ? 1 : 0;
assign detect_max[19][3] = (mid_1[167:160] > top_1[159:152]) ? 1 : 0;
assign detect_max[19][4] = (mid_1[167:160] > top_1[167:160]) ? 1 : 0;
assign detect_max[19][5] = (mid_1[167:160] > top_1[175:168]) ? 1 : 0;
assign detect_max[19][6] = (mid_1[167:160] > top_2[159:152]) ? 1 : 0;
assign detect_max[19][7] = (mid_1[167:160] > top_2[167:160]) ? 1 : 0;
assign detect_max[19][8] = (mid_1[167:160] > top_2[175:168]) ? 1 : 0;
assign detect_max[19][9] = (mid_1[167:160] > mid_0[159:152]) ? 1 : 0;
assign detect_max[19][10] = (mid_1[167:160] > mid_0[167:160]) ? 1 : 0;
assign detect_max[19][11] = (mid_1[167:160] > mid_0[175:168]) ? 1 : 0;
assign detect_max[19][12] = (mid_1[167:160] > mid_1[159:152]) ? 1 : 0;
assign detect_max[19][13] = (mid_1[167:160] > mid_1[175:168]) ? 1 : 0;
assign detect_max[19][14] = (mid_1[167:160] > mid_2[159:152]) ? 1 : 0;
assign detect_max[19][15] = (mid_1[167:160] > mid_2[167:160]) ? 1 : 0;
assign detect_max[19][16] = (mid_1[167:160] > mid_2[175:168]) ? 1 : 0;
assign detect_max[19][17] = (mid_1[167:160] > btm_0[159:152]) ? 1 : 0;
assign detect_max[19][18] = (mid_1[167:160] > btm_0[167:160]) ? 1 : 0;
assign detect_max[19][19] = (mid_1[167:160] > btm_0[175:168]) ? 1 : 0;
assign detect_max[19][20] = (mid_1[167:160] > btm_1[159:152]) ? 1 : 0;
assign detect_max[19][21] = (mid_1[167:160] > btm_1[167:160]) ? 1 : 0;
assign detect_max[19][22] = (mid_1[167:160] > btm_1[175:168]) ? 1 : 0;
assign detect_max[19][23] = (mid_1[167:160] > btm_2[159:152]) ? 1 : 0;
assign detect_max[19][24] = (mid_1[167:160] > btm_2[167:160]) ? 1 : 0;
assign detect_max[19][25] = (mid_1[167:160] > btm_2[175:168]) ? 1 : 0;

assign detect_max[20][0] = (mid_1[175:168] > top_0[167:160]) ? 1 : 0;
assign detect_max[20][1] = (mid_1[175:168] > top_0[175:168]) ? 1 : 0;
assign detect_max[20][2] = (mid_1[175:168] > top_0[183:176]) ? 1 : 0;
assign detect_max[20][3] = (mid_1[175:168] > top_1[167:160]) ? 1 : 0;
assign detect_max[20][4] = (mid_1[175:168] > top_1[175:168]) ? 1 : 0;
assign detect_max[20][5] = (mid_1[175:168] > top_1[183:176]) ? 1 : 0;
assign detect_max[20][6] = (mid_1[175:168] > top_2[167:160]) ? 1 : 0;
assign detect_max[20][7] = (mid_1[175:168] > top_2[175:168]) ? 1 : 0;
assign detect_max[20][8] = (mid_1[175:168] > top_2[183:176]) ? 1 : 0;
assign detect_max[20][9] = (mid_1[175:168] > mid_0[167:160]) ? 1 : 0;
assign detect_max[20][10] = (mid_1[175:168] > mid_0[175:168]) ? 1 : 0;
assign detect_max[20][11] = (mid_1[175:168] > mid_0[183:176]) ? 1 : 0;
assign detect_max[20][12] = (mid_1[175:168] > mid_1[167:160]) ? 1 : 0;
assign detect_max[20][13] = (mid_1[175:168] > mid_1[183:176]) ? 1 : 0;
assign detect_max[20][14] = (mid_1[175:168] > mid_2[167:160]) ? 1 : 0;
assign detect_max[20][15] = (mid_1[175:168] > mid_2[175:168]) ? 1 : 0;
assign detect_max[20][16] = (mid_1[175:168] > mid_2[183:176]) ? 1 : 0;
assign detect_max[20][17] = (mid_1[175:168] > btm_0[167:160]) ? 1 : 0;
assign detect_max[20][18] = (mid_1[175:168] > btm_0[175:168]) ? 1 : 0;
assign detect_max[20][19] = (mid_1[175:168] > btm_0[183:176]) ? 1 : 0;
assign detect_max[20][20] = (mid_1[175:168] > btm_1[167:160]) ? 1 : 0;
assign detect_max[20][21] = (mid_1[175:168] > btm_1[175:168]) ? 1 : 0;
assign detect_max[20][22] = (mid_1[175:168] > btm_1[183:176]) ? 1 : 0;
assign detect_max[20][23] = (mid_1[175:168] > btm_2[167:160]) ? 1 : 0;
assign detect_max[20][24] = (mid_1[175:168] > btm_2[175:168]) ? 1 : 0;
assign detect_max[20][25] = (mid_1[175:168] > btm_2[183:176]) ? 1 : 0;

assign detect_max[21][0] = (mid_1[183:176] > top_0[175:168]) ? 1 : 0;
assign detect_max[21][1] = (mid_1[183:176] > top_0[183:176]) ? 1 : 0;
assign detect_max[21][2] = (mid_1[183:176] > top_0[191:184]) ? 1 : 0;
assign detect_max[21][3] = (mid_1[183:176] > top_1[175:168]) ? 1 : 0;
assign detect_max[21][4] = (mid_1[183:176] > top_1[183:176]) ? 1 : 0;
assign detect_max[21][5] = (mid_1[183:176] > top_1[191:184]) ? 1 : 0;
assign detect_max[21][6] = (mid_1[183:176] > top_2[175:168]) ? 1 : 0;
assign detect_max[21][7] = (mid_1[183:176] > top_2[183:176]) ? 1 : 0;
assign detect_max[21][8] = (mid_1[183:176] > top_2[191:184]) ? 1 : 0;
assign detect_max[21][9] = (mid_1[183:176] > mid_0[175:168]) ? 1 : 0;
assign detect_max[21][10] = (mid_1[183:176] > mid_0[183:176]) ? 1 : 0;
assign detect_max[21][11] = (mid_1[183:176] > mid_0[191:184]) ? 1 : 0;
assign detect_max[21][12] = (mid_1[183:176] > mid_1[175:168]) ? 1 : 0;
assign detect_max[21][13] = (mid_1[183:176] > mid_1[191:184]) ? 1 : 0;
assign detect_max[21][14] = (mid_1[183:176] > mid_2[175:168]) ? 1 : 0;
assign detect_max[21][15] = (mid_1[183:176] > mid_2[183:176]) ? 1 : 0;
assign detect_max[21][16] = (mid_1[183:176] > mid_2[191:184]) ? 1 : 0;
assign detect_max[21][17] = (mid_1[183:176] > btm_0[175:168]) ? 1 : 0;
assign detect_max[21][18] = (mid_1[183:176] > btm_0[183:176]) ? 1 : 0;
assign detect_max[21][19] = (mid_1[183:176] > btm_0[191:184]) ? 1 : 0;
assign detect_max[21][20] = (mid_1[183:176] > btm_1[175:168]) ? 1 : 0;
assign detect_max[21][21] = (mid_1[183:176] > btm_1[183:176]) ? 1 : 0;
assign detect_max[21][22] = (mid_1[183:176] > btm_1[191:184]) ? 1 : 0;
assign detect_max[21][23] = (mid_1[183:176] > btm_2[175:168]) ? 1 : 0;
assign detect_max[21][24] = (mid_1[183:176] > btm_2[183:176]) ? 1 : 0;
assign detect_max[21][25] = (mid_1[183:176] > btm_2[191:184]) ? 1 : 0;

assign detect_max[22][0] = (mid_1[191:184] > top_0[183:176]) ? 1 : 0;
assign detect_max[22][1] = (mid_1[191:184] > top_0[191:184]) ? 1 : 0;
assign detect_max[22][2] = (mid_1[191:184] > top_0[199:192]) ? 1 : 0;
assign detect_max[22][3] = (mid_1[191:184] > top_1[183:176]) ? 1 : 0;
assign detect_max[22][4] = (mid_1[191:184] > top_1[191:184]) ? 1 : 0;
assign detect_max[22][5] = (mid_1[191:184] > top_1[199:192]) ? 1 : 0;
assign detect_max[22][6] = (mid_1[191:184] > top_2[183:176]) ? 1 : 0;
assign detect_max[22][7] = (mid_1[191:184] > top_2[191:184]) ? 1 : 0;
assign detect_max[22][8] = (mid_1[191:184] > top_2[199:192]) ? 1 : 0;
assign detect_max[22][9] = (mid_1[191:184] > mid_0[183:176]) ? 1 : 0;
assign detect_max[22][10] = (mid_1[191:184] > mid_0[191:184]) ? 1 : 0;
assign detect_max[22][11] = (mid_1[191:184] > mid_0[199:192]) ? 1 : 0;
assign detect_max[22][12] = (mid_1[191:184] > mid_1[183:176]) ? 1 : 0;
assign detect_max[22][13] = (mid_1[191:184] > mid_1[199:192]) ? 1 : 0;
assign detect_max[22][14] = (mid_1[191:184] > mid_2[183:176]) ? 1 : 0;
assign detect_max[22][15] = (mid_1[191:184] > mid_2[191:184]) ? 1 : 0;
assign detect_max[22][16] = (mid_1[191:184] > mid_2[199:192]) ? 1 : 0;
assign detect_max[22][17] = (mid_1[191:184] > btm_0[183:176]) ? 1 : 0;
assign detect_max[22][18] = (mid_1[191:184] > btm_0[191:184]) ? 1 : 0;
assign detect_max[22][19] = (mid_1[191:184] > btm_0[199:192]) ? 1 : 0;
assign detect_max[22][20] = (mid_1[191:184] > btm_1[183:176]) ? 1 : 0;
assign detect_max[22][21] = (mid_1[191:184] > btm_1[191:184]) ? 1 : 0;
assign detect_max[22][22] = (mid_1[191:184] > btm_1[199:192]) ? 1 : 0;
assign detect_max[22][23] = (mid_1[191:184] > btm_2[183:176]) ? 1 : 0;
assign detect_max[22][24] = (mid_1[191:184] > btm_2[191:184]) ? 1 : 0;
assign detect_max[22][25] = (mid_1[191:184] > btm_2[199:192]) ? 1 : 0;

assign detect_max[23][0] = (mid_1[199:192] > top_0[191:184]) ? 1 : 0;
assign detect_max[23][1] = (mid_1[199:192] > top_0[199:192]) ? 1 : 0;
assign detect_max[23][2] = (mid_1[199:192] > top_0[207:200]) ? 1 : 0;
assign detect_max[23][3] = (mid_1[199:192] > top_1[191:184]) ? 1 : 0;
assign detect_max[23][4] = (mid_1[199:192] > top_1[199:192]) ? 1 : 0;
assign detect_max[23][5] = (mid_1[199:192] > top_1[207:200]) ? 1 : 0;
assign detect_max[23][6] = (mid_1[199:192] > top_2[191:184]) ? 1 : 0;
assign detect_max[23][7] = (mid_1[199:192] > top_2[199:192]) ? 1 : 0;
assign detect_max[23][8] = (mid_1[199:192] > top_2[207:200]) ? 1 : 0;
assign detect_max[23][9] = (mid_1[199:192] > mid_0[191:184]) ? 1 : 0;
assign detect_max[23][10] = (mid_1[199:192] > mid_0[199:192]) ? 1 : 0;
assign detect_max[23][11] = (mid_1[199:192] > mid_0[207:200]) ? 1 : 0;
assign detect_max[23][12] = (mid_1[199:192] > mid_1[191:184]) ? 1 : 0;
assign detect_max[23][13] = (mid_1[199:192] > mid_1[207:200]) ? 1 : 0;
assign detect_max[23][14] = (mid_1[199:192] > mid_2[191:184]) ? 1 : 0;
assign detect_max[23][15] = (mid_1[199:192] > mid_2[199:192]) ? 1 : 0;
assign detect_max[23][16] = (mid_1[199:192] > mid_2[207:200]) ? 1 : 0;
assign detect_max[23][17] = (mid_1[199:192] > btm_0[191:184]) ? 1 : 0;
assign detect_max[23][18] = (mid_1[199:192] > btm_0[199:192]) ? 1 : 0;
assign detect_max[23][19] = (mid_1[199:192] > btm_0[207:200]) ? 1 : 0;
assign detect_max[23][20] = (mid_1[199:192] > btm_1[191:184]) ? 1 : 0;
assign detect_max[23][21] = (mid_1[199:192] > btm_1[199:192]) ? 1 : 0;
assign detect_max[23][22] = (mid_1[199:192] > btm_1[207:200]) ? 1 : 0;
assign detect_max[23][23] = (mid_1[199:192] > btm_2[191:184]) ? 1 : 0;
assign detect_max[23][24] = (mid_1[199:192] > btm_2[199:192]) ? 1 : 0;
assign detect_max[23][25] = (mid_1[199:192] > btm_2[207:200]) ? 1 : 0;

assign detect_max[24][0] = (mid_1[207:200] > top_0[199:192]) ? 1 : 0;
assign detect_max[24][1] = (mid_1[207:200] > top_0[207:200]) ? 1 : 0;
assign detect_max[24][2] = (mid_1[207:200] > top_0[215:208]) ? 1 : 0;
assign detect_max[24][3] = (mid_1[207:200] > top_1[199:192]) ? 1 : 0;
assign detect_max[24][4] = (mid_1[207:200] > top_1[207:200]) ? 1 : 0;
assign detect_max[24][5] = (mid_1[207:200] > top_1[215:208]) ? 1 : 0;
assign detect_max[24][6] = (mid_1[207:200] > top_2[199:192]) ? 1 : 0;
assign detect_max[24][7] = (mid_1[207:200] > top_2[207:200]) ? 1 : 0;
assign detect_max[24][8] = (mid_1[207:200] > top_2[215:208]) ? 1 : 0;
assign detect_max[24][9] = (mid_1[207:200] > mid_0[199:192]) ? 1 : 0;
assign detect_max[24][10] = (mid_1[207:200] > mid_0[207:200]) ? 1 : 0;
assign detect_max[24][11] = (mid_1[207:200] > mid_0[215:208]) ? 1 : 0;
assign detect_max[24][12] = (mid_1[207:200] > mid_1[199:192]) ? 1 : 0;
assign detect_max[24][13] = (mid_1[207:200] > mid_1[215:208]) ? 1 : 0;
assign detect_max[24][14] = (mid_1[207:200] > mid_2[199:192]) ? 1 : 0;
assign detect_max[24][15] = (mid_1[207:200] > mid_2[207:200]) ? 1 : 0;
assign detect_max[24][16] = (mid_1[207:200] > mid_2[215:208]) ? 1 : 0;
assign detect_max[24][17] = (mid_1[207:200] > btm_0[199:192]) ? 1 : 0;
assign detect_max[24][18] = (mid_1[207:200] > btm_0[207:200]) ? 1 : 0;
assign detect_max[24][19] = (mid_1[207:200] > btm_0[215:208]) ? 1 : 0;
assign detect_max[24][20] = (mid_1[207:200] > btm_1[199:192]) ? 1 : 0;
assign detect_max[24][21] = (mid_1[207:200] > btm_1[207:200]) ? 1 : 0;
assign detect_max[24][22] = (mid_1[207:200] > btm_1[215:208]) ? 1 : 0;
assign detect_max[24][23] = (mid_1[207:200] > btm_2[199:192]) ? 1 : 0;
assign detect_max[24][24] = (mid_1[207:200] > btm_2[207:200]) ? 1 : 0;
assign detect_max[24][25] = (mid_1[207:200] > btm_2[215:208]) ? 1 : 0;

assign detect_max[25][0] = (mid_1[215:208] > top_0[207:200]) ? 1 : 0;
assign detect_max[25][1] = (mid_1[215:208] > top_0[215:208]) ? 1 : 0;
assign detect_max[25][2] = (mid_1[215:208] > top_0[223:216]) ? 1 : 0;
assign detect_max[25][3] = (mid_1[215:208] > top_1[207:200]) ? 1 : 0;
assign detect_max[25][4] = (mid_1[215:208] > top_1[215:208]) ? 1 : 0;
assign detect_max[25][5] = (mid_1[215:208] > top_1[223:216]) ? 1 : 0;
assign detect_max[25][6] = (mid_1[215:208] > top_2[207:200]) ? 1 : 0;
assign detect_max[25][7] = (mid_1[215:208] > top_2[215:208]) ? 1 : 0;
assign detect_max[25][8] = (mid_1[215:208] > top_2[223:216]) ? 1 : 0;
assign detect_max[25][9] = (mid_1[215:208] > mid_0[207:200]) ? 1 : 0;
assign detect_max[25][10] = (mid_1[215:208] > mid_0[215:208]) ? 1 : 0;
assign detect_max[25][11] = (mid_1[215:208] > mid_0[223:216]) ? 1 : 0;
assign detect_max[25][12] = (mid_1[215:208] > mid_1[207:200]) ? 1 : 0;
assign detect_max[25][13] = (mid_1[215:208] > mid_1[223:216]) ? 1 : 0;
assign detect_max[25][14] = (mid_1[215:208] > mid_2[207:200]) ? 1 : 0;
assign detect_max[25][15] = (mid_1[215:208] > mid_2[215:208]) ? 1 : 0;
assign detect_max[25][16] = (mid_1[215:208] > mid_2[223:216]) ? 1 : 0;
assign detect_max[25][17] = (mid_1[215:208] > btm_0[207:200]) ? 1 : 0;
assign detect_max[25][18] = (mid_1[215:208] > btm_0[215:208]) ? 1 : 0;
assign detect_max[25][19] = (mid_1[215:208] > btm_0[223:216]) ? 1 : 0;
assign detect_max[25][20] = (mid_1[215:208] > btm_1[207:200]) ? 1 : 0;
assign detect_max[25][21] = (mid_1[215:208] > btm_1[215:208]) ? 1 : 0;
assign detect_max[25][22] = (mid_1[215:208] > btm_1[223:216]) ? 1 : 0;
assign detect_max[25][23] = (mid_1[215:208] > btm_2[207:200]) ? 1 : 0;
assign detect_max[25][24] = (mid_1[215:208] > btm_2[215:208]) ? 1 : 0;
assign detect_max[25][25] = (mid_1[215:208] > btm_2[223:216]) ? 1 : 0;

assign detect_max[26][0] = (mid_1[223:216] > top_0[215:208]) ? 1 : 0;
assign detect_max[26][1] = (mid_1[223:216] > top_0[223:216]) ? 1 : 0;
assign detect_max[26][2] = (mid_1[223:216] > top_0[231:224]) ? 1 : 0;
assign detect_max[26][3] = (mid_1[223:216] > top_1[215:208]) ? 1 : 0;
assign detect_max[26][4] = (mid_1[223:216] > top_1[223:216]) ? 1 : 0;
assign detect_max[26][5] = (mid_1[223:216] > top_1[231:224]) ? 1 : 0;
assign detect_max[26][6] = (mid_1[223:216] > top_2[215:208]) ? 1 : 0;
assign detect_max[26][7] = (mid_1[223:216] > top_2[223:216]) ? 1 : 0;
assign detect_max[26][8] = (mid_1[223:216] > top_2[231:224]) ? 1 : 0;
assign detect_max[26][9] = (mid_1[223:216] > mid_0[215:208]) ? 1 : 0;
assign detect_max[26][10] = (mid_1[223:216] > mid_0[223:216]) ? 1 : 0;
assign detect_max[26][11] = (mid_1[223:216] > mid_0[231:224]) ? 1 : 0;
assign detect_max[26][12] = (mid_1[223:216] > mid_1[215:208]) ? 1 : 0;
assign detect_max[26][13] = (mid_1[223:216] > mid_1[231:224]) ? 1 : 0;
assign detect_max[26][14] = (mid_1[223:216] > mid_2[215:208]) ? 1 : 0;
assign detect_max[26][15] = (mid_1[223:216] > mid_2[223:216]) ? 1 : 0;
assign detect_max[26][16] = (mid_1[223:216] > mid_2[231:224]) ? 1 : 0;
assign detect_max[26][17] = (mid_1[223:216] > btm_0[215:208]) ? 1 : 0;
assign detect_max[26][18] = (mid_1[223:216] > btm_0[223:216]) ? 1 : 0;
assign detect_max[26][19] = (mid_1[223:216] > btm_0[231:224]) ? 1 : 0;
assign detect_max[26][20] = (mid_1[223:216] > btm_1[215:208]) ? 1 : 0;
assign detect_max[26][21] = (mid_1[223:216] > btm_1[223:216]) ? 1 : 0;
assign detect_max[26][22] = (mid_1[223:216] > btm_1[231:224]) ? 1 : 0;
assign detect_max[26][23] = (mid_1[223:216] > btm_2[215:208]) ? 1 : 0;
assign detect_max[26][24] = (mid_1[223:216] > btm_2[223:216]) ? 1 : 0;
assign detect_max[26][25] = (mid_1[223:216] > btm_2[231:224]) ? 1 : 0;

assign detect_max[27][0] = (mid_1[231:224] > top_0[223:216]) ? 1 : 0;
assign detect_max[27][1] = (mid_1[231:224] > top_0[231:224]) ? 1 : 0;
assign detect_max[27][2] = (mid_1[231:224] > top_0[239:232]) ? 1 : 0;
assign detect_max[27][3] = (mid_1[231:224] > top_1[223:216]) ? 1 : 0;
assign detect_max[27][4] = (mid_1[231:224] > top_1[231:224]) ? 1 : 0;
assign detect_max[27][5] = (mid_1[231:224] > top_1[239:232]) ? 1 : 0;
assign detect_max[27][6] = (mid_1[231:224] > top_2[223:216]) ? 1 : 0;
assign detect_max[27][7] = (mid_1[231:224] > top_2[231:224]) ? 1 : 0;
assign detect_max[27][8] = (mid_1[231:224] > top_2[239:232]) ? 1 : 0;
assign detect_max[27][9] = (mid_1[231:224] > mid_0[223:216]) ? 1 : 0;
assign detect_max[27][10] = (mid_1[231:224] > mid_0[231:224]) ? 1 : 0;
assign detect_max[27][11] = (mid_1[231:224] > mid_0[239:232]) ? 1 : 0;
assign detect_max[27][12] = (mid_1[231:224] > mid_1[223:216]) ? 1 : 0;
assign detect_max[27][13] = (mid_1[231:224] > mid_1[239:232]) ? 1 : 0;
assign detect_max[27][14] = (mid_1[231:224] > mid_2[223:216]) ? 1 : 0;
assign detect_max[27][15] = (mid_1[231:224] > mid_2[231:224]) ? 1 : 0;
assign detect_max[27][16] = (mid_1[231:224] > mid_2[239:232]) ? 1 : 0;
assign detect_max[27][17] = (mid_1[231:224] > btm_0[223:216]) ? 1 : 0;
assign detect_max[27][18] = (mid_1[231:224] > btm_0[231:224]) ? 1 : 0;
assign detect_max[27][19] = (mid_1[231:224] > btm_0[239:232]) ? 1 : 0;
assign detect_max[27][20] = (mid_1[231:224] > btm_1[223:216]) ? 1 : 0;
assign detect_max[27][21] = (mid_1[231:224] > btm_1[231:224]) ? 1 : 0;
assign detect_max[27][22] = (mid_1[231:224] > btm_1[239:232]) ? 1 : 0;
assign detect_max[27][23] = (mid_1[231:224] > btm_2[223:216]) ? 1 : 0;
assign detect_max[27][24] = (mid_1[231:224] > btm_2[231:224]) ? 1 : 0;
assign detect_max[27][25] = (mid_1[231:224] > btm_2[239:232]) ? 1 : 0;

assign detect_max[28][0] = (mid_1[239:232] > top_0[231:224]) ? 1 : 0;
assign detect_max[28][1] = (mid_1[239:232] > top_0[239:232]) ? 1 : 0;
assign detect_max[28][2] = (mid_1[239:232] > top_0[247:240]) ? 1 : 0;
assign detect_max[28][3] = (mid_1[239:232] > top_1[231:224]) ? 1 : 0;
assign detect_max[28][4] = (mid_1[239:232] > top_1[239:232]) ? 1 : 0;
assign detect_max[28][5] = (mid_1[239:232] > top_1[247:240]) ? 1 : 0;
assign detect_max[28][6] = (mid_1[239:232] > top_2[231:224]) ? 1 : 0;
assign detect_max[28][7] = (mid_1[239:232] > top_2[239:232]) ? 1 : 0;
assign detect_max[28][8] = (mid_1[239:232] > top_2[247:240]) ? 1 : 0;
assign detect_max[28][9] = (mid_1[239:232] > mid_0[231:224]) ? 1 : 0;
assign detect_max[28][10] = (mid_1[239:232] > mid_0[239:232]) ? 1 : 0;
assign detect_max[28][11] = (mid_1[239:232] > mid_0[247:240]) ? 1 : 0;
assign detect_max[28][12] = (mid_1[239:232] > mid_1[231:224]) ? 1 : 0;
assign detect_max[28][13] = (mid_1[239:232] > mid_1[247:240]) ? 1 : 0;
assign detect_max[28][14] = (mid_1[239:232] > mid_2[231:224]) ? 1 : 0;
assign detect_max[28][15] = (mid_1[239:232] > mid_2[239:232]) ? 1 : 0;
assign detect_max[28][16] = (mid_1[239:232] > mid_2[247:240]) ? 1 : 0;
assign detect_max[28][17] = (mid_1[239:232] > btm_0[231:224]) ? 1 : 0;
assign detect_max[28][18] = (mid_1[239:232] > btm_0[239:232]) ? 1 : 0;
assign detect_max[28][19] = (mid_1[239:232] > btm_0[247:240]) ? 1 : 0;
assign detect_max[28][20] = (mid_1[239:232] > btm_1[231:224]) ? 1 : 0;
assign detect_max[28][21] = (mid_1[239:232] > btm_1[239:232]) ? 1 : 0;
assign detect_max[28][22] = (mid_1[239:232] > btm_1[247:240]) ? 1 : 0;
assign detect_max[28][23] = (mid_1[239:232] > btm_2[231:224]) ? 1 : 0;
assign detect_max[28][24] = (mid_1[239:232] > btm_2[239:232]) ? 1 : 0;
assign detect_max[28][25] = (mid_1[239:232] > btm_2[247:240]) ? 1 : 0;

assign detect_max[29][0] = (mid_1[247:240] > top_0[239:232]) ? 1 : 0;
assign detect_max[29][1] = (mid_1[247:240] > top_0[247:240]) ? 1 : 0;
assign detect_max[29][2] = (mid_1[247:240] > top_0[255:248]) ? 1 : 0;
assign detect_max[29][3] = (mid_1[247:240] > top_1[239:232]) ? 1 : 0;
assign detect_max[29][4] = (mid_1[247:240] > top_1[247:240]) ? 1 : 0;
assign detect_max[29][5] = (mid_1[247:240] > top_1[255:248]) ? 1 : 0;
assign detect_max[29][6] = (mid_1[247:240] > top_2[239:232]) ? 1 : 0;
assign detect_max[29][7] = (mid_1[247:240] > top_2[247:240]) ? 1 : 0;
assign detect_max[29][8] = (mid_1[247:240] > top_2[255:248]) ? 1 : 0;
assign detect_max[29][9] = (mid_1[247:240] > mid_0[239:232]) ? 1 : 0;
assign detect_max[29][10] = (mid_1[247:240] > mid_0[247:240]) ? 1 : 0;
assign detect_max[29][11] = (mid_1[247:240] > mid_0[255:248]) ? 1 : 0;
assign detect_max[29][12] = (mid_1[247:240] > mid_1[239:232]) ? 1 : 0;
assign detect_max[29][13] = (mid_1[247:240] > mid_1[255:248]) ? 1 : 0;
assign detect_max[29][14] = (mid_1[247:240] > mid_2[239:232]) ? 1 : 0;
assign detect_max[29][15] = (mid_1[247:240] > mid_2[247:240]) ? 1 : 0;
assign detect_max[29][16] = (mid_1[247:240] > mid_2[255:248]) ? 1 : 0;
assign detect_max[29][17] = (mid_1[247:240] > btm_0[239:232]) ? 1 : 0;
assign detect_max[29][18] = (mid_1[247:240] > btm_0[247:240]) ? 1 : 0;
assign detect_max[29][19] = (mid_1[247:240] > btm_0[255:248]) ? 1 : 0;
assign detect_max[29][20] = (mid_1[247:240] > btm_1[239:232]) ? 1 : 0;
assign detect_max[29][21] = (mid_1[247:240] > btm_1[247:240]) ? 1 : 0;
assign detect_max[29][22] = (mid_1[247:240] > btm_1[255:248]) ? 1 : 0;
assign detect_max[29][23] = (mid_1[247:240] > btm_2[239:232]) ? 1 : 0;
assign detect_max[29][24] = (mid_1[247:240] > btm_2[247:240]) ? 1 : 0;
assign detect_max[29][25] = (mid_1[247:240] > btm_2[255:248]) ? 1 : 0;

assign detect_max[30][0] = (mid_1[255:248] > top_0[247:240]) ? 1 : 0;
assign detect_max[30][1] = (mid_1[255:248] > top_0[255:248]) ? 1 : 0;
assign detect_max[30][2] = (mid_1[255:248] > top_0[263:256]) ? 1 : 0;
assign detect_max[30][3] = (mid_1[255:248] > top_1[247:240]) ? 1 : 0;
assign detect_max[30][4] = (mid_1[255:248] > top_1[255:248]) ? 1 : 0;
assign detect_max[30][5] = (mid_1[255:248] > top_1[263:256]) ? 1 : 0;
assign detect_max[30][6] = (mid_1[255:248] > top_2[247:240]) ? 1 : 0;
assign detect_max[30][7] = (mid_1[255:248] > top_2[255:248]) ? 1 : 0;
assign detect_max[30][8] = (mid_1[255:248] > top_2[263:256]) ? 1 : 0;
assign detect_max[30][9] = (mid_1[255:248] > mid_0[247:240]) ? 1 : 0;
assign detect_max[30][10] = (mid_1[255:248] > mid_0[255:248]) ? 1 : 0;
assign detect_max[30][11] = (mid_1[255:248] > mid_0[263:256]) ? 1 : 0;
assign detect_max[30][12] = (mid_1[255:248] > mid_1[247:240]) ? 1 : 0;
assign detect_max[30][13] = (mid_1[255:248] > mid_1[263:256]) ? 1 : 0;
assign detect_max[30][14] = (mid_1[255:248] > mid_2[247:240]) ? 1 : 0;
assign detect_max[30][15] = (mid_1[255:248] > mid_2[255:248]) ? 1 : 0;
assign detect_max[30][16] = (mid_1[255:248] > mid_2[263:256]) ? 1 : 0;
assign detect_max[30][17] = (mid_1[255:248] > btm_0[247:240]) ? 1 : 0;
assign detect_max[30][18] = (mid_1[255:248] > btm_0[255:248]) ? 1 : 0;
assign detect_max[30][19] = (mid_1[255:248] > btm_0[263:256]) ? 1 : 0;
assign detect_max[30][20] = (mid_1[255:248] > btm_1[247:240]) ? 1 : 0;
assign detect_max[30][21] = (mid_1[255:248] > btm_1[255:248]) ? 1 : 0;
assign detect_max[30][22] = (mid_1[255:248] > btm_1[263:256]) ? 1 : 0;
assign detect_max[30][23] = (mid_1[255:248] > btm_2[247:240]) ? 1 : 0;
assign detect_max[30][24] = (mid_1[255:248] > btm_2[255:248]) ? 1 : 0;
assign detect_max[30][25] = (mid_1[255:248] > btm_2[263:256]) ? 1 : 0;

assign detect_max[31][0] = (mid_1[263:256] > top_0[255:248]) ? 1 : 0;
assign detect_max[31][1] = (mid_1[263:256] > top_0[263:256]) ? 1 : 0;
assign detect_max[31][2] = (mid_1[263:256] > top_0[271:264]) ? 1 : 0;
assign detect_max[31][3] = (mid_1[263:256] > top_1[255:248]) ? 1 : 0;
assign detect_max[31][4] = (mid_1[263:256] > top_1[263:256]) ? 1 : 0;
assign detect_max[31][5] = (mid_1[263:256] > top_1[271:264]) ? 1 : 0;
assign detect_max[31][6] = (mid_1[263:256] > top_2[255:248]) ? 1 : 0;
assign detect_max[31][7] = (mid_1[263:256] > top_2[263:256]) ? 1 : 0;
assign detect_max[31][8] = (mid_1[263:256] > top_2[271:264]) ? 1 : 0;
assign detect_max[31][9] = (mid_1[263:256] > mid_0[255:248]) ? 1 : 0;
assign detect_max[31][10] = (mid_1[263:256] > mid_0[263:256]) ? 1 : 0;
assign detect_max[31][11] = (mid_1[263:256] > mid_0[271:264]) ? 1 : 0;
assign detect_max[31][12] = (mid_1[263:256] > mid_1[255:248]) ? 1 : 0;
assign detect_max[31][13] = (mid_1[263:256] > mid_1[271:264]) ? 1 : 0;
assign detect_max[31][14] = (mid_1[263:256] > mid_2[255:248]) ? 1 : 0;
assign detect_max[31][15] = (mid_1[263:256] > mid_2[263:256]) ? 1 : 0;
assign detect_max[31][16] = (mid_1[263:256] > mid_2[271:264]) ? 1 : 0;
assign detect_max[31][17] = (mid_1[263:256] > btm_0[255:248]) ? 1 : 0;
assign detect_max[31][18] = (mid_1[263:256] > btm_0[263:256]) ? 1 : 0;
assign detect_max[31][19] = (mid_1[263:256] > btm_0[271:264]) ? 1 : 0;
assign detect_max[31][20] = (mid_1[263:256] > btm_1[255:248]) ? 1 : 0;
assign detect_max[31][21] = (mid_1[263:256] > btm_1[263:256]) ? 1 : 0;
assign detect_max[31][22] = (mid_1[263:256] > btm_1[271:264]) ? 1 : 0;
assign detect_max[31][23] = (mid_1[263:256] > btm_2[255:248]) ? 1 : 0;
assign detect_max[31][24] = (mid_1[263:256] > btm_2[263:256]) ? 1 : 0;
assign detect_max[31][25] = (mid_1[263:256] > btm_2[271:264]) ? 1 : 0;

assign detect_max[32][0] = (mid_1[271:264] > top_0[263:256]) ? 1 : 0;
assign detect_max[32][1] = (mid_1[271:264] > top_0[271:264]) ? 1 : 0;
assign detect_max[32][2] = (mid_1[271:264] > top_0[279:272]) ? 1 : 0;
assign detect_max[32][3] = (mid_1[271:264] > top_1[263:256]) ? 1 : 0;
assign detect_max[32][4] = (mid_1[271:264] > top_1[271:264]) ? 1 : 0;
assign detect_max[32][5] = (mid_1[271:264] > top_1[279:272]) ? 1 : 0;
assign detect_max[32][6] = (mid_1[271:264] > top_2[263:256]) ? 1 : 0;
assign detect_max[32][7] = (mid_1[271:264] > top_2[271:264]) ? 1 : 0;
assign detect_max[32][8] = (mid_1[271:264] > top_2[279:272]) ? 1 : 0;
assign detect_max[32][9] = (mid_1[271:264] > mid_0[263:256]) ? 1 : 0;
assign detect_max[32][10] = (mid_1[271:264] > mid_0[271:264]) ? 1 : 0;
assign detect_max[32][11] = (mid_1[271:264] > mid_0[279:272]) ? 1 : 0;
assign detect_max[32][12] = (mid_1[271:264] > mid_1[263:256]) ? 1 : 0;
assign detect_max[32][13] = (mid_1[271:264] > mid_1[279:272]) ? 1 : 0;
assign detect_max[32][14] = (mid_1[271:264] > mid_2[263:256]) ? 1 : 0;
assign detect_max[32][15] = (mid_1[271:264] > mid_2[271:264]) ? 1 : 0;
assign detect_max[32][16] = (mid_1[271:264] > mid_2[279:272]) ? 1 : 0;
assign detect_max[32][17] = (mid_1[271:264] > btm_0[263:256]) ? 1 : 0;
assign detect_max[32][18] = (mid_1[271:264] > btm_0[271:264]) ? 1 : 0;
assign detect_max[32][19] = (mid_1[271:264] > btm_0[279:272]) ? 1 : 0;
assign detect_max[32][20] = (mid_1[271:264] > btm_1[263:256]) ? 1 : 0;
assign detect_max[32][21] = (mid_1[271:264] > btm_1[271:264]) ? 1 : 0;
assign detect_max[32][22] = (mid_1[271:264] > btm_1[279:272]) ? 1 : 0;
assign detect_max[32][23] = (mid_1[271:264] > btm_2[263:256]) ? 1 : 0;
assign detect_max[32][24] = (mid_1[271:264] > btm_2[271:264]) ? 1 : 0;
assign detect_max[32][25] = (mid_1[271:264] > btm_2[279:272]) ? 1 : 0;

assign detect_max[33][0] = (mid_1[279:272] > top_0[271:264]) ? 1 : 0;
assign detect_max[33][1] = (mid_1[279:272] > top_0[279:272]) ? 1 : 0;
assign detect_max[33][2] = (mid_1[279:272] > top_0[287:280]) ? 1 : 0;
assign detect_max[33][3] = (mid_1[279:272] > top_1[271:264]) ? 1 : 0;
assign detect_max[33][4] = (mid_1[279:272] > top_1[279:272]) ? 1 : 0;
assign detect_max[33][5] = (mid_1[279:272] > top_1[287:280]) ? 1 : 0;
assign detect_max[33][6] = (mid_1[279:272] > top_2[271:264]) ? 1 : 0;
assign detect_max[33][7] = (mid_1[279:272] > top_2[279:272]) ? 1 : 0;
assign detect_max[33][8] = (mid_1[279:272] > top_2[287:280]) ? 1 : 0;
assign detect_max[33][9] = (mid_1[279:272] > mid_0[271:264]) ? 1 : 0;
assign detect_max[33][10] = (mid_1[279:272] > mid_0[279:272]) ? 1 : 0;
assign detect_max[33][11] = (mid_1[279:272] > mid_0[287:280]) ? 1 : 0;
assign detect_max[33][12] = (mid_1[279:272] > mid_1[271:264]) ? 1 : 0;
assign detect_max[33][13] = (mid_1[279:272] > mid_1[287:280]) ? 1 : 0;
assign detect_max[33][14] = (mid_1[279:272] > mid_2[271:264]) ? 1 : 0;
assign detect_max[33][15] = (mid_1[279:272] > mid_2[279:272]) ? 1 : 0;
assign detect_max[33][16] = (mid_1[279:272] > mid_2[287:280]) ? 1 : 0;
assign detect_max[33][17] = (mid_1[279:272] > btm_0[271:264]) ? 1 : 0;
assign detect_max[33][18] = (mid_1[279:272] > btm_0[279:272]) ? 1 : 0;
assign detect_max[33][19] = (mid_1[279:272] > btm_0[287:280]) ? 1 : 0;
assign detect_max[33][20] = (mid_1[279:272] > btm_1[271:264]) ? 1 : 0;
assign detect_max[33][21] = (mid_1[279:272] > btm_1[279:272]) ? 1 : 0;
assign detect_max[33][22] = (mid_1[279:272] > btm_1[287:280]) ? 1 : 0;
assign detect_max[33][23] = (mid_1[279:272] > btm_2[271:264]) ? 1 : 0;
assign detect_max[33][24] = (mid_1[279:272] > btm_2[279:272]) ? 1 : 0;
assign detect_max[33][25] = (mid_1[279:272] > btm_2[287:280]) ? 1 : 0;

assign detect_max[34][0] = (mid_1[287:280] > top_0[279:272]) ? 1 : 0;
assign detect_max[34][1] = (mid_1[287:280] > top_0[287:280]) ? 1 : 0;
assign detect_max[34][2] = (mid_1[287:280] > top_0[295:288]) ? 1 : 0;
assign detect_max[34][3] = (mid_1[287:280] > top_1[279:272]) ? 1 : 0;
assign detect_max[34][4] = (mid_1[287:280] > top_1[287:280]) ? 1 : 0;
assign detect_max[34][5] = (mid_1[287:280] > top_1[295:288]) ? 1 : 0;
assign detect_max[34][6] = (mid_1[287:280] > top_2[279:272]) ? 1 : 0;
assign detect_max[34][7] = (mid_1[287:280] > top_2[287:280]) ? 1 : 0;
assign detect_max[34][8] = (mid_1[287:280] > top_2[295:288]) ? 1 : 0;
assign detect_max[34][9] = (mid_1[287:280] > mid_0[279:272]) ? 1 : 0;
assign detect_max[34][10] = (mid_1[287:280] > mid_0[287:280]) ? 1 : 0;
assign detect_max[34][11] = (mid_1[287:280] > mid_0[295:288]) ? 1 : 0;
assign detect_max[34][12] = (mid_1[287:280] > mid_1[279:272]) ? 1 : 0;
assign detect_max[34][13] = (mid_1[287:280] > mid_1[295:288]) ? 1 : 0;
assign detect_max[34][14] = (mid_1[287:280] > mid_2[279:272]) ? 1 : 0;
assign detect_max[34][15] = (mid_1[287:280] > mid_2[287:280]) ? 1 : 0;
assign detect_max[34][16] = (mid_1[287:280] > mid_2[295:288]) ? 1 : 0;
assign detect_max[34][17] = (mid_1[287:280] > btm_0[279:272]) ? 1 : 0;
assign detect_max[34][18] = (mid_1[287:280] > btm_0[287:280]) ? 1 : 0;
assign detect_max[34][19] = (mid_1[287:280] > btm_0[295:288]) ? 1 : 0;
assign detect_max[34][20] = (mid_1[287:280] > btm_1[279:272]) ? 1 : 0;
assign detect_max[34][21] = (mid_1[287:280] > btm_1[287:280]) ? 1 : 0;
assign detect_max[34][22] = (mid_1[287:280] > btm_1[295:288]) ? 1 : 0;
assign detect_max[34][23] = (mid_1[287:280] > btm_2[279:272]) ? 1 : 0;
assign detect_max[34][24] = (mid_1[287:280] > btm_2[287:280]) ? 1 : 0;
assign detect_max[34][25] = (mid_1[287:280] > btm_2[295:288]) ? 1 : 0;

assign detect_max[35][0] = (mid_1[295:288] > top_0[287:280]) ? 1 : 0;
assign detect_max[35][1] = (mid_1[295:288] > top_0[295:288]) ? 1 : 0;
assign detect_max[35][2] = (mid_1[295:288] > top_0[303:296]) ? 1 : 0;
assign detect_max[35][3] = (mid_1[295:288] > top_1[287:280]) ? 1 : 0;
assign detect_max[35][4] = (mid_1[295:288] > top_1[295:288]) ? 1 : 0;
assign detect_max[35][5] = (mid_1[295:288] > top_1[303:296]) ? 1 : 0;
assign detect_max[35][6] = (mid_1[295:288] > top_2[287:280]) ? 1 : 0;
assign detect_max[35][7] = (mid_1[295:288] > top_2[295:288]) ? 1 : 0;
assign detect_max[35][8] = (mid_1[295:288] > top_2[303:296]) ? 1 : 0;
assign detect_max[35][9] = (mid_1[295:288] > mid_0[287:280]) ? 1 : 0;
assign detect_max[35][10] = (mid_1[295:288] > mid_0[295:288]) ? 1 : 0;
assign detect_max[35][11] = (mid_1[295:288] > mid_0[303:296]) ? 1 : 0;
assign detect_max[35][12] = (mid_1[295:288] > mid_1[287:280]) ? 1 : 0;
assign detect_max[35][13] = (mid_1[295:288] > mid_1[303:296]) ? 1 : 0;
assign detect_max[35][14] = (mid_1[295:288] > mid_2[287:280]) ? 1 : 0;
assign detect_max[35][15] = (mid_1[295:288] > mid_2[295:288]) ? 1 : 0;
assign detect_max[35][16] = (mid_1[295:288] > mid_2[303:296]) ? 1 : 0;
assign detect_max[35][17] = (mid_1[295:288] > btm_0[287:280]) ? 1 : 0;
assign detect_max[35][18] = (mid_1[295:288] > btm_0[295:288]) ? 1 : 0;
assign detect_max[35][19] = (mid_1[295:288] > btm_0[303:296]) ? 1 : 0;
assign detect_max[35][20] = (mid_1[295:288] > btm_1[287:280]) ? 1 : 0;
assign detect_max[35][21] = (mid_1[295:288] > btm_1[295:288]) ? 1 : 0;
assign detect_max[35][22] = (mid_1[295:288] > btm_1[303:296]) ? 1 : 0;
assign detect_max[35][23] = (mid_1[295:288] > btm_2[287:280]) ? 1 : 0;
assign detect_max[35][24] = (mid_1[295:288] > btm_2[295:288]) ? 1 : 0;
assign detect_max[35][25] = (mid_1[295:288] > btm_2[303:296]) ? 1 : 0;

assign detect_max[36][0] = (mid_1[303:296] > top_0[295:288]) ? 1 : 0;
assign detect_max[36][1] = (mid_1[303:296] > top_0[303:296]) ? 1 : 0;
assign detect_max[36][2] = (mid_1[303:296] > top_0[311:304]) ? 1 : 0;
assign detect_max[36][3] = (mid_1[303:296] > top_1[295:288]) ? 1 : 0;
assign detect_max[36][4] = (mid_1[303:296] > top_1[303:296]) ? 1 : 0;
assign detect_max[36][5] = (mid_1[303:296] > top_1[311:304]) ? 1 : 0;
assign detect_max[36][6] = (mid_1[303:296] > top_2[295:288]) ? 1 : 0;
assign detect_max[36][7] = (mid_1[303:296] > top_2[303:296]) ? 1 : 0;
assign detect_max[36][8] = (mid_1[303:296] > top_2[311:304]) ? 1 : 0;
assign detect_max[36][9] = (mid_1[303:296] > mid_0[295:288]) ? 1 : 0;
assign detect_max[36][10] = (mid_1[303:296] > mid_0[303:296]) ? 1 : 0;
assign detect_max[36][11] = (mid_1[303:296] > mid_0[311:304]) ? 1 : 0;
assign detect_max[36][12] = (mid_1[303:296] > mid_1[295:288]) ? 1 : 0;
assign detect_max[36][13] = (mid_1[303:296] > mid_1[311:304]) ? 1 : 0;
assign detect_max[36][14] = (mid_1[303:296] > mid_2[295:288]) ? 1 : 0;
assign detect_max[36][15] = (mid_1[303:296] > mid_2[303:296]) ? 1 : 0;
assign detect_max[36][16] = (mid_1[303:296] > mid_2[311:304]) ? 1 : 0;
assign detect_max[36][17] = (mid_1[303:296] > btm_0[295:288]) ? 1 : 0;
assign detect_max[36][18] = (mid_1[303:296] > btm_0[303:296]) ? 1 : 0;
assign detect_max[36][19] = (mid_1[303:296] > btm_0[311:304]) ? 1 : 0;
assign detect_max[36][20] = (mid_1[303:296] > btm_1[295:288]) ? 1 : 0;
assign detect_max[36][21] = (mid_1[303:296] > btm_1[303:296]) ? 1 : 0;
assign detect_max[36][22] = (mid_1[303:296] > btm_1[311:304]) ? 1 : 0;
assign detect_max[36][23] = (mid_1[303:296] > btm_2[295:288]) ? 1 : 0;
assign detect_max[36][24] = (mid_1[303:296] > btm_2[303:296]) ? 1 : 0;
assign detect_max[36][25] = (mid_1[303:296] > btm_2[311:304]) ? 1 : 0;

assign detect_max[37][0] = (mid_1[311:304] > top_0[303:296]) ? 1 : 0;
assign detect_max[37][1] = (mid_1[311:304] > top_0[311:304]) ? 1 : 0;
assign detect_max[37][2] = (mid_1[311:304] > top_0[319:312]) ? 1 : 0;
assign detect_max[37][3] = (mid_1[311:304] > top_1[303:296]) ? 1 : 0;
assign detect_max[37][4] = (mid_1[311:304] > top_1[311:304]) ? 1 : 0;
assign detect_max[37][5] = (mid_1[311:304] > top_1[319:312]) ? 1 : 0;
assign detect_max[37][6] = (mid_1[311:304] > top_2[303:296]) ? 1 : 0;
assign detect_max[37][7] = (mid_1[311:304] > top_2[311:304]) ? 1 : 0;
assign detect_max[37][8] = (mid_1[311:304] > top_2[319:312]) ? 1 : 0;
assign detect_max[37][9] = (mid_1[311:304] > mid_0[303:296]) ? 1 : 0;
assign detect_max[37][10] = (mid_1[311:304] > mid_0[311:304]) ? 1 : 0;
assign detect_max[37][11] = (mid_1[311:304] > mid_0[319:312]) ? 1 : 0;
assign detect_max[37][12] = (mid_1[311:304] > mid_1[303:296]) ? 1 : 0;
assign detect_max[37][13] = (mid_1[311:304] > mid_1[319:312]) ? 1 : 0;
assign detect_max[37][14] = (mid_1[311:304] > mid_2[303:296]) ? 1 : 0;
assign detect_max[37][15] = (mid_1[311:304] > mid_2[311:304]) ? 1 : 0;
assign detect_max[37][16] = (mid_1[311:304] > mid_2[319:312]) ? 1 : 0;
assign detect_max[37][17] = (mid_1[311:304] > btm_0[303:296]) ? 1 : 0;
assign detect_max[37][18] = (mid_1[311:304] > btm_0[311:304]) ? 1 : 0;
assign detect_max[37][19] = (mid_1[311:304] > btm_0[319:312]) ? 1 : 0;
assign detect_max[37][20] = (mid_1[311:304] > btm_1[303:296]) ? 1 : 0;
assign detect_max[37][21] = (mid_1[311:304] > btm_1[311:304]) ? 1 : 0;
assign detect_max[37][22] = (mid_1[311:304] > btm_1[319:312]) ? 1 : 0;
assign detect_max[37][23] = (mid_1[311:304] > btm_2[303:296]) ? 1 : 0;
assign detect_max[37][24] = (mid_1[311:304] > btm_2[311:304]) ? 1 : 0;
assign detect_max[37][25] = (mid_1[311:304] > btm_2[319:312]) ? 1 : 0;

assign detect_max[38][0] = (mid_1[319:312] > top_0[311:304]) ? 1 : 0;
assign detect_max[38][1] = (mid_1[319:312] > top_0[319:312]) ? 1 : 0;
assign detect_max[38][2] = (mid_1[319:312] > top_0[327:320]) ? 1 : 0;
assign detect_max[38][3] = (mid_1[319:312] > top_1[311:304]) ? 1 : 0;
assign detect_max[38][4] = (mid_1[319:312] > top_1[319:312]) ? 1 : 0;
assign detect_max[38][5] = (mid_1[319:312] > top_1[327:320]) ? 1 : 0;
assign detect_max[38][6] = (mid_1[319:312] > top_2[311:304]) ? 1 : 0;
assign detect_max[38][7] = (mid_1[319:312] > top_2[319:312]) ? 1 : 0;
assign detect_max[38][8] = (mid_1[319:312] > top_2[327:320]) ? 1 : 0;
assign detect_max[38][9] = (mid_1[319:312] > mid_0[311:304]) ? 1 : 0;
assign detect_max[38][10] = (mid_1[319:312] > mid_0[319:312]) ? 1 : 0;
assign detect_max[38][11] = (mid_1[319:312] > mid_0[327:320]) ? 1 : 0;
assign detect_max[38][12] = (mid_1[319:312] > mid_1[311:304]) ? 1 : 0;
assign detect_max[38][13] = (mid_1[319:312] > mid_1[327:320]) ? 1 : 0;
assign detect_max[38][14] = (mid_1[319:312] > mid_2[311:304]) ? 1 : 0;
assign detect_max[38][15] = (mid_1[319:312] > mid_2[319:312]) ? 1 : 0;
assign detect_max[38][16] = (mid_1[319:312] > mid_2[327:320]) ? 1 : 0;
assign detect_max[38][17] = (mid_1[319:312] > btm_0[311:304]) ? 1 : 0;
assign detect_max[38][18] = (mid_1[319:312] > btm_0[319:312]) ? 1 : 0;
assign detect_max[38][19] = (mid_1[319:312] > btm_0[327:320]) ? 1 : 0;
assign detect_max[38][20] = (mid_1[319:312] > btm_1[311:304]) ? 1 : 0;
assign detect_max[38][21] = (mid_1[319:312] > btm_1[319:312]) ? 1 : 0;
assign detect_max[38][22] = (mid_1[319:312] > btm_1[327:320]) ? 1 : 0;
assign detect_max[38][23] = (mid_1[319:312] > btm_2[311:304]) ? 1 : 0;
assign detect_max[38][24] = (mid_1[319:312] > btm_2[319:312]) ? 1 : 0;
assign detect_max[38][25] = (mid_1[319:312] > btm_2[327:320]) ? 1 : 0;

assign detect_max[39][0] = (mid_1[327:320] > top_0[319:312]) ? 1 : 0;
assign detect_max[39][1] = (mid_1[327:320] > top_0[327:320]) ? 1 : 0;
assign detect_max[39][2] = (mid_1[327:320] > top_0[335:328]) ? 1 : 0;
assign detect_max[39][3] = (mid_1[327:320] > top_1[319:312]) ? 1 : 0;
assign detect_max[39][4] = (mid_1[327:320] > top_1[327:320]) ? 1 : 0;
assign detect_max[39][5] = (mid_1[327:320] > top_1[335:328]) ? 1 : 0;
assign detect_max[39][6] = (mid_1[327:320] > top_2[319:312]) ? 1 : 0;
assign detect_max[39][7] = (mid_1[327:320] > top_2[327:320]) ? 1 : 0;
assign detect_max[39][8] = (mid_1[327:320] > top_2[335:328]) ? 1 : 0;
assign detect_max[39][9] = (mid_1[327:320] > mid_0[319:312]) ? 1 : 0;
assign detect_max[39][10] = (mid_1[327:320] > mid_0[327:320]) ? 1 : 0;
assign detect_max[39][11] = (mid_1[327:320] > mid_0[335:328]) ? 1 : 0;
assign detect_max[39][12] = (mid_1[327:320] > mid_1[319:312]) ? 1 : 0;
assign detect_max[39][13] = (mid_1[327:320] > mid_1[335:328]) ? 1 : 0;
assign detect_max[39][14] = (mid_1[327:320] > mid_2[319:312]) ? 1 : 0;
assign detect_max[39][15] = (mid_1[327:320] > mid_2[327:320]) ? 1 : 0;
assign detect_max[39][16] = (mid_1[327:320] > mid_2[335:328]) ? 1 : 0;
assign detect_max[39][17] = (mid_1[327:320] > btm_0[319:312]) ? 1 : 0;
assign detect_max[39][18] = (mid_1[327:320] > btm_0[327:320]) ? 1 : 0;
assign detect_max[39][19] = (mid_1[327:320] > btm_0[335:328]) ? 1 : 0;
assign detect_max[39][20] = (mid_1[327:320] > btm_1[319:312]) ? 1 : 0;
assign detect_max[39][21] = (mid_1[327:320] > btm_1[327:320]) ? 1 : 0;
assign detect_max[39][22] = (mid_1[327:320] > btm_1[335:328]) ? 1 : 0;
assign detect_max[39][23] = (mid_1[327:320] > btm_2[319:312]) ? 1 : 0;
assign detect_max[39][24] = (mid_1[327:320] > btm_2[327:320]) ? 1 : 0;
assign detect_max[39][25] = (mid_1[327:320] > btm_2[335:328]) ? 1 : 0;

assign detect_max[40][0] = (mid_1[335:328] > top_0[327:320]) ? 1 : 0;
assign detect_max[40][1] = (mid_1[335:328] > top_0[335:328]) ? 1 : 0;
assign detect_max[40][2] = (mid_1[335:328] > top_0[343:336]) ? 1 : 0;
assign detect_max[40][3] = (mid_1[335:328] > top_1[327:320]) ? 1 : 0;
assign detect_max[40][4] = (mid_1[335:328] > top_1[335:328]) ? 1 : 0;
assign detect_max[40][5] = (mid_1[335:328] > top_1[343:336]) ? 1 : 0;
assign detect_max[40][6] = (mid_1[335:328] > top_2[327:320]) ? 1 : 0;
assign detect_max[40][7] = (mid_1[335:328] > top_2[335:328]) ? 1 : 0;
assign detect_max[40][8] = (mid_1[335:328] > top_2[343:336]) ? 1 : 0;
assign detect_max[40][9] = (mid_1[335:328] > mid_0[327:320]) ? 1 : 0;
assign detect_max[40][10] = (mid_1[335:328] > mid_0[335:328]) ? 1 : 0;
assign detect_max[40][11] = (mid_1[335:328] > mid_0[343:336]) ? 1 : 0;
assign detect_max[40][12] = (mid_1[335:328] > mid_1[327:320]) ? 1 : 0;
assign detect_max[40][13] = (mid_1[335:328] > mid_1[343:336]) ? 1 : 0;
assign detect_max[40][14] = (mid_1[335:328] > mid_2[327:320]) ? 1 : 0;
assign detect_max[40][15] = (mid_1[335:328] > mid_2[335:328]) ? 1 : 0;
assign detect_max[40][16] = (mid_1[335:328] > mid_2[343:336]) ? 1 : 0;
assign detect_max[40][17] = (mid_1[335:328] > btm_0[327:320]) ? 1 : 0;
assign detect_max[40][18] = (mid_1[335:328] > btm_0[335:328]) ? 1 : 0;
assign detect_max[40][19] = (mid_1[335:328] > btm_0[343:336]) ? 1 : 0;
assign detect_max[40][20] = (mid_1[335:328] > btm_1[327:320]) ? 1 : 0;
assign detect_max[40][21] = (mid_1[335:328] > btm_1[335:328]) ? 1 : 0;
assign detect_max[40][22] = (mid_1[335:328] > btm_1[343:336]) ? 1 : 0;
assign detect_max[40][23] = (mid_1[335:328] > btm_2[327:320]) ? 1 : 0;
assign detect_max[40][24] = (mid_1[335:328] > btm_2[335:328]) ? 1 : 0;
assign detect_max[40][25] = (mid_1[335:328] > btm_2[343:336]) ? 1 : 0;

assign detect_max[41][0] = (mid_1[343:336] > top_0[335:328]) ? 1 : 0;
assign detect_max[41][1] = (mid_1[343:336] > top_0[343:336]) ? 1 : 0;
assign detect_max[41][2] = (mid_1[343:336] > top_0[351:344]) ? 1 : 0;
assign detect_max[41][3] = (mid_1[343:336] > top_1[335:328]) ? 1 : 0;
assign detect_max[41][4] = (mid_1[343:336] > top_1[343:336]) ? 1 : 0;
assign detect_max[41][5] = (mid_1[343:336] > top_1[351:344]) ? 1 : 0;
assign detect_max[41][6] = (mid_1[343:336] > top_2[335:328]) ? 1 : 0;
assign detect_max[41][7] = (mid_1[343:336] > top_2[343:336]) ? 1 : 0;
assign detect_max[41][8] = (mid_1[343:336] > top_2[351:344]) ? 1 : 0;
assign detect_max[41][9] = (mid_1[343:336] > mid_0[335:328]) ? 1 : 0;
assign detect_max[41][10] = (mid_1[343:336] > mid_0[343:336]) ? 1 : 0;
assign detect_max[41][11] = (mid_1[343:336] > mid_0[351:344]) ? 1 : 0;
assign detect_max[41][12] = (mid_1[343:336] > mid_1[335:328]) ? 1 : 0;
assign detect_max[41][13] = (mid_1[343:336] > mid_1[351:344]) ? 1 : 0;
assign detect_max[41][14] = (mid_1[343:336] > mid_2[335:328]) ? 1 : 0;
assign detect_max[41][15] = (mid_1[343:336] > mid_2[343:336]) ? 1 : 0;
assign detect_max[41][16] = (mid_1[343:336] > mid_2[351:344]) ? 1 : 0;
assign detect_max[41][17] = (mid_1[343:336] > btm_0[335:328]) ? 1 : 0;
assign detect_max[41][18] = (mid_1[343:336] > btm_0[343:336]) ? 1 : 0;
assign detect_max[41][19] = (mid_1[343:336] > btm_0[351:344]) ? 1 : 0;
assign detect_max[41][20] = (mid_1[343:336] > btm_1[335:328]) ? 1 : 0;
assign detect_max[41][21] = (mid_1[343:336] > btm_1[343:336]) ? 1 : 0;
assign detect_max[41][22] = (mid_1[343:336] > btm_1[351:344]) ? 1 : 0;
assign detect_max[41][23] = (mid_1[343:336] > btm_2[335:328]) ? 1 : 0;
assign detect_max[41][24] = (mid_1[343:336] > btm_2[343:336]) ? 1 : 0;
assign detect_max[41][25] = (mid_1[343:336] > btm_2[351:344]) ? 1 : 0;

assign detect_max[42][0] = (mid_1[351:344] > top_0[343:336]) ? 1 : 0;
assign detect_max[42][1] = (mid_1[351:344] > top_0[351:344]) ? 1 : 0;
assign detect_max[42][2] = (mid_1[351:344] > top_0[359:352]) ? 1 : 0;
assign detect_max[42][3] = (mid_1[351:344] > top_1[343:336]) ? 1 : 0;
assign detect_max[42][4] = (mid_1[351:344] > top_1[351:344]) ? 1 : 0;
assign detect_max[42][5] = (mid_1[351:344] > top_1[359:352]) ? 1 : 0;
assign detect_max[42][6] = (mid_1[351:344] > top_2[343:336]) ? 1 : 0;
assign detect_max[42][7] = (mid_1[351:344] > top_2[351:344]) ? 1 : 0;
assign detect_max[42][8] = (mid_1[351:344] > top_2[359:352]) ? 1 : 0;
assign detect_max[42][9] = (mid_1[351:344] > mid_0[343:336]) ? 1 : 0;
assign detect_max[42][10] = (mid_1[351:344] > mid_0[351:344]) ? 1 : 0;
assign detect_max[42][11] = (mid_1[351:344] > mid_0[359:352]) ? 1 : 0;
assign detect_max[42][12] = (mid_1[351:344] > mid_1[343:336]) ? 1 : 0;
assign detect_max[42][13] = (mid_1[351:344] > mid_1[359:352]) ? 1 : 0;
assign detect_max[42][14] = (mid_1[351:344] > mid_2[343:336]) ? 1 : 0;
assign detect_max[42][15] = (mid_1[351:344] > mid_2[351:344]) ? 1 : 0;
assign detect_max[42][16] = (mid_1[351:344] > mid_2[359:352]) ? 1 : 0;
assign detect_max[42][17] = (mid_1[351:344] > btm_0[343:336]) ? 1 : 0;
assign detect_max[42][18] = (mid_1[351:344] > btm_0[351:344]) ? 1 : 0;
assign detect_max[42][19] = (mid_1[351:344] > btm_0[359:352]) ? 1 : 0;
assign detect_max[42][20] = (mid_1[351:344] > btm_1[343:336]) ? 1 : 0;
assign detect_max[42][21] = (mid_1[351:344] > btm_1[351:344]) ? 1 : 0;
assign detect_max[42][22] = (mid_1[351:344] > btm_1[359:352]) ? 1 : 0;
assign detect_max[42][23] = (mid_1[351:344] > btm_2[343:336]) ? 1 : 0;
assign detect_max[42][24] = (mid_1[351:344] > btm_2[351:344]) ? 1 : 0;
assign detect_max[42][25] = (mid_1[351:344] > btm_2[359:352]) ? 1 : 0;

assign detect_max[43][0] = (mid_1[359:352] > top_0[351:344]) ? 1 : 0;
assign detect_max[43][1] = (mid_1[359:352] > top_0[359:352]) ? 1 : 0;
assign detect_max[43][2] = (mid_1[359:352] > top_0[367:360]) ? 1 : 0;
assign detect_max[43][3] = (mid_1[359:352] > top_1[351:344]) ? 1 : 0;
assign detect_max[43][4] = (mid_1[359:352] > top_1[359:352]) ? 1 : 0;
assign detect_max[43][5] = (mid_1[359:352] > top_1[367:360]) ? 1 : 0;
assign detect_max[43][6] = (mid_1[359:352] > top_2[351:344]) ? 1 : 0;
assign detect_max[43][7] = (mid_1[359:352] > top_2[359:352]) ? 1 : 0;
assign detect_max[43][8] = (mid_1[359:352] > top_2[367:360]) ? 1 : 0;
assign detect_max[43][9] = (mid_1[359:352] > mid_0[351:344]) ? 1 : 0;
assign detect_max[43][10] = (mid_1[359:352] > mid_0[359:352]) ? 1 : 0;
assign detect_max[43][11] = (mid_1[359:352] > mid_0[367:360]) ? 1 : 0;
assign detect_max[43][12] = (mid_1[359:352] > mid_1[351:344]) ? 1 : 0;
assign detect_max[43][13] = (mid_1[359:352] > mid_1[367:360]) ? 1 : 0;
assign detect_max[43][14] = (mid_1[359:352] > mid_2[351:344]) ? 1 : 0;
assign detect_max[43][15] = (mid_1[359:352] > mid_2[359:352]) ? 1 : 0;
assign detect_max[43][16] = (mid_1[359:352] > mid_2[367:360]) ? 1 : 0;
assign detect_max[43][17] = (mid_1[359:352] > btm_0[351:344]) ? 1 : 0;
assign detect_max[43][18] = (mid_1[359:352] > btm_0[359:352]) ? 1 : 0;
assign detect_max[43][19] = (mid_1[359:352] > btm_0[367:360]) ? 1 : 0;
assign detect_max[43][20] = (mid_1[359:352] > btm_1[351:344]) ? 1 : 0;
assign detect_max[43][21] = (mid_1[359:352] > btm_1[359:352]) ? 1 : 0;
assign detect_max[43][22] = (mid_1[359:352] > btm_1[367:360]) ? 1 : 0;
assign detect_max[43][23] = (mid_1[359:352] > btm_2[351:344]) ? 1 : 0;
assign detect_max[43][24] = (mid_1[359:352] > btm_2[359:352]) ? 1 : 0;
assign detect_max[43][25] = (mid_1[359:352] > btm_2[367:360]) ? 1 : 0;

assign detect_max[44][0] = (mid_1[367:360] > top_0[359:352]) ? 1 : 0;
assign detect_max[44][1] = (mid_1[367:360] > top_0[367:360]) ? 1 : 0;
assign detect_max[44][2] = (mid_1[367:360] > top_0[375:368]) ? 1 : 0;
assign detect_max[44][3] = (mid_1[367:360] > top_1[359:352]) ? 1 : 0;
assign detect_max[44][4] = (mid_1[367:360] > top_1[367:360]) ? 1 : 0;
assign detect_max[44][5] = (mid_1[367:360] > top_1[375:368]) ? 1 : 0;
assign detect_max[44][6] = (mid_1[367:360] > top_2[359:352]) ? 1 : 0;
assign detect_max[44][7] = (mid_1[367:360] > top_2[367:360]) ? 1 : 0;
assign detect_max[44][8] = (mid_1[367:360] > top_2[375:368]) ? 1 : 0;
assign detect_max[44][9] = (mid_1[367:360] > mid_0[359:352]) ? 1 : 0;
assign detect_max[44][10] = (mid_1[367:360] > mid_0[367:360]) ? 1 : 0;
assign detect_max[44][11] = (mid_1[367:360] > mid_0[375:368]) ? 1 : 0;
assign detect_max[44][12] = (mid_1[367:360] > mid_1[359:352]) ? 1 : 0;
assign detect_max[44][13] = (mid_1[367:360] > mid_1[375:368]) ? 1 : 0;
assign detect_max[44][14] = (mid_1[367:360] > mid_2[359:352]) ? 1 : 0;
assign detect_max[44][15] = (mid_1[367:360] > mid_2[367:360]) ? 1 : 0;
assign detect_max[44][16] = (mid_1[367:360] > mid_2[375:368]) ? 1 : 0;
assign detect_max[44][17] = (mid_1[367:360] > btm_0[359:352]) ? 1 : 0;
assign detect_max[44][18] = (mid_1[367:360] > btm_0[367:360]) ? 1 : 0;
assign detect_max[44][19] = (mid_1[367:360] > btm_0[375:368]) ? 1 : 0;
assign detect_max[44][20] = (mid_1[367:360] > btm_1[359:352]) ? 1 : 0;
assign detect_max[44][21] = (mid_1[367:360] > btm_1[367:360]) ? 1 : 0;
assign detect_max[44][22] = (mid_1[367:360] > btm_1[375:368]) ? 1 : 0;
assign detect_max[44][23] = (mid_1[367:360] > btm_2[359:352]) ? 1 : 0;
assign detect_max[44][24] = (mid_1[367:360] > btm_2[367:360]) ? 1 : 0;
assign detect_max[44][25] = (mid_1[367:360] > btm_2[375:368]) ? 1 : 0;

assign detect_max[45][0] = (mid_1[375:368] > top_0[367:360]) ? 1 : 0;
assign detect_max[45][1] = (mid_1[375:368] > top_0[375:368]) ? 1 : 0;
assign detect_max[45][2] = (mid_1[375:368] > top_0[383:376]) ? 1 : 0;
assign detect_max[45][3] = (mid_1[375:368] > top_1[367:360]) ? 1 : 0;
assign detect_max[45][4] = (mid_1[375:368] > top_1[375:368]) ? 1 : 0;
assign detect_max[45][5] = (mid_1[375:368] > top_1[383:376]) ? 1 : 0;
assign detect_max[45][6] = (mid_1[375:368] > top_2[367:360]) ? 1 : 0;
assign detect_max[45][7] = (mid_1[375:368] > top_2[375:368]) ? 1 : 0;
assign detect_max[45][8] = (mid_1[375:368] > top_2[383:376]) ? 1 : 0;
assign detect_max[45][9] = (mid_1[375:368] > mid_0[367:360]) ? 1 : 0;
assign detect_max[45][10] = (mid_1[375:368] > mid_0[375:368]) ? 1 : 0;
assign detect_max[45][11] = (mid_1[375:368] > mid_0[383:376]) ? 1 : 0;
assign detect_max[45][12] = (mid_1[375:368] > mid_1[367:360]) ? 1 : 0;
assign detect_max[45][13] = (mid_1[375:368] > mid_1[383:376]) ? 1 : 0;
assign detect_max[45][14] = (mid_1[375:368] > mid_2[367:360]) ? 1 : 0;
assign detect_max[45][15] = (mid_1[375:368] > mid_2[375:368]) ? 1 : 0;
assign detect_max[45][16] = (mid_1[375:368] > mid_2[383:376]) ? 1 : 0;
assign detect_max[45][17] = (mid_1[375:368] > btm_0[367:360]) ? 1 : 0;
assign detect_max[45][18] = (mid_1[375:368] > btm_0[375:368]) ? 1 : 0;
assign detect_max[45][19] = (mid_1[375:368] > btm_0[383:376]) ? 1 : 0;
assign detect_max[45][20] = (mid_1[375:368] > btm_1[367:360]) ? 1 : 0;
assign detect_max[45][21] = (mid_1[375:368] > btm_1[375:368]) ? 1 : 0;
assign detect_max[45][22] = (mid_1[375:368] > btm_1[383:376]) ? 1 : 0;
assign detect_max[45][23] = (mid_1[375:368] > btm_2[367:360]) ? 1 : 0;
assign detect_max[45][24] = (mid_1[375:368] > btm_2[375:368]) ? 1 : 0;
assign detect_max[45][25] = (mid_1[375:368] > btm_2[383:376]) ? 1 : 0;

assign detect_max[46][0] = (mid_1[383:376] > top_0[375:368]) ? 1 : 0;
assign detect_max[46][1] = (mid_1[383:376] > top_0[383:376]) ? 1 : 0;
assign detect_max[46][2] = (mid_1[383:376] > top_0[391:384]) ? 1 : 0;
assign detect_max[46][3] = (mid_1[383:376] > top_1[375:368]) ? 1 : 0;
assign detect_max[46][4] = (mid_1[383:376] > top_1[383:376]) ? 1 : 0;
assign detect_max[46][5] = (mid_1[383:376] > top_1[391:384]) ? 1 : 0;
assign detect_max[46][6] = (mid_1[383:376] > top_2[375:368]) ? 1 : 0;
assign detect_max[46][7] = (mid_1[383:376] > top_2[383:376]) ? 1 : 0;
assign detect_max[46][8] = (mid_1[383:376] > top_2[391:384]) ? 1 : 0;
assign detect_max[46][9] = (mid_1[383:376] > mid_0[375:368]) ? 1 : 0;
assign detect_max[46][10] = (mid_1[383:376] > mid_0[383:376]) ? 1 : 0;
assign detect_max[46][11] = (mid_1[383:376] > mid_0[391:384]) ? 1 : 0;
assign detect_max[46][12] = (mid_1[383:376] > mid_1[375:368]) ? 1 : 0;
assign detect_max[46][13] = (mid_1[383:376] > mid_1[391:384]) ? 1 : 0;
assign detect_max[46][14] = (mid_1[383:376] > mid_2[375:368]) ? 1 : 0;
assign detect_max[46][15] = (mid_1[383:376] > mid_2[383:376]) ? 1 : 0;
assign detect_max[46][16] = (mid_1[383:376] > mid_2[391:384]) ? 1 : 0;
assign detect_max[46][17] = (mid_1[383:376] > btm_0[375:368]) ? 1 : 0;
assign detect_max[46][18] = (mid_1[383:376] > btm_0[383:376]) ? 1 : 0;
assign detect_max[46][19] = (mid_1[383:376] > btm_0[391:384]) ? 1 : 0;
assign detect_max[46][20] = (mid_1[383:376] > btm_1[375:368]) ? 1 : 0;
assign detect_max[46][21] = (mid_1[383:376] > btm_1[383:376]) ? 1 : 0;
assign detect_max[46][22] = (mid_1[383:376] > btm_1[391:384]) ? 1 : 0;
assign detect_max[46][23] = (mid_1[383:376] > btm_2[375:368]) ? 1 : 0;
assign detect_max[46][24] = (mid_1[383:376] > btm_2[383:376]) ? 1 : 0;
assign detect_max[46][25] = (mid_1[383:376] > btm_2[391:384]) ? 1 : 0;

assign detect_max[47][0] = (mid_1[391:384] > top_0[383:376]) ? 1 : 0;
assign detect_max[47][1] = (mid_1[391:384] > top_0[391:384]) ? 1 : 0;
assign detect_max[47][2] = (mid_1[391:384] > top_0[399:392]) ? 1 : 0;
assign detect_max[47][3] = (mid_1[391:384] > top_1[383:376]) ? 1 : 0;
assign detect_max[47][4] = (mid_1[391:384] > top_1[391:384]) ? 1 : 0;
assign detect_max[47][5] = (mid_1[391:384] > top_1[399:392]) ? 1 : 0;
assign detect_max[47][6] = (mid_1[391:384] > top_2[383:376]) ? 1 : 0;
assign detect_max[47][7] = (mid_1[391:384] > top_2[391:384]) ? 1 : 0;
assign detect_max[47][8] = (mid_1[391:384] > top_2[399:392]) ? 1 : 0;
assign detect_max[47][9] = (mid_1[391:384] > mid_0[383:376]) ? 1 : 0;
assign detect_max[47][10] = (mid_1[391:384] > mid_0[391:384]) ? 1 : 0;
assign detect_max[47][11] = (mid_1[391:384] > mid_0[399:392]) ? 1 : 0;
assign detect_max[47][12] = (mid_1[391:384] > mid_1[383:376]) ? 1 : 0;
assign detect_max[47][13] = (mid_1[391:384] > mid_1[399:392]) ? 1 : 0;
assign detect_max[47][14] = (mid_1[391:384] > mid_2[383:376]) ? 1 : 0;
assign detect_max[47][15] = (mid_1[391:384] > mid_2[391:384]) ? 1 : 0;
assign detect_max[47][16] = (mid_1[391:384] > mid_2[399:392]) ? 1 : 0;
assign detect_max[47][17] = (mid_1[391:384] > btm_0[383:376]) ? 1 : 0;
assign detect_max[47][18] = (mid_1[391:384] > btm_0[391:384]) ? 1 : 0;
assign detect_max[47][19] = (mid_1[391:384] > btm_0[399:392]) ? 1 : 0;
assign detect_max[47][20] = (mid_1[391:384] > btm_1[383:376]) ? 1 : 0;
assign detect_max[47][21] = (mid_1[391:384] > btm_1[391:384]) ? 1 : 0;
assign detect_max[47][22] = (mid_1[391:384] > btm_1[399:392]) ? 1 : 0;
assign detect_max[47][23] = (mid_1[391:384] > btm_2[383:376]) ? 1 : 0;
assign detect_max[47][24] = (mid_1[391:384] > btm_2[391:384]) ? 1 : 0;
assign detect_max[47][25] = (mid_1[391:384] > btm_2[399:392]) ? 1 : 0;

assign detect_max[48][0] = (mid_1[399:392] > top_0[391:384]) ? 1 : 0;
assign detect_max[48][1] = (mid_1[399:392] > top_0[399:392]) ? 1 : 0;
assign detect_max[48][2] = (mid_1[399:392] > top_0[407:400]) ? 1 : 0;
assign detect_max[48][3] = (mid_1[399:392] > top_1[391:384]) ? 1 : 0;
assign detect_max[48][4] = (mid_1[399:392] > top_1[399:392]) ? 1 : 0;
assign detect_max[48][5] = (mid_1[399:392] > top_1[407:400]) ? 1 : 0;
assign detect_max[48][6] = (mid_1[399:392] > top_2[391:384]) ? 1 : 0;
assign detect_max[48][7] = (mid_1[399:392] > top_2[399:392]) ? 1 : 0;
assign detect_max[48][8] = (mid_1[399:392] > top_2[407:400]) ? 1 : 0;
assign detect_max[48][9] = (mid_1[399:392] > mid_0[391:384]) ? 1 : 0;
assign detect_max[48][10] = (mid_1[399:392] > mid_0[399:392]) ? 1 : 0;
assign detect_max[48][11] = (mid_1[399:392] > mid_0[407:400]) ? 1 : 0;
assign detect_max[48][12] = (mid_1[399:392] > mid_1[391:384]) ? 1 : 0;
assign detect_max[48][13] = (mid_1[399:392] > mid_1[407:400]) ? 1 : 0;
assign detect_max[48][14] = (mid_1[399:392] > mid_2[391:384]) ? 1 : 0;
assign detect_max[48][15] = (mid_1[399:392] > mid_2[399:392]) ? 1 : 0;
assign detect_max[48][16] = (mid_1[399:392] > mid_2[407:400]) ? 1 : 0;
assign detect_max[48][17] = (mid_1[399:392] > btm_0[391:384]) ? 1 : 0;
assign detect_max[48][18] = (mid_1[399:392] > btm_0[399:392]) ? 1 : 0;
assign detect_max[48][19] = (mid_1[399:392] > btm_0[407:400]) ? 1 : 0;
assign detect_max[48][20] = (mid_1[399:392] > btm_1[391:384]) ? 1 : 0;
assign detect_max[48][21] = (mid_1[399:392] > btm_1[399:392]) ? 1 : 0;
assign detect_max[48][22] = (mid_1[399:392] > btm_1[407:400]) ? 1 : 0;
assign detect_max[48][23] = (mid_1[399:392] > btm_2[391:384]) ? 1 : 0;
assign detect_max[48][24] = (mid_1[399:392] > btm_2[399:392]) ? 1 : 0;
assign detect_max[48][25] = (mid_1[399:392] > btm_2[407:400]) ? 1 : 0;

assign detect_max[49][0] = (mid_1[407:400] > top_0[399:392]) ? 1 : 0;
assign detect_max[49][1] = (mid_1[407:400] > top_0[407:400]) ? 1 : 0;
assign detect_max[49][2] = (mid_1[407:400] > top_0[415:408]) ? 1 : 0;
assign detect_max[49][3] = (mid_1[407:400] > top_1[399:392]) ? 1 : 0;
assign detect_max[49][4] = (mid_1[407:400] > top_1[407:400]) ? 1 : 0;
assign detect_max[49][5] = (mid_1[407:400] > top_1[415:408]) ? 1 : 0;
assign detect_max[49][6] = (mid_1[407:400] > top_2[399:392]) ? 1 : 0;
assign detect_max[49][7] = (mid_1[407:400] > top_2[407:400]) ? 1 : 0;
assign detect_max[49][8] = (mid_1[407:400] > top_2[415:408]) ? 1 : 0;
assign detect_max[49][9] = (mid_1[407:400] > mid_0[399:392]) ? 1 : 0;
assign detect_max[49][10] = (mid_1[407:400] > mid_0[407:400]) ? 1 : 0;
assign detect_max[49][11] = (mid_1[407:400] > mid_0[415:408]) ? 1 : 0;
assign detect_max[49][12] = (mid_1[407:400] > mid_1[399:392]) ? 1 : 0;
assign detect_max[49][13] = (mid_1[407:400] > mid_1[415:408]) ? 1 : 0;
assign detect_max[49][14] = (mid_1[407:400] > mid_2[399:392]) ? 1 : 0;
assign detect_max[49][15] = (mid_1[407:400] > mid_2[407:400]) ? 1 : 0;
assign detect_max[49][16] = (mid_1[407:400] > mid_2[415:408]) ? 1 : 0;
assign detect_max[49][17] = (mid_1[407:400] > btm_0[399:392]) ? 1 : 0;
assign detect_max[49][18] = (mid_1[407:400] > btm_0[407:400]) ? 1 : 0;
assign detect_max[49][19] = (mid_1[407:400] > btm_0[415:408]) ? 1 : 0;
assign detect_max[49][20] = (mid_1[407:400] > btm_1[399:392]) ? 1 : 0;
assign detect_max[49][21] = (mid_1[407:400] > btm_1[407:400]) ? 1 : 0;
assign detect_max[49][22] = (mid_1[407:400] > btm_1[415:408]) ? 1 : 0;
assign detect_max[49][23] = (mid_1[407:400] > btm_2[399:392]) ? 1 : 0;
assign detect_max[49][24] = (mid_1[407:400] > btm_2[407:400]) ? 1 : 0;
assign detect_max[49][25] = (mid_1[407:400] > btm_2[415:408]) ? 1 : 0;

assign detect_max[50][0] = (mid_1[415:408] > top_0[407:400]) ? 1 : 0;
assign detect_max[50][1] = (mid_1[415:408] > top_0[415:408]) ? 1 : 0;
assign detect_max[50][2] = (mid_1[415:408] > top_0[423:416]) ? 1 : 0;
assign detect_max[50][3] = (mid_1[415:408] > top_1[407:400]) ? 1 : 0;
assign detect_max[50][4] = (mid_1[415:408] > top_1[415:408]) ? 1 : 0;
assign detect_max[50][5] = (mid_1[415:408] > top_1[423:416]) ? 1 : 0;
assign detect_max[50][6] = (mid_1[415:408] > top_2[407:400]) ? 1 : 0;
assign detect_max[50][7] = (mid_1[415:408] > top_2[415:408]) ? 1 : 0;
assign detect_max[50][8] = (mid_1[415:408] > top_2[423:416]) ? 1 : 0;
assign detect_max[50][9] = (mid_1[415:408] > mid_0[407:400]) ? 1 : 0;
assign detect_max[50][10] = (mid_1[415:408] > mid_0[415:408]) ? 1 : 0;
assign detect_max[50][11] = (mid_1[415:408] > mid_0[423:416]) ? 1 : 0;
assign detect_max[50][12] = (mid_1[415:408] > mid_1[407:400]) ? 1 : 0;
assign detect_max[50][13] = (mid_1[415:408] > mid_1[423:416]) ? 1 : 0;
assign detect_max[50][14] = (mid_1[415:408] > mid_2[407:400]) ? 1 : 0;
assign detect_max[50][15] = (mid_1[415:408] > mid_2[415:408]) ? 1 : 0;
assign detect_max[50][16] = (mid_1[415:408] > mid_2[423:416]) ? 1 : 0;
assign detect_max[50][17] = (mid_1[415:408] > btm_0[407:400]) ? 1 : 0;
assign detect_max[50][18] = (mid_1[415:408] > btm_0[415:408]) ? 1 : 0;
assign detect_max[50][19] = (mid_1[415:408] > btm_0[423:416]) ? 1 : 0;
assign detect_max[50][20] = (mid_1[415:408] > btm_1[407:400]) ? 1 : 0;
assign detect_max[50][21] = (mid_1[415:408] > btm_1[415:408]) ? 1 : 0;
assign detect_max[50][22] = (mid_1[415:408] > btm_1[423:416]) ? 1 : 0;
assign detect_max[50][23] = (mid_1[415:408] > btm_2[407:400]) ? 1 : 0;
assign detect_max[50][24] = (mid_1[415:408] > btm_2[415:408]) ? 1 : 0;
assign detect_max[50][25] = (mid_1[415:408] > btm_2[423:416]) ? 1 : 0;

assign detect_max[51][0] = (mid_1[423:416] > top_0[415:408]) ? 1 : 0;
assign detect_max[51][1] = (mid_1[423:416] > top_0[423:416]) ? 1 : 0;
assign detect_max[51][2] = (mid_1[423:416] > top_0[431:424]) ? 1 : 0;
assign detect_max[51][3] = (mid_1[423:416] > top_1[415:408]) ? 1 : 0;
assign detect_max[51][4] = (mid_1[423:416] > top_1[423:416]) ? 1 : 0;
assign detect_max[51][5] = (mid_1[423:416] > top_1[431:424]) ? 1 : 0;
assign detect_max[51][6] = (mid_1[423:416] > top_2[415:408]) ? 1 : 0;
assign detect_max[51][7] = (mid_1[423:416] > top_2[423:416]) ? 1 : 0;
assign detect_max[51][8] = (mid_1[423:416] > top_2[431:424]) ? 1 : 0;
assign detect_max[51][9] = (mid_1[423:416] > mid_0[415:408]) ? 1 : 0;
assign detect_max[51][10] = (mid_1[423:416] > mid_0[423:416]) ? 1 : 0;
assign detect_max[51][11] = (mid_1[423:416] > mid_0[431:424]) ? 1 : 0;
assign detect_max[51][12] = (mid_1[423:416] > mid_1[415:408]) ? 1 : 0;
assign detect_max[51][13] = (mid_1[423:416] > mid_1[431:424]) ? 1 : 0;
assign detect_max[51][14] = (mid_1[423:416] > mid_2[415:408]) ? 1 : 0;
assign detect_max[51][15] = (mid_1[423:416] > mid_2[423:416]) ? 1 : 0;
assign detect_max[51][16] = (mid_1[423:416] > mid_2[431:424]) ? 1 : 0;
assign detect_max[51][17] = (mid_1[423:416] > btm_0[415:408]) ? 1 : 0;
assign detect_max[51][18] = (mid_1[423:416] > btm_0[423:416]) ? 1 : 0;
assign detect_max[51][19] = (mid_1[423:416] > btm_0[431:424]) ? 1 : 0;
assign detect_max[51][20] = (mid_1[423:416] > btm_1[415:408]) ? 1 : 0;
assign detect_max[51][21] = (mid_1[423:416] > btm_1[423:416]) ? 1 : 0;
assign detect_max[51][22] = (mid_1[423:416] > btm_1[431:424]) ? 1 : 0;
assign detect_max[51][23] = (mid_1[423:416] > btm_2[415:408]) ? 1 : 0;
assign detect_max[51][24] = (mid_1[423:416] > btm_2[423:416]) ? 1 : 0;
assign detect_max[51][25] = (mid_1[423:416] > btm_2[431:424]) ? 1 : 0;

assign detect_max[52][0] = (mid_1[431:424] > top_0[423:416]) ? 1 : 0;
assign detect_max[52][1] = (mid_1[431:424] > top_0[431:424]) ? 1 : 0;
assign detect_max[52][2] = (mid_1[431:424] > top_0[439:432]) ? 1 : 0;
assign detect_max[52][3] = (mid_1[431:424] > top_1[423:416]) ? 1 : 0;
assign detect_max[52][4] = (mid_1[431:424] > top_1[431:424]) ? 1 : 0;
assign detect_max[52][5] = (mid_1[431:424] > top_1[439:432]) ? 1 : 0;
assign detect_max[52][6] = (mid_1[431:424] > top_2[423:416]) ? 1 : 0;
assign detect_max[52][7] = (mid_1[431:424] > top_2[431:424]) ? 1 : 0;
assign detect_max[52][8] = (mid_1[431:424] > top_2[439:432]) ? 1 : 0;
assign detect_max[52][9] = (mid_1[431:424] > mid_0[423:416]) ? 1 : 0;
assign detect_max[52][10] = (mid_1[431:424] > mid_0[431:424]) ? 1 : 0;
assign detect_max[52][11] = (mid_1[431:424] > mid_0[439:432]) ? 1 : 0;
assign detect_max[52][12] = (mid_1[431:424] > mid_1[423:416]) ? 1 : 0;
assign detect_max[52][13] = (mid_1[431:424] > mid_1[439:432]) ? 1 : 0;
assign detect_max[52][14] = (mid_1[431:424] > mid_2[423:416]) ? 1 : 0;
assign detect_max[52][15] = (mid_1[431:424] > mid_2[431:424]) ? 1 : 0;
assign detect_max[52][16] = (mid_1[431:424] > mid_2[439:432]) ? 1 : 0;
assign detect_max[52][17] = (mid_1[431:424] > btm_0[423:416]) ? 1 : 0;
assign detect_max[52][18] = (mid_1[431:424] > btm_0[431:424]) ? 1 : 0;
assign detect_max[52][19] = (mid_1[431:424] > btm_0[439:432]) ? 1 : 0;
assign detect_max[52][20] = (mid_1[431:424] > btm_1[423:416]) ? 1 : 0;
assign detect_max[52][21] = (mid_1[431:424] > btm_1[431:424]) ? 1 : 0;
assign detect_max[52][22] = (mid_1[431:424] > btm_1[439:432]) ? 1 : 0;
assign detect_max[52][23] = (mid_1[431:424] > btm_2[423:416]) ? 1 : 0;
assign detect_max[52][24] = (mid_1[431:424] > btm_2[431:424]) ? 1 : 0;
assign detect_max[52][25] = (mid_1[431:424] > btm_2[439:432]) ? 1 : 0;

assign detect_max[53][0] = (mid_1[439:432] > top_0[431:424]) ? 1 : 0;
assign detect_max[53][1] = (mid_1[439:432] > top_0[439:432]) ? 1 : 0;
assign detect_max[53][2] = (mid_1[439:432] > top_0[447:440]) ? 1 : 0;
assign detect_max[53][3] = (mid_1[439:432] > top_1[431:424]) ? 1 : 0;
assign detect_max[53][4] = (mid_1[439:432] > top_1[439:432]) ? 1 : 0;
assign detect_max[53][5] = (mid_1[439:432] > top_1[447:440]) ? 1 : 0;
assign detect_max[53][6] = (mid_1[439:432] > top_2[431:424]) ? 1 : 0;
assign detect_max[53][7] = (mid_1[439:432] > top_2[439:432]) ? 1 : 0;
assign detect_max[53][8] = (mid_1[439:432] > top_2[447:440]) ? 1 : 0;
assign detect_max[53][9] = (mid_1[439:432] > mid_0[431:424]) ? 1 : 0;
assign detect_max[53][10] = (mid_1[439:432] > mid_0[439:432]) ? 1 : 0;
assign detect_max[53][11] = (mid_1[439:432] > mid_0[447:440]) ? 1 : 0;
assign detect_max[53][12] = (mid_1[439:432] > mid_1[431:424]) ? 1 : 0;
assign detect_max[53][13] = (mid_1[439:432] > mid_1[447:440]) ? 1 : 0;
assign detect_max[53][14] = (mid_1[439:432] > mid_2[431:424]) ? 1 : 0;
assign detect_max[53][15] = (mid_1[439:432] > mid_2[439:432]) ? 1 : 0;
assign detect_max[53][16] = (mid_1[439:432] > mid_2[447:440]) ? 1 : 0;
assign detect_max[53][17] = (mid_1[439:432] > btm_0[431:424]) ? 1 : 0;
assign detect_max[53][18] = (mid_1[439:432] > btm_0[439:432]) ? 1 : 0;
assign detect_max[53][19] = (mid_1[439:432] > btm_0[447:440]) ? 1 : 0;
assign detect_max[53][20] = (mid_1[439:432] > btm_1[431:424]) ? 1 : 0;
assign detect_max[53][21] = (mid_1[439:432] > btm_1[439:432]) ? 1 : 0;
assign detect_max[53][22] = (mid_1[439:432] > btm_1[447:440]) ? 1 : 0;
assign detect_max[53][23] = (mid_1[439:432] > btm_2[431:424]) ? 1 : 0;
assign detect_max[53][24] = (mid_1[439:432] > btm_2[439:432]) ? 1 : 0;
assign detect_max[53][25] = (mid_1[439:432] > btm_2[447:440]) ? 1 : 0;

assign detect_max[54][0] = (mid_1[447:440] > top_0[439:432]) ? 1 : 0;
assign detect_max[54][1] = (mid_1[447:440] > top_0[447:440]) ? 1 : 0;
assign detect_max[54][2] = (mid_1[447:440] > top_0[455:448]) ? 1 : 0;
assign detect_max[54][3] = (mid_1[447:440] > top_1[439:432]) ? 1 : 0;
assign detect_max[54][4] = (mid_1[447:440] > top_1[447:440]) ? 1 : 0;
assign detect_max[54][5] = (mid_1[447:440] > top_1[455:448]) ? 1 : 0;
assign detect_max[54][6] = (mid_1[447:440] > top_2[439:432]) ? 1 : 0;
assign detect_max[54][7] = (mid_1[447:440] > top_2[447:440]) ? 1 : 0;
assign detect_max[54][8] = (mid_1[447:440] > top_2[455:448]) ? 1 : 0;
assign detect_max[54][9] = (mid_1[447:440] > mid_0[439:432]) ? 1 : 0;
assign detect_max[54][10] = (mid_1[447:440] > mid_0[447:440]) ? 1 : 0;
assign detect_max[54][11] = (mid_1[447:440] > mid_0[455:448]) ? 1 : 0;
assign detect_max[54][12] = (mid_1[447:440] > mid_1[439:432]) ? 1 : 0;
assign detect_max[54][13] = (mid_1[447:440] > mid_1[455:448]) ? 1 : 0;
assign detect_max[54][14] = (mid_1[447:440] > mid_2[439:432]) ? 1 : 0;
assign detect_max[54][15] = (mid_1[447:440] > mid_2[447:440]) ? 1 : 0;
assign detect_max[54][16] = (mid_1[447:440] > mid_2[455:448]) ? 1 : 0;
assign detect_max[54][17] = (mid_1[447:440] > btm_0[439:432]) ? 1 : 0;
assign detect_max[54][18] = (mid_1[447:440] > btm_0[447:440]) ? 1 : 0;
assign detect_max[54][19] = (mid_1[447:440] > btm_0[455:448]) ? 1 : 0;
assign detect_max[54][20] = (mid_1[447:440] > btm_1[439:432]) ? 1 : 0;
assign detect_max[54][21] = (mid_1[447:440] > btm_1[447:440]) ? 1 : 0;
assign detect_max[54][22] = (mid_1[447:440] > btm_1[455:448]) ? 1 : 0;
assign detect_max[54][23] = (mid_1[447:440] > btm_2[439:432]) ? 1 : 0;
assign detect_max[54][24] = (mid_1[447:440] > btm_2[447:440]) ? 1 : 0;
assign detect_max[54][25] = (mid_1[447:440] > btm_2[455:448]) ? 1 : 0;

assign detect_max[55][0] = (mid_1[455:448] > top_0[447:440]) ? 1 : 0;
assign detect_max[55][1] = (mid_1[455:448] > top_0[455:448]) ? 1 : 0;
assign detect_max[55][2] = (mid_1[455:448] > top_0[463:456]) ? 1 : 0;
assign detect_max[55][3] = (mid_1[455:448] > top_1[447:440]) ? 1 : 0;
assign detect_max[55][4] = (mid_1[455:448] > top_1[455:448]) ? 1 : 0;
assign detect_max[55][5] = (mid_1[455:448] > top_1[463:456]) ? 1 : 0;
assign detect_max[55][6] = (mid_1[455:448] > top_2[447:440]) ? 1 : 0;
assign detect_max[55][7] = (mid_1[455:448] > top_2[455:448]) ? 1 : 0;
assign detect_max[55][8] = (mid_1[455:448] > top_2[463:456]) ? 1 : 0;
assign detect_max[55][9] = (mid_1[455:448] > mid_0[447:440]) ? 1 : 0;
assign detect_max[55][10] = (mid_1[455:448] > mid_0[455:448]) ? 1 : 0;
assign detect_max[55][11] = (mid_1[455:448] > mid_0[463:456]) ? 1 : 0;
assign detect_max[55][12] = (mid_1[455:448] > mid_1[447:440]) ? 1 : 0;
assign detect_max[55][13] = (mid_1[455:448] > mid_1[463:456]) ? 1 : 0;
assign detect_max[55][14] = (mid_1[455:448] > mid_2[447:440]) ? 1 : 0;
assign detect_max[55][15] = (mid_1[455:448] > mid_2[455:448]) ? 1 : 0;
assign detect_max[55][16] = (mid_1[455:448] > mid_2[463:456]) ? 1 : 0;
assign detect_max[55][17] = (mid_1[455:448] > btm_0[447:440]) ? 1 : 0;
assign detect_max[55][18] = (mid_1[455:448] > btm_0[455:448]) ? 1 : 0;
assign detect_max[55][19] = (mid_1[455:448] > btm_0[463:456]) ? 1 : 0;
assign detect_max[55][20] = (mid_1[455:448] > btm_1[447:440]) ? 1 : 0;
assign detect_max[55][21] = (mid_1[455:448] > btm_1[455:448]) ? 1 : 0;
assign detect_max[55][22] = (mid_1[455:448] > btm_1[463:456]) ? 1 : 0;
assign detect_max[55][23] = (mid_1[455:448] > btm_2[447:440]) ? 1 : 0;
assign detect_max[55][24] = (mid_1[455:448] > btm_2[455:448]) ? 1 : 0;
assign detect_max[55][25] = (mid_1[455:448] > btm_2[463:456]) ? 1 : 0;

assign detect_max[56][0] = (mid_1[463:456] > top_0[455:448]) ? 1 : 0;
assign detect_max[56][1] = (mid_1[463:456] > top_0[463:456]) ? 1 : 0;
assign detect_max[56][2] = (mid_1[463:456] > top_0[471:464]) ? 1 : 0;
assign detect_max[56][3] = (mid_1[463:456] > top_1[455:448]) ? 1 : 0;
assign detect_max[56][4] = (mid_1[463:456] > top_1[463:456]) ? 1 : 0;
assign detect_max[56][5] = (mid_1[463:456] > top_1[471:464]) ? 1 : 0;
assign detect_max[56][6] = (mid_1[463:456] > top_2[455:448]) ? 1 : 0;
assign detect_max[56][7] = (mid_1[463:456] > top_2[463:456]) ? 1 : 0;
assign detect_max[56][8] = (mid_1[463:456] > top_2[471:464]) ? 1 : 0;
assign detect_max[56][9] = (mid_1[463:456] > mid_0[455:448]) ? 1 : 0;
assign detect_max[56][10] = (mid_1[463:456] > mid_0[463:456]) ? 1 : 0;
assign detect_max[56][11] = (mid_1[463:456] > mid_0[471:464]) ? 1 : 0;
assign detect_max[56][12] = (mid_1[463:456] > mid_1[455:448]) ? 1 : 0;
assign detect_max[56][13] = (mid_1[463:456] > mid_1[471:464]) ? 1 : 0;
assign detect_max[56][14] = (mid_1[463:456] > mid_2[455:448]) ? 1 : 0;
assign detect_max[56][15] = (mid_1[463:456] > mid_2[463:456]) ? 1 : 0;
assign detect_max[56][16] = (mid_1[463:456] > mid_2[471:464]) ? 1 : 0;
assign detect_max[56][17] = (mid_1[463:456] > btm_0[455:448]) ? 1 : 0;
assign detect_max[56][18] = (mid_1[463:456] > btm_0[463:456]) ? 1 : 0;
assign detect_max[56][19] = (mid_1[463:456] > btm_0[471:464]) ? 1 : 0;
assign detect_max[56][20] = (mid_1[463:456] > btm_1[455:448]) ? 1 : 0;
assign detect_max[56][21] = (mid_1[463:456] > btm_1[463:456]) ? 1 : 0;
assign detect_max[56][22] = (mid_1[463:456] > btm_1[471:464]) ? 1 : 0;
assign detect_max[56][23] = (mid_1[463:456] > btm_2[455:448]) ? 1 : 0;
assign detect_max[56][24] = (mid_1[463:456] > btm_2[463:456]) ? 1 : 0;
assign detect_max[56][25] = (mid_1[463:456] > btm_2[471:464]) ? 1 : 0;

assign detect_max[57][0] = (mid_1[471:464] > top_0[463:456]) ? 1 : 0;
assign detect_max[57][1] = (mid_1[471:464] > top_0[471:464]) ? 1 : 0;
assign detect_max[57][2] = (mid_1[471:464] > top_0[479:472]) ? 1 : 0;
assign detect_max[57][3] = (mid_1[471:464] > top_1[463:456]) ? 1 : 0;
assign detect_max[57][4] = (mid_1[471:464] > top_1[471:464]) ? 1 : 0;
assign detect_max[57][5] = (mid_1[471:464] > top_1[479:472]) ? 1 : 0;
assign detect_max[57][6] = (mid_1[471:464] > top_2[463:456]) ? 1 : 0;
assign detect_max[57][7] = (mid_1[471:464] > top_2[471:464]) ? 1 : 0;
assign detect_max[57][8] = (mid_1[471:464] > top_2[479:472]) ? 1 : 0;
assign detect_max[57][9] = (mid_1[471:464] > mid_0[463:456]) ? 1 : 0;
assign detect_max[57][10] = (mid_1[471:464] > mid_0[471:464]) ? 1 : 0;
assign detect_max[57][11] = (mid_1[471:464] > mid_0[479:472]) ? 1 : 0;
assign detect_max[57][12] = (mid_1[471:464] > mid_1[463:456]) ? 1 : 0;
assign detect_max[57][13] = (mid_1[471:464] > mid_1[479:472]) ? 1 : 0;
assign detect_max[57][14] = (mid_1[471:464] > mid_2[463:456]) ? 1 : 0;
assign detect_max[57][15] = (mid_1[471:464] > mid_2[471:464]) ? 1 : 0;
assign detect_max[57][16] = (mid_1[471:464] > mid_2[479:472]) ? 1 : 0;
assign detect_max[57][17] = (mid_1[471:464] > btm_0[463:456]) ? 1 : 0;
assign detect_max[57][18] = (mid_1[471:464] > btm_0[471:464]) ? 1 : 0;
assign detect_max[57][19] = (mid_1[471:464] > btm_0[479:472]) ? 1 : 0;
assign detect_max[57][20] = (mid_1[471:464] > btm_1[463:456]) ? 1 : 0;
assign detect_max[57][21] = (mid_1[471:464] > btm_1[471:464]) ? 1 : 0;
assign detect_max[57][22] = (mid_1[471:464] > btm_1[479:472]) ? 1 : 0;
assign detect_max[57][23] = (mid_1[471:464] > btm_2[463:456]) ? 1 : 0;
assign detect_max[57][24] = (mid_1[471:464] > btm_2[471:464]) ? 1 : 0;
assign detect_max[57][25] = (mid_1[471:464] > btm_2[479:472]) ? 1 : 0;

assign detect_max[58][0] = (mid_1[479:472] > top_0[471:464]) ? 1 : 0;
assign detect_max[58][1] = (mid_1[479:472] > top_0[479:472]) ? 1 : 0;
assign detect_max[58][2] = (mid_1[479:472] > top_0[487:480]) ? 1 : 0;
assign detect_max[58][3] = (mid_1[479:472] > top_1[471:464]) ? 1 : 0;
assign detect_max[58][4] = (mid_1[479:472] > top_1[479:472]) ? 1 : 0;
assign detect_max[58][5] = (mid_1[479:472] > top_1[487:480]) ? 1 : 0;
assign detect_max[58][6] = (mid_1[479:472] > top_2[471:464]) ? 1 : 0;
assign detect_max[58][7] = (mid_1[479:472] > top_2[479:472]) ? 1 : 0;
assign detect_max[58][8] = (mid_1[479:472] > top_2[487:480]) ? 1 : 0;
assign detect_max[58][9] = (mid_1[479:472] > mid_0[471:464]) ? 1 : 0;
assign detect_max[58][10] = (mid_1[479:472] > mid_0[479:472]) ? 1 : 0;
assign detect_max[58][11] = (mid_1[479:472] > mid_0[487:480]) ? 1 : 0;
assign detect_max[58][12] = (mid_1[479:472] > mid_1[471:464]) ? 1 : 0;
assign detect_max[58][13] = (mid_1[479:472] > mid_1[487:480]) ? 1 : 0;
assign detect_max[58][14] = (mid_1[479:472] > mid_2[471:464]) ? 1 : 0;
assign detect_max[58][15] = (mid_1[479:472] > mid_2[479:472]) ? 1 : 0;
assign detect_max[58][16] = (mid_1[479:472] > mid_2[487:480]) ? 1 : 0;
assign detect_max[58][17] = (mid_1[479:472] > btm_0[471:464]) ? 1 : 0;
assign detect_max[58][18] = (mid_1[479:472] > btm_0[479:472]) ? 1 : 0;
assign detect_max[58][19] = (mid_1[479:472] > btm_0[487:480]) ? 1 : 0;
assign detect_max[58][20] = (mid_1[479:472] > btm_1[471:464]) ? 1 : 0;
assign detect_max[58][21] = (mid_1[479:472] > btm_1[479:472]) ? 1 : 0;
assign detect_max[58][22] = (mid_1[479:472] > btm_1[487:480]) ? 1 : 0;
assign detect_max[58][23] = (mid_1[479:472] > btm_2[471:464]) ? 1 : 0;
assign detect_max[58][24] = (mid_1[479:472] > btm_2[479:472]) ? 1 : 0;
assign detect_max[58][25] = (mid_1[479:472] > btm_2[487:480]) ? 1 : 0;

assign detect_max[59][0] = (mid_1[487:480] > top_0[479:472]) ? 1 : 0;
assign detect_max[59][1] = (mid_1[487:480] > top_0[487:480]) ? 1 : 0;
assign detect_max[59][2] = (mid_1[487:480] > top_0[495:488]) ? 1 : 0;
assign detect_max[59][3] = (mid_1[487:480] > top_1[479:472]) ? 1 : 0;
assign detect_max[59][4] = (mid_1[487:480] > top_1[487:480]) ? 1 : 0;
assign detect_max[59][5] = (mid_1[487:480] > top_1[495:488]) ? 1 : 0;
assign detect_max[59][6] = (mid_1[487:480] > top_2[479:472]) ? 1 : 0;
assign detect_max[59][7] = (mid_1[487:480] > top_2[487:480]) ? 1 : 0;
assign detect_max[59][8] = (mid_1[487:480] > top_2[495:488]) ? 1 : 0;
assign detect_max[59][9] = (mid_1[487:480] > mid_0[479:472]) ? 1 : 0;
assign detect_max[59][10] = (mid_1[487:480] > mid_0[487:480]) ? 1 : 0;
assign detect_max[59][11] = (mid_1[487:480] > mid_0[495:488]) ? 1 : 0;
assign detect_max[59][12] = (mid_1[487:480] > mid_1[479:472]) ? 1 : 0;
assign detect_max[59][13] = (mid_1[487:480] > mid_1[495:488]) ? 1 : 0;
assign detect_max[59][14] = (mid_1[487:480] > mid_2[479:472]) ? 1 : 0;
assign detect_max[59][15] = (mid_1[487:480] > mid_2[487:480]) ? 1 : 0;
assign detect_max[59][16] = (mid_1[487:480] > mid_2[495:488]) ? 1 : 0;
assign detect_max[59][17] = (mid_1[487:480] > btm_0[479:472]) ? 1 : 0;
assign detect_max[59][18] = (mid_1[487:480] > btm_0[487:480]) ? 1 : 0;
assign detect_max[59][19] = (mid_1[487:480] > btm_0[495:488]) ? 1 : 0;
assign detect_max[59][20] = (mid_1[487:480] > btm_1[479:472]) ? 1 : 0;
assign detect_max[59][21] = (mid_1[487:480] > btm_1[487:480]) ? 1 : 0;
assign detect_max[59][22] = (mid_1[487:480] > btm_1[495:488]) ? 1 : 0;
assign detect_max[59][23] = (mid_1[487:480] > btm_2[479:472]) ? 1 : 0;
assign detect_max[59][24] = (mid_1[487:480] > btm_2[487:480]) ? 1 : 0;
assign detect_max[59][25] = (mid_1[487:480] > btm_2[495:488]) ? 1 : 0;

assign detect_max[60][0] = (mid_1[495:488] > top_0[487:480]) ? 1 : 0;
assign detect_max[60][1] = (mid_1[495:488] > top_0[495:488]) ? 1 : 0;
assign detect_max[60][2] = (mid_1[495:488] > top_0[503:496]) ? 1 : 0;
assign detect_max[60][3] = (mid_1[495:488] > top_1[487:480]) ? 1 : 0;
assign detect_max[60][4] = (mid_1[495:488] > top_1[495:488]) ? 1 : 0;
assign detect_max[60][5] = (mid_1[495:488] > top_1[503:496]) ? 1 : 0;
assign detect_max[60][6] = (mid_1[495:488] > top_2[487:480]) ? 1 : 0;
assign detect_max[60][7] = (mid_1[495:488] > top_2[495:488]) ? 1 : 0;
assign detect_max[60][8] = (mid_1[495:488] > top_2[503:496]) ? 1 : 0;
assign detect_max[60][9] = (mid_1[495:488] > mid_0[487:480]) ? 1 : 0;
assign detect_max[60][10] = (mid_1[495:488] > mid_0[495:488]) ? 1 : 0;
assign detect_max[60][11] = (mid_1[495:488] > mid_0[503:496]) ? 1 : 0;
assign detect_max[60][12] = (mid_1[495:488] > mid_1[487:480]) ? 1 : 0;
assign detect_max[60][13] = (mid_1[495:488] > mid_1[503:496]) ? 1 : 0;
assign detect_max[60][14] = (mid_1[495:488] > mid_2[487:480]) ? 1 : 0;
assign detect_max[60][15] = (mid_1[495:488] > mid_2[495:488]) ? 1 : 0;
assign detect_max[60][16] = (mid_1[495:488] > mid_2[503:496]) ? 1 : 0;
assign detect_max[60][17] = (mid_1[495:488] > btm_0[487:480]) ? 1 : 0;
assign detect_max[60][18] = (mid_1[495:488] > btm_0[495:488]) ? 1 : 0;
assign detect_max[60][19] = (mid_1[495:488] > btm_0[503:496]) ? 1 : 0;
assign detect_max[60][20] = (mid_1[495:488] > btm_1[487:480]) ? 1 : 0;
assign detect_max[60][21] = (mid_1[495:488] > btm_1[495:488]) ? 1 : 0;
assign detect_max[60][22] = (mid_1[495:488] > btm_1[503:496]) ? 1 : 0;
assign detect_max[60][23] = (mid_1[495:488] > btm_2[487:480]) ? 1 : 0;
assign detect_max[60][24] = (mid_1[495:488] > btm_2[495:488]) ? 1 : 0;
assign detect_max[60][25] = (mid_1[495:488] > btm_2[503:496]) ? 1 : 0;

assign detect_max[61][0] = (mid_1[503:496] > top_0[495:488]) ? 1 : 0;
assign detect_max[61][1] = (mid_1[503:496] > top_0[503:496]) ? 1 : 0;
assign detect_max[61][2] = (mid_1[503:496] > top_0[511:504]) ? 1 : 0;
assign detect_max[61][3] = (mid_1[503:496] > top_1[495:488]) ? 1 : 0;
assign detect_max[61][4] = (mid_1[503:496] > top_1[503:496]) ? 1 : 0;
assign detect_max[61][5] = (mid_1[503:496] > top_1[511:504]) ? 1 : 0;
assign detect_max[61][6] = (mid_1[503:496] > top_2[495:488]) ? 1 : 0;
assign detect_max[61][7] = (mid_1[503:496] > top_2[503:496]) ? 1 : 0;
assign detect_max[61][8] = (mid_1[503:496] > top_2[511:504]) ? 1 : 0;
assign detect_max[61][9] = (mid_1[503:496] > mid_0[495:488]) ? 1 : 0;
assign detect_max[61][10] = (mid_1[503:496] > mid_0[503:496]) ? 1 : 0;
assign detect_max[61][11] = (mid_1[503:496] > mid_0[511:504]) ? 1 : 0;
assign detect_max[61][12] = (mid_1[503:496] > mid_1[495:488]) ? 1 : 0;
assign detect_max[61][13] = (mid_1[503:496] > mid_1[511:504]) ? 1 : 0;
assign detect_max[61][14] = (mid_1[503:496] > mid_2[495:488]) ? 1 : 0;
assign detect_max[61][15] = (mid_1[503:496] > mid_2[503:496]) ? 1 : 0;
assign detect_max[61][16] = (mid_1[503:496] > mid_2[511:504]) ? 1 : 0;
assign detect_max[61][17] = (mid_1[503:496] > btm_0[495:488]) ? 1 : 0;
assign detect_max[61][18] = (mid_1[503:496] > btm_0[503:496]) ? 1 : 0;
assign detect_max[61][19] = (mid_1[503:496] > btm_0[511:504]) ? 1 : 0;
assign detect_max[61][20] = (mid_1[503:496] > btm_1[495:488]) ? 1 : 0;
assign detect_max[61][21] = (mid_1[503:496] > btm_1[503:496]) ? 1 : 0;
assign detect_max[61][22] = (mid_1[503:496] > btm_1[511:504]) ? 1 : 0;
assign detect_max[61][23] = (mid_1[503:496] > btm_2[495:488]) ? 1 : 0;
assign detect_max[61][24] = (mid_1[503:496] > btm_2[503:496]) ? 1 : 0;
assign detect_max[61][25] = (mid_1[503:496] > btm_2[511:504]) ? 1 : 0;

assign detect_max[62][0] = (mid_1[511:504] > top_0[503:496]) ? 1 : 0;
assign detect_max[62][1] = (mid_1[511:504] > top_0[511:504]) ? 1 : 0;
assign detect_max[62][2] = (mid_1[511:504] > top_0[519:512]) ? 1 : 0;
assign detect_max[62][3] = (mid_1[511:504] > top_1[503:496]) ? 1 : 0;
assign detect_max[62][4] = (mid_1[511:504] > top_1[511:504]) ? 1 : 0;
assign detect_max[62][5] = (mid_1[511:504] > top_1[519:512]) ? 1 : 0;
assign detect_max[62][6] = (mid_1[511:504] > top_2[503:496]) ? 1 : 0;
assign detect_max[62][7] = (mid_1[511:504] > top_2[511:504]) ? 1 : 0;
assign detect_max[62][8] = (mid_1[511:504] > top_2[519:512]) ? 1 : 0;
assign detect_max[62][9] = (mid_1[511:504] > mid_0[503:496]) ? 1 : 0;
assign detect_max[62][10] = (mid_1[511:504] > mid_0[511:504]) ? 1 : 0;
assign detect_max[62][11] = (mid_1[511:504] > mid_0[519:512]) ? 1 : 0;
assign detect_max[62][12] = (mid_1[511:504] > mid_1[503:496]) ? 1 : 0;
assign detect_max[62][13] = (mid_1[511:504] > mid_1[519:512]) ? 1 : 0;
assign detect_max[62][14] = (mid_1[511:504] > mid_2[503:496]) ? 1 : 0;
assign detect_max[62][15] = (mid_1[511:504] > mid_2[511:504]) ? 1 : 0;
assign detect_max[62][16] = (mid_1[511:504] > mid_2[519:512]) ? 1 : 0;
assign detect_max[62][17] = (mid_1[511:504] > btm_0[503:496]) ? 1 : 0;
assign detect_max[62][18] = (mid_1[511:504] > btm_0[511:504]) ? 1 : 0;
assign detect_max[62][19] = (mid_1[511:504] > btm_0[519:512]) ? 1 : 0;
assign detect_max[62][20] = (mid_1[511:504] > btm_1[503:496]) ? 1 : 0;
assign detect_max[62][21] = (mid_1[511:504] > btm_1[511:504]) ? 1 : 0;
assign detect_max[62][22] = (mid_1[511:504] > btm_1[519:512]) ? 1 : 0;
assign detect_max[62][23] = (mid_1[511:504] > btm_2[503:496]) ? 1 : 0;
assign detect_max[62][24] = (mid_1[511:504] > btm_2[511:504]) ? 1 : 0;
assign detect_max[62][25] = (mid_1[511:504] > btm_2[519:512]) ? 1 : 0;

assign detect_max[63][0] = (mid_1[519:512] > top_0[511:504]) ? 1 : 0;
assign detect_max[63][1] = (mid_1[519:512] > top_0[519:512]) ? 1 : 0;
assign detect_max[63][2] = (mid_1[519:512] > top_0[527:520]) ? 1 : 0;
assign detect_max[63][3] = (mid_1[519:512] > top_1[511:504]) ? 1 : 0;
assign detect_max[63][4] = (mid_1[519:512] > top_1[519:512]) ? 1 : 0;
assign detect_max[63][5] = (mid_1[519:512] > top_1[527:520]) ? 1 : 0;
assign detect_max[63][6] = (mid_1[519:512] > top_2[511:504]) ? 1 : 0;
assign detect_max[63][7] = (mid_1[519:512] > top_2[519:512]) ? 1 : 0;
assign detect_max[63][8] = (mid_1[519:512] > top_2[527:520]) ? 1 : 0;
assign detect_max[63][9] = (mid_1[519:512] > mid_0[511:504]) ? 1 : 0;
assign detect_max[63][10] = (mid_1[519:512] > mid_0[519:512]) ? 1 : 0;
assign detect_max[63][11] = (mid_1[519:512] > mid_0[527:520]) ? 1 : 0;
assign detect_max[63][12] = (mid_1[519:512] > mid_1[511:504]) ? 1 : 0;
assign detect_max[63][13] = (mid_1[519:512] > mid_1[527:520]) ? 1 : 0;
assign detect_max[63][14] = (mid_1[519:512] > mid_2[511:504]) ? 1 : 0;
assign detect_max[63][15] = (mid_1[519:512] > mid_2[519:512]) ? 1 : 0;
assign detect_max[63][16] = (mid_1[519:512] > mid_2[527:520]) ? 1 : 0;
assign detect_max[63][17] = (mid_1[519:512] > btm_0[511:504]) ? 1 : 0;
assign detect_max[63][18] = (mid_1[519:512] > btm_0[519:512]) ? 1 : 0;
assign detect_max[63][19] = (mid_1[519:512] > btm_0[527:520]) ? 1 : 0;
assign detect_max[63][20] = (mid_1[519:512] > btm_1[511:504]) ? 1 : 0;
assign detect_max[63][21] = (mid_1[519:512] > btm_1[519:512]) ? 1 : 0;
assign detect_max[63][22] = (mid_1[519:512] > btm_1[527:520]) ? 1 : 0;
assign detect_max[63][23] = (mid_1[519:512] > btm_2[511:504]) ? 1 : 0;
assign detect_max[63][24] = (mid_1[519:512] > btm_2[519:512]) ? 1 : 0;
assign detect_max[63][25] = (mid_1[519:512] > btm_2[527:520]) ? 1 : 0;

assign detect_max[64][0] = (mid_1[527:520] > top_0[519:512]) ? 1 : 0;
assign detect_max[64][1] = (mid_1[527:520] > top_0[527:520]) ? 1 : 0;
assign detect_max[64][2] = (mid_1[527:520] > top_0[535:528]) ? 1 : 0;
assign detect_max[64][3] = (mid_1[527:520] > top_1[519:512]) ? 1 : 0;
assign detect_max[64][4] = (mid_1[527:520] > top_1[527:520]) ? 1 : 0;
assign detect_max[64][5] = (mid_1[527:520] > top_1[535:528]) ? 1 : 0;
assign detect_max[64][6] = (mid_1[527:520] > top_2[519:512]) ? 1 : 0;
assign detect_max[64][7] = (mid_1[527:520] > top_2[527:520]) ? 1 : 0;
assign detect_max[64][8] = (mid_1[527:520] > top_2[535:528]) ? 1 : 0;
assign detect_max[64][9] = (mid_1[527:520] > mid_0[519:512]) ? 1 : 0;
assign detect_max[64][10] = (mid_1[527:520] > mid_0[527:520]) ? 1 : 0;
assign detect_max[64][11] = (mid_1[527:520] > mid_0[535:528]) ? 1 : 0;
assign detect_max[64][12] = (mid_1[527:520] > mid_1[519:512]) ? 1 : 0;
assign detect_max[64][13] = (mid_1[527:520] > mid_1[535:528]) ? 1 : 0;
assign detect_max[64][14] = (mid_1[527:520] > mid_2[519:512]) ? 1 : 0;
assign detect_max[64][15] = (mid_1[527:520] > mid_2[527:520]) ? 1 : 0;
assign detect_max[64][16] = (mid_1[527:520] > mid_2[535:528]) ? 1 : 0;
assign detect_max[64][17] = (mid_1[527:520] > btm_0[519:512]) ? 1 : 0;
assign detect_max[64][18] = (mid_1[527:520] > btm_0[527:520]) ? 1 : 0;
assign detect_max[64][19] = (mid_1[527:520] > btm_0[535:528]) ? 1 : 0;
assign detect_max[64][20] = (mid_1[527:520] > btm_1[519:512]) ? 1 : 0;
assign detect_max[64][21] = (mid_1[527:520] > btm_1[527:520]) ? 1 : 0;
assign detect_max[64][22] = (mid_1[527:520] > btm_1[535:528]) ? 1 : 0;
assign detect_max[64][23] = (mid_1[527:520] > btm_2[519:512]) ? 1 : 0;
assign detect_max[64][24] = (mid_1[527:520] > btm_2[527:520]) ? 1 : 0;
assign detect_max[64][25] = (mid_1[527:520] > btm_2[535:528]) ? 1 : 0;

assign detect_max[65][0] = (mid_1[535:528] > top_0[527:520]) ? 1 : 0;
assign detect_max[65][1] = (mid_1[535:528] > top_0[535:528]) ? 1 : 0;
assign detect_max[65][2] = (mid_1[535:528] > top_0[543:536]) ? 1 : 0;
assign detect_max[65][3] = (mid_1[535:528] > top_1[527:520]) ? 1 : 0;
assign detect_max[65][4] = (mid_1[535:528] > top_1[535:528]) ? 1 : 0;
assign detect_max[65][5] = (mid_1[535:528] > top_1[543:536]) ? 1 : 0;
assign detect_max[65][6] = (mid_1[535:528] > top_2[527:520]) ? 1 : 0;
assign detect_max[65][7] = (mid_1[535:528] > top_2[535:528]) ? 1 : 0;
assign detect_max[65][8] = (mid_1[535:528] > top_2[543:536]) ? 1 : 0;
assign detect_max[65][9] = (mid_1[535:528] > mid_0[527:520]) ? 1 : 0;
assign detect_max[65][10] = (mid_1[535:528] > mid_0[535:528]) ? 1 : 0;
assign detect_max[65][11] = (mid_1[535:528] > mid_0[543:536]) ? 1 : 0;
assign detect_max[65][12] = (mid_1[535:528] > mid_1[527:520]) ? 1 : 0;
assign detect_max[65][13] = (mid_1[535:528] > mid_1[543:536]) ? 1 : 0;
assign detect_max[65][14] = (mid_1[535:528] > mid_2[527:520]) ? 1 : 0;
assign detect_max[65][15] = (mid_1[535:528] > mid_2[535:528]) ? 1 : 0;
assign detect_max[65][16] = (mid_1[535:528] > mid_2[543:536]) ? 1 : 0;
assign detect_max[65][17] = (mid_1[535:528] > btm_0[527:520]) ? 1 : 0;
assign detect_max[65][18] = (mid_1[535:528] > btm_0[535:528]) ? 1 : 0;
assign detect_max[65][19] = (mid_1[535:528] > btm_0[543:536]) ? 1 : 0;
assign detect_max[65][20] = (mid_1[535:528] > btm_1[527:520]) ? 1 : 0;
assign detect_max[65][21] = (mid_1[535:528] > btm_1[535:528]) ? 1 : 0;
assign detect_max[65][22] = (mid_1[535:528] > btm_1[543:536]) ? 1 : 0;
assign detect_max[65][23] = (mid_1[535:528] > btm_2[527:520]) ? 1 : 0;
assign detect_max[65][24] = (mid_1[535:528] > btm_2[535:528]) ? 1 : 0;
assign detect_max[65][25] = (mid_1[535:528] > btm_2[543:536]) ? 1 : 0;

assign detect_max[66][0] = (mid_1[543:536] > top_0[535:528]) ? 1 : 0;
assign detect_max[66][1] = (mid_1[543:536] > top_0[543:536]) ? 1 : 0;
assign detect_max[66][2] = (mid_1[543:536] > top_0[551:544]) ? 1 : 0;
assign detect_max[66][3] = (mid_1[543:536] > top_1[535:528]) ? 1 : 0;
assign detect_max[66][4] = (mid_1[543:536] > top_1[543:536]) ? 1 : 0;
assign detect_max[66][5] = (mid_1[543:536] > top_1[551:544]) ? 1 : 0;
assign detect_max[66][6] = (mid_1[543:536] > top_2[535:528]) ? 1 : 0;
assign detect_max[66][7] = (mid_1[543:536] > top_2[543:536]) ? 1 : 0;
assign detect_max[66][8] = (mid_1[543:536] > top_2[551:544]) ? 1 : 0;
assign detect_max[66][9] = (mid_1[543:536] > mid_0[535:528]) ? 1 : 0;
assign detect_max[66][10] = (mid_1[543:536] > mid_0[543:536]) ? 1 : 0;
assign detect_max[66][11] = (mid_1[543:536] > mid_0[551:544]) ? 1 : 0;
assign detect_max[66][12] = (mid_1[543:536] > mid_1[535:528]) ? 1 : 0;
assign detect_max[66][13] = (mid_1[543:536] > mid_1[551:544]) ? 1 : 0;
assign detect_max[66][14] = (mid_1[543:536] > mid_2[535:528]) ? 1 : 0;
assign detect_max[66][15] = (mid_1[543:536] > mid_2[543:536]) ? 1 : 0;
assign detect_max[66][16] = (mid_1[543:536] > mid_2[551:544]) ? 1 : 0;
assign detect_max[66][17] = (mid_1[543:536] > btm_0[535:528]) ? 1 : 0;
assign detect_max[66][18] = (mid_1[543:536] > btm_0[543:536]) ? 1 : 0;
assign detect_max[66][19] = (mid_1[543:536] > btm_0[551:544]) ? 1 : 0;
assign detect_max[66][20] = (mid_1[543:536] > btm_1[535:528]) ? 1 : 0;
assign detect_max[66][21] = (mid_1[543:536] > btm_1[543:536]) ? 1 : 0;
assign detect_max[66][22] = (mid_1[543:536] > btm_1[551:544]) ? 1 : 0;
assign detect_max[66][23] = (mid_1[543:536] > btm_2[535:528]) ? 1 : 0;
assign detect_max[66][24] = (mid_1[543:536] > btm_2[543:536]) ? 1 : 0;
assign detect_max[66][25] = (mid_1[543:536] > btm_2[551:544]) ? 1 : 0;

assign detect_max[67][0] = (mid_1[551:544] > top_0[543:536]) ? 1 : 0;
assign detect_max[67][1] = (mid_1[551:544] > top_0[551:544]) ? 1 : 0;
assign detect_max[67][2] = (mid_1[551:544] > top_0[559:552]) ? 1 : 0;
assign detect_max[67][3] = (mid_1[551:544] > top_1[543:536]) ? 1 : 0;
assign detect_max[67][4] = (mid_1[551:544] > top_1[551:544]) ? 1 : 0;
assign detect_max[67][5] = (mid_1[551:544] > top_1[559:552]) ? 1 : 0;
assign detect_max[67][6] = (mid_1[551:544] > top_2[543:536]) ? 1 : 0;
assign detect_max[67][7] = (mid_1[551:544] > top_2[551:544]) ? 1 : 0;
assign detect_max[67][8] = (mid_1[551:544] > top_2[559:552]) ? 1 : 0;
assign detect_max[67][9] = (mid_1[551:544] > mid_0[543:536]) ? 1 : 0;
assign detect_max[67][10] = (mid_1[551:544] > mid_0[551:544]) ? 1 : 0;
assign detect_max[67][11] = (mid_1[551:544] > mid_0[559:552]) ? 1 : 0;
assign detect_max[67][12] = (mid_1[551:544] > mid_1[543:536]) ? 1 : 0;
assign detect_max[67][13] = (mid_1[551:544] > mid_1[559:552]) ? 1 : 0;
assign detect_max[67][14] = (mid_1[551:544] > mid_2[543:536]) ? 1 : 0;
assign detect_max[67][15] = (mid_1[551:544] > mid_2[551:544]) ? 1 : 0;
assign detect_max[67][16] = (mid_1[551:544] > mid_2[559:552]) ? 1 : 0;
assign detect_max[67][17] = (mid_1[551:544] > btm_0[543:536]) ? 1 : 0;
assign detect_max[67][18] = (mid_1[551:544] > btm_0[551:544]) ? 1 : 0;
assign detect_max[67][19] = (mid_1[551:544] > btm_0[559:552]) ? 1 : 0;
assign detect_max[67][20] = (mid_1[551:544] > btm_1[543:536]) ? 1 : 0;
assign detect_max[67][21] = (mid_1[551:544] > btm_1[551:544]) ? 1 : 0;
assign detect_max[67][22] = (mid_1[551:544] > btm_1[559:552]) ? 1 : 0;
assign detect_max[67][23] = (mid_1[551:544] > btm_2[543:536]) ? 1 : 0;
assign detect_max[67][24] = (mid_1[551:544] > btm_2[551:544]) ? 1 : 0;
assign detect_max[67][25] = (mid_1[551:544] > btm_2[559:552]) ? 1 : 0;

assign detect_max[68][0] = (mid_1[559:552] > top_0[551:544]) ? 1 : 0;
assign detect_max[68][1] = (mid_1[559:552] > top_0[559:552]) ? 1 : 0;
assign detect_max[68][2] = (mid_1[559:552] > top_0[567:560]) ? 1 : 0;
assign detect_max[68][3] = (mid_1[559:552] > top_1[551:544]) ? 1 : 0;
assign detect_max[68][4] = (mid_1[559:552] > top_1[559:552]) ? 1 : 0;
assign detect_max[68][5] = (mid_1[559:552] > top_1[567:560]) ? 1 : 0;
assign detect_max[68][6] = (mid_1[559:552] > top_2[551:544]) ? 1 : 0;
assign detect_max[68][7] = (mid_1[559:552] > top_2[559:552]) ? 1 : 0;
assign detect_max[68][8] = (mid_1[559:552] > top_2[567:560]) ? 1 : 0;
assign detect_max[68][9] = (mid_1[559:552] > mid_0[551:544]) ? 1 : 0;
assign detect_max[68][10] = (mid_1[559:552] > mid_0[559:552]) ? 1 : 0;
assign detect_max[68][11] = (mid_1[559:552] > mid_0[567:560]) ? 1 : 0;
assign detect_max[68][12] = (mid_1[559:552] > mid_1[551:544]) ? 1 : 0;
assign detect_max[68][13] = (mid_1[559:552] > mid_1[567:560]) ? 1 : 0;
assign detect_max[68][14] = (mid_1[559:552] > mid_2[551:544]) ? 1 : 0;
assign detect_max[68][15] = (mid_1[559:552] > mid_2[559:552]) ? 1 : 0;
assign detect_max[68][16] = (mid_1[559:552] > mid_2[567:560]) ? 1 : 0;
assign detect_max[68][17] = (mid_1[559:552] > btm_0[551:544]) ? 1 : 0;
assign detect_max[68][18] = (mid_1[559:552] > btm_0[559:552]) ? 1 : 0;
assign detect_max[68][19] = (mid_1[559:552] > btm_0[567:560]) ? 1 : 0;
assign detect_max[68][20] = (mid_1[559:552] > btm_1[551:544]) ? 1 : 0;
assign detect_max[68][21] = (mid_1[559:552] > btm_1[559:552]) ? 1 : 0;
assign detect_max[68][22] = (mid_1[559:552] > btm_1[567:560]) ? 1 : 0;
assign detect_max[68][23] = (mid_1[559:552] > btm_2[551:544]) ? 1 : 0;
assign detect_max[68][24] = (mid_1[559:552] > btm_2[559:552]) ? 1 : 0;
assign detect_max[68][25] = (mid_1[559:552] > btm_2[567:560]) ? 1 : 0;

assign detect_max[69][0] = (mid_1[567:560] > top_0[559:552]) ? 1 : 0;
assign detect_max[69][1] = (mid_1[567:560] > top_0[567:560]) ? 1 : 0;
assign detect_max[69][2] = (mid_1[567:560] > top_0[575:568]) ? 1 : 0;
assign detect_max[69][3] = (mid_1[567:560] > top_1[559:552]) ? 1 : 0;
assign detect_max[69][4] = (mid_1[567:560] > top_1[567:560]) ? 1 : 0;
assign detect_max[69][5] = (mid_1[567:560] > top_1[575:568]) ? 1 : 0;
assign detect_max[69][6] = (mid_1[567:560] > top_2[559:552]) ? 1 : 0;
assign detect_max[69][7] = (mid_1[567:560] > top_2[567:560]) ? 1 : 0;
assign detect_max[69][8] = (mid_1[567:560] > top_2[575:568]) ? 1 : 0;
assign detect_max[69][9] = (mid_1[567:560] > mid_0[559:552]) ? 1 : 0;
assign detect_max[69][10] = (mid_1[567:560] > mid_0[567:560]) ? 1 : 0;
assign detect_max[69][11] = (mid_1[567:560] > mid_0[575:568]) ? 1 : 0;
assign detect_max[69][12] = (mid_1[567:560] > mid_1[559:552]) ? 1 : 0;
assign detect_max[69][13] = (mid_1[567:560] > mid_1[575:568]) ? 1 : 0;
assign detect_max[69][14] = (mid_1[567:560] > mid_2[559:552]) ? 1 : 0;
assign detect_max[69][15] = (mid_1[567:560] > mid_2[567:560]) ? 1 : 0;
assign detect_max[69][16] = (mid_1[567:560] > mid_2[575:568]) ? 1 : 0;
assign detect_max[69][17] = (mid_1[567:560] > btm_0[559:552]) ? 1 : 0;
assign detect_max[69][18] = (mid_1[567:560] > btm_0[567:560]) ? 1 : 0;
assign detect_max[69][19] = (mid_1[567:560] > btm_0[575:568]) ? 1 : 0;
assign detect_max[69][20] = (mid_1[567:560] > btm_1[559:552]) ? 1 : 0;
assign detect_max[69][21] = (mid_1[567:560] > btm_1[567:560]) ? 1 : 0;
assign detect_max[69][22] = (mid_1[567:560] > btm_1[575:568]) ? 1 : 0;
assign detect_max[69][23] = (mid_1[567:560] > btm_2[559:552]) ? 1 : 0;
assign detect_max[69][24] = (mid_1[567:560] > btm_2[567:560]) ? 1 : 0;
assign detect_max[69][25] = (mid_1[567:560] > btm_2[575:568]) ? 1 : 0;

assign detect_max[70][0] = (mid_1[575:568] > top_0[567:560]) ? 1 : 0;
assign detect_max[70][1] = (mid_1[575:568] > top_0[575:568]) ? 1 : 0;
assign detect_max[70][2] = (mid_1[575:568] > top_0[583:576]) ? 1 : 0;
assign detect_max[70][3] = (mid_1[575:568] > top_1[567:560]) ? 1 : 0;
assign detect_max[70][4] = (mid_1[575:568] > top_1[575:568]) ? 1 : 0;
assign detect_max[70][5] = (mid_1[575:568] > top_1[583:576]) ? 1 : 0;
assign detect_max[70][6] = (mid_1[575:568] > top_2[567:560]) ? 1 : 0;
assign detect_max[70][7] = (mid_1[575:568] > top_2[575:568]) ? 1 : 0;
assign detect_max[70][8] = (mid_1[575:568] > top_2[583:576]) ? 1 : 0;
assign detect_max[70][9] = (mid_1[575:568] > mid_0[567:560]) ? 1 : 0;
assign detect_max[70][10] = (mid_1[575:568] > mid_0[575:568]) ? 1 : 0;
assign detect_max[70][11] = (mid_1[575:568] > mid_0[583:576]) ? 1 : 0;
assign detect_max[70][12] = (mid_1[575:568] > mid_1[567:560]) ? 1 : 0;
assign detect_max[70][13] = (mid_1[575:568] > mid_1[583:576]) ? 1 : 0;
assign detect_max[70][14] = (mid_1[575:568] > mid_2[567:560]) ? 1 : 0;
assign detect_max[70][15] = (mid_1[575:568] > mid_2[575:568]) ? 1 : 0;
assign detect_max[70][16] = (mid_1[575:568] > mid_2[583:576]) ? 1 : 0;
assign detect_max[70][17] = (mid_1[575:568] > btm_0[567:560]) ? 1 : 0;
assign detect_max[70][18] = (mid_1[575:568] > btm_0[575:568]) ? 1 : 0;
assign detect_max[70][19] = (mid_1[575:568] > btm_0[583:576]) ? 1 : 0;
assign detect_max[70][20] = (mid_1[575:568] > btm_1[567:560]) ? 1 : 0;
assign detect_max[70][21] = (mid_1[575:568] > btm_1[575:568]) ? 1 : 0;
assign detect_max[70][22] = (mid_1[575:568] > btm_1[583:576]) ? 1 : 0;
assign detect_max[70][23] = (mid_1[575:568] > btm_2[567:560]) ? 1 : 0;
assign detect_max[70][24] = (mid_1[575:568] > btm_2[575:568]) ? 1 : 0;
assign detect_max[70][25] = (mid_1[575:568] > btm_2[583:576]) ? 1 : 0;

assign detect_max[71][0] = (mid_1[583:576] > top_0[575:568]) ? 1 : 0;
assign detect_max[71][1] = (mid_1[583:576] > top_0[583:576]) ? 1 : 0;
assign detect_max[71][2] = (mid_1[583:576] > top_0[591:584]) ? 1 : 0;
assign detect_max[71][3] = (mid_1[583:576] > top_1[575:568]) ? 1 : 0;
assign detect_max[71][4] = (mid_1[583:576] > top_1[583:576]) ? 1 : 0;
assign detect_max[71][5] = (mid_1[583:576] > top_1[591:584]) ? 1 : 0;
assign detect_max[71][6] = (mid_1[583:576] > top_2[575:568]) ? 1 : 0;
assign detect_max[71][7] = (mid_1[583:576] > top_2[583:576]) ? 1 : 0;
assign detect_max[71][8] = (mid_1[583:576] > top_2[591:584]) ? 1 : 0;
assign detect_max[71][9] = (mid_1[583:576] > mid_0[575:568]) ? 1 : 0;
assign detect_max[71][10] = (mid_1[583:576] > mid_0[583:576]) ? 1 : 0;
assign detect_max[71][11] = (mid_1[583:576] > mid_0[591:584]) ? 1 : 0;
assign detect_max[71][12] = (mid_1[583:576] > mid_1[575:568]) ? 1 : 0;
assign detect_max[71][13] = (mid_1[583:576] > mid_1[591:584]) ? 1 : 0;
assign detect_max[71][14] = (mid_1[583:576] > mid_2[575:568]) ? 1 : 0;
assign detect_max[71][15] = (mid_1[583:576] > mid_2[583:576]) ? 1 : 0;
assign detect_max[71][16] = (mid_1[583:576] > mid_2[591:584]) ? 1 : 0;
assign detect_max[71][17] = (mid_1[583:576] > btm_0[575:568]) ? 1 : 0;
assign detect_max[71][18] = (mid_1[583:576] > btm_0[583:576]) ? 1 : 0;
assign detect_max[71][19] = (mid_1[583:576] > btm_0[591:584]) ? 1 : 0;
assign detect_max[71][20] = (mid_1[583:576] > btm_1[575:568]) ? 1 : 0;
assign detect_max[71][21] = (mid_1[583:576] > btm_1[583:576]) ? 1 : 0;
assign detect_max[71][22] = (mid_1[583:576] > btm_1[591:584]) ? 1 : 0;
assign detect_max[71][23] = (mid_1[583:576] > btm_2[575:568]) ? 1 : 0;
assign detect_max[71][24] = (mid_1[583:576] > btm_2[583:576]) ? 1 : 0;
assign detect_max[71][25] = (mid_1[583:576] > btm_2[591:584]) ? 1 : 0;

assign detect_max[72][0] = (mid_1[591:584] > top_0[583:576]) ? 1 : 0;
assign detect_max[72][1] = (mid_1[591:584] > top_0[591:584]) ? 1 : 0;
assign detect_max[72][2] = (mid_1[591:584] > top_0[599:592]) ? 1 : 0;
assign detect_max[72][3] = (mid_1[591:584] > top_1[583:576]) ? 1 : 0;
assign detect_max[72][4] = (mid_1[591:584] > top_1[591:584]) ? 1 : 0;
assign detect_max[72][5] = (mid_1[591:584] > top_1[599:592]) ? 1 : 0;
assign detect_max[72][6] = (mid_1[591:584] > top_2[583:576]) ? 1 : 0;
assign detect_max[72][7] = (mid_1[591:584] > top_2[591:584]) ? 1 : 0;
assign detect_max[72][8] = (mid_1[591:584] > top_2[599:592]) ? 1 : 0;
assign detect_max[72][9] = (mid_1[591:584] > mid_0[583:576]) ? 1 : 0;
assign detect_max[72][10] = (mid_1[591:584] > mid_0[591:584]) ? 1 : 0;
assign detect_max[72][11] = (mid_1[591:584] > mid_0[599:592]) ? 1 : 0;
assign detect_max[72][12] = (mid_1[591:584] > mid_1[583:576]) ? 1 : 0;
assign detect_max[72][13] = (mid_1[591:584] > mid_1[599:592]) ? 1 : 0;
assign detect_max[72][14] = (mid_1[591:584] > mid_2[583:576]) ? 1 : 0;
assign detect_max[72][15] = (mid_1[591:584] > mid_2[591:584]) ? 1 : 0;
assign detect_max[72][16] = (mid_1[591:584] > mid_2[599:592]) ? 1 : 0;
assign detect_max[72][17] = (mid_1[591:584] > btm_0[583:576]) ? 1 : 0;
assign detect_max[72][18] = (mid_1[591:584] > btm_0[591:584]) ? 1 : 0;
assign detect_max[72][19] = (mid_1[591:584] > btm_0[599:592]) ? 1 : 0;
assign detect_max[72][20] = (mid_1[591:584] > btm_1[583:576]) ? 1 : 0;
assign detect_max[72][21] = (mid_1[591:584] > btm_1[591:584]) ? 1 : 0;
assign detect_max[72][22] = (mid_1[591:584] > btm_1[599:592]) ? 1 : 0;
assign detect_max[72][23] = (mid_1[591:584] > btm_2[583:576]) ? 1 : 0;
assign detect_max[72][24] = (mid_1[591:584] > btm_2[591:584]) ? 1 : 0;
assign detect_max[72][25] = (mid_1[591:584] > btm_2[599:592]) ? 1 : 0;

assign detect_max[73][0] = (mid_1[599:592] > top_0[591:584]) ? 1 : 0;
assign detect_max[73][1] = (mid_1[599:592] > top_0[599:592]) ? 1 : 0;
assign detect_max[73][2] = (mid_1[599:592] > top_0[607:600]) ? 1 : 0;
assign detect_max[73][3] = (mid_1[599:592] > top_1[591:584]) ? 1 : 0;
assign detect_max[73][4] = (mid_1[599:592] > top_1[599:592]) ? 1 : 0;
assign detect_max[73][5] = (mid_1[599:592] > top_1[607:600]) ? 1 : 0;
assign detect_max[73][6] = (mid_1[599:592] > top_2[591:584]) ? 1 : 0;
assign detect_max[73][7] = (mid_1[599:592] > top_2[599:592]) ? 1 : 0;
assign detect_max[73][8] = (mid_1[599:592] > top_2[607:600]) ? 1 : 0;
assign detect_max[73][9] = (mid_1[599:592] > mid_0[591:584]) ? 1 : 0;
assign detect_max[73][10] = (mid_1[599:592] > mid_0[599:592]) ? 1 : 0;
assign detect_max[73][11] = (mid_1[599:592] > mid_0[607:600]) ? 1 : 0;
assign detect_max[73][12] = (mid_1[599:592] > mid_1[591:584]) ? 1 : 0;
assign detect_max[73][13] = (mid_1[599:592] > mid_1[607:600]) ? 1 : 0;
assign detect_max[73][14] = (mid_1[599:592] > mid_2[591:584]) ? 1 : 0;
assign detect_max[73][15] = (mid_1[599:592] > mid_2[599:592]) ? 1 : 0;
assign detect_max[73][16] = (mid_1[599:592] > mid_2[607:600]) ? 1 : 0;
assign detect_max[73][17] = (mid_1[599:592] > btm_0[591:584]) ? 1 : 0;
assign detect_max[73][18] = (mid_1[599:592] > btm_0[599:592]) ? 1 : 0;
assign detect_max[73][19] = (mid_1[599:592] > btm_0[607:600]) ? 1 : 0;
assign detect_max[73][20] = (mid_1[599:592] > btm_1[591:584]) ? 1 : 0;
assign detect_max[73][21] = (mid_1[599:592] > btm_1[599:592]) ? 1 : 0;
assign detect_max[73][22] = (mid_1[599:592] > btm_1[607:600]) ? 1 : 0;
assign detect_max[73][23] = (mid_1[599:592] > btm_2[591:584]) ? 1 : 0;
assign detect_max[73][24] = (mid_1[599:592] > btm_2[599:592]) ? 1 : 0;
assign detect_max[73][25] = (mid_1[599:592] > btm_2[607:600]) ? 1 : 0;

assign detect_max[74][0] = (mid_1[607:600] > top_0[599:592]) ? 1 : 0;
assign detect_max[74][1] = (mid_1[607:600] > top_0[607:600]) ? 1 : 0;
assign detect_max[74][2] = (mid_1[607:600] > top_0[615:608]) ? 1 : 0;
assign detect_max[74][3] = (mid_1[607:600] > top_1[599:592]) ? 1 : 0;
assign detect_max[74][4] = (mid_1[607:600] > top_1[607:600]) ? 1 : 0;
assign detect_max[74][5] = (mid_1[607:600] > top_1[615:608]) ? 1 : 0;
assign detect_max[74][6] = (mid_1[607:600] > top_2[599:592]) ? 1 : 0;
assign detect_max[74][7] = (mid_1[607:600] > top_2[607:600]) ? 1 : 0;
assign detect_max[74][8] = (mid_1[607:600] > top_2[615:608]) ? 1 : 0;
assign detect_max[74][9] = (mid_1[607:600] > mid_0[599:592]) ? 1 : 0;
assign detect_max[74][10] = (mid_1[607:600] > mid_0[607:600]) ? 1 : 0;
assign detect_max[74][11] = (mid_1[607:600] > mid_0[615:608]) ? 1 : 0;
assign detect_max[74][12] = (mid_1[607:600] > mid_1[599:592]) ? 1 : 0;
assign detect_max[74][13] = (mid_1[607:600] > mid_1[615:608]) ? 1 : 0;
assign detect_max[74][14] = (mid_1[607:600] > mid_2[599:592]) ? 1 : 0;
assign detect_max[74][15] = (mid_1[607:600] > mid_2[607:600]) ? 1 : 0;
assign detect_max[74][16] = (mid_1[607:600] > mid_2[615:608]) ? 1 : 0;
assign detect_max[74][17] = (mid_1[607:600] > btm_0[599:592]) ? 1 : 0;
assign detect_max[74][18] = (mid_1[607:600] > btm_0[607:600]) ? 1 : 0;
assign detect_max[74][19] = (mid_1[607:600] > btm_0[615:608]) ? 1 : 0;
assign detect_max[74][20] = (mid_1[607:600] > btm_1[599:592]) ? 1 : 0;
assign detect_max[74][21] = (mid_1[607:600] > btm_1[607:600]) ? 1 : 0;
assign detect_max[74][22] = (mid_1[607:600] > btm_1[615:608]) ? 1 : 0;
assign detect_max[74][23] = (mid_1[607:600] > btm_2[599:592]) ? 1 : 0;
assign detect_max[74][24] = (mid_1[607:600] > btm_2[607:600]) ? 1 : 0;
assign detect_max[74][25] = (mid_1[607:600] > btm_2[615:608]) ? 1 : 0;

assign detect_max[75][0] = (mid_1[615:608] > top_0[607:600]) ? 1 : 0;
assign detect_max[75][1] = (mid_1[615:608] > top_0[615:608]) ? 1 : 0;
assign detect_max[75][2] = (mid_1[615:608] > top_0[623:616]) ? 1 : 0;
assign detect_max[75][3] = (mid_1[615:608] > top_1[607:600]) ? 1 : 0;
assign detect_max[75][4] = (mid_1[615:608] > top_1[615:608]) ? 1 : 0;
assign detect_max[75][5] = (mid_1[615:608] > top_1[623:616]) ? 1 : 0;
assign detect_max[75][6] = (mid_1[615:608] > top_2[607:600]) ? 1 : 0;
assign detect_max[75][7] = (mid_1[615:608] > top_2[615:608]) ? 1 : 0;
assign detect_max[75][8] = (mid_1[615:608] > top_2[623:616]) ? 1 : 0;
assign detect_max[75][9] = (mid_1[615:608] > mid_0[607:600]) ? 1 : 0;
assign detect_max[75][10] = (mid_1[615:608] > mid_0[615:608]) ? 1 : 0;
assign detect_max[75][11] = (mid_1[615:608] > mid_0[623:616]) ? 1 : 0;
assign detect_max[75][12] = (mid_1[615:608] > mid_1[607:600]) ? 1 : 0;
assign detect_max[75][13] = (mid_1[615:608] > mid_1[623:616]) ? 1 : 0;
assign detect_max[75][14] = (mid_1[615:608] > mid_2[607:600]) ? 1 : 0;
assign detect_max[75][15] = (mid_1[615:608] > mid_2[615:608]) ? 1 : 0;
assign detect_max[75][16] = (mid_1[615:608] > mid_2[623:616]) ? 1 : 0;
assign detect_max[75][17] = (mid_1[615:608] > btm_0[607:600]) ? 1 : 0;
assign detect_max[75][18] = (mid_1[615:608] > btm_0[615:608]) ? 1 : 0;
assign detect_max[75][19] = (mid_1[615:608] > btm_0[623:616]) ? 1 : 0;
assign detect_max[75][20] = (mid_1[615:608] > btm_1[607:600]) ? 1 : 0;
assign detect_max[75][21] = (mid_1[615:608] > btm_1[615:608]) ? 1 : 0;
assign detect_max[75][22] = (mid_1[615:608] > btm_1[623:616]) ? 1 : 0;
assign detect_max[75][23] = (mid_1[615:608] > btm_2[607:600]) ? 1 : 0;
assign detect_max[75][24] = (mid_1[615:608] > btm_2[615:608]) ? 1 : 0;
assign detect_max[75][25] = (mid_1[615:608] > btm_2[623:616]) ? 1 : 0;

assign detect_max[76][0] = (mid_1[623:616] > top_0[615:608]) ? 1 : 0;
assign detect_max[76][1] = (mid_1[623:616] > top_0[623:616]) ? 1 : 0;
assign detect_max[76][2] = (mid_1[623:616] > top_0[631:624]) ? 1 : 0;
assign detect_max[76][3] = (mid_1[623:616] > top_1[615:608]) ? 1 : 0;
assign detect_max[76][4] = (mid_1[623:616] > top_1[623:616]) ? 1 : 0;
assign detect_max[76][5] = (mid_1[623:616] > top_1[631:624]) ? 1 : 0;
assign detect_max[76][6] = (mid_1[623:616] > top_2[615:608]) ? 1 : 0;
assign detect_max[76][7] = (mid_1[623:616] > top_2[623:616]) ? 1 : 0;
assign detect_max[76][8] = (mid_1[623:616] > top_2[631:624]) ? 1 : 0;
assign detect_max[76][9] = (mid_1[623:616] > mid_0[615:608]) ? 1 : 0;
assign detect_max[76][10] = (mid_1[623:616] > mid_0[623:616]) ? 1 : 0;
assign detect_max[76][11] = (mid_1[623:616] > mid_0[631:624]) ? 1 : 0;
assign detect_max[76][12] = (mid_1[623:616] > mid_1[615:608]) ? 1 : 0;
assign detect_max[76][13] = (mid_1[623:616] > mid_1[631:624]) ? 1 : 0;
assign detect_max[76][14] = (mid_1[623:616] > mid_2[615:608]) ? 1 : 0;
assign detect_max[76][15] = (mid_1[623:616] > mid_2[623:616]) ? 1 : 0;
assign detect_max[76][16] = (mid_1[623:616] > mid_2[631:624]) ? 1 : 0;
assign detect_max[76][17] = (mid_1[623:616] > btm_0[615:608]) ? 1 : 0;
assign detect_max[76][18] = (mid_1[623:616] > btm_0[623:616]) ? 1 : 0;
assign detect_max[76][19] = (mid_1[623:616] > btm_0[631:624]) ? 1 : 0;
assign detect_max[76][20] = (mid_1[623:616] > btm_1[615:608]) ? 1 : 0;
assign detect_max[76][21] = (mid_1[623:616] > btm_1[623:616]) ? 1 : 0;
assign detect_max[76][22] = (mid_1[623:616] > btm_1[631:624]) ? 1 : 0;
assign detect_max[76][23] = (mid_1[623:616] > btm_2[615:608]) ? 1 : 0;
assign detect_max[76][24] = (mid_1[623:616] > btm_2[623:616]) ? 1 : 0;
assign detect_max[76][25] = (mid_1[623:616] > btm_2[631:624]) ? 1 : 0;

assign detect_max[77][0] = (mid_1[631:624] > top_0[623:616]) ? 1 : 0;
assign detect_max[77][1] = (mid_1[631:624] > top_0[631:624]) ? 1 : 0;
assign detect_max[77][2] = (mid_1[631:624] > top_0[639:632]) ? 1 : 0;
assign detect_max[77][3] = (mid_1[631:624] > top_1[623:616]) ? 1 : 0;
assign detect_max[77][4] = (mid_1[631:624] > top_1[631:624]) ? 1 : 0;
assign detect_max[77][5] = (mid_1[631:624] > top_1[639:632]) ? 1 : 0;
assign detect_max[77][6] = (mid_1[631:624] > top_2[623:616]) ? 1 : 0;
assign detect_max[77][7] = (mid_1[631:624] > top_2[631:624]) ? 1 : 0;
assign detect_max[77][8] = (mid_1[631:624] > top_2[639:632]) ? 1 : 0;
assign detect_max[77][9] = (mid_1[631:624] > mid_0[623:616]) ? 1 : 0;
assign detect_max[77][10] = (mid_1[631:624] > mid_0[631:624]) ? 1 : 0;
assign detect_max[77][11] = (mid_1[631:624] > mid_0[639:632]) ? 1 : 0;
assign detect_max[77][12] = (mid_1[631:624] > mid_1[623:616]) ? 1 : 0;
assign detect_max[77][13] = (mid_1[631:624] > mid_1[639:632]) ? 1 : 0;
assign detect_max[77][14] = (mid_1[631:624] > mid_2[623:616]) ? 1 : 0;
assign detect_max[77][15] = (mid_1[631:624] > mid_2[631:624]) ? 1 : 0;
assign detect_max[77][16] = (mid_1[631:624] > mid_2[639:632]) ? 1 : 0;
assign detect_max[77][17] = (mid_1[631:624] > btm_0[623:616]) ? 1 : 0;
assign detect_max[77][18] = (mid_1[631:624] > btm_0[631:624]) ? 1 : 0;
assign detect_max[77][19] = (mid_1[631:624] > btm_0[639:632]) ? 1 : 0;
assign detect_max[77][20] = (mid_1[631:624] > btm_1[623:616]) ? 1 : 0;
assign detect_max[77][21] = (mid_1[631:624] > btm_1[631:624]) ? 1 : 0;
assign detect_max[77][22] = (mid_1[631:624] > btm_1[639:632]) ? 1 : 0;
assign detect_max[77][23] = (mid_1[631:624] > btm_2[623:616]) ? 1 : 0;
assign detect_max[77][24] = (mid_1[631:624] > btm_2[631:624]) ? 1 : 0;
assign detect_max[77][25] = (mid_1[631:624] > btm_2[639:632]) ? 1 : 0;

assign detect_max[78][0] = (mid_1[639:632] > top_0[631:624]) ? 1 : 0;
assign detect_max[78][1] = (mid_1[639:632] > top_0[639:632]) ? 1 : 0;
assign detect_max[78][2] = (mid_1[639:632] > top_0[647:640]) ? 1 : 0;
assign detect_max[78][3] = (mid_1[639:632] > top_1[631:624]) ? 1 : 0;
assign detect_max[78][4] = (mid_1[639:632] > top_1[639:632]) ? 1 : 0;
assign detect_max[78][5] = (mid_1[639:632] > top_1[647:640]) ? 1 : 0;
assign detect_max[78][6] = (mid_1[639:632] > top_2[631:624]) ? 1 : 0;
assign detect_max[78][7] = (mid_1[639:632] > top_2[639:632]) ? 1 : 0;
assign detect_max[78][8] = (mid_1[639:632] > top_2[647:640]) ? 1 : 0;
assign detect_max[78][9] = (mid_1[639:632] > mid_0[631:624]) ? 1 : 0;
assign detect_max[78][10] = (mid_1[639:632] > mid_0[639:632]) ? 1 : 0;
assign detect_max[78][11] = (mid_1[639:632] > mid_0[647:640]) ? 1 : 0;
assign detect_max[78][12] = (mid_1[639:632] > mid_1[631:624]) ? 1 : 0;
assign detect_max[78][13] = (mid_1[639:632] > mid_1[647:640]) ? 1 : 0;
assign detect_max[78][14] = (mid_1[639:632] > mid_2[631:624]) ? 1 : 0;
assign detect_max[78][15] = (mid_1[639:632] > mid_2[639:632]) ? 1 : 0;
assign detect_max[78][16] = (mid_1[639:632] > mid_2[647:640]) ? 1 : 0;
assign detect_max[78][17] = (mid_1[639:632] > btm_0[631:624]) ? 1 : 0;
assign detect_max[78][18] = (mid_1[639:632] > btm_0[639:632]) ? 1 : 0;
assign detect_max[78][19] = (mid_1[639:632] > btm_0[647:640]) ? 1 : 0;
assign detect_max[78][20] = (mid_1[639:632] > btm_1[631:624]) ? 1 : 0;
assign detect_max[78][21] = (mid_1[639:632] > btm_1[639:632]) ? 1 : 0;
assign detect_max[78][22] = (mid_1[639:632] > btm_1[647:640]) ? 1 : 0;
assign detect_max[78][23] = (mid_1[639:632] > btm_2[631:624]) ? 1 : 0;
assign detect_max[78][24] = (mid_1[639:632] > btm_2[639:632]) ? 1 : 0;
assign detect_max[78][25] = (mid_1[639:632] > btm_2[647:640]) ? 1 : 0;

assign detect_max[79][0] = (mid_1[647:640] > top_0[639:632]) ? 1 : 0;
assign detect_max[79][1] = (mid_1[647:640] > top_0[647:640]) ? 1 : 0;
assign detect_max[79][2] = (mid_1[647:640] > top_0[655:648]) ? 1 : 0;
assign detect_max[79][3] = (mid_1[647:640] > top_1[639:632]) ? 1 : 0;
assign detect_max[79][4] = (mid_1[647:640] > top_1[647:640]) ? 1 : 0;
assign detect_max[79][5] = (mid_1[647:640] > top_1[655:648]) ? 1 : 0;
assign detect_max[79][6] = (mid_1[647:640] > top_2[639:632]) ? 1 : 0;
assign detect_max[79][7] = (mid_1[647:640] > top_2[647:640]) ? 1 : 0;
assign detect_max[79][8] = (mid_1[647:640] > top_2[655:648]) ? 1 : 0;
assign detect_max[79][9] = (mid_1[647:640] > mid_0[639:632]) ? 1 : 0;
assign detect_max[79][10] = (mid_1[647:640] > mid_0[647:640]) ? 1 : 0;
assign detect_max[79][11] = (mid_1[647:640] > mid_0[655:648]) ? 1 : 0;
assign detect_max[79][12] = (mid_1[647:640] > mid_1[639:632]) ? 1 : 0;
assign detect_max[79][13] = (mid_1[647:640] > mid_1[655:648]) ? 1 : 0;
assign detect_max[79][14] = (mid_1[647:640] > mid_2[639:632]) ? 1 : 0;
assign detect_max[79][15] = (mid_1[647:640] > mid_2[647:640]) ? 1 : 0;
assign detect_max[79][16] = (mid_1[647:640] > mid_2[655:648]) ? 1 : 0;
assign detect_max[79][17] = (mid_1[647:640] > btm_0[639:632]) ? 1 : 0;
assign detect_max[79][18] = (mid_1[647:640] > btm_0[647:640]) ? 1 : 0;
assign detect_max[79][19] = (mid_1[647:640] > btm_0[655:648]) ? 1 : 0;
assign detect_max[79][20] = (mid_1[647:640] > btm_1[639:632]) ? 1 : 0;
assign detect_max[79][21] = (mid_1[647:640] > btm_1[647:640]) ? 1 : 0;
assign detect_max[79][22] = (mid_1[647:640] > btm_1[655:648]) ? 1 : 0;
assign detect_max[79][23] = (mid_1[647:640] > btm_2[639:632]) ? 1 : 0;
assign detect_max[79][24] = (mid_1[647:640] > btm_2[647:640]) ? 1 : 0;
assign detect_max[79][25] = (mid_1[647:640] > btm_2[655:648]) ? 1 : 0;

assign detect_max[80][0] = (mid_1[655:648] > top_0[647:640]) ? 1 : 0;
assign detect_max[80][1] = (mid_1[655:648] > top_0[655:648]) ? 1 : 0;
assign detect_max[80][2] = (mid_1[655:648] > top_0[663:656]) ? 1 : 0;
assign detect_max[80][3] = (mid_1[655:648] > top_1[647:640]) ? 1 : 0;
assign detect_max[80][4] = (mid_1[655:648] > top_1[655:648]) ? 1 : 0;
assign detect_max[80][5] = (mid_1[655:648] > top_1[663:656]) ? 1 : 0;
assign detect_max[80][6] = (mid_1[655:648] > top_2[647:640]) ? 1 : 0;
assign detect_max[80][7] = (mid_1[655:648] > top_2[655:648]) ? 1 : 0;
assign detect_max[80][8] = (mid_1[655:648] > top_2[663:656]) ? 1 : 0;
assign detect_max[80][9] = (mid_1[655:648] > mid_0[647:640]) ? 1 : 0;
assign detect_max[80][10] = (mid_1[655:648] > mid_0[655:648]) ? 1 : 0;
assign detect_max[80][11] = (mid_1[655:648] > mid_0[663:656]) ? 1 : 0;
assign detect_max[80][12] = (mid_1[655:648] > mid_1[647:640]) ? 1 : 0;
assign detect_max[80][13] = (mid_1[655:648] > mid_1[663:656]) ? 1 : 0;
assign detect_max[80][14] = (mid_1[655:648] > mid_2[647:640]) ? 1 : 0;
assign detect_max[80][15] = (mid_1[655:648] > mid_2[655:648]) ? 1 : 0;
assign detect_max[80][16] = (mid_1[655:648] > mid_2[663:656]) ? 1 : 0;
assign detect_max[80][17] = (mid_1[655:648] > btm_0[647:640]) ? 1 : 0;
assign detect_max[80][18] = (mid_1[655:648] > btm_0[655:648]) ? 1 : 0;
assign detect_max[80][19] = (mid_1[655:648] > btm_0[663:656]) ? 1 : 0;
assign detect_max[80][20] = (mid_1[655:648] > btm_1[647:640]) ? 1 : 0;
assign detect_max[80][21] = (mid_1[655:648] > btm_1[655:648]) ? 1 : 0;
assign detect_max[80][22] = (mid_1[655:648] > btm_1[663:656]) ? 1 : 0;
assign detect_max[80][23] = (mid_1[655:648] > btm_2[647:640]) ? 1 : 0;
assign detect_max[80][24] = (mid_1[655:648] > btm_2[655:648]) ? 1 : 0;
assign detect_max[80][25] = (mid_1[655:648] > btm_2[663:656]) ? 1 : 0;

assign detect_max[81][0] = (mid_1[663:656] > top_0[655:648]) ? 1 : 0;
assign detect_max[81][1] = (mid_1[663:656] > top_0[663:656]) ? 1 : 0;
assign detect_max[81][2] = (mid_1[663:656] > top_0[671:664]) ? 1 : 0;
assign detect_max[81][3] = (mid_1[663:656] > top_1[655:648]) ? 1 : 0;
assign detect_max[81][4] = (mid_1[663:656] > top_1[663:656]) ? 1 : 0;
assign detect_max[81][5] = (mid_1[663:656] > top_1[671:664]) ? 1 : 0;
assign detect_max[81][6] = (mid_1[663:656] > top_2[655:648]) ? 1 : 0;
assign detect_max[81][7] = (mid_1[663:656] > top_2[663:656]) ? 1 : 0;
assign detect_max[81][8] = (mid_1[663:656] > top_2[671:664]) ? 1 : 0;
assign detect_max[81][9] = (mid_1[663:656] > mid_0[655:648]) ? 1 : 0;
assign detect_max[81][10] = (mid_1[663:656] > mid_0[663:656]) ? 1 : 0;
assign detect_max[81][11] = (mid_1[663:656] > mid_0[671:664]) ? 1 : 0;
assign detect_max[81][12] = (mid_1[663:656] > mid_1[655:648]) ? 1 : 0;
assign detect_max[81][13] = (mid_1[663:656] > mid_1[671:664]) ? 1 : 0;
assign detect_max[81][14] = (mid_1[663:656] > mid_2[655:648]) ? 1 : 0;
assign detect_max[81][15] = (mid_1[663:656] > mid_2[663:656]) ? 1 : 0;
assign detect_max[81][16] = (mid_1[663:656] > mid_2[671:664]) ? 1 : 0;
assign detect_max[81][17] = (mid_1[663:656] > btm_0[655:648]) ? 1 : 0;
assign detect_max[81][18] = (mid_1[663:656] > btm_0[663:656]) ? 1 : 0;
assign detect_max[81][19] = (mid_1[663:656] > btm_0[671:664]) ? 1 : 0;
assign detect_max[81][20] = (mid_1[663:656] > btm_1[655:648]) ? 1 : 0;
assign detect_max[81][21] = (mid_1[663:656] > btm_1[663:656]) ? 1 : 0;
assign detect_max[81][22] = (mid_1[663:656] > btm_1[671:664]) ? 1 : 0;
assign detect_max[81][23] = (mid_1[663:656] > btm_2[655:648]) ? 1 : 0;
assign detect_max[81][24] = (mid_1[663:656] > btm_2[663:656]) ? 1 : 0;
assign detect_max[81][25] = (mid_1[663:656] > btm_2[671:664]) ? 1 : 0;

assign detect_max[82][0] = (mid_1[671:664] > top_0[663:656]) ? 1 : 0;
assign detect_max[82][1] = (mid_1[671:664] > top_0[671:664]) ? 1 : 0;
assign detect_max[82][2] = (mid_1[671:664] > top_0[679:672]) ? 1 : 0;
assign detect_max[82][3] = (mid_1[671:664] > top_1[663:656]) ? 1 : 0;
assign detect_max[82][4] = (mid_1[671:664] > top_1[671:664]) ? 1 : 0;
assign detect_max[82][5] = (mid_1[671:664] > top_1[679:672]) ? 1 : 0;
assign detect_max[82][6] = (mid_1[671:664] > top_2[663:656]) ? 1 : 0;
assign detect_max[82][7] = (mid_1[671:664] > top_2[671:664]) ? 1 : 0;
assign detect_max[82][8] = (mid_1[671:664] > top_2[679:672]) ? 1 : 0;
assign detect_max[82][9] = (mid_1[671:664] > mid_0[663:656]) ? 1 : 0;
assign detect_max[82][10] = (mid_1[671:664] > mid_0[671:664]) ? 1 : 0;
assign detect_max[82][11] = (mid_1[671:664] > mid_0[679:672]) ? 1 : 0;
assign detect_max[82][12] = (mid_1[671:664] > mid_1[663:656]) ? 1 : 0;
assign detect_max[82][13] = (mid_1[671:664] > mid_1[679:672]) ? 1 : 0;
assign detect_max[82][14] = (mid_1[671:664] > mid_2[663:656]) ? 1 : 0;
assign detect_max[82][15] = (mid_1[671:664] > mid_2[671:664]) ? 1 : 0;
assign detect_max[82][16] = (mid_1[671:664] > mid_2[679:672]) ? 1 : 0;
assign detect_max[82][17] = (mid_1[671:664] > btm_0[663:656]) ? 1 : 0;
assign detect_max[82][18] = (mid_1[671:664] > btm_0[671:664]) ? 1 : 0;
assign detect_max[82][19] = (mid_1[671:664] > btm_0[679:672]) ? 1 : 0;
assign detect_max[82][20] = (mid_1[671:664] > btm_1[663:656]) ? 1 : 0;
assign detect_max[82][21] = (mid_1[671:664] > btm_1[671:664]) ? 1 : 0;
assign detect_max[82][22] = (mid_1[671:664] > btm_1[679:672]) ? 1 : 0;
assign detect_max[82][23] = (mid_1[671:664] > btm_2[663:656]) ? 1 : 0;
assign detect_max[82][24] = (mid_1[671:664] > btm_2[671:664]) ? 1 : 0;
assign detect_max[82][25] = (mid_1[671:664] > btm_2[679:672]) ? 1 : 0;

assign detect_max[83][0] = (mid_1[679:672] > top_0[671:664]) ? 1 : 0;
assign detect_max[83][1] = (mid_1[679:672] > top_0[679:672]) ? 1 : 0;
assign detect_max[83][2] = (mid_1[679:672] > top_0[687:680]) ? 1 : 0;
assign detect_max[83][3] = (mid_1[679:672] > top_1[671:664]) ? 1 : 0;
assign detect_max[83][4] = (mid_1[679:672] > top_1[679:672]) ? 1 : 0;
assign detect_max[83][5] = (mid_1[679:672] > top_1[687:680]) ? 1 : 0;
assign detect_max[83][6] = (mid_1[679:672] > top_2[671:664]) ? 1 : 0;
assign detect_max[83][7] = (mid_1[679:672] > top_2[679:672]) ? 1 : 0;
assign detect_max[83][8] = (mid_1[679:672] > top_2[687:680]) ? 1 : 0;
assign detect_max[83][9] = (mid_1[679:672] > mid_0[671:664]) ? 1 : 0;
assign detect_max[83][10] = (mid_1[679:672] > mid_0[679:672]) ? 1 : 0;
assign detect_max[83][11] = (mid_1[679:672] > mid_0[687:680]) ? 1 : 0;
assign detect_max[83][12] = (mid_1[679:672] > mid_1[671:664]) ? 1 : 0;
assign detect_max[83][13] = (mid_1[679:672] > mid_1[687:680]) ? 1 : 0;
assign detect_max[83][14] = (mid_1[679:672] > mid_2[671:664]) ? 1 : 0;
assign detect_max[83][15] = (mid_1[679:672] > mid_2[679:672]) ? 1 : 0;
assign detect_max[83][16] = (mid_1[679:672] > mid_2[687:680]) ? 1 : 0;
assign detect_max[83][17] = (mid_1[679:672] > btm_0[671:664]) ? 1 : 0;
assign detect_max[83][18] = (mid_1[679:672] > btm_0[679:672]) ? 1 : 0;
assign detect_max[83][19] = (mid_1[679:672] > btm_0[687:680]) ? 1 : 0;
assign detect_max[83][20] = (mid_1[679:672] > btm_1[671:664]) ? 1 : 0;
assign detect_max[83][21] = (mid_1[679:672] > btm_1[679:672]) ? 1 : 0;
assign detect_max[83][22] = (mid_1[679:672] > btm_1[687:680]) ? 1 : 0;
assign detect_max[83][23] = (mid_1[679:672] > btm_2[671:664]) ? 1 : 0;
assign detect_max[83][24] = (mid_1[679:672] > btm_2[679:672]) ? 1 : 0;
assign detect_max[83][25] = (mid_1[679:672] > btm_2[687:680]) ? 1 : 0;

assign detect_max[84][0] = (mid_1[687:680] > top_0[679:672]) ? 1 : 0;
assign detect_max[84][1] = (mid_1[687:680] > top_0[687:680]) ? 1 : 0;
assign detect_max[84][2] = (mid_1[687:680] > top_0[695:688]) ? 1 : 0;
assign detect_max[84][3] = (mid_1[687:680] > top_1[679:672]) ? 1 : 0;
assign detect_max[84][4] = (mid_1[687:680] > top_1[687:680]) ? 1 : 0;
assign detect_max[84][5] = (mid_1[687:680] > top_1[695:688]) ? 1 : 0;
assign detect_max[84][6] = (mid_1[687:680] > top_2[679:672]) ? 1 : 0;
assign detect_max[84][7] = (mid_1[687:680] > top_2[687:680]) ? 1 : 0;
assign detect_max[84][8] = (mid_1[687:680] > top_2[695:688]) ? 1 : 0;
assign detect_max[84][9] = (mid_1[687:680] > mid_0[679:672]) ? 1 : 0;
assign detect_max[84][10] = (mid_1[687:680] > mid_0[687:680]) ? 1 : 0;
assign detect_max[84][11] = (mid_1[687:680] > mid_0[695:688]) ? 1 : 0;
assign detect_max[84][12] = (mid_1[687:680] > mid_1[679:672]) ? 1 : 0;
assign detect_max[84][13] = (mid_1[687:680] > mid_1[695:688]) ? 1 : 0;
assign detect_max[84][14] = (mid_1[687:680] > mid_2[679:672]) ? 1 : 0;
assign detect_max[84][15] = (mid_1[687:680] > mid_2[687:680]) ? 1 : 0;
assign detect_max[84][16] = (mid_1[687:680] > mid_2[695:688]) ? 1 : 0;
assign detect_max[84][17] = (mid_1[687:680] > btm_0[679:672]) ? 1 : 0;
assign detect_max[84][18] = (mid_1[687:680] > btm_0[687:680]) ? 1 : 0;
assign detect_max[84][19] = (mid_1[687:680] > btm_0[695:688]) ? 1 : 0;
assign detect_max[84][20] = (mid_1[687:680] > btm_1[679:672]) ? 1 : 0;
assign detect_max[84][21] = (mid_1[687:680] > btm_1[687:680]) ? 1 : 0;
assign detect_max[84][22] = (mid_1[687:680] > btm_1[695:688]) ? 1 : 0;
assign detect_max[84][23] = (mid_1[687:680] > btm_2[679:672]) ? 1 : 0;
assign detect_max[84][24] = (mid_1[687:680] > btm_2[687:680]) ? 1 : 0;
assign detect_max[84][25] = (mid_1[687:680] > btm_2[695:688]) ? 1 : 0;

assign detect_max[85][0] = (mid_1[695:688] > top_0[687:680]) ? 1 : 0;
assign detect_max[85][1] = (mid_1[695:688] > top_0[695:688]) ? 1 : 0;
assign detect_max[85][2] = (mid_1[695:688] > top_0[703:696]) ? 1 : 0;
assign detect_max[85][3] = (mid_1[695:688] > top_1[687:680]) ? 1 : 0;
assign detect_max[85][4] = (mid_1[695:688] > top_1[695:688]) ? 1 : 0;
assign detect_max[85][5] = (mid_1[695:688] > top_1[703:696]) ? 1 : 0;
assign detect_max[85][6] = (mid_1[695:688] > top_2[687:680]) ? 1 : 0;
assign detect_max[85][7] = (mid_1[695:688] > top_2[695:688]) ? 1 : 0;
assign detect_max[85][8] = (mid_1[695:688] > top_2[703:696]) ? 1 : 0;
assign detect_max[85][9] = (mid_1[695:688] > mid_0[687:680]) ? 1 : 0;
assign detect_max[85][10] = (mid_1[695:688] > mid_0[695:688]) ? 1 : 0;
assign detect_max[85][11] = (mid_1[695:688] > mid_0[703:696]) ? 1 : 0;
assign detect_max[85][12] = (mid_1[695:688] > mid_1[687:680]) ? 1 : 0;
assign detect_max[85][13] = (mid_1[695:688] > mid_1[703:696]) ? 1 : 0;
assign detect_max[85][14] = (mid_1[695:688] > mid_2[687:680]) ? 1 : 0;
assign detect_max[85][15] = (mid_1[695:688] > mid_2[695:688]) ? 1 : 0;
assign detect_max[85][16] = (mid_1[695:688] > mid_2[703:696]) ? 1 : 0;
assign detect_max[85][17] = (mid_1[695:688] > btm_0[687:680]) ? 1 : 0;
assign detect_max[85][18] = (mid_1[695:688] > btm_0[695:688]) ? 1 : 0;
assign detect_max[85][19] = (mid_1[695:688] > btm_0[703:696]) ? 1 : 0;
assign detect_max[85][20] = (mid_1[695:688] > btm_1[687:680]) ? 1 : 0;
assign detect_max[85][21] = (mid_1[695:688] > btm_1[695:688]) ? 1 : 0;
assign detect_max[85][22] = (mid_1[695:688] > btm_1[703:696]) ? 1 : 0;
assign detect_max[85][23] = (mid_1[695:688] > btm_2[687:680]) ? 1 : 0;
assign detect_max[85][24] = (mid_1[695:688] > btm_2[695:688]) ? 1 : 0;
assign detect_max[85][25] = (mid_1[695:688] > btm_2[703:696]) ? 1 : 0;

assign detect_max[86][0] = (mid_1[703:696] > top_0[695:688]) ? 1 : 0;
assign detect_max[86][1] = (mid_1[703:696] > top_0[703:696]) ? 1 : 0;
assign detect_max[86][2] = (mid_1[703:696] > top_0[711:704]) ? 1 : 0;
assign detect_max[86][3] = (mid_1[703:696] > top_1[695:688]) ? 1 : 0;
assign detect_max[86][4] = (mid_1[703:696] > top_1[703:696]) ? 1 : 0;
assign detect_max[86][5] = (mid_1[703:696] > top_1[711:704]) ? 1 : 0;
assign detect_max[86][6] = (mid_1[703:696] > top_2[695:688]) ? 1 : 0;
assign detect_max[86][7] = (mid_1[703:696] > top_2[703:696]) ? 1 : 0;
assign detect_max[86][8] = (mid_1[703:696] > top_2[711:704]) ? 1 : 0;
assign detect_max[86][9] = (mid_1[703:696] > mid_0[695:688]) ? 1 : 0;
assign detect_max[86][10] = (mid_1[703:696] > mid_0[703:696]) ? 1 : 0;
assign detect_max[86][11] = (mid_1[703:696] > mid_0[711:704]) ? 1 : 0;
assign detect_max[86][12] = (mid_1[703:696] > mid_1[695:688]) ? 1 : 0;
assign detect_max[86][13] = (mid_1[703:696] > mid_1[711:704]) ? 1 : 0;
assign detect_max[86][14] = (mid_1[703:696] > mid_2[695:688]) ? 1 : 0;
assign detect_max[86][15] = (mid_1[703:696] > mid_2[703:696]) ? 1 : 0;
assign detect_max[86][16] = (mid_1[703:696] > mid_2[711:704]) ? 1 : 0;
assign detect_max[86][17] = (mid_1[703:696] > btm_0[695:688]) ? 1 : 0;
assign detect_max[86][18] = (mid_1[703:696] > btm_0[703:696]) ? 1 : 0;
assign detect_max[86][19] = (mid_1[703:696] > btm_0[711:704]) ? 1 : 0;
assign detect_max[86][20] = (mid_1[703:696] > btm_1[695:688]) ? 1 : 0;
assign detect_max[86][21] = (mid_1[703:696] > btm_1[703:696]) ? 1 : 0;
assign detect_max[86][22] = (mid_1[703:696] > btm_1[711:704]) ? 1 : 0;
assign detect_max[86][23] = (mid_1[703:696] > btm_2[695:688]) ? 1 : 0;
assign detect_max[86][24] = (mid_1[703:696] > btm_2[703:696]) ? 1 : 0;
assign detect_max[86][25] = (mid_1[703:696] > btm_2[711:704]) ? 1 : 0;

assign detect_max[87][0] = (mid_1[711:704] > top_0[703:696]) ? 1 : 0;
assign detect_max[87][1] = (mid_1[711:704] > top_0[711:704]) ? 1 : 0;
assign detect_max[87][2] = (mid_1[711:704] > top_0[719:712]) ? 1 : 0;
assign detect_max[87][3] = (mid_1[711:704] > top_1[703:696]) ? 1 : 0;
assign detect_max[87][4] = (mid_1[711:704] > top_1[711:704]) ? 1 : 0;
assign detect_max[87][5] = (mid_1[711:704] > top_1[719:712]) ? 1 : 0;
assign detect_max[87][6] = (mid_1[711:704] > top_2[703:696]) ? 1 : 0;
assign detect_max[87][7] = (mid_1[711:704] > top_2[711:704]) ? 1 : 0;
assign detect_max[87][8] = (mid_1[711:704] > top_2[719:712]) ? 1 : 0;
assign detect_max[87][9] = (mid_1[711:704] > mid_0[703:696]) ? 1 : 0;
assign detect_max[87][10] = (mid_1[711:704] > mid_0[711:704]) ? 1 : 0;
assign detect_max[87][11] = (mid_1[711:704] > mid_0[719:712]) ? 1 : 0;
assign detect_max[87][12] = (mid_1[711:704] > mid_1[703:696]) ? 1 : 0;
assign detect_max[87][13] = (mid_1[711:704] > mid_1[719:712]) ? 1 : 0;
assign detect_max[87][14] = (mid_1[711:704] > mid_2[703:696]) ? 1 : 0;
assign detect_max[87][15] = (mid_1[711:704] > mid_2[711:704]) ? 1 : 0;
assign detect_max[87][16] = (mid_1[711:704] > mid_2[719:712]) ? 1 : 0;
assign detect_max[87][17] = (mid_1[711:704] > btm_0[703:696]) ? 1 : 0;
assign detect_max[87][18] = (mid_1[711:704] > btm_0[711:704]) ? 1 : 0;
assign detect_max[87][19] = (mid_1[711:704] > btm_0[719:712]) ? 1 : 0;
assign detect_max[87][20] = (mid_1[711:704] > btm_1[703:696]) ? 1 : 0;
assign detect_max[87][21] = (mid_1[711:704] > btm_1[711:704]) ? 1 : 0;
assign detect_max[87][22] = (mid_1[711:704] > btm_1[719:712]) ? 1 : 0;
assign detect_max[87][23] = (mid_1[711:704] > btm_2[703:696]) ? 1 : 0;
assign detect_max[87][24] = (mid_1[711:704] > btm_2[711:704]) ? 1 : 0;
assign detect_max[87][25] = (mid_1[711:704] > btm_2[719:712]) ? 1 : 0;

assign detect_max[88][0] = (mid_1[719:712] > top_0[711:704]) ? 1 : 0;
assign detect_max[88][1] = (mid_1[719:712] > top_0[719:712]) ? 1 : 0;
assign detect_max[88][2] = (mid_1[719:712] > top_0[727:720]) ? 1 : 0;
assign detect_max[88][3] = (mid_1[719:712] > top_1[711:704]) ? 1 : 0;
assign detect_max[88][4] = (mid_1[719:712] > top_1[719:712]) ? 1 : 0;
assign detect_max[88][5] = (mid_1[719:712] > top_1[727:720]) ? 1 : 0;
assign detect_max[88][6] = (mid_1[719:712] > top_2[711:704]) ? 1 : 0;
assign detect_max[88][7] = (mid_1[719:712] > top_2[719:712]) ? 1 : 0;
assign detect_max[88][8] = (mid_1[719:712] > top_2[727:720]) ? 1 : 0;
assign detect_max[88][9] = (mid_1[719:712] > mid_0[711:704]) ? 1 : 0;
assign detect_max[88][10] = (mid_1[719:712] > mid_0[719:712]) ? 1 : 0;
assign detect_max[88][11] = (mid_1[719:712] > mid_0[727:720]) ? 1 : 0;
assign detect_max[88][12] = (mid_1[719:712] > mid_1[711:704]) ? 1 : 0;
assign detect_max[88][13] = (mid_1[719:712] > mid_1[727:720]) ? 1 : 0;
assign detect_max[88][14] = (mid_1[719:712] > mid_2[711:704]) ? 1 : 0;
assign detect_max[88][15] = (mid_1[719:712] > mid_2[719:712]) ? 1 : 0;
assign detect_max[88][16] = (mid_1[719:712] > mid_2[727:720]) ? 1 : 0;
assign detect_max[88][17] = (mid_1[719:712] > btm_0[711:704]) ? 1 : 0;
assign detect_max[88][18] = (mid_1[719:712] > btm_0[719:712]) ? 1 : 0;
assign detect_max[88][19] = (mid_1[719:712] > btm_0[727:720]) ? 1 : 0;
assign detect_max[88][20] = (mid_1[719:712] > btm_1[711:704]) ? 1 : 0;
assign detect_max[88][21] = (mid_1[719:712] > btm_1[719:712]) ? 1 : 0;
assign detect_max[88][22] = (mid_1[719:712] > btm_1[727:720]) ? 1 : 0;
assign detect_max[88][23] = (mid_1[719:712] > btm_2[711:704]) ? 1 : 0;
assign detect_max[88][24] = (mid_1[719:712] > btm_2[719:712]) ? 1 : 0;
assign detect_max[88][25] = (mid_1[719:712] > btm_2[727:720]) ? 1 : 0;

assign detect_max[89][0] = (mid_1[727:720] > top_0[719:712]) ? 1 : 0;
assign detect_max[89][1] = (mid_1[727:720] > top_0[727:720]) ? 1 : 0;
assign detect_max[89][2] = (mid_1[727:720] > top_0[735:728]) ? 1 : 0;
assign detect_max[89][3] = (mid_1[727:720] > top_1[719:712]) ? 1 : 0;
assign detect_max[89][4] = (mid_1[727:720] > top_1[727:720]) ? 1 : 0;
assign detect_max[89][5] = (mid_1[727:720] > top_1[735:728]) ? 1 : 0;
assign detect_max[89][6] = (mid_1[727:720] > top_2[719:712]) ? 1 : 0;
assign detect_max[89][7] = (mid_1[727:720] > top_2[727:720]) ? 1 : 0;
assign detect_max[89][8] = (mid_1[727:720] > top_2[735:728]) ? 1 : 0;
assign detect_max[89][9] = (mid_1[727:720] > mid_0[719:712]) ? 1 : 0;
assign detect_max[89][10] = (mid_1[727:720] > mid_0[727:720]) ? 1 : 0;
assign detect_max[89][11] = (mid_1[727:720] > mid_0[735:728]) ? 1 : 0;
assign detect_max[89][12] = (mid_1[727:720] > mid_1[719:712]) ? 1 : 0;
assign detect_max[89][13] = (mid_1[727:720] > mid_1[735:728]) ? 1 : 0;
assign detect_max[89][14] = (mid_1[727:720] > mid_2[719:712]) ? 1 : 0;
assign detect_max[89][15] = (mid_1[727:720] > mid_2[727:720]) ? 1 : 0;
assign detect_max[89][16] = (mid_1[727:720] > mid_2[735:728]) ? 1 : 0;
assign detect_max[89][17] = (mid_1[727:720] > btm_0[719:712]) ? 1 : 0;
assign detect_max[89][18] = (mid_1[727:720] > btm_0[727:720]) ? 1 : 0;
assign detect_max[89][19] = (mid_1[727:720] > btm_0[735:728]) ? 1 : 0;
assign detect_max[89][20] = (mid_1[727:720] > btm_1[719:712]) ? 1 : 0;
assign detect_max[89][21] = (mid_1[727:720] > btm_1[727:720]) ? 1 : 0;
assign detect_max[89][22] = (mid_1[727:720] > btm_1[735:728]) ? 1 : 0;
assign detect_max[89][23] = (mid_1[727:720] > btm_2[719:712]) ? 1 : 0;
assign detect_max[89][24] = (mid_1[727:720] > btm_2[727:720]) ? 1 : 0;
assign detect_max[89][25] = (mid_1[727:720] > btm_2[735:728]) ? 1 : 0;

assign detect_max[90][0] = (mid_1[735:728] > top_0[727:720]) ? 1 : 0;
assign detect_max[90][1] = (mid_1[735:728] > top_0[735:728]) ? 1 : 0;
assign detect_max[90][2] = (mid_1[735:728] > top_0[743:736]) ? 1 : 0;
assign detect_max[90][3] = (mid_1[735:728] > top_1[727:720]) ? 1 : 0;
assign detect_max[90][4] = (mid_1[735:728] > top_1[735:728]) ? 1 : 0;
assign detect_max[90][5] = (mid_1[735:728] > top_1[743:736]) ? 1 : 0;
assign detect_max[90][6] = (mid_1[735:728] > top_2[727:720]) ? 1 : 0;
assign detect_max[90][7] = (mid_1[735:728] > top_2[735:728]) ? 1 : 0;
assign detect_max[90][8] = (mid_1[735:728] > top_2[743:736]) ? 1 : 0;
assign detect_max[90][9] = (mid_1[735:728] > mid_0[727:720]) ? 1 : 0;
assign detect_max[90][10] = (mid_1[735:728] > mid_0[735:728]) ? 1 : 0;
assign detect_max[90][11] = (mid_1[735:728] > mid_0[743:736]) ? 1 : 0;
assign detect_max[90][12] = (mid_1[735:728] > mid_1[727:720]) ? 1 : 0;
assign detect_max[90][13] = (mid_1[735:728] > mid_1[743:736]) ? 1 : 0;
assign detect_max[90][14] = (mid_1[735:728] > mid_2[727:720]) ? 1 : 0;
assign detect_max[90][15] = (mid_1[735:728] > mid_2[735:728]) ? 1 : 0;
assign detect_max[90][16] = (mid_1[735:728] > mid_2[743:736]) ? 1 : 0;
assign detect_max[90][17] = (mid_1[735:728] > btm_0[727:720]) ? 1 : 0;
assign detect_max[90][18] = (mid_1[735:728] > btm_0[735:728]) ? 1 : 0;
assign detect_max[90][19] = (mid_1[735:728] > btm_0[743:736]) ? 1 : 0;
assign detect_max[90][20] = (mid_1[735:728] > btm_1[727:720]) ? 1 : 0;
assign detect_max[90][21] = (mid_1[735:728] > btm_1[735:728]) ? 1 : 0;
assign detect_max[90][22] = (mid_1[735:728] > btm_1[743:736]) ? 1 : 0;
assign detect_max[90][23] = (mid_1[735:728] > btm_2[727:720]) ? 1 : 0;
assign detect_max[90][24] = (mid_1[735:728] > btm_2[735:728]) ? 1 : 0;
assign detect_max[90][25] = (mid_1[735:728] > btm_2[743:736]) ? 1 : 0;

assign detect_max[91][0] = (mid_1[743:736] > top_0[735:728]) ? 1 : 0;
assign detect_max[91][1] = (mid_1[743:736] > top_0[743:736]) ? 1 : 0;
assign detect_max[91][2] = (mid_1[743:736] > top_0[751:744]) ? 1 : 0;
assign detect_max[91][3] = (mid_1[743:736] > top_1[735:728]) ? 1 : 0;
assign detect_max[91][4] = (mid_1[743:736] > top_1[743:736]) ? 1 : 0;
assign detect_max[91][5] = (mid_1[743:736] > top_1[751:744]) ? 1 : 0;
assign detect_max[91][6] = (mid_1[743:736] > top_2[735:728]) ? 1 : 0;
assign detect_max[91][7] = (mid_1[743:736] > top_2[743:736]) ? 1 : 0;
assign detect_max[91][8] = (mid_1[743:736] > top_2[751:744]) ? 1 : 0;
assign detect_max[91][9] = (mid_1[743:736] > mid_0[735:728]) ? 1 : 0;
assign detect_max[91][10] = (mid_1[743:736] > mid_0[743:736]) ? 1 : 0;
assign detect_max[91][11] = (mid_1[743:736] > mid_0[751:744]) ? 1 : 0;
assign detect_max[91][12] = (mid_1[743:736] > mid_1[735:728]) ? 1 : 0;
assign detect_max[91][13] = (mid_1[743:736] > mid_1[751:744]) ? 1 : 0;
assign detect_max[91][14] = (mid_1[743:736] > mid_2[735:728]) ? 1 : 0;
assign detect_max[91][15] = (mid_1[743:736] > mid_2[743:736]) ? 1 : 0;
assign detect_max[91][16] = (mid_1[743:736] > mid_2[751:744]) ? 1 : 0;
assign detect_max[91][17] = (mid_1[743:736] > btm_0[735:728]) ? 1 : 0;
assign detect_max[91][18] = (mid_1[743:736] > btm_0[743:736]) ? 1 : 0;
assign detect_max[91][19] = (mid_1[743:736] > btm_0[751:744]) ? 1 : 0;
assign detect_max[91][20] = (mid_1[743:736] > btm_1[735:728]) ? 1 : 0;
assign detect_max[91][21] = (mid_1[743:736] > btm_1[743:736]) ? 1 : 0;
assign detect_max[91][22] = (mid_1[743:736] > btm_1[751:744]) ? 1 : 0;
assign detect_max[91][23] = (mid_1[743:736] > btm_2[735:728]) ? 1 : 0;
assign detect_max[91][24] = (mid_1[743:736] > btm_2[743:736]) ? 1 : 0;
assign detect_max[91][25] = (mid_1[743:736] > btm_2[751:744]) ? 1 : 0;

assign detect_max[92][0] = (mid_1[751:744] > top_0[743:736]) ? 1 : 0;
assign detect_max[92][1] = (mid_1[751:744] > top_0[751:744]) ? 1 : 0;
assign detect_max[92][2] = (mid_1[751:744] > top_0[759:752]) ? 1 : 0;
assign detect_max[92][3] = (mid_1[751:744] > top_1[743:736]) ? 1 : 0;
assign detect_max[92][4] = (mid_1[751:744] > top_1[751:744]) ? 1 : 0;
assign detect_max[92][5] = (mid_1[751:744] > top_1[759:752]) ? 1 : 0;
assign detect_max[92][6] = (mid_1[751:744] > top_2[743:736]) ? 1 : 0;
assign detect_max[92][7] = (mid_1[751:744] > top_2[751:744]) ? 1 : 0;
assign detect_max[92][8] = (mid_1[751:744] > top_2[759:752]) ? 1 : 0;
assign detect_max[92][9] = (mid_1[751:744] > mid_0[743:736]) ? 1 : 0;
assign detect_max[92][10] = (mid_1[751:744] > mid_0[751:744]) ? 1 : 0;
assign detect_max[92][11] = (mid_1[751:744] > mid_0[759:752]) ? 1 : 0;
assign detect_max[92][12] = (mid_1[751:744] > mid_1[743:736]) ? 1 : 0;
assign detect_max[92][13] = (mid_1[751:744] > mid_1[759:752]) ? 1 : 0;
assign detect_max[92][14] = (mid_1[751:744] > mid_2[743:736]) ? 1 : 0;
assign detect_max[92][15] = (mid_1[751:744] > mid_2[751:744]) ? 1 : 0;
assign detect_max[92][16] = (mid_1[751:744] > mid_2[759:752]) ? 1 : 0;
assign detect_max[92][17] = (mid_1[751:744] > btm_0[743:736]) ? 1 : 0;
assign detect_max[92][18] = (mid_1[751:744] > btm_0[751:744]) ? 1 : 0;
assign detect_max[92][19] = (mid_1[751:744] > btm_0[759:752]) ? 1 : 0;
assign detect_max[92][20] = (mid_1[751:744] > btm_1[743:736]) ? 1 : 0;
assign detect_max[92][21] = (mid_1[751:744] > btm_1[751:744]) ? 1 : 0;
assign detect_max[92][22] = (mid_1[751:744] > btm_1[759:752]) ? 1 : 0;
assign detect_max[92][23] = (mid_1[751:744] > btm_2[743:736]) ? 1 : 0;
assign detect_max[92][24] = (mid_1[751:744] > btm_2[751:744]) ? 1 : 0;
assign detect_max[92][25] = (mid_1[751:744] > btm_2[759:752]) ? 1 : 0;

assign detect_max[93][0] = (mid_1[759:752] > top_0[751:744]) ? 1 : 0;
assign detect_max[93][1] = (mid_1[759:752] > top_0[759:752]) ? 1 : 0;
assign detect_max[93][2] = (mid_1[759:752] > top_0[767:760]) ? 1 : 0;
assign detect_max[93][3] = (mid_1[759:752] > top_1[751:744]) ? 1 : 0;
assign detect_max[93][4] = (mid_1[759:752] > top_1[759:752]) ? 1 : 0;
assign detect_max[93][5] = (mid_1[759:752] > top_1[767:760]) ? 1 : 0;
assign detect_max[93][6] = (mid_1[759:752] > top_2[751:744]) ? 1 : 0;
assign detect_max[93][7] = (mid_1[759:752] > top_2[759:752]) ? 1 : 0;
assign detect_max[93][8] = (mid_1[759:752] > top_2[767:760]) ? 1 : 0;
assign detect_max[93][9] = (mid_1[759:752] > mid_0[751:744]) ? 1 : 0;
assign detect_max[93][10] = (mid_1[759:752] > mid_0[759:752]) ? 1 : 0;
assign detect_max[93][11] = (mid_1[759:752] > mid_0[767:760]) ? 1 : 0;
assign detect_max[93][12] = (mid_1[759:752] > mid_1[751:744]) ? 1 : 0;
assign detect_max[93][13] = (mid_1[759:752] > mid_1[767:760]) ? 1 : 0;
assign detect_max[93][14] = (mid_1[759:752] > mid_2[751:744]) ? 1 : 0;
assign detect_max[93][15] = (mid_1[759:752] > mid_2[759:752]) ? 1 : 0;
assign detect_max[93][16] = (mid_1[759:752] > mid_2[767:760]) ? 1 : 0;
assign detect_max[93][17] = (mid_1[759:752] > btm_0[751:744]) ? 1 : 0;
assign detect_max[93][18] = (mid_1[759:752] > btm_0[759:752]) ? 1 : 0;
assign detect_max[93][19] = (mid_1[759:752] > btm_0[767:760]) ? 1 : 0;
assign detect_max[93][20] = (mid_1[759:752] > btm_1[751:744]) ? 1 : 0;
assign detect_max[93][21] = (mid_1[759:752] > btm_1[759:752]) ? 1 : 0;
assign detect_max[93][22] = (mid_1[759:752] > btm_1[767:760]) ? 1 : 0;
assign detect_max[93][23] = (mid_1[759:752] > btm_2[751:744]) ? 1 : 0;
assign detect_max[93][24] = (mid_1[759:752] > btm_2[759:752]) ? 1 : 0;
assign detect_max[93][25] = (mid_1[759:752] > btm_2[767:760]) ? 1 : 0;

assign detect_max[94][0] = (mid_1[767:760] > top_0[759:752]) ? 1 : 0;
assign detect_max[94][1] = (mid_1[767:760] > top_0[767:760]) ? 1 : 0;
assign detect_max[94][2] = (mid_1[767:760] > top_0[775:768]) ? 1 : 0;
assign detect_max[94][3] = (mid_1[767:760] > top_1[759:752]) ? 1 : 0;
assign detect_max[94][4] = (mid_1[767:760] > top_1[767:760]) ? 1 : 0;
assign detect_max[94][5] = (mid_1[767:760] > top_1[775:768]) ? 1 : 0;
assign detect_max[94][6] = (mid_1[767:760] > top_2[759:752]) ? 1 : 0;
assign detect_max[94][7] = (mid_1[767:760] > top_2[767:760]) ? 1 : 0;
assign detect_max[94][8] = (mid_1[767:760] > top_2[775:768]) ? 1 : 0;
assign detect_max[94][9] = (mid_1[767:760] > mid_0[759:752]) ? 1 : 0;
assign detect_max[94][10] = (mid_1[767:760] > mid_0[767:760]) ? 1 : 0;
assign detect_max[94][11] = (mid_1[767:760] > mid_0[775:768]) ? 1 : 0;
assign detect_max[94][12] = (mid_1[767:760] > mid_1[759:752]) ? 1 : 0;
assign detect_max[94][13] = (mid_1[767:760] > mid_1[775:768]) ? 1 : 0;
assign detect_max[94][14] = (mid_1[767:760] > mid_2[759:752]) ? 1 : 0;
assign detect_max[94][15] = (mid_1[767:760] > mid_2[767:760]) ? 1 : 0;
assign detect_max[94][16] = (mid_1[767:760] > mid_2[775:768]) ? 1 : 0;
assign detect_max[94][17] = (mid_1[767:760] > btm_0[759:752]) ? 1 : 0;
assign detect_max[94][18] = (mid_1[767:760] > btm_0[767:760]) ? 1 : 0;
assign detect_max[94][19] = (mid_1[767:760] > btm_0[775:768]) ? 1 : 0;
assign detect_max[94][20] = (mid_1[767:760] > btm_1[759:752]) ? 1 : 0;
assign detect_max[94][21] = (mid_1[767:760] > btm_1[767:760]) ? 1 : 0;
assign detect_max[94][22] = (mid_1[767:760] > btm_1[775:768]) ? 1 : 0;
assign detect_max[94][23] = (mid_1[767:760] > btm_2[759:752]) ? 1 : 0;
assign detect_max[94][24] = (mid_1[767:760] > btm_2[767:760]) ? 1 : 0;
assign detect_max[94][25] = (mid_1[767:760] > btm_2[775:768]) ? 1 : 0;

assign detect_max[95][0] = (mid_1[775:768] > top_0[767:760]) ? 1 : 0;
assign detect_max[95][1] = (mid_1[775:768] > top_0[775:768]) ? 1 : 0;
assign detect_max[95][2] = (mid_1[775:768] > top_0[783:776]) ? 1 : 0;
assign detect_max[95][3] = (mid_1[775:768] > top_1[767:760]) ? 1 : 0;
assign detect_max[95][4] = (mid_1[775:768] > top_1[775:768]) ? 1 : 0;
assign detect_max[95][5] = (mid_1[775:768] > top_1[783:776]) ? 1 : 0;
assign detect_max[95][6] = (mid_1[775:768] > top_2[767:760]) ? 1 : 0;
assign detect_max[95][7] = (mid_1[775:768] > top_2[775:768]) ? 1 : 0;
assign detect_max[95][8] = (mid_1[775:768] > top_2[783:776]) ? 1 : 0;
assign detect_max[95][9] = (mid_1[775:768] > mid_0[767:760]) ? 1 : 0;
assign detect_max[95][10] = (mid_1[775:768] > mid_0[775:768]) ? 1 : 0;
assign detect_max[95][11] = (mid_1[775:768] > mid_0[783:776]) ? 1 : 0;
assign detect_max[95][12] = (mid_1[775:768] > mid_1[767:760]) ? 1 : 0;
assign detect_max[95][13] = (mid_1[775:768] > mid_1[783:776]) ? 1 : 0;
assign detect_max[95][14] = (mid_1[775:768] > mid_2[767:760]) ? 1 : 0;
assign detect_max[95][15] = (mid_1[775:768] > mid_2[775:768]) ? 1 : 0;
assign detect_max[95][16] = (mid_1[775:768] > mid_2[783:776]) ? 1 : 0;
assign detect_max[95][17] = (mid_1[775:768] > btm_0[767:760]) ? 1 : 0;
assign detect_max[95][18] = (mid_1[775:768] > btm_0[775:768]) ? 1 : 0;
assign detect_max[95][19] = (mid_1[775:768] > btm_0[783:776]) ? 1 : 0;
assign detect_max[95][20] = (mid_1[775:768] > btm_1[767:760]) ? 1 : 0;
assign detect_max[95][21] = (mid_1[775:768] > btm_1[775:768]) ? 1 : 0;
assign detect_max[95][22] = (mid_1[775:768] > btm_1[783:776]) ? 1 : 0;
assign detect_max[95][23] = (mid_1[775:768] > btm_2[767:760]) ? 1 : 0;
assign detect_max[95][24] = (mid_1[775:768] > btm_2[775:768]) ? 1 : 0;
assign detect_max[95][25] = (mid_1[775:768] > btm_2[783:776]) ? 1 : 0;

assign detect_max[96][0] = (mid_1[783:776] > top_0[775:768]) ? 1 : 0;
assign detect_max[96][1] = (mid_1[783:776] > top_0[783:776]) ? 1 : 0;
assign detect_max[96][2] = (mid_1[783:776] > top_0[791:784]) ? 1 : 0;
assign detect_max[96][3] = (mid_1[783:776] > top_1[775:768]) ? 1 : 0;
assign detect_max[96][4] = (mid_1[783:776] > top_1[783:776]) ? 1 : 0;
assign detect_max[96][5] = (mid_1[783:776] > top_1[791:784]) ? 1 : 0;
assign detect_max[96][6] = (mid_1[783:776] > top_2[775:768]) ? 1 : 0;
assign detect_max[96][7] = (mid_1[783:776] > top_2[783:776]) ? 1 : 0;
assign detect_max[96][8] = (mid_1[783:776] > top_2[791:784]) ? 1 : 0;
assign detect_max[96][9] = (mid_1[783:776] > mid_0[775:768]) ? 1 : 0;
assign detect_max[96][10] = (mid_1[783:776] > mid_0[783:776]) ? 1 : 0;
assign detect_max[96][11] = (mid_1[783:776] > mid_0[791:784]) ? 1 : 0;
assign detect_max[96][12] = (mid_1[783:776] > mid_1[775:768]) ? 1 : 0;
assign detect_max[96][13] = (mid_1[783:776] > mid_1[791:784]) ? 1 : 0;
assign detect_max[96][14] = (mid_1[783:776] > mid_2[775:768]) ? 1 : 0;
assign detect_max[96][15] = (mid_1[783:776] > mid_2[783:776]) ? 1 : 0;
assign detect_max[96][16] = (mid_1[783:776] > mid_2[791:784]) ? 1 : 0;
assign detect_max[96][17] = (mid_1[783:776] > btm_0[775:768]) ? 1 : 0;
assign detect_max[96][18] = (mid_1[783:776] > btm_0[783:776]) ? 1 : 0;
assign detect_max[96][19] = (mid_1[783:776] > btm_0[791:784]) ? 1 : 0;
assign detect_max[96][20] = (mid_1[783:776] > btm_1[775:768]) ? 1 : 0;
assign detect_max[96][21] = (mid_1[783:776] > btm_1[783:776]) ? 1 : 0;
assign detect_max[96][22] = (mid_1[783:776] > btm_1[791:784]) ? 1 : 0;
assign detect_max[96][23] = (mid_1[783:776] > btm_2[775:768]) ? 1 : 0;
assign detect_max[96][24] = (mid_1[783:776] > btm_2[783:776]) ? 1 : 0;
assign detect_max[96][25] = (mid_1[783:776] > btm_2[791:784]) ? 1 : 0;

assign detect_max[97][0] = (mid_1[791:784] > top_0[783:776]) ? 1 : 0;
assign detect_max[97][1] = (mid_1[791:784] > top_0[791:784]) ? 1 : 0;
assign detect_max[97][2] = (mid_1[791:784] > top_0[799:792]) ? 1 : 0;
assign detect_max[97][3] = (mid_1[791:784] > top_1[783:776]) ? 1 : 0;
assign detect_max[97][4] = (mid_1[791:784] > top_1[791:784]) ? 1 : 0;
assign detect_max[97][5] = (mid_1[791:784] > top_1[799:792]) ? 1 : 0;
assign detect_max[97][6] = (mid_1[791:784] > top_2[783:776]) ? 1 : 0;
assign detect_max[97][7] = (mid_1[791:784] > top_2[791:784]) ? 1 : 0;
assign detect_max[97][8] = (mid_1[791:784] > top_2[799:792]) ? 1 : 0;
assign detect_max[97][9] = (mid_1[791:784] > mid_0[783:776]) ? 1 : 0;
assign detect_max[97][10] = (mid_1[791:784] > mid_0[791:784]) ? 1 : 0;
assign detect_max[97][11] = (mid_1[791:784] > mid_0[799:792]) ? 1 : 0;
assign detect_max[97][12] = (mid_1[791:784] > mid_1[783:776]) ? 1 : 0;
assign detect_max[97][13] = (mid_1[791:784] > mid_1[799:792]) ? 1 : 0;
assign detect_max[97][14] = (mid_1[791:784] > mid_2[783:776]) ? 1 : 0;
assign detect_max[97][15] = (mid_1[791:784] > mid_2[791:784]) ? 1 : 0;
assign detect_max[97][16] = (mid_1[791:784] > mid_2[799:792]) ? 1 : 0;
assign detect_max[97][17] = (mid_1[791:784] > btm_0[783:776]) ? 1 : 0;
assign detect_max[97][18] = (mid_1[791:784] > btm_0[791:784]) ? 1 : 0;
assign detect_max[97][19] = (mid_1[791:784] > btm_0[799:792]) ? 1 : 0;
assign detect_max[97][20] = (mid_1[791:784] > btm_1[783:776]) ? 1 : 0;
assign detect_max[97][21] = (mid_1[791:784] > btm_1[791:784]) ? 1 : 0;
assign detect_max[97][22] = (mid_1[791:784] > btm_1[799:792]) ? 1 : 0;
assign detect_max[97][23] = (mid_1[791:784] > btm_2[783:776]) ? 1 : 0;
assign detect_max[97][24] = (mid_1[791:784] > btm_2[791:784]) ? 1 : 0;
assign detect_max[97][25] = (mid_1[791:784] > btm_2[799:792]) ? 1 : 0;

assign detect_max[98][0] = (mid_1[799:792] > top_0[791:784]) ? 1 : 0;
assign detect_max[98][1] = (mid_1[799:792] > top_0[799:792]) ? 1 : 0;
assign detect_max[98][2] = (mid_1[799:792] > top_0[807:800]) ? 1 : 0;
assign detect_max[98][3] = (mid_1[799:792] > top_1[791:784]) ? 1 : 0;
assign detect_max[98][4] = (mid_1[799:792] > top_1[799:792]) ? 1 : 0;
assign detect_max[98][5] = (mid_1[799:792] > top_1[807:800]) ? 1 : 0;
assign detect_max[98][6] = (mid_1[799:792] > top_2[791:784]) ? 1 : 0;
assign detect_max[98][7] = (mid_1[799:792] > top_2[799:792]) ? 1 : 0;
assign detect_max[98][8] = (mid_1[799:792] > top_2[807:800]) ? 1 : 0;
assign detect_max[98][9] = (mid_1[799:792] > mid_0[791:784]) ? 1 : 0;
assign detect_max[98][10] = (mid_1[799:792] > mid_0[799:792]) ? 1 : 0;
assign detect_max[98][11] = (mid_1[799:792] > mid_0[807:800]) ? 1 : 0;
assign detect_max[98][12] = (mid_1[799:792] > mid_1[791:784]) ? 1 : 0;
assign detect_max[98][13] = (mid_1[799:792] > mid_1[807:800]) ? 1 : 0;
assign detect_max[98][14] = (mid_1[799:792] > mid_2[791:784]) ? 1 : 0;
assign detect_max[98][15] = (mid_1[799:792] > mid_2[799:792]) ? 1 : 0;
assign detect_max[98][16] = (mid_1[799:792] > mid_2[807:800]) ? 1 : 0;
assign detect_max[98][17] = (mid_1[799:792] > btm_0[791:784]) ? 1 : 0;
assign detect_max[98][18] = (mid_1[799:792] > btm_0[799:792]) ? 1 : 0;
assign detect_max[98][19] = (mid_1[799:792] > btm_0[807:800]) ? 1 : 0;
assign detect_max[98][20] = (mid_1[799:792] > btm_1[791:784]) ? 1 : 0;
assign detect_max[98][21] = (mid_1[799:792] > btm_1[799:792]) ? 1 : 0;
assign detect_max[98][22] = (mid_1[799:792] > btm_1[807:800]) ? 1 : 0;
assign detect_max[98][23] = (mid_1[799:792] > btm_2[791:784]) ? 1 : 0;
assign detect_max[98][24] = (mid_1[799:792] > btm_2[799:792]) ? 1 : 0;
assign detect_max[98][25] = (mid_1[799:792] > btm_2[807:800]) ? 1 : 0;

assign detect_max[99][0] = (mid_1[807:800] > top_0[799:792]) ? 1 : 0;
assign detect_max[99][1] = (mid_1[807:800] > top_0[807:800]) ? 1 : 0;
assign detect_max[99][2] = (mid_1[807:800] > top_0[815:808]) ? 1 : 0;
assign detect_max[99][3] = (mid_1[807:800] > top_1[799:792]) ? 1 : 0;
assign detect_max[99][4] = (mid_1[807:800] > top_1[807:800]) ? 1 : 0;
assign detect_max[99][5] = (mid_1[807:800] > top_1[815:808]) ? 1 : 0;
assign detect_max[99][6] = (mid_1[807:800] > top_2[799:792]) ? 1 : 0;
assign detect_max[99][7] = (mid_1[807:800] > top_2[807:800]) ? 1 : 0;
assign detect_max[99][8] = (mid_1[807:800] > top_2[815:808]) ? 1 : 0;
assign detect_max[99][9] = (mid_1[807:800] > mid_0[799:792]) ? 1 : 0;
assign detect_max[99][10] = (mid_1[807:800] > mid_0[807:800]) ? 1 : 0;
assign detect_max[99][11] = (mid_1[807:800] > mid_0[815:808]) ? 1 : 0;
assign detect_max[99][12] = (mid_1[807:800] > mid_1[799:792]) ? 1 : 0;
assign detect_max[99][13] = (mid_1[807:800] > mid_1[815:808]) ? 1 : 0;
assign detect_max[99][14] = (mid_1[807:800] > mid_2[799:792]) ? 1 : 0;
assign detect_max[99][15] = (mid_1[807:800] > mid_2[807:800]) ? 1 : 0;
assign detect_max[99][16] = (mid_1[807:800] > mid_2[815:808]) ? 1 : 0;
assign detect_max[99][17] = (mid_1[807:800] > btm_0[799:792]) ? 1 : 0;
assign detect_max[99][18] = (mid_1[807:800] > btm_0[807:800]) ? 1 : 0;
assign detect_max[99][19] = (mid_1[807:800] > btm_0[815:808]) ? 1 : 0;
assign detect_max[99][20] = (mid_1[807:800] > btm_1[799:792]) ? 1 : 0;
assign detect_max[99][21] = (mid_1[807:800] > btm_1[807:800]) ? 1 : 0;
assign detect_max[99][22] = (mid_1[807:800] > btm_1[815:808]) ? 1 : 0;
assign detect_max[99][23] = (mid_1[807:800] > btm_2[799:792]) ? 1 : 0;
assign detect_max[99][24] = (mid_1[807:800] > btm_2[807:800]) ? 1 : 0;
assign detect_max[99][25] = (mid_1[807:800] > btm_2[815:808]) ? 1 : 0;

assign detect_max[100][0] = (mid_1[815:808] > top_0[807:800]) ? 1 : 0;
assign detect_max[100][1] = (mid_1[815:808] > top_0[815:808]) ? 1 : 0;
assign detect_max[100][2] = (mid_1[815:808] > top_0[823:816]) ? 1 : 0;
assign detect_max[100][3] = (mid_1[815:808] > top_1[807:800]) ? 1 : 0;
assign detect_max[100][4] = (mid_1[815:808] > top_1[815:808]) ? 1 : 0;
assign detect_max[100][5] = (mid_1[815:808] > top_1[823:816]) ? 1 : 0;
assign detect_max[100][6] = (mid_1[815:808] > top_2[807:800]) ? 1 : 0;
assign detect_max[100][7] = (mid_1[815:808] > top_2[815:808]) ? 1 : 0;
assign detect_max[100][8] = (mid_1[815:808] > top_2[823:816]) ? 1 : 0;
assign detect_max[100][9] = (mid_1[815:808] > mid_0[807:800]) ? 1 : 0;
assign detect_max[100][10] = (mid_1[815:808] > mid_0[815:808]) ? 1 : 0;
assign detect_max[100][11] = (mid_1[815:808] > mid_0[823:816]) ? 1 : 0;
assign detect_max[100][12] = (mid_1[815:808] > mid_1[807:800]) ? 1 : 0;
assign detect_max[100][13] = (mid_1[815:808] > mid_1[823:816]) ? 1 : 0;
assign detect_max[100][14] = (mid_1[815:808] > mid_2[807:800]) ? 1 : 0;
assign detect_max[100][15] = (mid_1[815:808] > mid_2[815:808]) ? 1 : 0;
assign detect_max[100][16] = (mid_1[815:808] > mid_2[823:816]) ? 1 : 0;
assign detect_max[100][17] = (mid_1[815:808] > btm_0[807:800]) ? 1 : 0;
assign detect_max[100][18] = (mid_1[815:808] > btm_0[815:808]) ? 1 : 0;
assign detect_max[100][19] = (mid_1[815:808] > btm_0[823:816]) ? 1 : 0;
assign detect_max[100][20] = (mid_1[815:808] > btm_1[807:800]) ? 1 : 0;
assign detect_max[100][21] = (mid_1[815:808] > btm_1[815:808]) ? 1 : 0;
assign detect_max[100][22] = (mid_1[815:808] > btm_1[823:816]) ? 1 : 0;
assign detect_max[100][23] = (mid_1[815:808] > btm_2[807:800]) ? 1 : 0;
assign detect_max[100][24] = (mid_1[815:808] > btm_2[815:808]) ? 1 : 0;
assign detect_max[100][25] = (mid_1[815:808] > btm_2[823:816]) ? 1 : 0;

assign detect_max[101][0] = (mid_1[823:816] > top_0[815:808]) ? 1 : 0;
assign detect_max[101][1] = (mid_1[823:816] > top_0[823:816]) ? 1 : 0;
assign detect_max[101][2] = (mid_1[823:816] > top_0[831:824]) ? 1 : 0;
assign detect_max[101][3] = (mid_1[823:816] > top_1[815:808]) ? 1 : 0;
assign detect_max[101][4] = (mid_1[823:816] > top_1[823:816]) ? 1 : 0;
assign detect_max[101][5] = (mid_1[823:816] > top_1[831:824]) ? 1 : 0;
assign detect_max[101][6] = (mid_1[823:816] > top_2[815:808]) ? 1 : 0;
assign detect_max[101][7] = (mid_1[823:816] > top_2[823:816]) ? 1 : 0;
assign detect_max[101][8] = (mid_1[823:816] > top_2[831:824]) ? 1 : 0;
assign detect_max[101][9] = (mid_1[823:816] > mid_0[815:808]) ? 1 : 0;
assign detect_max[101][10] = (mid_1[823:816] > mid_0[823:816]) ? 1 : 0;
assign detect_max[101][11] = (mid_1[823:816] > mid_0[831:824]) ? 1 : 0;
assign detect_max[101][12] = (mid_1[823:816] > mid_1[815:808]) ? 1 : 0;
assign detect_max[101][13] = (mid_1[823:816] > mid_1[831:824]) ? 1 : 0;
assign detect_max[101][14] = (mid_1[823:816] > mid_2[815:808]) ? 1 : 0;
assign detect_max[101][15] = (mid_1[823:816] > mid_2[823:816]) ? 1 : 0;
assign detect_max[101][16] = (mid_1[823:816] > mid_2[831:824]) ? 1 : 0;
assign detect_max[101][17] = (mid_1[823:816] > btm_0[815:808]) ? 1 : 0;
assign detect_max[101][18] = (mid_1[823:816] > btm_0[823:816]) ? 1 : 0;
assign detect_max[101][19] = (mid_1[823:816] > btm_0[831:824]) ? 1 : 0;
assign detect_max[101][20] = (mid_1[823:816] > btm_1[815:808]) ? 1 : 0;
assign detect_max[101][21] = (mid_1[823:816] > btm_1[823:816]) ? 1 : 0;
assign detect_max[101][22] = (mid_1[823:816] > btm_1[831:824]) ? 1 : 0;
assign detect_max[101][23] = (mid_1[823:816] > btm_2[815:808]) ? 1 : 0;
assign detect_max[101][24] = (mid_1[823:816] > btm_2[823:816]) ? 1 : 0;
assign detect_max[101][25] = (mid_1[823:816] > btm_2[831:824]) ? 1 : 0;

assign detect_max[102][0] = (mid_1[831:824] > top_0[823:816]) ? 1 : 0;
assign detect_max[102][1] = (mid_1[831:824] > top_0[831:824]) ? 1 : 0;
assign detect_max[102][2] = (mid_1[831:824] > top_0[839:832]) ? 1 : 0;
assign detect_max[102][3] = (mid_1[831:824] > top_1[823:816]) ? 1 : 0;
assign detect_max[102][4] = (mid_1[831:824] > top_1[831:824]) ? 1 : 0;
assign detect_max[102][5] = (mid_1[831:824] > top_1[839:832]) ? 1 : 0;
assign detect_max[102][6] = (mid_1[831:824] > top_2[823:816]) ? 1 : 0;
assign detect_max[102][7] = (mid_1[831:824] > top_2[831:824]) ? 1 : 0;
assign detect_max[102][8] = (mid_1[831:824] > top_2[839:832]) ? 1 : 0;
assign detect_max[102][9] = (mid_1[831:824] > mid_0[823:816]) ? 1 : 0;
assign detect_max[102][10] = (mid_1[831:824] > mid_0[831:824]) ? 1 : 0;
assign detect_max[102][11] = (mid_1[831:824] > mid_0[839:832]) ? 1 : 0;
assign detect_max[102][12] = (mid_1[831:824] > mid_1[823:816]) ? 1 : 0;
assign detect_max[102][13] = (mid_1[831:824] > mid_1[839:832]) ? 1 : 0;
assign detect_max[102][14] = (mid_1[831:824] > mid_2[823:816]) ? 1 : 0;
assign detect_max[102][15] = (mid_1[831:824] > mid_2[831:824]) ? 1 : 0;
assign detect_max[102][16] = (mid_1[831:824] > mid_2[839:832]) ? 1 : 0;
assign detect_max[102][17] = (mid_1[831:824] > btm_0[823:816]) ? 1 : 0;
assign detect_max[102][18] = (mid_1[831:824] > btm_0[831:824]) ? 1 : 0;
assign detect_max[102][19] = (mid_1[831:824] > btm_0[839:832]) ? 1 : 0;
assign detect_max[102][20] = (mid_1[831:824] > btm_1[823:816]) ? 1 : 0;
assign detect_max[102][21] = (mid_1[831:824] > btm_1[831:824]) ? 1 : 0;
assign detect_max[102][22] = (mid_1[831:824] > btm_1[839:832]) ? 1 : 0;
assign detect_max[102][23] = (mid_1[831:824] > btm_2[823:816]) ? 1 : 0;
assign detect_max[102][24] = (mid_1[831:824] > btm_2[831:824]) ? 1 : 0;
assign detect_max[102][25] = (mid_1[831:824] > btm_2[839:832]) ? 1 : 0;

assign detect_max[103][0] = (mid_1[839:832] > top_0[831:824]) ? 1 : 0;
assign detect_max[103][1] = (mid_1[839:832] > top_0[839:832]) ? 1 : 0;
assign detect_max[103][2] = (mid_1[839:832] > top_0[847:840]) ? 1 : 0;
assign detect_max[103][3] = (mid_1[839:832] > top_1[831:824]) ? 1 : 0;
assign detect_max[103][4] = (mid_1[839:832] > top_1[839:832]) ? 1 : 0;
assign detect_max[103][5] = (mid_1[839:832] > top_1[847:840]) ? 1 : 0;
assign detect_max[103][6] = (mid_1[839:832] > top_2[831:824]) ? 1 : 0;
assign detect_max[103][7] = (mid_1[839:832] > top_2[839:832]) ? 1 : 0;
assign detect_max[103][8] = (mid_1[839:832] > top_2[847:840]) ? 1 : 0;
assign detect_max[103][9] = (mid_1[839:832] > mid_0[831:824]) ? 1 : 0;
assign detect_max[103][10] = (mid_1[839:832] > mid_0[839:832]) ? 1 : 0;
assign detect_max[103][11] = (mid_1[839:832] > mid_0[847:840]) ? 1 : 0;
assign detect_max[103][12] = (mid_1[839:832] > mid_1[831:824]) ? 1 : 0;
assign detect_max[103][13] = (mid_1[839:832] > mid_1[847:840]) ? 1 : 0;
assign detect_max[103][14] = (mid_1[839:832] > mid_2[831:824]) ? 1 : 0;
assign detect_max[103][15] = (mid_1[839:832] > mid_2[839:832]) ? 1 : 0;
assign detect_max[103][16] = (mid_1[839:832] > mid_2[847:840]) ? 1 : 0;
assign detect_max[103][17] = (mid_1[839:832] > btm_0[831:824]) ? 1 : 0;
assign detect_max[103][18] = (mid_1[839:832] > btm_0[839:832]) ? 1 : 0;
assign detect_max[103][19] = (mid_1[839:832] > btm_0[847:840]) ? 1 : 0;
assign detect_max[103][20] = (mid_1[839:832] > btm_1[831:824]) ? 1 : 0;
assign detect_max[103][21] = (mid_1[839:832] > btm_1[839:832]) ? 1 : 0;
assign detect_max[103][22] = (mid_1[839:832] > btm_1[847:840]) ? 1 : 0;
assign detect_max[103][23] = (mid_1[839:832] > btm_2[831:824]) ? 1 : 0;
assign detect_max[103][24] = (mid_1[839:832] > btm_2[839:832]) ? 1 : 0;
assign detect_max[103][25] = (mid_1[839:832] > btm_2[847:840]) ? 1 : 0;

assign detect_max[104][0] = (mid_1[847:840] > top_0[839:832]) ? 1 : 0;
assign detect_max[104][1] = (mid_1[847:840] > top_0[847:840]) ? 1 : 0;
assign detect_max[104][2] = (mid_1[847:840] > top_0[855:848]) ? 1 : 0;
assign detect_max[104][3] = (mid_1[847:840] > top_1[839:832]) ? 1 : 0;
assign detect_max[104][4] = (mid_1[847:840] > top_1[847:840]) ? 1 : 0;
assign detect_max[104][5] = (mid_1[847:840] > top_1[855:848]) ? 1 : 0;
assign detect_max[104][6] = (mid_1[847:840] > top_2[839:832]) ? 1 : 0;
assign detect_max[104][7] = (mid_1[847:840] > top_2[847:840]) ? 1 : 0;
assign detect_max[104][8] = (mid_1[847:840] > top_2[855:848]) ? 1 : 0;
assign detect_max[104][9] = (mid_1[847:840] > mid_0[839:832]) ? 1 : 0;
assign detect_max[104][10] = (mid_1[847:840] > mid_0[847:840]) ? 1 : 0;
assign detect_max[104][11] = (mid_1[847:840] > mid_0[855:848]) ? 1 : 0;
assign detect_max[104][12] = (mid_1[847:840] > mid_1[839:832]) ? 1 : 0;
assign detect_max[104][13] = (mid_1[847:840] > mid_1[855:848]) ? 1 : 0;
assign detect_max[104][14] = (mid_1[847:840] > mid_2[839:832]) ? 1 : 0;
assign detect_max[104][15] = (mid_1[847:840] > mid_2[847:840]) ? 1 : 0;
assign detect_max[104][16] = (mid_1[847:840] > mid_2[855:848]) ? 1 : 0;
assign detect_max[104][17] = (mid_1[847:840] > btm_0[839:832]) ? 1 : 0;
assign detect_max[104][18] = (mid_1[847:840] > btm_0[847:840]) ? 1 : 0;
assign detect_max[104][19] = (mid_1[847:840] > btm_0[855:848]) ? 1 : 0;
assign detect_max[104][20] = (mid_1[847:840] > btm_1[839:832]) ? 1 : 0;
assign detect_max[104][21] = (mid_1[847:840] > btm_1[847:840]) ? 1 : 0;
assign detect_max[104][22] = (mid_1[847:840] > btm_1[855:848]) ? 1 : 0;
assign detect_max[104][23] = (mid_1[847:840] > btm_2[839:832]) ? 1 : 0;
assign detect_max[104][24] = (mid_1[847:840] > btm_2[847:840]) ? 1 : 0;
assign detect_max[104][25] = (mid_1[847:840] > btm_2[855:848]) ? 1 : 0;

assign detect_max[105][0] = (mid_1[855:848] > top_0[847:840]) ? 1 : 0;
assign detect_max[105][1] = (mid_1[855:848] > top_0[855:848]) ? 1 : 0;
assign detect_max[105][2] = (mid_1[855:848] > top_0[863:856]) ? 1 : 0;
assign detect_max[105][3] = (mid_1[855:848] > top_1[847:840]) ? 1 : 0;
assign detect_max[105][4] = (mid_1[855:848] > top_1[855:848]) ? 1 : 0;
assign detect_max[105][5] = (mid_1[855:848] > top_1[863:856]) ? 1 : 0;
assign detect_max[105][6] = (mid_1[855:848] > top_2[847:840]) ? 1 : 0;
assign detect_max[105][7] = (mid_1[855:848] > top_2[855:848]) ? 1 : 0;
assign detect_max[105][8] = (mid_1[855:848] > top_2[863:856]) ? 1 : 0;
assign detect_max[105][9] = (mid_1[855:848] > mid_0[847:840]) ? 1 : 0;
assign detect_max[105][10] = (mid_1[855:848] > mid_0[855:848]) ? 1 : 0;
assign detect_max[105][11] = (mid_1[855:848] > mid_0[863:856]) ? 1 : 0;
assign detect_max[105][12] = (mid_1[855:848] > mid_1[847:840]) ? 1 : 0;
assign detect_max[105][13] = (mid_1[855:848] > mid_1[863:856]) ? 1 : 0;
assign detect_max[105][14] = (mid_1[855:848] > mid_2[847:840]) ? 1 : 0;
assign detect_max[105][15] = (mid_1[855:848] > mid_2[855:848]) ? 1 : 0;
assign detect_max[105][16] = (mid_1[855:848] > mid_2[863:856]) ? 1 : 0;
assign detect_max[105][17] = (mid_1[855:848] > btm_0[847:840]) ? 1 : 0;
assign detect_max[105][18] = (mid_1[855:848] > btm_0[855:848]) ? 1 : 0;
assign detect_max[105][19] = (mid_1[855:848] > btm_0[863:856]) ? 1 : 0;
assign detect_max[105][20] = (mid_1[855:848] > btm_1[847:840]) ? 1 : 0;
assign detect_max[105][21] = (mid_1[855:848] > btm_1[855:848]) ? 1 : 0;
assign detect_max[105][22] = (mid_1[855:848] > btm_1[863:856]) ? 1 : 0;
assign detect_max[105][23] = (mid_1[855:848] > btm_2[847:840]) ? 1 : 0;
assign detect_max[105][24] = (mid_1[855:848] > btm_2[855:848]) ? 1 : 0;
assign detect_max[105][25] = (mid_1[855:848] > btm_2[863:856]) ? 1 : 0;

assign detect_max[106][0] = (mid_1[863:856] > top_0[855:848]) ? 1 : 0;
assign detect_max[106][1] = (mid_1[863:856] > top_0[863:856]) ? 1 : 0;
assign detect_max[106][2] = (mid_1[863:856] > top_0[871:864]) ? 1 : 0;
assign detect_max[106][3] = (mid_1[863:856] > top_1[855:848]) ? 1 : 0;
assign detect_max[106][4] = (mid_1[863:856] > top_1[863:856]) ? 1 : 0;
assign detect_max[106][5] = (mid_1[863:856] > top_1[871:864]) ? 1 : 0;
assign detect_max[106][6] = (mid_1[863:856] > top_2[855:848]) ? 1 : 0;
assign detect_max[106][7] = (mid_1[863:856] > top_2[863:856]) ? 1 : 0;
assign detect_max[106][8] = (mid_1[863:856] > top_2[871:864]) ? 1 : 0;
assign detect_max[106][9] = (mid_1[863:856] > mid_0[855:848]) ? 1 : 0;
assign detect_max[106][10] = (mid_1[863:856] > mid_0[863:856]) ? 1 : 0;
assign detect_max[106][11] = (mid_1[863:856] > mid_0[871:864]) ? 1 : 0;
assign detect_max[106][12] = (mid_1[863:856] > mid_1[855:848]) ? 1 : 0;
assign detect_max[106][13] = (mid_1[863:856] > mid_1[871:864]) ? 1 : 0;
assign detect_max[106][14] = (mid_1[863:856] > mid_2[855:848]) ? 1 : 0;
assign detect_max[106][15] = (mid_1[863:856] > mid_2[863:856]) ? 1 : 0;
assign detect_max[106][16] = (mid_1[863:856] > mid_2[871:864]) ? 1 : 0;
assign detect_max[106][17] = (mid_1[863:856] > btm_0[855:848]) ? 1 : 0;
assign detect_max[106][18] = (mid_1[863:856] > btm_0[863:856]) ? 1 : 0;
assign detect_max[106][19] = (mid_1[863:856] > btm_0[871:864]) ? 1 : 0;
assign detect_max[106][20] = (mid_1[863:856] > btm_1[855:848]) ? 1 : 0;
assign detect_max[106][21] = (mid_1[863:856] > btm_1[863:856]) ? 1 : 0;
assign detect_max[106][22] = (mid_1[863:856] > btm_1[871:864]) ? 1 : 0;
assign detect_max[106][23] = (mid_1[863:856] > btm_2[855:848]) ? 1 : 0;
assign detect_max[106][24] = (mid_1[863:856] > btm_2[863:856]) ? 1 : 0;
assign detect_max[106][25] = (mid_1[863:856] > btm_2[871:864]) ? 1 : 0;

assign detect_max[107][0] = (mid_1[871:864] > top_0[863:856]) ? 1 : 0;
assign detect_max[107][1] = (mid_1[871:864] > top_0[871:864]) ? 1 : 0;
assign detect_max[107][2] = (mid_1[871:864] > top_0[879:872]) ? 1 : 0;
assign detect_max[107][3] = (mid_1[871:864] > top_1[863:856]) ? 1 : 0;
assign detect_max[107][4] = (mid_1[871:864] > top_1[871:864]) ? 1 : 0;
assign detect_max[107][5] = (mid_1[871:864] > top_1[879:872]) ? 1 : 0;
assign detect_max[107][6] = (mid_1[871:864] > top_2[863:856]) ? 1 : 0;
assign detect_max[107][7] = (mid_1[871:864] > top_2[871:864]) ? 1 : 0;
assign detect_max[107][8] = (mid_1[871:864] > top_2[879:872]) ? 1 : 0;
assign detect_max[107][9] = (mid_1[871:864] > mid_0[863:856]) ? 1 : 0;
assign detect_max[107][10] = (mid_1[871:864] > mid_0[871:864]) ? 1 : 0;
assign detect_max[107][11] = (mid_1[871:864] > mid_0[879:872]) ? 1 : 0;
assign detect_max[107][12] = (mid_1[871:864] > mid_1[863:856]) ? 1 : 0;
assign detect_max[107][13] = (mid_1[871:864] > mid_1[879:872]) ? 1 : 0;
assign detect_max[107][14] = (mid_1[871:864] > mid_2[863:856]) ? 1 : 0;
assign detect_max[107][15] = (mid_1[871:864] > mid_2[871:864]) ? 1 : 0;
assign detect_max[107][16] = (mid_1[871:864] > mid_2[879:872]) ? 1 : 0;
assign detect_max[107][17] = (mid_1[871:864] > btm_0[863:856]) ? 1 : 0;
assign detect_max[107][18] = (mid_1[871:864] > btm_0[871:864]) ? 1 : 0;
assign detect_max[107][19] = (mid_1[871:864] > btm_0[879:872]) ? 1 : 0;
assign detect_max[107][20] = (mid_1[871:864] > btm_1[863:856]) ? 1 : 0;
assign detect_max[107][21] = (mid_1[871:864] > btm_1[871:864]) ? 1 : 0;
assign detect_max[107][22] = (mid_1[871:864] > btm_1[879:872]) ? 1 : 0;
assign detect_max[107][23] = (mid_1[871:864] > btm_2[863:856]) ? 1 : 0;
assign detect_max[107][24] = (mid_1[871:864] > btm_2[871:864]) ? 1 : 0;
assign detect_max[107][25] = (mid_1[871:864] > btm_2[879:872]) ? 1 : 0;

assign detect_max[108][0] = (mid_1[879:872] > top_0[871:864]) ? 1 : 0;
assign detect_max[108][1] = (mid_1[879:872] > top_0[879:872]) ? 1 : 0;
assign detect_max[108][2] = (mid_1[879:872] > top_0[887:880]) ? 1 : 0;
assign detect_max[108][3] = (mid_1[879:872] > top_1[871:864]) ? 1 : 0;
assign detect_max[108][4] = (mid_1[879:872] > top_1[879:872]) ? 1 : 0;
assign detect_max[108][5] = (mid_1[879:872] > top_1[887:880]) ? 1 : 0;
assign detect_max[108][6] = (mid_1[879:872] > top_2[871:864]) ? 1 : 0;
assign detect_max[108][7] = (mid_1[879:872] > top_2[879:872]) ? 1 : 0;
assign detect_max[108][8] = (mid_1[879:872] > top_2[887:880]) ? 1 : 0;
assign detect_max[108][9] = (mid_1[879:872] > mid_0[871:864]) ? 1 : 0;
assign detect_max[108][10] = (mid_1[879:872] > mid_0[879:872]) ? 1 : 0;
assign detect_max[108][11] = (mid_1[879:872] > mid_0[887:880]) ? 1 : 0;
assign detect_max[108][12] = (mid_1[879:872] > mid_1[871:864]) ? 1 : 0;
assign detect_max[108][13] = (mid_1[879:872] > mid_1[887:880]) ? 1 : 0;
assign detect_max[108][14] = (mid_1[879:872] > mid_2[871:864]) ? 1 : 0;
assign detect_max[108][15] = (mid_1[879:872] > mid_2[879:872]) ? 1 : 0;
assign detect_max[108][16] = (mid_1[879:872] > mid_2[887:880]) ? 1 : 0;
assign detect_max[108][17] = (mid_1[879:872] > btm_0[871:864]) ? 1 : 0;
assign detect_max[108][18] = (mid_1[879:872] > btm_0[879:872]) ? 1 : 0;
assign detect_max[108][19] = (mid_1[879:872] > btm_0[887:880]) ? 1 : 0;
assign detect_max[108][20] = (mid_1[879:872] > btm_1[871:864]) ? 1 : 0;
assign detect_max[108][21] = (mid_1[879:872] > btm_1[879:872]) ? 1 : 0;
assign detect_max[108][22] = (mid_1[879:872] > btm_1[887:880]) ? 1 : 0;
assign detect_max[108][23] = (mid_1[879:872] > btm_2[871:864]) ? 1 : 0;
assign detect_max[108][24] = (mid_1[879:872] > btm_2[879:872]) ? 1 : 0;
assign detect_max[108][25] = (mid_1[879:872] > btm_2[887:880]) ? 1 : 0;

assign detect_max[109][0] = (mid_1[887:880] > top_0[879:872]) ? 1 : 0;
assign detect_max[109][1] = (mid_1[887:880] > top_0[887:880]) ? 1 : 0;
assign detect_max[109][2] = (mid_1[887:880] > top_0[895:888]) ? 1 : 0;
assign detect_max[109][3] = (mid_1[887:880] > top_1[879:872]) ? 1 : 0;
assign detect_max[109][4] = (mid_1[887:880] > top_1[887:880]) ? 1 : 0;
assign detect_max[109][5] = (mid_1[887:880] > top_1[895:888]) ? 1 : 0;
assign detect_max[109][6] = (mid_1[887:880] > top_2[879:872]) ? 1 : 0;
assign detect_max[109][7] = (mid_1[887:880] > top_2[887:880]) ? 1 : 0;
assign detect_max[109][8] = (mid_1[887:880] > top_2[895:888]) ? 1 : 0;
assign detect_max[109][9] = (mid_1[887:880] > mid_0[879:872]) ? 1 : 0;
assign detect_max[109][10] = (mid_1[887:880] > mid_0[887:880]) ? 1 : 0;
assign detect_max[109][11] = (mid_1[887:880] > mid_0[895:888]) ? 1 : 0;
assign detect_max[109][12] = (mid_1[887:880] > mid_1[879:872]) ? 1 : 0;
assign detect_max[109][13] = (mid_1[887:880] > mid_1[895:888]) ? 1 : 0;
assign detect_max[109][14] = (mid_1[887:880] > mid_2[879:872]) ? 1 : 0;
assign detect_max[109][15] = (mid_1[887:880] > mid_2[887:880]) ? 1 : 0;
assign detect_max[109][16] = (mid_1[887:880] > mid_2[895:888]) ? 1 : 0;
assign detect_max[109][17] = (mid_1[887:880] > btm_0[879:872]) ? 1 : 0;
assign detect_max[109][18] = (mid_1[887:880] > btm_0[887:880]) ? 1 : 0;
assign detect_max[109][19] = (mid_1[887:880] > btm_0[895:888]) ? 1 : 0;
assign detect_max[109][20] = (mid_1[887:880] > btm_1[879:872]) ? 1 : 0;
assign detect_max[109][21] = (mid_1[887:880] > btm_1[887:880]) ? 1 : 0;
assign detect_max[109][22] = (mid_1[887:880] > btm_1[895:888]) ? 1 : 0;
assign detect_max[109][23] = (mid_1[887:880] > btm_2[879:872]) ? 1 : 0;
assign detect_max[109][24] = (mid_1[887:880] > btm_2[887:880]) ? 1 : 0;
assign detect_max[109][25] = (mid_1[887:880] > btm_2[895:888]) ? 1 : 0;

assign detect_max[110][0] = (mid_1[895:888] > top_0[887:880]) ? 1 : 0;
assign detect_max[110][1] = (mid_1[895:888] > top_0[895:888]) ? 1 : 0;
assign detect_max[110][2] = (mid_1[895:888] > top_0[903:896]) ? 1 : 0;
assign detect_max[110][3] = (mid_1[895:888] > top_1[887:880]) ? 1 : 0;
assign detect_max[110][4] = (mid_1[895:888] > top_1[895:888]) ? 1 : 0;
assign detect_max[110][5] = (mid_1[895:888] > top_1[903:896]) ? 1 : 0;
assign detect_max[110][6] = (mid_1[895:888] > top_2[887:880]) ? 1 : 0;
assign detect_max[110][7] = (mid_1[895:888] > top_2[895:888]) ? 1 : 0;
assign detect_max[110][8] = (mid_1[895:888] > top_2[903:896]) ? 1 : 0;
assign detect_max[110][9] = (mid_1[895:888] > mid_0[887:880]) ? 1 : 0;
assign detect_max[110][10] = (mid_1[895:888] > mid_0[895:888]) ? 1 : 0;
assign detect_max[110][11] = (mid_1[895:888] > mid_0[903:896]) ? 1 : 0;
assign detect_max[110][12] = (mid_1[895:888] > mid_1[887:880]) ? 1 : 0;
assign detect_max[110][13] = (mid_1[895:888] > mid_1[903:896]) ? 1 : 0;
assign detect_max[110][14] = (mid_1[895:888] > mid_2[887:880]) ? 1 : 0;
assign detect_max[110][15] = (mid_1[895:888] > mid_2[895:888]) ? 1 : 0;
assign detect_max[110][16] = (mid_1[895:888] > mid_2[903:896]) ? 1 : 0;
assign detect_max[110][17] = (mid_1[895:888] > btm_0[887:880]) ? 1 : 0;
assign detect_max[110][18] = (mid_1[895:888] > btm_0[895:888]) ? 1 : 0;
assign detect_max[110][19] = (mid_1[895:888] > btm_0[903:896]) ? 1 : 0;
assign detect_max[110][20] = (mid_1[895:888] > btm_1[887:880]) ? 1 : 0;
assign detect_max[110][21] = (mid_1[895:888] > btm_1[895:888]) ? 1 : 0;
assign detect_max[110][22] = (mid_1[895:888] > btm_1[903:896]) ? 1 : 0;
assign detect_max[110][23] = (mid_1[895:888] > btm_2[887:880]) ? 1 : 0;
assign detect_max[110][24] = (mid_1[895:888] > btm_2[895:888]) ? 1 : 0;
assign detect_max[110][25] = (mid_1[895:888] > btm_2[903:896]) ? 1 : 0;

assign detect_max[111][0] = (mid_1[903:896] > top_0[895:888]) ? 1 : 0;
assign detect_max[111][1] = (mid_1[903:896] > top_0[903:896]) ? 1 : 0;
assign detect_max[111][2] = (mid_1[903:896] > top_0[911:904]) ? 1 : 0;
assign detect_max[111][3] = (mid_1[903:896] > top_1[895:888]) ? 1 : 0;
assign detect_max[111][4] = (mid_1[903:896] > top_1[903:896]) ? 1 : 0;
assign detect_max[111][5] = (mid_1[903:896] > top_1[911:904]) ? 1 : 0;
assign detect_max[111][6] = (mid_1[903:896] > top_2[895:888]) ? 1 : 0;
assign detect_max[111][7] = (mid_1[903:896] > top_2[903:896]) ? 1 : 0;
assign detect_max[111][8] = (mid_1[903:896] > top_2[911:904]) ? 1 : 0;
assign detect_max[111][9] = (mid_1[903:896] > mid_0[895:888]) ? 1 : 0;
assign detect_max[111][10] = (mid_1[903:896] > mid_0[903:896]) ? 1 : 0;
assign detect_max[111][11] = (mid_1[903:896] > mid_0[911:904]) ? 1 : 0;
assign detect_max[111][12] = (mid_1[903:896] > mid_1[895:888]) ? 1 : 0;
assign detect_max[111][13] = (mid_1[903:896] > mid_1[911:904]) ? 1 : 0;
assign detect_max[111][14] = (mid_1[903:896] > mid_2[895:888]) ? 1 : 0;
assign detect_max[111][15] = (mid_1[903:896] > mid_2[903:896]) ? 1 : 0;
assign detect_max[111][16] = (mid_1[903:896] > mid_2[911:904]) ? 1 : 0;
assign detect_max[111][17] = (mid_1[903:896] > btm_0[895:888]) ? 1 : 0;
assign detect_max[111][18] = (mid_1[903:896] > btm_0[903:896]) ? 1 : 0;
assign detect_max[111][19] = (mid_1[903:896] > btm_0[911:904]) ? 1 : 0;
assign detect_max[111][20] = (mid_1[903:896] > btm_1[895:888]) ? 1 : 0;
assign detect_max[111][21] = (mid_1[903:896] > btm_1[903:896]) ? 1 : 0;
assign detect_max[111][22] = (mid_1[903:896] > btm_1[911:904]) ? 1 : 0;
assign detect_max[111][23] = (mid_1[903:896] > btm_2[895:888]) ? 1 : 0;
assign detect_max[111][24] = (mid_1[903:896] > btm_2[903:896]) ? 1 : 0;
assign detect_max[111][25] = (mid_1[903:896] > btm_2[911:904]) ? 1 : 0;

assign detect_max[112][0] = (mid_1[911:904] > top_0[903:896]) ? 1 : 0;
assign detect_max[112][1] = (mid_1[911:904] > top_0[911:904]) ? 1 : 0;
assign detect_max[112][2] = (mid_1[911:904] > top_0[919:912]) ? 1 : 0;
assign detect_max[112][3] = (mid_1[911:904] > top_1[903:896]) ? 1 : 0;
assign detect_max[112][4] = (mid_1[911:904] > top_1[911:904]) ? 1 : 0;
assign detect_max[112][5] = (mid_1[911:904] > top_1[919:912]) ? 1 : 0;
assign detect_max[112][6] = (mid_1[911:904] > top_2[903:896]) ? 1 : 0;
assign detect_max[112][7] = (mid_1[911:904] > top_2[911:904]) ? 1 : 0;
assign detect_max[112][8] = (mid_1[911:904] > top_2[919:912]) ? 1 : 0;
assign detect_max[112][9] = (mid_1[911:904] > mid_0[903:896]) ? 1 : 0;
assign detect_max[112][10] = (mid_1[911:904] > mid_0[911:904]) ? 1 : 0;
assign detect_max[112][11] = (mid_1[911:904] > mid_0[919:912]) ? 1 : 0;
assign detect_max[112][12] = (mid_1[911:904] > mid_1[903:896]) ? 1 : 0;
assign detect_max[112][13] = (mid_1[911:904] > mid_1[919:912]) ? 1 : 0;
assign detect_max[112][14] = (mid_1[911:904] > mid_2[903:896]) ? 1 : 0;
assign detect_max[112][15] = (mid_1[911:904] > mid_2[911:904]) ? 1 : 0;
assign detect_max[112][16] = (mid_1[911:904] > mid_2[919:912]) ? 1 : 0;
assign detect_max[112][17] = (mid_1[911:904] > btm_0[903:896]) ? 1 : 0;
assign detect_max[112][18] = (mid_1[911:904] > btm_0[911:904]) ? 1 : 0;
assign detect_max[112][19] = (mid_1[911:904] > btm_0[919:912]) ? 1 : 0;
assign detect_max[112][20] = (mid_1[911:904] > btm_1[903:896]) ? 1 : 0;
assign detect_max[112][21] = (mid_1[911:904] > btm_1[911:904]) ? 1 : 0;
assign detect_max[112][22] = (mid_1[911:904] > btm_1[919:912]) ? 1 : 0;
assign detect_max[112][23] = (mid_1[911:904] > btm_2[903:896]) ? 1 : 0;
assign detect_max[112][24] = (mid_1[911:904] > btm_2[911:904]) ? 1 : 0;
assign detect_max[112][25] = (mid_1[911:904] > btm_2[919:912]) ? 1 : 0;

assign detect_max[113][0] = (mid_1[919:912] > top_0[911:904]) ? 1 : 0;
assign detect_max[113][1] = (mid_1[919:912] > top_0[919:912]) ? 1 : 0;
assign detect_max[113][2] = (mid_1[919:912] > top_0[927:920]) ? 1 : 0;
assign detect_max[113][3] = (mid_1[919:912] > top_1[911:904]) ? 1 : 0;
assign detect_max[113][4] = (mid_1[919:912] > top_1[919:912]) ? 1 : 0;
assign detect_max[113][5] = (mid_1[919:912] > top_1[927:920]) ? 1 : 0;
assign detect_max[113][6] = (mid_1[919:912] > top_2[911:904]) ? 1 : 0;
assign detect_max[113][7] = (mid_1[919:912] > top_2[919:912]) ? 1 : 0;
assign detect_max[113][8] = (mid_1[919:912] > top_2[927:920]) ? 1 : 0;
assign detect_max[113][9] = (mid_1[919:912] > mid_0[911:904]) ? 1 : 0;
assign detect_max[113][10] = (mid_1[919:912] > mid_0[919:912]) ? 1 : 0;
assign detect_max[113][11] = (mid_1[919:912] > mid_0[927:920]) ? 1 : 0;
assign detect_max[113][12] = (mid_1[919:912] > mid_1[911:904]) ? 1 : 0;
assign detect_max[113][13] = (mid_1[919:912] > mid_1[927:920]) ? 1 : 0;
assign detect_max[113][14] = (mid_1[919:912] > mid_2[911:904]) ? 1 : 0;
assign detect_max[113][15] = (mid_1[919:912] > mid_2[919:912]) ? 1 : 0;
assign detect_max[113][16] = (mid_1[919:912] > mid_2[927:920]) ? 1 : 0;
assign detect_max[113][17] = (mid_1[919:912] > btm_0[911:904]) ? 1 : 0;
assign detect_max[113][18] = (mid_1[919:912] > btm_0[919:912]) ? 1 : 0;
assign detect_max[113][19] = (mid_1[919:912] > btm_0[927:920]) ? 1 : 0;
assign detect_max[113][20] = (mid_1[919:912] > btm_1[911:904]) ? 1 : 0;
assign detect_max[113][21] = (mid_1[919:912] > btm_1[919:912]) ? 1 : 0;
assign detect_max[113][22] = (mid_1[919:912] > btm_1[927:920]) ? 1 : 0;
assign detect_max[113][23] = (mid_1[919:912] > btm_2[911:904]) ? 1 : 0;
assign detect_max[113][24] = (mid_1[919:912] > btm_2[919:912]) ? 1 : 0;
assign detect_max[113][25] = (mid_1[919:912] > btm_2[927:920]) ? 1 : 0;

assign detect_max[114][0] = (mid_1[927:920] > top_0[919:912]) ? 1 : 0;
assign detect_max[114][1] = (mid_1[927:920] > top_0[927:920]) ? 1 : 0;
assign detect_max[114][2] = (mid_1[927:920] > top_0[935:928]) ? 1 : 0;
assign detect_max[114][3] = (mid_1[927:920] > top_1[919:912]) ? 1 : 0;
assign detect_max[114][4] = (mid_1[927:920] > top_1[927:920]) ? 1 : 0;
assign detect_max[114][5] = (mid_1[927:920] > top_1[935:928]) ? 1 : 0;
assign detect_max[114][6] = (mid_1[927:920] > top_2[919:912]) ? 1 : 0;
assign detect_max[114][7] = (mid_1[927:920] > top_2[927:920]) ? 1 : 0;
assign detect_max[114][8] = (mid_1[927:920] > top_2[935:928]) ? 1 : 0;
assign detect_max[114][9] = (mid_1[927:920] > mid_0[919:912]) ? 1 : 0;
assign detect_max[114][10] = (mid_1[927:920] > mid_0[927:920]) ? 1 : 0;
assign detect_max[114][11] = (mid_1[927:920] > mid_0[935:928]) ? 1 : 0;
assign detect_max[114][12] = (mid_1[927:920] > mid_1[919:912]) ? 1 : 0;
assign detect_max[114][13] = (mid_1[927:920] > mid_1[935:928]) ? 1 : 0;
assign detect_max[114][14] = (mid_1[927:920] > mid_2[919:912]) ? 1 : 0;
assign detect_max[114][15] = (mid_1[927:920] > mid_2[927:920]) ? 1 : 0;
assign detect_max[114][16] = (mid_1[927:920] > mid_2[935:928]) ? 1 : 0;
assign detect_max[114][17] = (mid_1[927:920] > btm_0[919:912]) ? 1 : 0;
assign detect_max[114][18] = (mid_1[927:920] > btm_0[927:920]) ? 1 : 0;
assign detect_max[114][19] = (mid_1[927:920] > btm_0[935:928]) ? 1 : 0;
assign detect_max[114][20] = (mid_1[927:920] > btm_1[919:912]) ? 1 : 0;
assign detect_max[114][21] = (mid_1[927:920] > btm_1[927:920]) ? 1 : 0;
assign detect_max[114][22] = (mid_1[927:920] > btm_1[935:928]) ? 1 : 0;
assign detect_max[114][23] = (mid_1[927:920] > btm_2[919:912]) ? 1 : 0;
assign detect_max[114][24] = (mid_1[927:920] > btm_2[927:920]) ? 1 : 0;
assign detect_max[114][25] = (mid_1[927:920] > btm_2[935:928]) ? 1 : 0;

assign detect_max[115][0] = (mid_1[935:928] > top_0[927:920]) ? 1 : 0;
assign detect_max[115][1] = (mid_1[935:928] > top_0[935:928]) ? 1 : 0;
assign detect_max[115][2] = (mid_1[935:928] > top_0[943:936]) ? 1 : 0;
assign detect_max[115][3] = (mid_1[935:928] > top_1[927:920]) ? 1 : 0;
assign detect_max[115][4] = (mid_1[935:928] > top_1[935:928]) ? 1 : 0;
assign detect_max[115][5] = (mid_1[935:928] > top_1[943:936]) ? 1 : 0;
assign detect_max[115][6] = (mid_1[935:928] > top_2[927:920]) ? 1 : 0;
assign detect_max[115][7] = (mid_1[935:928] > top_2[935:928]) ? 1 : 0;
assign detect_max[115][8] = (mid_1[935:928] > top_2[943:936]) ? 1 : 0;
assign detect_max[115][9] = (mid_1[935:928] > mid_0[927:920]) ? 1 : 0;
assign detect_max[115][10] = (mid_1[935:928] > mid_0[935:928]) ? 1 : 0;
assign detect_max[115][11] = (mid_1[935:928] > mid_0[943:936]) ? 1 : 0;
assign detect_max[115][12] = (mid_1[935:928] > mid_1[927:920]) ? 1 : 0;
assign detect_max[115][13] = (mid_1[935:928] > mid_1[943:936]) ? 1 : 0;
assign detect_max[115][14] = (mid_1[935:928] > mid_2[927:920]) ? 1 : 0;
assign detect_max[115][15] = (mid_1[935:928] > mid_2[935:928]) ? 1 : 0;
assign detect_max[115][16] = (mid_1[935:928] > mid_2[943:936]) ? 1 : 0;
assign detect_max[115][17] = (mid_1[935:928] > btm_0[927:920]) ? 1 : 0;
assign detect_max[115][18] = (mid_1[935:928] > btm_0[935:928]) ? 1 : 0;
assign detect_max[115][19] = (mid_1[935:928] > btm_0[943:936]) ? 1 : 0;
assign detect_max[115][20] = (mid_1[935:928] > btm_1[927:920]) ? 1 : 0;
assign detect_max[115][21] = (mid_1[935:928] > btm_1[935:928]) ? 1 : 0;
assign detect_max[115][22] = (mid_1[935:928] > btm_1[943:936]) ? 1 : 0;
assign detect_max[115][23] = (mid_1[935:928] > btm_2[927:920]) ? 1 : 0;
assign detect_max[115][24] = (mid_1[935:928] > btm_2[935:928]) ? 1 : 0;
assign detect_max[115][25] = (mid_1[935:928] > btm_2[943:936]) ? 1 : 0;

assign detect_max[116][0] = (mid_1[943:936] > top_0[935:928]) ? 1 : 0;
assign detect_max[116][1] = (mid_1[943:936] > top_0[943:936]) ? 1 : 0;
assign detect_max[116][2] = (mid_1[943:936] > top_0[951:944]) ? 1 : 0;
assign detect_max[116][3] = (mid_1[943:936] > top_1[935:928]) ? 1 : 0;
assign detect_max[116][4] = (mid_1[943:936] > top_1[943:936]) ? 1 : 0;
assign detect_max[116][5] = (mid_1[943:936] > top_1[951:944]) ? 1 : 0;
assign detect_max[116][6] = (mid_1[943:936] > top_2[935:928]) ? 1 : 0;
assign detect_max[116][7] = (mid_1[943:936] > top_2[943:936]) ? 1 : 0;
assign detect_max[116][8] = (mid_1[943:936] > top_2[951:944]) ? 1 : 0;
assign detect_max[116][9] = (mid_1[943:936] > mid_0[935:928]) ? 1 : 0;
assign detect_max[116][10] = (mid_1[943:936] > mid_0[943:936]) ? 1 : 0;
assign detect_max[116][11] = (mid_1[943:936] > mid_0[951:944]) ? 1 : 0;
assign detect_max[116][12] = (mid_1[943:936] > mid_1[935:928]) ? 1 : 0;
assign detect_max[116][13] = (mid_1[943:936] > mid_1[951:944]) ? 1 : 0;
assign detect_max[116][14] = (mid_1[943:936] > mid_2[935:928]) ? 1 : 0;
assign detect_max[116][15] = (mid_1[943:936] > mid_2[943:936]) ? 1 : 0;
assign detect_max[116][16] = (mid_1[943:936] > mid_2[951:944]) ? 1 : 0;
assign detect_max[116][17] = (mid_1[943:936] > btm_0[935:928]) ? 1 : 0;
assign detect_max[116][18] = (mid_1[943:936] > btm_0[943:936]) ? 1 : 0;
assign detect_max[116][19] = (mid_1[943:936] > btm_0[951:944]) ? 1 : 0;
assign detect_max[116][20] = (mid_1[943:936] > btm_1[935:928]) ? 1 : 0;
assign detect_max[116][21] = (mid_1[943:936] > btm_1[943:936]) ? 1 : 0;
assign detect_max[116][22] = (mid_1[943:936] > btm_1[951:944]) ? 1 : 0;
assign detect_max[116][23] = (mid_1[943:936] > btm_2[935:928]) ? 1 : 0;
assign detect_max[116][24] = (mid_1[943:936] > btm_2[943:936]) ? 1 : 0;
assign detect_max[116][25] = (mid_1[943:936] > btm_2[951:944]) ? 1 : 0;

assign detect_max[117][0] = (mid_1[951:944] > top_0[943:936]) ? 1 : 0;
assign detect_max[117][1] = (mid_1[951:944] > top_0[951:944]) ? 1 : 0;
assign detect_max[117][2] = (mid_1[951:944] > top_0[959:952]) ? 1 : 0;
assign detect_max[117][3] = (mid_1[951:944] > top_1[943:936]) ? 1 : 0;
assign detect_max[117][4] = (mid_1[951:944] > top_1[951:944]) ? 1 : 0;
assign detect_max[117][5] = (mid_1[951:944] > top_1[959:952]) ? 1 : 0;
assign detect_max[117][6] = (mid_1[951:944] > top_2[943:936]) ? 1 : 0;
assign detect_max[117][7] = (mid_1[951:944] > top_2[951:944]) ? 1 : 0;
assign detect_max[117][8] = (mid_1[951:944] > top_2[959:952]) ? 1 : 0;
assign detect_max[117][9] = (mid_1[951:944] > mid_0[943:936]) ? 1 : 0;
assign detect_max[117][10] = (mid_1[951:944] > mid_0[951:944]) ? 1 : 0;
assign detect_max[117][11] = (mid_1[951:944] > mid_0[959:952]) ? 1 : 0;
assign detect_max[117][12] = (mid_1[951:944] > mid_1[943:936]) ? 1 : 0;
assign detect_max[117][13] = (mid_1[951:944] > mid_1[959:952]) ? 1 : 0;
assign detect_max[117][14] = (mid_1[951:944] > mid_2[943:936]) ? 1 : 0;
assign detect_max[117][15] = (mid_1[951:944] > mid_2[951:944]) ? 1 : 0;
assign detect_max[117][16] = (mid_1[951:944] > mid_2[959:952]) ? 1 : 0;
assign detect_max[117][17] = (mid_1[951:944] > btm_0[943:936]) ? 1 : 0;
assign detect_max[117][18] = (mid_1[951:944] > btm_0[951:944]) ? 1 : 0;
assign detect_max[117][19] = (mid_1[951:944] > btm_0[959:952]) ? 1 : 0;
assign detect_max[117][20] = (mid_1[951:944] > btm_1[943:936]) ? 1 : 0;
assign detect_max[117][21] = (mid_1[951:944] > btm_1[951:944]) ? 1 : 0;
assign detect_max[117][22] = (mid_1[951:944] > btm_1[959:952]) ? 1 : 0;
assign detect_max[117][23] = (mid_1[951:944] > btm_2[943:936]) ? 1 : 0;
assign detect_max[117][24] = (mid_1[951:944] > btm_2[951:944]) ? 1 : 0;
assign detect_max[117][25] = (mid_1[951:944] > btm_2[959:952]) ? 1 : 0;

assign detect_max[118][0] = (mid_1[959:952] > top_0[951:944]) ? 1 : 0;
assign detect_max[118][1] = (mid_1[959:952] > top_0[959:952]) ? 1 : 0;
assign detect_max[118][2] = (mid_1[959:952] > top_0[967:960]) ? 1 : 0;
assign detect_max[118][3] = (mid_1[959:952] > top_1[951:944]) ? 1 : 0;
assign detect_max[118][4] = (mid_1[959:952] > top_1[959:952]) ? 1 : 0;
assign detect_max[118][5] = (mid_1[959:952] > top_1[967:960]) ? 1 : 0;
assign detect_max[118][6] = (mid_1[959:952] > top_2[951:944]) ? 1 : 0;
assign detect_max[118][7] = (mid_1[959:952] > top_2[959:952]) ? 1 : 0;
assign detect_max[118][8] = (mid_1[959:952] > top_2[967:960]) ? 1 : 0;
assign detect_max[118][9] = (mid_1[959:952] > mid_0[951:944]) ? 1 : 0;
assign detect_max[118][10] = (mid_1[959:952] > mid_0[959:952]) ? 1 : 0;
assign detect_max[118][11] = (mid_1[959:952] > mid_0[967:960]) ? 1 : 0;
assign detect_max[118][12] = (mid_1[959:952] > mid_1[951:944]) ? 1 : 0;
assign detect_max[118][13] = (mid_1[959:952] > mid_1[967:960]) ? 1 : 0;
assign detect_max[118][14] = (mid_1[959:952] > mid_2[951:944]) ? 1 : 0;
assign detect_max[118][15] = (mid_1[959:952] > mid_2[959:952]) ? 1 : 0;
assign detect_max[118][16] = (mid_1[959:952] > mid_2[967:960]) ? 1 : 0;
assign detect_max[118][17] = (mid_1[959:952] > btm_0[951:944]) ? 1 : 0;
assign detect_max[118][18] = (mid_1[959:952] > btm_0[959:952]) ? 1 : 0;
assign detect_max[118][19] = (mid_1[959:952] > btm_0[967:960]) ? 1 : 0;
assign detect_max[118][20] = (mid_1[959:952] > btm_1[951:944]) ? 1 : 0;
assign detect_max[118][21] = (mid_1[959:952] > btm_1[959:952]) ? 1 : 0;
assign detect_max[118][22] = (mid_1[959:952] > btm_1[967:960]) ? 1 : 0;
assign detect_max[118][23] = (mid_1[959:952] > btm_2[951:944]) ? 1 : 0;
assign detect_max[118][24] = (mid_1[959:952] > btm_2[959:952]) ? 1 : 0;
assign detect_max[118][25] = (mid_1[959:952] > btm_2[967:960]) ? 1 : 0;

assign detect_max[119][0] = (mid_1[967:960] > top_0[959:952]) ? 1 : 0;
assign detect_max[119][1] = (mid_1[967:960] > top_0[967:960]) ? 1 : 0;
assign detect_max[119][2] = (mid_1[967:960] > top_0[975:968]) ? 1 : 0;
assign detect_max[119][3] = (mid_1[967:960] > top_1[959:952]) ? 1 : 0;
assign detect_max[119][4] = (mid_1[967:960] > top_1[967:960]) ? 1 : 0;
assign detect_max[119][5] = (mid_1[967:960] > top_1[975:968]) ? 1 : 0;
assign detect_max[119][6] = (mid_1[967:960] > top_2[959:952]) ? 1 : 0;
assign detect_max[119][7] = (mid_1[967:960] > top_2[967:960]) ? 1 : 0;
assign detect_max[119][8] = (mid_1[967:960] > top_2[975:968]) ? 1 : 0;
assign detect_max[119][9] = (mid_1[967:960] > mid_0[959:952]) ? 1 : 0;
assign detect_max[119][10] = (mid_1[967:960] > mid_0[967:960]) ? 1 : 0;
assign detect_max[119][11] = (mid_1[967:960] > mid_0[975:968]) ? 1 : 0;
assign detect_max[119][12] = (mid_1[967:960] > mid_1[959:952]) ? 1 : 0;
assign detect_max[119][13] = (mid_1[967:960] > mid_1[975:968]) ? 1 : 0;
assign detect_max[119][14] = (mid_1[967:960] > mid_2[959:952]) ? 1 : 0;
assign detect_max[119][15] = (mid_1[967:960] > mid_2[967:960]) ? 1 : 0;
assign detect_max[119][16] = (mid_1[967:960] > mid_2[975:968]) ? 1 : 0;
assign detect_max[119][17] = (mid_1[967:960] > btm_0[959:952]) ? 1 : 0;
assign detect_max[119][18] = (mid_1[967:960] > btm_0[967:960]) ? 1 : 0;
assign detect_max[119][19] = (mid_1[967:960] > btm_0[975:968]) ? 1 : 0;
assign detect_max[119][20] = (mid_1[967:960] > btm_1[959:952]) ? 1 : 0;
assign detect_max[119][21] = (mid_1[967:960] > btm_1[967:960]) ? 1 : 0;
assign detect_max[119][22] = (mid_1[967:960] > btm_1[975:968]) ? 1 : 0;
assign detect_max[119][23] = (mid_1[967:960] > btm_2[959:952]) ? 1 : 0;
assign detect_max[119][24] = (mid_1[967:960] > btm_2[967:960]) ? 1 : 0;
assign detect_max[119][25] = (mid_1[967:960] > btm_2[975:968]) ? 1 : 0;

assign detect_max[120][0] = (mid_1[975:968] > top_0[967:960]) ? 1 : 0;
assign detect_max[120][1] = (mid_1[975:968] > top_0[975:968]) ? 1 : 0;
assign detect_max[120][2] = (mid_1[975:968] > top_0[983:976]) ? 1 : 0;
assign detect_max[120][3] = (mid_1[975:968] > top_1[967:960]) ? 1 : 0;
assign detect_max[120][4] = (mid_1[975:968] > top_1[975:968]) ? 1 : 0;
assign detect_max[120][5] = (mid_1[975:968] > top_1[983:976]) ? 1 : 0;
assign detect_max[120][6] = (mid_1[975:968] > top_2[967:960]) ? 1 : 0;
assign detect_max[120][7] = (mid_1[975:968] > top_2[975:968]) ? 1 : 0;
assign detect_max[120][8] = (mid_1[975:968] > top_2[983:976]) ? 1 : 0;
assign detect_max[120][9] = (mid_1[975:968] > mid_0[967:960]) ? 1 : 0;
assign detect_max[120][10] = (mid_1[975:968] > mid_0[975:968]) ? 1 : 0;
assign detect_max[120][11] = (mid_1[975:968] > mid_0[983:976]) ? 1 : 0;
assign detect_max[120][12] = (mid_1[975:968] > mid_1[967:960]) ? 1 : 0;
assign detect_max[120][13] = (mid_1[975:968] > mid_1[983:976]) ? 1 : 0;
assign detect_max[120][14] = (mid_1[975:968] > mid_2[967:960]) ? 1 : 0;
assign detect_max[120][15] = (mid_1[975:968] > mid_2[975:968]) ? 1 : 0;
assign detect_max[120][16] = (mid_1[975:968] > mid_2[983:976]) ? 1 : 0;
assign detect_max[120][17] = (mid_1[975:968] > btm_0[967:960]) ? 1 : 0;
assign detect_max[120][18] = (mid_1[975:968] > btm_0[975:968]) ? 1 : 0;
assign detect_max[120][19] = (mid_1[975:968] > btm_0[983:976]) ? 1 : 0;
assign detect_max[120][20] = (mid_1[975:968] > btm_1[967:960]) ? 1 : 0;
assign detect_max[120][21] = (mid_1[975:968] > btm_1[975:968]) ? 1 : 0;
assign detect_max[120][22] = (mid_1[975:968] > btm_1[983:976]) ? 1 : 0;
assign detect_max[120][23] = (mid_1[975:968] > btm_2[967:960]) ? 1 : 0;
assign detect_max[120][24] = (mid_1[975:968] > btm_2[975:968]) ? 1 : 0;
assign detect_max[120][25] = (mid_1[975:968] > btm_2[983:976]) ? 1 : 0;

assign detect_max[121][0] = (mid_1[983:976] > top_0[975:968]) ? 1 : 0;
assign detect_max[121][1] = (mid_1[983:976] > top_0[983:976]) ? 1 : 0;
assign detect_max[121][2] = (mid_1[983:976] > top_0[991:984]) ? 1 : 0;
assign detect_max[121][3] = (mid_1[983:976] > top_1[975:968]) ? 1 : 0;
assign detect_max[121][4] = (mid_1[983:976] > top_1[983:976]) ? 1 : 0;
assign detect_max[121][5] = (mid_1[983:976] > top_1[991:984]) ? 1 : 0;
assign detect_max[121][6] = (mid_1[983:976] > top_2[975:968]) ? 1 : 0;
assign detect_max[121][7] = (mid_1[983:976] > top_2[983:976]) ? 1 : 0;
assign detect_max[121][8] = (mid_1[983:976] > top_2[991:984]) ? 1 : 0;
assign detect_max[121][9] = (mid_1[983:976] > mid_0[975:968]) ? 1 : 0;
assign detect_max[121][10] = (mid_1[983:976] > mid_0[983:976]) ? 1 : 0;
assign detect_max[121][11] = (mid_1[983:976] > mid_0[991:984]) ? 1 : 0;
assign detect_max[121][12] = (mid_1[983:976] > mid_1[975:968]) ? 1 : 0;
assign detect_max[121][13] = (mid_1[983:976] > mid_1[991:984]) ? 1 : 0;
assign detect_max[121][14] = (mid_1[983:976] > mid_2[975:968]) ? 1 : 0;
assign detect_max[121][15] = (mid_1[983:976] > mid_2[983:976]) ? 1 : 0;
assign detect_max[121][16] = (mid_1[983:976] > mid_2[991:984]) ? 1 : 0;
assign detect_max[121][17] = (mid_1[983:976] > btm_0[975:968]) ? 1 : 0;
assign detect_max[121][18] = (mid_1[983:976] > btm_0[983:976]) ? 1 : 0;
assign detect_max[121][19] = (mid_1[983:976] > btm_0[991:984]) ? 1 : 0;
assign detect_max[121][20] = (mid_1[983:976] > btm_1[975:968]) ? 1 : 0;
assign detect_max[121][21] = (mid_1[983:976] > btm_1[983:976]) ? 1 : 0;
assign detect_max[121][22] = (mid_1[983:976] > btm_1[991:984]) ? 1 : 0;
assign detect_max[121][23] = (mid_1[983:976] > btm_2[975:968]) ? 1 : 0;
assign detect_max[121][24] = (mid_1[983:976] > btm_2[983:976]) ? 1 : 0;
assign detect_max[121][25] = (mid_1[983:976] > btm_2[991:984]) ? 1 : 0;

assign detect_max[122][0] = (mid_1[991:984] > top_0[983:976]) ? 1 : 0;
assign detect_max[122][1] = (mid_1[991:984] > top_0[991:984]) ? 1 : 0;
assign detect_max[122][2] = (mid_1[991:984] > top_0[999:992]) ? 1 : 0;
assign detect_max[122][3] = (mid_1[991:984] > top_1[983:976]) ? 1 : 0;
assign detect_max[122][4] = (mid_1[991:984] > top_1[991:984]) ? 1 : 0;
assign detect_max[122][5] = (mid_1[991:984] > top_1[999:992]) ? 1 : 0;
assign detect_max[122][6] = (mid_1[991:984] > top_2[983:976]) ? 1 : 0;
assign detect_max[122][7] = (mid_1[991:984] > top_2[991:984]) ? 1 : 0;
assign detect_max[122][8] = (mid_1[991:984] > top_2[999:992]) ? 1 : 0;
assign detect_max[122][9] = (mid_1[991:984] > mid_0[983:976]) ? 1 : 0;
assign detect_max[122][10] = (mid_1[991:984] > mid_0[991:984]) ? 1 : 0;
assign detect_max[122][11] = (mid_1[991:984] > mid_0[999:992]) ? 1 : 0;
assign detect_max[122][12] = (mid_1[991:984] > mid_1[983:976]) ? 1 : 0;
assign detect_max[122][13] = (mid_1[991:984] > mid_1[999:992]) ? 1 : 0;
assign detect_max[122][14] = (mid_1[991:984] > mid_2[983:976]) ? 1 : 0;
assign detect_max[122][15] = (mid_1[991:984] > mid_2[991:984]) ? 1 : 0;
assign detect_max[122][16] = (mid_1[991:984] > mid_2[999:992]) ? 1 : 0;
assign detect_max[122][17] = (mid_1[991:984] > btm_0[983:976]) ? 1 : 0;
assign detect_max[122][18] = (mid_1[991:984] > btm_0[991:984]) ? 1 : 0;
assign detect_max[122][19] = (mid_1[991:984] > btm_0[999:992]) ? 1 : 0;
assign detect_max[122][20] = (mid_1[991:984] > btm_1[983:976]) ? 1 : 0;
assign detect_max[122][21] = (mid_1[991:984] > btm_1[991:984]) ? 1 : 0;
assign detect_max[122][22] = (mid_1[991:984] > btm_1[999:992]) ? 1 : 0;
assign detect_max[122][23] = (mid_1[991:984] > btm_2[983:976]) ? 1 : 0;
assign detect_max[122][24] = (mid_1[991:984] > btm_2[991:984]) ? 1 : 0;
assign detect_max[122][25] = (mid_1[991:984] > btm_2[999:992]) ? 1 : 0;

assign detect_max[123][0] = (mid_1[999:992] > top_0[991:984]) ? 1 : 0;
assign detect_max[123][1] = (mid_1[999:992] > top_0[999:992]) ? 1 : 0;
assign detect_max[123][2] = (mid_1[999:992] > top_0[1007:1000]) ? 1 : 0;
assign detect_max[123][3] = (mid_1[999:992] > top_1[991:984]) ? 1 : 0;
assign detect_max[123][4] = (mid_1[999:992] > top_1[999:992]) ? 1 : 0;
assign detect_max[123][5] = (mid_1[999:992] > top_1[1007:1000]) ? 1 : 0;
assign detect_max[123][6] = (mid_1[999:992] > top_2[991:984]) ? 1 : 0;
assign detect_max[123][7] = (mid_1[999:992] > top_2[999:992]) ? 1 : 0;
assign detect_max[123][8] = (mid_1[999:992] > top_2[1007:1000]) ? 1 : 0;
assign detect_max[123][9] = (mid_1[999:992] > mid_0[991:984]) ? 1 : 0;
assign detect_max[123][10] = (mid_1[999:992] > mid_0[999:992]) ? 1 : 0;
assign detect_max[123][11] = (mid_1[999:992] > mid_0[1007:1000]) ? 1 : 0;
assign detect_max[123][12] = (mid_1[999:992] > mid_1[991:984]) ? 1 : 0;
assign detect_max[123][13] = (mid_1[999:992] > mid_1[1007:1000]) ? 1 : 0;
assign detect_max[123][14] = (mid_1[999:992] > mid_2[991:984]) ? 1 : 0;
assign detect_max[123][15] = (mid_1[999:992] > mid_2[999:992]) ? 1 : 0;
assign detect_max[123][16] = (mid_1[999:992] > mid_2[1007:1000]) ? 1 : 0;
assign detect_max[123][17] = (mid_1[999:992] > btm_0[991:984]) ? 1 : 0;
assign detect_max[123][18] = (mid_1[999:992] > btm_0[999:992]) ? 1 : 0;
assign detect_max[123][19] = (mid_1[999:992] > btm_0[1007:1000]) ? 1 : 0;
assign detect_max[123][20] = (mid_1[999:992] > btm_1[991:984]) ? 1 : 0;
assign detect_max[123][21] = (mid_1[999:992] > btm_1[999:992]) ? 1 : 0;
assign detect_max[123][22] = (mid_1[999:992] > btm_1[1007:1000]) ? 1 : 0;
assign detect_max[123][23] = (mid_1[999:992] > btm_2[991:984]) ? 1 : 0;
assign detect_max[123][24] = (mid_1[999:992] > btm_2[999:992]) ? 1 : 0;
assign detect_max[123][25] = (mid_1[999:992] > btm_2[1007:1000]) ? 1 : 0;

assign detect_max[124][0] = (mid_1[1007:1000] > top_0[999:992]) ? 1 : 0;
assign detect_max[124][1] = (mid_1[1007:1000] > top_0[1007:1000]) ? 1 : 0;
assign detect_max[124][2] = (mid_1[1007:1000] > top_0[1015:1008]) ? 1 : 0;
assign detect_max[124][3] = (mid_1[1007:1000] > top_1[999:992]) ? 1 : 0;
assign detect_max[124][4] = (mid_1[1007:1000] > top_1[1007:1000]) ? 1 : 0;
assign detect_max[124][5] = (mid_1[1007:1000] > top_1[1015:1008]) ? 1 : 0;
assign detect_max[124][6] = (mid_1[1007:1000] > top_2[999:992]) ? 1 : 0;
assign detect_max[124][7] = (mid_1[1007:1000] > top_2[1007:1000]) ? 1 : 0;
assign detect_max[124][8] = (mid_1[1007:1000] > top_2[1015:1008]) ? 1 : 0;
assign detect_max[124][9] = (mid_1[1007:1000] > mid_0[999:992]) ? 1 : 0;
assign detect_max[124][10] = (mid_1[1007:1000] > mid_0[1007:1000]) ? 1 : 0;
assign detect_max[124][11] = (mid_1[1007:1000] > mid_0[1015:1008]) ? 1 : 0;
assign detect_max[124][12] = (mid_1[1007:1000] > mid_1[999:992]) ? 1 : 0;
assign detect_max[124][13] = (mid_1[1007:1000] > mid_1[1015:1008]) ? 1 : 0;
assign detect_max[124][14] = (mid_1[1007:1000] > mid_2[999:992]) ? 1 : 0;
assign detect_max[124][15] = (mid_1[1007:1000] > mid_2[1007:1000]) ? 1 : 0;
assign detect_max[124][16] = (mid_1[1007:1000] > mid_2[1015:1008]) ? 1 : 0;
assign detect_max[124][17] = (mid_1[1007:1000] > btm_0[999:992]) ? 1 : 0;
assign detect_max[124][18] = (mid_1[1007:1000] > btm_0[1007:1000]) ? 1 : 0;
assign detect_max[124][19] = (mid_1[1007:1000] > btm_0[1015:1008]) ? 1 : 0;
assign detect_max[124][20] = (mid_1[1007:1000] > btm_1[999:992]) ? 1 : 0;
assign detect_max[124][21] = (mid_1[1007:1000] > btm_1[1007:1000]) ? 1 : 0;
assign detect_max[124][22] = (mid_1[1007:1000] > btm_1[1015:1008]) ? 1 : 0;
assign detect_max[124][23] = (mid_1[1007:1000] > btm_2[999:992]) ? 1 : 0;
assign detect_max[124][24] = (mid_1[1007:1000] > btm_2[1007:1000]) ? 1 : 0;
assign detect_max[124][25] = (mid_1[1007:1000] > btm_2[1015:1008]) ? 1 : 0;

assign detect_max[125][0] = (mid_1[1015:1008] > top_0[1007:1000]) ? 1 : 0;
assign detect_max[125][1] = (mid_1[1015:1008] > top_0[1015:1008]) ? 1 : 0;
assign detect_max[125][2] = (mid_1[1015:1008] > top_0[1023:1016]) ? 1 : 0;
assign detect_max[125][3] = (mid_1[1015:1008] > top_1[1007:1000]) ? 1 : 0;
assign detect_max[125][4] = (mid_1[1015:1008] > top_1[1015:1008]) ? 1 : 0;
assign detect_max[125][5] = (mid_1[1015:1008] > top_1[1023:1016]) ? 1 : 0;
assign detect_max[125][6] = (mid_1[1015:1008] > top_2[1007:1000]) ? 1 : 0;
assign detect_max[125][7] = (mid_1[1015:1008] > top_2[1015:1008]) ? 1 : 0;
assign detect_max[125][8] = (mid_1[1015:1008] > top_2[1023:1016]) ? 1 : 0;
assign detect_max[125][9] = (mid_1[1015:1008] > mid_0[1007:1000]) ? 1 : 0;
assign detect_max[125][10] = (mid_1[1015:1008] > mid_0[1015:1008]) ? 1 : 0;
assign detect_max[125][11] = (mid_1[1015:1008] > mid_0[1023:1016]) ? 1 : 0;
assign detect_max[125][12] = (mid_1[1015:1008] > mid_1[1007:1000]) ? 1 : 0;
assign detect_max[125][13] = (mid_1[1015:1008] > mid_1[1023:1016]) ? 1 : 0;
assign detect_max[125][14] = (mid_1[1015:1008] > mid_2[1007:1000]) ? 1 : 0;
assign detect_max[125][15] = (mid_1[1015:1008] > mid_2[1015:1008]) ? 1 : 0;
assign detect_max[125][16] = (mid_1[1015:1008] > mid_2[1023:1016]) ? 1 : 0;
assign detect_max[125][17] = (mid_1[1015:1008] > btm_0[1007:1000]) ? 1 : 0;
assign detect_max[125][18] = (mid_1[1015:1008] > btm_0[1015:1008]) ? 1 : 0;
assign detect_max[125][19] = (mid_1[1015:1008] > btm_0[1023:1016]) ? 1 : 0;
assign detect_max[125][20] = (mid_1[1015:1008] > btm_1[1007:1000]) ? 1 : 0;
assign detect_max[125][21] = (mid_1[1015:1008] > btm_1[1015:1008]) ? 1 : 0;
assign detect_max[125][22] = (mid_1[1015:1008] > btm_1[1023:1016]) ? 1 : 0;
assign detect_max[125][23] = (mid_1[1015:1008] > btm_2[1007:1000]) ? 1 : 0;
assign detect_max[125][24] = (mid_1[1015:1008] > btm_2[1015:1008]) ? 1 : 0;
assign detect_max[125][25] = (mid_1[1015:1008] > btm_2[1023:1016]) ? 1 : 0;

assign detect_max[126][0] = (mid_1[1023:1016] > top_0[1015:1008]) ? 1 : 0;
assign detect_max[126][1] = (mid_1[1023:1016] > top_0[1023:1016]) ? 1 : 0;
assign detect_max[126][2] = (mid_1[1023:1016] > top_0[1031:1024]) ? 1 : 0;
assign detect_max[126][3] = (mid_1[1023:1016] > top_1[1015:1008]) ? 1 : 0;
assign detect_max[126][4] = (mid_1[1023:1016] > top_1[1023:1016]) ? 1 : 0;
assign detect_max[126][5] = (mid_1[1023:1016] > top_1[1031:1024]) ? 1 : 0;
assign detect_max[126][6] = (mid_1[1023:1016] > top_2[1015:1008]) ? 1 : 0;
assign detect_max[126][7] = (mid_1[1023:1016] > top_2[1023:1016]) ? 1 : 0;
assign detect_max[126][8] = (mid_1[1023:1016] > top_2[1031:1024]) ? 1 : 0;
assign detect_max[126][9] = (mid_1[1023:1016] > mid_0[1015:1008]) ? 1 : 0;
assign detect_max[126][10] = (mid_1[1023:1016] > mid_0[1023:1016]) ? 1 : 0;
assign detect_max[126][11] = (mid_1[1023:1016] > mid_0[1031:1024]) ? 1 : 0;
assign detect_max[126][12] = (mid_1[1023:1016] > mid_1[1015:1008]) ? 1 : 0;
assign detect_max[126][13] = (mid_1[1023:1016] > mid_1[1031:1024]) ? 1 : 0;
assign detect_max[126][14] = (mid_1[1023:1016] > mid_2[1015:1008]) ? 1 : 0;
assign detect_max[126][15] = (mid_1[1023:1016] > mid_2[1023:1016]) ? 1 : 0;
assign detect_max[126][16] = (mid_1[1023:1016] > mid_2[1031:1024]) ? 1 : 0;
assign detect_max[126][17] = (mid_1[1023:1016] > btm_0[1015:1008]) ? 1 : 0;
assign detect_max[126][18] = (mid_1[1023:1016] > btm_0[1023:1016]) ? 1 : 0;
assign detect_max[126][19] = (mid_1[1023:1016] > btm_0[1031:1024]) ? 1 : 0;
assign detect_max[126][20] = (mid_1[1023:1016] > btm_1[1015:1008]) ? 1 : 0;
assign detect_max[126][21] = (mid_1[1023:1016] > btm_1[1023:1016]) ? 1 : 0;
assign detect_max[126][22] = (mid_1[1023:1016] > btm_1[1031:1024]) ? 1 : 0;
assign detect_max[126][23] = (mid_1[1023:1016] > btm_2[1015:1008]) ? 1 : 0;
assign detect_max[126][24] = (mid_1[1023:1016] > btm_2[1023:1016]) ? 1 : 0;
assign detect_max[126][25] = (mid_1[1023:1016] > btm_2[1031:1024]) ? 1 : 0;

assign detect_max[127][0] = (mid_1[1031:1024] > top_0[1023:1016]) ? 1 : 0;
assign detect_max[127][1] = (mid_1[1031:1024] > top_0[1031:1024]) ? 1 : 0;
assign detect_max[127][2] = (mid_1[1031:1024] > top_0[1039:1032]) ? 1 : 0;
assign detect_max[127][3] = (mid_1[1031:1024] > top_1[1023:1016]) ? 1 : 0;
assign detect_max[127][4] = (mid_1[1031:1024] > top_1[1031:1024]) ? 1 : 0;
assign detect_max[127][5] = (mid_1[1031:1024] > top_1[1039:1032]) ? 1 : 0;
assign detect_max[127][6] = (mid_1[1031:1024] > top_2[1023:1016]) ? 1 : 0;
assign detect_max[127][7] = (mid_1[1031:1024] > top_2[1031:1024]) ? 1 : 0;
assign detect_max[127][8] = (mid_1[1031:1024] > top_2[1039:1032]) ? 1 : 0;
assign detect_max[127][9] = (mid_1[1031:1024] > mid_0[1023:1016]) ? 1 : 0;
assign detect_max[127][10] = (mid_1[1031:1024] > mid_0[1031:1024]) ? 1 : 0;
assign detect_max[127][11] = (mid_1[1031:1024] > mid_0[1039:1032]) ? 1 : 0;
assign detect_max[127][12] = (mid_1[1031:1024] > mid_1[1023:1016]) ? 1 : 0;
assign detect_max[127][13] = (mid_1[1031:1024] > mid_1[1039:1032]) ? 1 : 0;
assign detect_max[127][14] = (mid_1[1031:1024] > mid_2[1023:1016]) ? 1 : 0;
assign detect_max[127][15] = (mid_1[1031:1024] > mid_2[1031:1024]) ? 1 : 0;
assign detect_max[127][16] = (mid_1[1031:1024] > mid_2[1039:1032]) ? 1 : 0;
assign detect_max[127][17] = (mid_1[1031:1024] > btm_0[1023:1016]) ? 1 : 0;
assign detect_max[127][18] = (mid_1[1031:1024] > btm_0[1031:1024]) ? 1 : 0;
assign detect_max[127][19] = (mid_1[1031:1024] > btm_0[1039:1032]) ? 1 : 0;
assign detect_max[127][20] = (mid_1[1031:1024] > btm_1[1023:1016]) ? 1 : 0;
assign detect_max[127][21] = (mid_1[1031:1024] > btm_1[1031:1024]) ? 1 : 0;
assign detect_max[127][22] = (mid_1[1031:1024] > btm_1[1039:1032]) ? 1 : 0;
assign detect_max[127][23] = (mid_1[1031:1024] > btm_2[1023:1016]) ? 1 : 0;
assign detect_max[127][24] = (mid_1[1031:1024] > btm_2[1031:1024]) ? 1 : 0;
assign detect_max[127][25] = (mid_1[1031:1024] > btm_2[1039:1032]) ? 1 : 0;

assign detect_max[128][0] = (mid_1[1039:1032] > top_0[1031:1024]) ? 1 : 0;
assign detect_max[128][1] = (mid_1[1039:1032] > top_0[1039:1032]) ? 1 : 0;
assign detect_max[128][2] = (mid_1[1039:1032] > top_0[1047:1040]) ? 1 : 0;
assign detect_max[128][3] = (mid_1[1039:1032] > top_1[1031:1024]) ? 1 : 0;
assign detect_max[128][4] = (mid_1[1039:1032] > top_1[1039:1032]) ? 1 : 0;
assign detect_max[128][5] = (mid_1[1039:1032] > top_1[1047:1040]) ? 1 : 0;
assign detect_max[128][6] = (mid_1[1039:1032] > top_2[1031:1024]) ? 1 : 0;
assign detect_max[128][7] = (mid_1[1039:1032] > top_2[1039:1032]) ? 1 : 0;
assign detect_max[128][8] = (mid_1[1039:1032] > top_2[1047:1040]) ? 1 : 0;
assign detect_max[128][9] = (mid_1[1039:1032] > mid_0[1031:1024]) ? 1 : 0;
assign detect_max[128][10] = (mid_1[1039:1032] > mid_0[1039:1032]) ? 1 : 0;
assign detect_max[128][11] = (mid_1[1039:1032] > mid_0[1047:1040]) ? 1 : 0;
assign detect_max[128][12] = (mid_1[1039:1032] > mid_1[1031:1024]) ? 1 : 0;
assign detect_max[128][13] = (mid_1[1039:1032] > mid_1[1047:1040]) ? 1 : 0;
assign detect_max[128][14] = (mid_1[1039:1032] > mid_2[1031:1024]) ? 1 : 0;
assign detect_max[128][15] = (mid_1[1039:1032] > mid_2[1039:1032]) ? 1 : 0;
assign detect_max[128][16] = (mid_1[1039:1032] > mid_2[1047:1040]) ? 1 : 0;
assign detect_max[128][17] = (mid_1[1039:1032] > btm_0[1031:1024]) ? 1 : 0;
assign detect_max[128][18] = (mid_1[1039:1032] > btm_0[1039:1032]) ? 1 : 0;
assign detect_max[128][19] = (mid_1[1039:1032] > btm_0[1047:1040]) ? 1 : 0;
assign detect_max[128][20] = (mid_1[1039:1032] > btm_1[1031:1024]) ? 1 : 0;
assign detect_max[128][21] = (mid_1[1039:1032] > btm_1[1039:1032]) ? 1 : 0;
assign detect_max[128][22] = (mid_1[1039:1032] > btm_1[1047:1040]) ? 1 : 0;
assign detect_max[128][23] = (mid_1[1039:1032] > btm_2[1031:1024]) ? 1 : 0;
assign detect_max[128][24] = (mid_1[1039:1032] > btm_2[1039:1032]) ? 1 : 0;
assign detect_max[128][25] = (mid_1[1039:1032] > btm_2[1047:1040]) ? 1 : 0;

assign detect_max[129][0] = (mid_1[1047:1040] > top_0[1039:1032]) ? 1 : 0;
assign detect_max[129][1] = (mid_1[1047:1040] > top_0[1047:1040]) ? 1 : 0;
assign detect_max[129][2] = (mid_1[1047:1040] > top_0[1055:1048]) ? 1 : 0;
assign detect_max[129][3] = (mid_1[1047:1040] > top_1[1039:1032]) ? 1 : 0;
assign detect_max[129][4] = (mid_1[1047:1040] > top_1[1047:1040]) ? 1 : 0;
assign detect_max[129][5] = (mid_1[1047:1040] > top_1[1055:1048]) ? 1 : 0;
assign detect_max[129][6] = (mid_1[1047:1040] > top_2[1039:1032]) ? 1 : 0;
assign detect_max[129][7] = (mid_1[1047:1040] > top_2[1047:1040]) ? 1 : 0;
assign detect_max[129][8] = (mid_1[1047:1040] > top_2[1055:1048]) ? 1 : 0;
assign detect_max[129][9] = (mid_1[1047:1040] > mid_0[1039:1032]) ? 1 : 0;
assign detect_max[129][10] = (mid_1[1047:1040] > mid_0[1047:1040]) ? 1 : 0;
assign detect_max[129][11] = (mid_1[1047:1040] > mid_0[1055:1048]) ? 1 : 0;
assign detect_max[129][12] = (mid_1[1047:1040] > mid_1[1039:1032]) ? 1 : 0;
assign detect_max[129][13] = (mid_1[1047:1040] > mid_1[1055:1048]) ? 1 : 0;
assign detect_max[129][14] = (mid_1[1047:1040] > mid_2[1039:1032]) ? 1 : 0;
assign detect_max[129][15] = (mid_1[1047:1040] > mid_2[1047:1040]) ? 1 : 0;
assign detect_max[129][16] = (mid_1[1047:1040] > mid_2[1055:1048]) ? 1 : 0;
assign detect_max[129][17] = (mid_1[1047:1040] > btm_0[1039:1032]) ? 1 : 0;
assign detect_max[129][18] = (mid_1[1047:1040] > btm_0[1047:1040]) ? 1 : 0;
assign detect_max[129][19] = (mid_1[1047:1040] > btm_0[1055:1048]) ? 1 : 0;
assign detect_max[129][20] = (mid_1[1047:1040] > btm_1[1039:1032]) ? 1 : 0;
assign detect_max[129][21] = (mid_1[1047:1040] > btm_1[1047:1040]) ? 1 : 0;
assign detect_max[129][22] = (mid_1[1047:1040] > btm_1[1055:1048]) ? 1 : 0;
assign detect_max[129][23] = (mid_1[1047:1040] > btm_2[1039:1032]) ? 1 : 0;
assign detect_max[129][24] = (mid_1[1047:1040] > btm_2[1047:1040]) ? 1 : 0;
assign detect_max[129][25] = (mid_1[1047:1040] > btm_2[1055:1048]) ? 1 : 0;

assign detect_max[130][0] = (mid_1[1055:1048] > top_0[1047:1040]) ? 1 : 0;
assign detect_max[130][1] = (mid_1[1055:1048] > top_0[1055:1048]) ? 1 : 0;
assign detect_max[130][2] = (mid_1[1055:1048] > top_0[1063:1056]) ? 1 : 0;
assign detect_max[130][3] = (mid_1[1055:1048] > top_1[1047:1040]) ? 1 : 0;
assign detect_max[130][4] = (mid_1[1055:1048] > top_1[1055:1048]) ? 1 : 0;
assign detect_max[130][5] = (mid_1[1055:1048] > top_1[1063:1056]) ? 1 : 0;
assign detect_max[130][6] = (mid_1[1055:1048] > top_2[1047:1040]) ? 1 : 0;
assign detect_max[130][7] = (mid_1[1055:1048] > top_2[1055:1048]) ? 1 : 0;
assign detect_max[130][8] = (mid_1[1055:1048] > top_2[1063:1056]) ? 1 : 0;
assign detect_max[130][9] = (mid_1[1055:1048] > mid_0[1047:1040]) ? 1 : 0;
assign detect_max[130][10] = (mid_1[1055:1048] > mid_0[1055:1048]) ? 1 : 0;
assign detect_max[130][11] = (mid_1[1055:1048] > mid_0[1063:1056]) ? 1 : 0;
assign detect_max[130][12] = (mid_1[1055:1048] > mid_1[1047:1040]) ? 1 : 0;
assign detect_max[130][13] = (mid_1[1055:1048] > mid_1[1063:1056]) ? 1 : 0;
assign detect_max[130][14] = (mid_1[1055:1048] > mid_2[1047:1040]) ? 1 : 0;
assign detect_max[130][15] = (mid_1[1055:1048] > mid_2[1055:1048]) ? 1 : 0;
assign detect_max[130][16] = (mid_1[1055:1048] > mid_2[1063:1056]) ? 1 : 0;
assign detect_max[130][17] = (mid_1[1055:1048] > btm_0[1047:1040]) ? 1 : 0;
assign detect_max[130][18] = (mid_1[1055:1048] > btm_0[1055:1048]) ? 1 : 0;
assign detect_max[130][19] = (mid_1[1055:1048] > btm_0[1063:1056]) ? 1 : 0;
assign detect_max[130][20] = (mid_1[1055:1048] > btm_1[1047:1040]) ? 1 : 0;
assign detect_max[130][21] = (mid_1[1055:1048] > btm_1[1055:1048]) ? 1 : 0;
assign detect_max[130][22] = (mid_1[1055:1048] > btm_1[1063:1056]) ? 1 : 0;
assign detect_max[130][23] = (mid_1[1055:1048] > btm_2[1047:1040]) ? 1 : 0;
assign detect_max[130][24] = (mid_1[1055:1048] > btm_2[1055:1048]) ? 1 : 0;
assign detect_max[130][25] = (mid_1[1055:1048] > btm_2[1063:1056]) ? 1 : 0;

assign detect_max[131][0] = (mid_1[1063:1056] > top_0[1055:1048]) ? 1 : 0;
assign detect_max[131][1] = (mid_1[1063:1056] > top_0[1063:1056]) ? 1 : 0;
assign detect_max[131][2] = (mid_1[1063:1056] > top_0[1071:1064]) ? 1 : 0;
assign detect_max[131][3] = (mid_1[1063:1056] > top_1[1055:1048]) ? 1 : 0;
assign detect_max[131][4] = (mid_1[1063:1056] > top_1[1063:1056]) ? 1 : 0;
assign detect_max[131][5] = (mid_1[1063:1056] > top_1[1071:1064]) ? 1 : 0;
assign detect_max[131][6] = (mid_1[1063:1056] > top_2[1055:1048]) ? 1 : 0;
assign detect_max[131][7] = (mid_1[1063:1056] > top_2[1063:1056]) ? 1 : 0;
assign detect_max[131][8] = (mid_1[1063:1056] > top_2[1071:1064]) ? 1 : 0;
assign detect_max[131][9] = (mid_1[1063:1056] > mid_0[1055:1048]) ? 1 : 0;
assign detect_max[131][10] = (mid_1[1063:1056] > mid_0[1063:1056]) ? 1 : 0;
assign detect_max[131][11] = (mid_1[1063:1056] > mid_0[1071:1064]) ? 1 : 0;
assign detect_max[131][12] = (mid_1[1063:1056] > mid_1[1055:1048]) ? 1 : 0;
assign detect_max[131][13] = (mid_1[1063:1056] > mid_1[1071:1064]) ? 1 : 0;
assign detect_max[131][14] = (mid_1[1063:1056] > mid_2[1055:1048]) ? 1 : 0;
assign detect_max[131][15] = (mid_1[1063:1056] > mid_2[1063:1056]) ? 1 : 0;
assign detect_max[131][16] = (mid_1[1063:1056] > mid_2[1071:1064]) ? 1 : 0;
assign detect_max[131][17] = (mid_1[1063:1056] > btm_0[1055:1048]) ? 1 : 0;
assign detect_max[131][18] = (mid_1[1063:1056] > btm_0[1063:1056]) ? 1 : 0;
assign detect_max[131][19] = (mid_1[1063:1056] > btm_0[1071:1064]) ? 1 : 0;
assign detect_max[131][20] = (mid_1[1063:1056] > btm_1[1055:1048]) ? 1 : 0;
assign detect_max[131][21] = (mid_1[1063:1056] > btm_1[1063:1056]) ? 1 : 0;
assign detect_max[131][22] = (mid_1[1063:1056] > btm_1[1071:1064]) ? 1 : 0;
assign detect_max[131][23] = (mid_1[1063:1056] > btm_2[1055:1048]) ? 1 : 0;
assign detect_max[131][24] = (mid_1[1063:1056] > btm_2[1063:1056]) ? 1 : 0;
assign detect_max[131][25] = (mid_1[1063:1056] > btm_2[1071:1064]) ? 1 : 0;

assign detect_max[132][0] = (mid_1[1071:1064] > top_0[1063:1056]) ? 1 : 0;
assign detect_max[132][1] = (mid_1[1071:1064] > top_0[1071:1064]) ? 1 : 0;
assign detect_max[132][2] = (mid_1[1071:1064] > top_0[1079:1072]) ? 1 : 0;
assign detect_max[132][3] = (mid_1[1071:1064] > top_1[1063:1056]) ? 1 : 0;
assign detect_max[132][4] = (mid_1[1071:1064] > top_1[1071:1064]) ? 1 : 0;
assign detect_max[132][5] = (mid_1[1071:1064] > top_1[1079:1072]) ? 1 : 0;
assign detect_max[132][6] = (mid_1[1071:1064] > top_2[1063:1056]) ? 1 : 0;
assign detect_max[132][7] = (mid_1[1071:1064] > top_2[1071:1064]) ? 1 : 0;
assign detect_max[132][8] = (mid_1[1071:1064] > top_2[1079:1072]) ? 1 : 0;
assign detect_max[132][9] = (mid_1[1071:1064] > mid_0[1063:1056]) ? 1 : 0;
assign detect_max[132][10] = (mid_1[1071:1064] > mid_0[1071:1064]) ? 1 : 0;
assign detect_max[132][11] = (mid_1[1071:1064] > mid_0[1079:1072]) ? 1 : 0;
assign detect_max[132][12] = (mid_1[1071:1064] > mid_1[1063:1056]) ? 1 : 0;
assign detect_max[132][13] = (mid_1[1071:1064] > mid_1[1079:1072]) ? 1 : 0;
assign detect_max[132][14] = (mid_1[1071:1064] > mid_2[1063:1056]) ? 1 : 0;
assign detect_max[132][15] = (mid_1[1071:1064] > mid_2[1071:1064]) ? 1 : 0;
assign detect_max[132][16] = (mid_1[1071:1064] > mid_2[1079:1072]) ? 1 : 0;
assign detect_max[132][17] = (mid_1[1071:1064] > btm_0[1063:1056]) ? 1 : 0;
assign detect_max[132][18] = (mid_1[1071:1064] > btm_0[1071:1064]) ? 1 : 0;
assign detect_max[132][19] = (mid_1[1071:1064] > btm_0[1079:1072]) ? 1 : 0;
assign detect_max[132][20] = (mid_1[1071:1064] > btm_1[1063:1056]) ? 1 : 0;
assign detect_max[132][21] = (mid_1[1071:1064] > btm_1[1071:1064]) ? 1 : 0;
assign detect_max[132][22] = (mid_1[1071:1064] > btm_1[1079:1072]) ? 1 : 0;
assign detect_max[132][23] = (mid_1[1071:1064] > btm_2[1063:1056]) ? 1 : 0;
assign detect_max[132][24] = (mid_1[1071:1064] > btm_2[1071:1064]) ? 1 : 0;
assign detect_max[132][25] = (mid_1[1071:1064] > btm_2[1079:1072]) ? 1 : 0;

assign detect_max[133][0] = (mid_1[1079:1072] > top_0[1071:1064]) ? 1 : 0;
assign detect_max[133][1] = (mid_1[1079:1072] > top_0[1079:1072]) ? 1 : 0;
assign detect_max[133][2] = (mid_1[1079:1072] > top_0[1087:1080]) ? 1 : 0;
assign detect_max[133][3] = (mid_1[1079:1072] > top_1[1071:1064]) ? 1 : 0;
assign detect_max[133][4] = (mid_1[1079:1072] > top_1[1079:1072]) ? 1 : 0;
assign detect_max[133][5] = (mid_1[1079:1072] > top_1[1087:1080]) ? 1 : 0;
assign detect_max[133][6] = (mid_1[1079:1072] > top_2[1071:1064]) ? 1 : 0;
assign detect_max[133][7] = (mid_1[1079:1072] > top_2[1079:1072]) ? 1 : 0;
assign detect_max[133][8] = (mid_1[1079:1072] > top_2[1087:1080]) ? 1 : 0;
assign detect_max[133][9] = (mid_1[1079:1072] > mid_0[1071:1064]) ? 1 : 0;
assign detect_max[133][10] = (mid_1[1079:1072] > mid_0[1079:1072]) ? 1 : 0;
assign detect_max[133][11] = (mid_1[1079:1072] > mid_0[1087:1080]) ? 1 : 0;
assign detect_max[133][12] = (mid_1[1079:1072] > mid_1[1071:1064]) ? 1 : 0;
assign detect_max[133][13] = (mid_1[1079:1072] > mid_1[1087:1080]) ? 1 : 0;
assign detect_max[133][14] = (mid_1[1079:1072] > mid_2[1071:1064]) ? 1 : 0;
assign detect_max[133][15] = (mid_1[1079:1072] > mid_2[1079:1072]) ? 1 : 0;
assign detect_max[133][16] = (mid_1[1079:1072] > mid_2[1087:1080]) ? 1 : 0;
assign detect_max[133][17] = (mid_1[1079:1072] > btm_0[1071:1064]) ? 1 : 0;
assign detect_max[133][18] = (mid_1[1079:1072] > btm_0[1079:1072]) ? 1 : 0;
assign detect_max[133][19] = (mid_1[1079:1072] > btm_0[1087:1080]) ? 1 : 0;
assign detect_max[133][20] = (mid_1[1079:1072] > btm_1[1071:1064]) ? 1 : 0;
assign detect_max[133][21] = (mid_1[1079:1072] > btm_1[1079:1072]) ? 1 : 0;
assign detect_max[133][22] = (mid_1[1079:1072] > btm_1[1087:1080]) ? 1 : 0;
assign detect_max[133][23] = (mid_1[1079:1072] > btm_2[1071:1064]) ? 1 : 0;
assign detect_max[133][24] = (mid_1[1079:1072] > btm_2[1079:1072]) ? 1 : 0;
assign detect_max[133][25] = (mid_1[1079:1072] > btm_2[1087:1080]) ? 1 : 0;

assign detect_max[134][0] = (mid_1[1087:1080] > top_0[1079:1072]) ? 1 : 0;
assign detect_max[134][1] = (mid_1[1087:1080] > top_0[1087:1080]) ? 1 : 0;
assign detect_max[134][2] = (mid_1[1087:1080] > top_0[1095:1088]) ? 1 : 0;
assign detect_max[134][3] = (mid_1[1087:1080] > top_1[1079:1072]) ? 1 : 0;
assign detect_max[134][4] = (mid_1[1087:1080] > top_1[1087:1080]) ? 1 : 0;
assign detect_max[134][5] = (mid_1[1087:1080] > top_1[1095:1088]) ? 1 : 0;
assign detect_max[134][6] = (mid_1[1087:1080] > top_2[1079:1072]) ? 1 : 0;
assign detect_max[134][7] = (mid_1[1087:1080] > top_2[1087:1080]) ? 1 : 0;
assign detect_max[134][8] = (mid_1[1087:1080] > top_2[1095:1088]) ? 1 : 0;
assign detect_max[134][9] = (mid_1[1087:1080] > mid_0[1079:1072]) ? 1 : 0;
assign detect_max[134][10] = (mid_1[1087:1080] > mid_0[1087:1080]) ? 1 : 0;
assign detect_max[134][11] = (mid_1[1087:1080] > mid_0[1095:1088]) ? 1 : 0;
assign detect_max[134][12] = (mid_1[1087:1080] > mid_1[1079:1072]) ? 1 : 0;
assign detect_max[134][13] = (mid_1[1087:1080] > mid_1[1095:1088]) ? 1 : 0;
assign detect_max[134][14] = (mid_1[1087:1080] > mid_2[1079:1072]) ? 1 : 0;
assign detect_max[134][15] = (mid_1[1087:1080] > mid_2[1087:1080]) ? 1 : 0;
assign detect_max[134][16] = (mid_1[1087:1080] > mid_2[1095:1088]) ? 1 : 0;
assign detect_max[134][17] = (mid_1[1087:1080] > btm_0[1079:1072]) ? 1 : 0;
assign detect_max[134][18] = (mid_1[1087:1080] > btm_0[1087:1080]) ? 1 : 0;
assign detect_max[134][19] = (mid_1[1087:1080] > btm_0[1095:1088]) ? 1 : 0;
assign detect_max[134][20] = (mid_1[1087:1080] > btm_1[1079:1072]) ? 1 : 0;
assign detect_max[134][21] = (mid_1[1087:1080] > btm_1[1087:1080]) ? 1 : 0;
assign detect_max[134][22] = (mid_1[1087:1080] > btm_1[1095:1088]) ? 1 : 0;
assign detect_max[134][23] = (mid_1[1087:1080] > btm_2[1079:1072]) ? 1 : 0;
assign detect_max[134][24] = (mid_1[1087:1080] > btm_2[1087:1080]) ? 1 : 0;
assign detect_max[134][25] = (mid_1[1087:1080] > btm_2[1095:1088]) ? 1 : 0;

assign detect_max[135][0] = (mid_1[1095:1088] > top_0[1087:1080]) ? 1 : 0;
assign detect_max[135][1] = (mid_1[1095:1088] > top_0[1095:1088]) ? 1 : 0;
assign detect_max[135][2] = (mid_1[1095:1088] > top_0[1103:1096]) ? 1 : 0;
assign detect_max[135][3] = (mid_1[1095:1088] > top_1[1087:1080]) ? 1 : 0;
assign detect_max[135][4] = (mid_1[1095:1088] > top_1[1095:1088]) ? 1 : 0;
assign detect_max[135][5] = (mid_1[1095:1088] > top_1[1103:1096]) ? 1 : 0;
assign detect_max[135][6] = (mid_1[1095:1088] > top_2[1087:1080]) ? 1 : 0;
assign detect_max[135][7] = (mid_1[1095:1088] > top_2[1095:1088]) ? 1 : 0;
assign detect_max[135][8] = (mid_1[1095:1088] > top_2[1103:1096]) ? 1 : 0;
assign detect_max[135][9] = (mid_1[1095:1088] > mid_0[1087:1080]) ? 1 : 0;
assign detect_max[135][10] = (mid_1[1095:1088] > mid_0[1095:1088]) ? 1 : 0;
assign detect_max[135][11] = (mid_1[1095:1088] > mid_0[1103:1096]) ? 1 : 0;
assign detect_max[135][12] = (mid_1[1095:1088] > mid_1[1087:1080]) ? 1 : 0;
assign detect_max[135][13] = (mid_1[1095:1088] > mid_1[1103:1096]) ? 1 : 0;
assign detect_max[135][14] = (mid_1[1095:1088] > mid_2[1087:1080]) ? 1 : 0;
assign detect_max[135][15] = (mid_1[1095:1088] > mid_2[1095:1088]) ? 1 : 0;
assign detect_max[135][16] = (mid_1[1095:1088] > mid_2[1103:1096]) ? 1 : 0;
assign detect_max[135][17] = (mid_1[1095:1088] > btm_0[1087:1080]) ? 1 : 0;
assign detect_max[135][18] = (mid_1[1095:1088] > btm_0[1095:1088]) ? 1 : 0;
assign detect_max[135][19] = (mid_1[1095:1088] > btm_0[1103:1096]) ? 1 : 0;
assign detect_max[135][20] = (mid_1[1095:1088] > btm_1[1087:1080]) ? 1 : 0;
assign detect_max[135][21] = (mid_1[1095:1088] > btm_1[1095:1088]) ? 1 : 0;
assign detect_max[135][22] = (mid_1[1095:1088] > btm_1[1103:1096]) ? 1 : 0;
assign detect_max[135][23] = (mid_1[1095:1088] > btm_2[1087:1080]) ? 1 : 0;
assign detect_max[135][24] = (mid_1[1095:1088] > btm_2[1095:1088]) ? 1 : 0;
assign detect_max[135][25] = (mid_1[1095:1088] > btm_2[1103:1096]) ? 1 : 0;

assign detect_max[136][0] = (mid_1[1103:1096] > top_0[1095:1088]) ? 1 : 0;
assign detect_max[136][1] = (mid_1[1103:1096] > top_0[1103:1096]) ? 1 : 0;
assign detect_max[136][2] = (mid_1[1103:1096] > top_0[1111:1104]) ? 1 : 0;
assign detect_max[136][3] = (mid_1[1103:1096] > top_1[1095:1088]) ? 1 : 0;
assign detect_max[136][4] = (mid_1[1103:1096] > top_1[1103:1096]) ? 1 : 0;
assign detect_max[136][5] = (mid_1[1103:1096] > top_1[1111:1104]) ? 1 : 0;
assign detect_max[136][6] = (mid_1[1103:1096] > top_2[1095:1088]) ? 1 : 0;
assign detect_max[136][7] = (mid_1[1103:1096] > top_2[1103:1096]) ? 1 : 0;
assign detect_max[136][8] = (mid_1[1103:1096] > top_2[1111:1104]) ? 1 : 0;
assign detect_max[136][9] = (mid_1[1103:1096] > mid_0[1095:1088]) ? 1 : 0;
assign detect_max[136][10] = (mid_1[1103:1096] > mid_0[1103:1096]) ? 1 : 0;
assign detect_max[136][11] = (mid_1[1103:1096] > mid_0[1111:1104]) ? 1 : 0;
assign detect_max[136][12] = (mid_1[1103:1096] > mid_1[1095:1088]) ? 1 : 0;
assign detect_max[136][13] = (mid_1[1103:1096] > mid_1[1111:1104]) ? 1 : 0;
assign detect_max[136][14] = (mid_1[1103:1096] > mid_2[1095:1088]) ? 1 : 0;
assign detect_max[136][15] = (mid_1[1103:1096] > mid_2[1103:1096]) ? 1 : 0;
assign detect_max[136][16] = (mid_1[1103:1096] > mid_2[1111:1104]) ? 1 : 0;
assign detect_max[136][17] = (mid_1[1103:1096] > btm_0[1095:1088]) ? 1 : 0;
assign detect_max[136][18] = (mid_1[1103:1096] > btm_0[1103:1096]) ? 1 : 0;
assign detect_max[136][19] = (mid_1[1103:1096] > btm_0[1111:1104]) ? 1 : 0;
assign detect_max[136][20] = (mid_1[1103:1096] > btm_1[1095:1088]) ? 1 : 0;
assign detect_max[136][21] = (mid_1[1103:1096] > btm_1[1103:1096]) ? 1 : 0;
assign detect_max[136][22] = (mid_1[1103:1096] > btm_1[1111:1104]) ? 1 : 0;
assign detect_max[136][23] = (mid_1[1103:1096] > btm_2[1095:1088]) ? 1 : 0;
assign detect_max[136][24] = (mid_1[1103:1096] > btm_2[1103:1096]) ? 1 : 0;
assign detect_max[136][25] = (mid_1[1103:1096] > btm_2[1111:1104]) ? 1 : 0;

assign detect_max[137][0] = (mid_1[1111:1104] > top_0[1103:1096]) ? 1 : 0;
assign detect_max[137][1] = (mid_1[1111:1104] > top_0[1111:1104]) ? 1 : 0;
assign detect_max[137][2] = (mid_1[1111:1104] > top_0[1119:1112]) ? 1 : 0;
assign detect_max[137][3] = (mid_1[1111:1104] > top_1[1103:1096]) ? 1 : 0;
assign detect_max[137][4] = (mid_1[1111:1104] > top_1[1111:1104]) ? 1 : 0;
assign detect_max[137][5] = (mid_1[1111:1104] > top_1[1119:1112]) ? 1 : 0;
assign detect_max[137][6] = (mid_1[1111:1104] > top_2[1103:1096]) ? 1 : 0;
assign detect_max[137][7] = (mid_1[1111:1104] > top_2[1111:1104]) ? 1 : 0;
assign detect_max[137][8] = (mid_1[1111:1104] > top_2[1119:1112]) ? 1 : 0;
assign detect_max[137][9] = (mid_1[1111:1104] > mid_0[1103:1096]) ? 1 : 0;
assign detect_max[137][10] = (mid_1[1111:1104] > mid_0[1111:1104]) ? 1 : 0;
assign detect_max[137][11] = (mid_1[1111:1104] > mid_0[1119:1112]) ? 1 : 0;
assign detect_max[137][12] = (mid_1[1111:1104] > mid_1[1103:1096]) ? 1 : 0;
assign detect_max[137][13] = (mid_1[1111:1104] > mid_1[1119:1112]) ? 1 : 0;
assign detect_max[137][14] = (mid_1[1111:1104] > mid_2[1103:1096]) ? 1 : 0;
assign detect_max[137][15] = (mid_1[1111:1104] > mid_2[1111:1104]) ? 1 : 0;
assign detect_max[137][16] = (mid_1[1111:1104] > mid_2[1119:1112]) ? 1 : 0;
assign detect_max[137][17] = (mid_1[1111:1104] > btm_0[1103:1096]) ? 1 : 0;
assign detect_max[137][18] = (mid_1[1111:1104] > btm_0[1111:1104]) ? 1 : 0;
assign detect_max[137][19] = (mid_1[1111:1104] > btm_0[1119:1112]) ? 1 : 0;
assign detect_max[137][20] = (mid_1[1111:1104] > btm_1[1103:1096]) ? 1 : 0;
assign detect_max[137][21] = (mid_1[1111:1104] > btm_1[1111:1104]) ? 1 : 0;
assign detect_max[137][22] = (mid_1[1111:1104] > btm_1[1119:1112]) ? 1 : 0;
assign detect_max[137][23] = (mid_1[1111:1104] > btm_2[1103:1096]) ? 1 : 0;
assign detect_max[137][24] = (mid_1[1111:1104] > btm_2[1111:1104]) ? 1 : 0;
assign detect_max[137][25] = (mid_1[1111:1104] > btm_2[1119:1112]) ? 1 : 0;

assign detect_max[138][0] = (mid_1[1119:1112] > top_0[1111:1104]) ? 1 : 0;
assign detect_max[138][1] = (mid_1[1119:1112] > top_0[1119:1112]) ? 1 : 0;
assign detect_max[138][2] = (mid_1[1119:1112] > top_0[1127:1120]) ? 1 : 0;
assign detect_max[138][3] = (mid_1[1119:1112] > top_1[1111:1104]) ? 1 : 0;
assign detect_max[138][4] = (mid_1[1119:1112] > top_1[1119:1112]) ? 1 : 0;
assign detect_max[138][5] = (mid_1[1119:1112] > top_1[1127:1120]) ? 1 : 0;
assign detect_max[138][6] = (mid_1[1119:1112] > top_2[1111:1104]) ? 1 : 0;
assign detect_max[138][7] = (mid_1[1119:1112] > top_2[1119:1112]) ? 1 : 0;
assign detect_max[138][8] = (mid_1[1119:1112] > top_2[1127:1120]) ? 1 : 0;
assign detect_max[138][9] = (mid_1[1119:1112] > mid_0[1111:1104]) ? 1 : 0;
assign detect_max[138][10] = (mid_1[1119:1112] > mid_0[1119:1112]) ? 1 : 0;
assign detect_max[138][11] = (mid_1[1119:1112] > mid_0[1127:1120]) ? 1 : 0;
assign detect_max[138][12] = (mid_1[1119:1112] > mid_1[1111:1104]) ? 1 : 0;
assign detect_max[138][13] = (mid_1[1119:1112] > mid_1[1127:1120]) ? 1 : 0;
assign detect_max[138][14] = (mid_1[1119:1112] > mid_2[1111:1104]) ? 1 : 0;
assign detect_max[138][15] = (mid_1[1119:1112] > mid_2[1119:1112]) ? 1 : 0;
assign detect_max[138][16] = (mid_1[1119:1112] > mid_2[1127:1120]) ? 1 : 0;
assign detect_max[138][17] = (mid_1[1119:1112] > btm_0[1111:1104]) ? 1 : 0;
assign detect_max[138][18] = (mid_1[1119:1112] > btm_0[1119:1112]) ? 1 : 0;
assign detect_max[138][19] = (mid_1[1119:1112] > btm_0[1127:1120]) ? 1 : 0;
assign detect_max[138][20] = (mid_1[1119:1112] > btm_1[1111:1104]) ? 1 : 0;
assign detect_max[138][21] = (mid_1[1119:1112] > btm_1[1119:1112]) ? 1 : 0;
assign detect_max[138][22] = (mid_1[1119:1112] > btm_1[1127:1120]) ? 1 : 0;
assign detect_max[138][23] = (mid_1[1119:1112] > btm_2[1111:1104]) ? 1 : 0;
assign detect_max[138][24] = (mid_1[1119:1112] > btm_2[1119:1112]) ? 1 : 0;
assign detect_max[138][25] = (mid_1[1119:1112] > btm_2[1127:1120]) ? 1 : 0;

assign detect_max[139][0] = (mid_1[1127:1120] > top_0[1119:1112]) ? 1 : 0;
assign detect_max[139][1] = (mid_1[1127:1120] > top_0[1127:1120]) ? 1 : 0;
assign detect_max[139][2] = (mid_1[1127:1120] > top_0[1135:1128]) ? 1 : 0;
assign detect_max[139][3] = (mid_1[1127:1120] > top_1[1119:1112]) ? 1 : 0;
assign detect_max[139][4] = (mid_1[1127:1120] > top_1[1127:1120]) ? 1 : 0;
assign detect_max[139][5] = (mid_1[1127:1120] > top_1[1135:1128]) ? 1 : 0;
assign detect_max[139][6] = (mid_1[1127:1120] > top_2[1119:1112]) ? 1 : 0;
assign detect_max[139][7] = (mid_1[1127:1120] > top_2[1127:1120]) ? 1 : 0;
assign detect_max[139][8] = (mid_1[1127:1120] > top_2[1135:1128]) ? 1 : 0;
assign detect_max[139][9] = (mid_1[1127:1120] > mid_0[1119:1112]) ? 1 : 0;
assign detect_max[139][10] = (mid_1[1127:1120] > mid_0[1127:1120]) ? 1 : 0;
assign detect_max[139][11] = (mid_1[1127:1120] > mid_0[1135:1128]) ? 1 : 0;
assign detect_max[139][12] = (mid_1[1127:1120] > mid_1[1119:1112]) ? 1 : 0;
assign detect_max[139][13] = (mid_1[1127:1120] > mid_1[1135:1128]) ? 1 : 0;
assign detect_max[139][14] = (mid_1[1127:1120] > mid_2[1119:1112]) ? 1 : 0;
assign detect_max[139][15] = (mid_1[1127:1120] > mid_2[1127:1120]) ? 1 : 0;
assign detect_max[139][16] = (mid_1[1127:1120] > mid_2[1135:1128]) ? 1 : 0;
assign detect_max[139][17] = (mid_1[1127:1120] > btm_0[1119:1112]) ? 1 : 0;
assign detect_max[139][18] = (mid_1[1127:1120] > btm_0[1127:1120]) ? 1 : 0;
assign detect_max[139][19] = (mid_1[1127:1120] > btm_0[1135:1128]) ? 1 : 0;
assign detect_max[139][20] = (mid_1[1127:1120] > btm_1[1119:1112]) ? 1 : 0;
assign detect_max[139][21] = (mid_1[1127:1120] > btm_1[1127:1120]) ? 1 : 0;
assign detect_max[139][22] = (mid_1[1127:1120] > btm_1[1135:1128]) ? 1 : 0;
assign detect_max[139][23] = (mid_1[1127:1120] > btm_2[1119:1112]) ? 1 : 0;
assign detect_max[139][24] = (mid_1[1127:1120] > btm_2[1127:1120]) ? 1 : 0;
assign detect_max[139][25] = (mid_1[1127:1120] > btm_2[1135:1128]) ? 1 : 0;

assign detect_max[140][0] = (mid_1[1135:1128] > top_0[1127:1120]) ? 1 : 0;
assign detect_max[140][1] = (mid_1[1135:1128] > top_0[1135:1128]) ? 1 : 0;
assign detect_max[140][2] = (mid_1[1135:1128] > top_0[1143:1136]) ? 1 : 0;
assign detect_max[140][3] = (mid_1[1135:1128] > top_1[1127:1120]) ? 1 : 0;
assign detect_max[140][4] = (mid_1[1135:1128] > top_1[1135:1128]) ? 1 : 0;
assign detect_max[140][5] = (mid_1[1135:1128] > top_1[1143:1136]) ? 1 : 0;
assign detect_max[140][6] = (mid_1[1135:1128] > top_2[1127:1120]) ? 1 : 0;
assign detect_max[140][7] = (mid_1[1135:1128] > top_2[1135:1128]) ? 1 : 0;
assign detect_max[140][8] = (mid_1[1135:1128] > top_2[1143:1136]) ? 1 : 0;
assign detect_max[140][9] = (mid_1[1135:1128] > mid_0[1127:1120]) ? 1 : 0;
assign detect_max[140][10] = (mid_1[1135:1128] > mid_0[1135:1128]) ? 1 : 0;
assign detect_max[140][11] = (mid_1[1135:1128] > mid_0[1143:1136]) ? 1 : 0;
assign detect_max[140][12] = (mid_1[1135:1128] > mid_1[1127:1120]) ? 1 : 0;
assign detect_max[140][13] = (mid_1[1135:1128] > mid_1[1143:1136]) ? 1 : 0;
assign detect_max[140][14] = (mid_1[1135:1128] > mid_2[1127:1120]) ? 1 : 0;
assign detect_max[140][15] = (mid_1[1135:1128] > mid_2[1135:1128]) ? 1 : 0;
assign detect_max[140][16] = (mid_1[1135:1128] > mid_2[1143:1136]) ? 1 : 0;
assign detect_max[140][17] = (mid_1[1135:1128] > btm_0[1127:1120]) ? 1 : 0;
assign detect_max[140][18] = (mid_1[1135:1128] > btm_0[1135:1128]) ? 1 : 0;
assign detect_max[140][19] = (mid_1[1135:1128] > btm_0[1143:1136]) ? 1 : 0;
assign detect_max[140][20] = (mid_1[1135:1128] > btm_1[1127:1120]) ? 1 : 0;
assign detect_max[140][21] = (mid_1[1135:1128] > btm_1[1135:1128]) ? 1 : 0;
assign detect_max[140][22] = (mid_1[1135:1128] > btm_1[1143:1136]) ? 1 : 0;
assign detect_max[140][23] = (mid_1[1135:1128] > btm_2[1127:1120]) ? 1 : 0;
assign detect_max[140][24] = (mid_1[1135:1128] > btm_2[1135:1128]) ? 1 : 0;
assign detect_max[140][25] = (mid_1[1135:1128] > btm_2[1143:1136]) ? 1 : 0;

assign detect_max[141][0] = (mid_1[1143:1136] > top_0[1135:1128]) ? 1 : 0;
assign detect_max[141][1] = (mid_1[1143:1136] > top_0[1143:1136]) ? 1 : 0;
assign detect_max[141][2] = (mid_1[1143:1136] > top_0[1151:1144]) ? 1 : 0;
assign detect_max[141][3] = (mid_1[1143:1136] > top_1[1135:1128]) ? 1 : 0;
assign detect_max[141][4] = (mid_1[1143:1136] > top_1[1143:1136]) ? 1 : 0;
assign detect_max[141][5] = (mid_1[1143:1136] > top_1[1151:1144]) ? 1 : 0;
assign detect_max[141][6] = (mid_1[1143:1136] > top_2[1135:1128]) ? 1 : 0;
assign detect_max[141][7] = (mid_1[1143:1136] > top_2[1143:1136]) ? 1 : 0;
assign detect_max[141][8] = (mid_1[1143:1136] > top_2[1151:1144]) ? 1 : 0;
assign detect_max[141][9] = (mid_1[1143:1136] > mid_0[1135:1128]) ? 1 : 0;
assign detect_max[141][10] = (mid_1[1143:1136] > mid_0[1143:1136]) ? 1 : 0;
assign detect_max[141][11] = (mid_1[1143:1136] > mid_0[1151:1144]) ? 1 : 0;
assign detect_max[141][12] = (mid_1[1143:1136] > mid_1[1135:1128]) ? 1 : 0;
assign detect_max[141][13] = (mid_1[1143:1136] > mid_1[1151:1144]) ? 1 : 0;
assign detect_max[141][14] = (mid_1[1143:1136] > mid_2[1135:1128]) ? 1 : 0;
assign detect_max[141][15] = (mid_1[1143:1136] > mid_2[1143:1136]) ? 1 : 0;
assign detect_max[141][16] = (mid_1[1143:1136] > mid_2[1151:1144]) ? 1 : 0;
assign detect_max[141][17] = (mid_1[1143:1136] > btm_0[1135:1128]) ? 1 : 0;
assign detect_max[141][18] = (mid_1[1143:1136] > btm_0[1143:1136]) ? 1 : 0;
assign detect_max[141][19] = (mid_1[1143:1136] > btm_0[1151:1144]) ? 1 : 0;
assign detect_max[141][20] = (mid_1[1143:1136] > btm_1[1135:1128]) ? 1 : 0;
assign detect_max[141][21] = (mid_1[1143:1136] > btm_1[1143:1136]) ? 1 : 0;
assign detect_max[141][22] = (mid_1[1143:1136] > btm_1[1151:1144]) ? 1 : 0;
assign detect_max[141][23] = (mid_1[1143:1136] > btm_2[1135:1128]) ? 1 : 0;
assign detect_max[141][24] = (mid_1[1143:1136] > btm_2[1143:1136]) ? 1 : 0;
assign detect_max[141][25] = (mid_1[1143:1136] > btm_2[1151:1144]) ? 1 : 0;

assign detect_max[142][0] = (mid_1[1151:1144] > top_0[1143:1136]) ? 1 : 0;
assign detect_max[142][1] = (mid_1[1151:1144] > top_0[1151:1144]) ? 1 : 0;
assign detect_max[142][2] = (mid_1[1151:1144] > top_0[1159:1152]) ? 1 : 0;
assign detect_max[142][3] = (mid_1[1151:1144] > top_1[1143:1136]) ? 1 : 0;
assign detect_max[142][4] = (mid_1[1151:1144] > top_1[1151:1144]) ? 1 : 0;
assign detect_max[142][5] = (mid_1[1151:1144] > top_1[1159:1152]) ? 1 : 0;
assign detect_max[142][6] = (mid_1[1151:1144] > top_2[1143:1136]) ? 1 : 0;
assign detect_max[142][7] = (mid_1[1151:1144] > top_2[1151:1144]) ? 1 : 0;
assign detect_max[142][8] = (mid_1[1151:1144] > top_2[1159:1152]) ? 1 : 0;
assign detect_max[142][9] = (mid_1[1151:1144] > mid_0[1143:1136]) ? 1 : 0;
assign detect_max[142][10] = (mid_1[1151:1144] > mid_0[1151:1144]) ? 1 : 0;
assign detect_max[142][11] = (mid_1[1151:1144] > mid_0[1159:1152]) ? 1 : 0;
assign detect_max[142][12] = (mid_1[1151:1144] > mid_1[1143:1136]) ? 1 : 0;
assign detect_max[142][13] = (mid_1[1151:1144] > mid_1[1159:1152]) ? 1 : 0;
assign detect_max[142][14] = (mid_1[1151:1144] > mid_2[1143:1136]) ? 1 : 0;
assign detect_max[142][15] = (mid_1[1151:1144] > mid_2[1151:1144]) ? 1 : 0;
assign detect_max[142][16] = (mid_1[1151:1144] > mid_2[1159:1152]) ? 1 : 0;
assign detect_max[142][17] = (mid_1[1151:1144] > btm_0[1143:1136]) ? 1 : 0;
assign detect_max[142][18] = (mid_1[1151:1144] > btm_0[1151:1144]) ? 1 : 0;
assign detect_max[142][19] = (mid_1[1151:1144] > btm_0[1159:1152]) ? 1 : 0;
assign detect_max[142][20] = (mid_1[1151:1144] > btm_1[1143:1136]) ? 1 : 0;
assign detect_max[142][21] = (mid_1[1151:1144] > btm_1[1151:1144]) ? 1 : 0;
assign detect_max[142][22] = (mid_1[1151:1144] > btm_1[1159:1152]) ? 1 : 0;
assign detect_max[142][23] = (mid_1[1151:1144] > btm_2[1143:1136]) ? 1 : 0;
assign detect_max[142][24] = (mid_1[1151:1144] > btm_2[1151:1144]) ? 1 : 0;
assign detect_max[142][25] = (mid_1[1151:1144] > btm_2[1159:1152]) ? 1 : 0;

assign detect_max[143][0] = (mid_1[1159:1152] > top_0[1151:1144]) ? 1 : 0;
assign detect_max[143][1] = (mid_1[1159:1152] > top_0[1159:1152]) ? 1 : 0;
assign detect_max[143][2] = (mid_1[1159:1152] > top_0[1167:1160]) ? 1 : 0;
assign detect_max[143][3] = (mid_1[1159:1152] > top_1[1151:1144]) ? 1 : 0;
assign detect_max[143][4] = (mid_1[1159:1152] > top_1[1159:1152]) ? 1 : 0;
assign detect_max[143][5] = (mid_1[1159:1152] > top_1[1167:1160]) ? 1 : 0;
assign detect_max[143][6] = (mid_1[1159:1152] > top_2[1151:1144]) ? 1 : 0;
assign detect_max[143][7] = (mid_1[1159:1152] > top_2[1159:1152]) ? 1 : 0;
assign detect_max[143][8] = (mid_1[1159:1152] > top_2[1167:1160]) ? 1 : 0;
assign detect_max[143][9] = (mid_1[1159:1152] > mid_0[1151:1144]) ? 1 : 0;
assign detect_max[143][10] = (mid_1[1159:1152] > mid_0[1159:1152]) ? 1 : 0;
assign detect_max[143][11] = (mid_1[1159:1152] > mid_0[1167:1160]) ? 1 : 0;
assign detect_max[143][12] = (mid_1[1159:1152] > mid_1[1151:1144]) ? 1 : 0;
assign detect_max[143][13] = (mid_1[1159:1152] > mid_1[1167:1160]) ? 1 : 0;
assign detect_max[143][14] = (mid_1[1159:1152] > mid_2[1151:1144]) ? 1 : 0;
assign detect_max[143][15] = (mid_1[1159:1152] > mid_2[1159:1152]) ? 1 : 0;
assign detect_max[143][16] = (mid_1[1159:1152] > mid_2[1167:1160]) ? 1 : 0;
assign detect_max[143][17] = (mid_1[1159:1152] > btm_0[1151:1144]) ? 1 : 0;
assign detect_max[143][18] = (mid_1[1159:1152] > btm_0[1159:1152]) ? 1 : 0;
assign detect_max[143][19] = (mid_1[1159:1152] > btm_0[1167:1160]) ? 1 : 0;
assign detect_max[143][20] = (mid_1[1159:1152] > btm_1[1151:1144]) ? 1 : 0;
assign detect_max[143][21] = (mid_1[1159:1152] > btm_1[1159:1152]) ? 1 : 0;
assign detect_max[143][22] = (mid_1[1159:1152] > btm_1[1167:1160]) ? 1 : 0;
assign detect_max[143][23] = (mid_1[1159:1152] > btm_2[1151:1144]) ? 1 : 0;
assign detect_max[143][24] = (mid_1[1159:1152] > btm_2[1159:1152]) ? 1 : 0;
assign detect_max[143][25] = (mid_1[1159:1152] > btm_2[1167:1160]) ? 1 : 0;

assign detect_max[144][0] = (mid_1[1167:1160] > top_0[1159:1152]) ? 1 : 0;
assign detect_max[144][1] = (mid_1[1167:1160] > top_0[1167:1160]) ? 1 : 0;
assign detect_max[144][2] = (mid_1[1167:1160] > top_0[1175:1168]) ? 1 : 0;
assign detect_max[144][3] = (mid_1[1167:1160] > top_1[1159:1152]) ? 1 : 0;
assign detect_max[144][4] = (mid_1[1167:1160] > top_1[1167:1160]) ? 1 : 0;
assign detect_max[144][5] = (mid_1[1167:1160] > top_1[1175:1168]) ? 1 : 0;
assign detect_max[144][6] = (mid_1[1167:1160] > top_2[1159:1152]) ? 1 : 0;
assign detect_max[144][7] = (mid_1[1167:1160] > top_2[1167:1160]) ? 1 : 0;
assign detect_max[144][8] = (mid_1[1167:1160] > top_2[1175:1168]) ? 1 : 0;
assign detect_max[144][9] = (mid_1[1167:1160] > mid_0[1159:1152]) ? 1 : 0;
assign detect_max[144][10] = (mid_1[1167:1160] > mid_0[1167:1160]) ? 1 : 0;
assign detect_max[144][11] = (mid_1[1167:1160] > mid_0[1175:1168]) ? 1 : 0;
assign detect_max[144][12] = (mid_1[1167:1160] > mid_1[1159:1152]) ? 1 : 0;
assign detect_max[144][13] = (mid_1[1167:1160] > mid_1[1175:1168]) ? 1 : 0;
assign detect_max[144][14] = (mid_1[1167:1160] > mid_2[1159:1152]) ? 1 : 0;
assign detect_max[144][15] = (mid_1[1167:1160] > mid_2[1167:1160]) ? 1 : 0;
assign detect_max[144][16] = (mid_1[1167:1160] > mid_2[1175:1168]) ? 1 : 0;
assign detect_max[144][17] = (mid_1[1167:1160] > btm_0[1159:1152]) ? 1 : 0;
assign detect_max[144][18] = (mid_1[1167:1160] > btm_0[1167:1160]) ? 1 : 0;
assign detect_max[144][19] = (mid_1[1167:1160] > btm_0[1175:1168]) ? 1 : 0;
assign detect_max[144][20] = (mid_1[1167:1160] > btm_1[1159:1152]) ? 1 : 0;
assign detect_max[144][21] = (mid_1[1167:1160] > btm_1[1167:1160]) ? 1 : 0;
assign detect_max[144][22] = (mid_1[1167:1160] > btm_1[1175:1168]) ? 1 : 0;
assign detect_max[144][23] = (mid_1[1167:1160] > btm_2[1159:1152]) ? 1 : 0;
assign detect_max[144][24] = (mid_1[1167:1160] > btm_2[1167:1160]) ? 1 : 0;
assign detect_max[144][25] = (mid_1[1167:1160] > btm_2[1175:1168]) ? 1 : 0;

assign detect_max[145][0] = (mid_1[1175:1168] > top_0[1167:1160]) ? 1 : 0;
assign detect_max[145][1] = (mid_1[1175:1168] > top_0[1175:1168]) ? 1 : 0;
assign detect_max[145][2] = (mid_1[1175:1168] > top_0[1183:1176]) ? 1 : 0;
assign detect_max[145][3] = (mid_1[1175:1168] > top_1[1167:1160]) ? 1 : 0;
assign detect_max[145][4] = (mid_1[1175:1168] > top_1[1175:1168]) ? 1 : 0;
assign detect_max[145][5] = (mid_1[1175:1168] > top_1[1183:1176]) ? 1 : 0;
assign detect_max[145][6] = (mid_1[1175:1168] > top_2[1167:1160]) ? 1 : 0;
assign detect_max[145][7] = (mid_1[1175:1168] > top_2[1175:1168]) ? 1 : 0;
assign detect_max[145][8] = (mid_1[1175:1168] > top_2[1183:1176]) ? 1 : 0;
assign detect_max[145][9] = (mid_1[1175:1168] > mid_0[1167:1160]) ? 1 : 0;
assign detect_max[145][10] = (mid_1[1175:1168] > mid_0[1175:1168]) ? 1 : 0;
assign detect_max[145][11] = (mid_1[1175:1168] > mid_0[1183:1176]) ? 1 : 0;
assign detect_max[145][12] = (mid_1[1175:1168] > mid_1[1167:1160]) ? 1 : 0;
assign detect_max[145][13] = (mid_1[1175:1168] > mid_1[1183:1176]) ? 1 : 0;
assign detect_max[145][14] = (mid_1[1175:1168] > mid_2[1167:1160]) ? 1 : 0;
assign detect_max[145][15] = (mid_1[1175:1168] > mid_2[1175:1168]) ? 1 : 0;
assign detect_max[145][16] = (mid_1[1175:1168] > mid_2[1183:1176]) ? 1 : 0;
assign detect_max[145][17] = (mid_1[1175:1168] > btm_0[1167:1160]) ? 1 : 0;
assign detect_max[145][18] = (mid_1[1175:1168] > btm_0[1175:1168]) ? 1 : 0;
assign detect_max[145][19] = (mid_1[1175:1168] > btm_0[1183:1176]) ? 1 : 0;
assign detect_max[145][20] = (mid_1[1175:1168] > btm_1[1167:1160]) ? 1 : 0;
assign detect_max[145][21] = (mid_1[1175:1168] > btm_1[1175:1168]) ? 1 : 0;
assign detect_max[145][22] = (mid_1[1175:1168] > btm_1[1183:1176]) ? 1 : 0;
assign detect_max[145][23] = (mid_1[1175:1168] > btm_2[1167:1160]) ? 1 : 0;
assign detect_max[145][24] = (mid_1[1175:1168] > btm_2[1175:1168]) ? 1 : 0;
assign detect_max[145][25] = (mid_1[1175:1168] > btm_2[1183:1176]) ? 1 : 0;

assign detect_max[146][0] = (mid_1[1183:1176] > top_0[1175:1168]) ? 1 : 0;
assign detect_max[146][1] = (mid_1[1183:1176] > top_0[1183:1176]) ? 1 : 0;
assign detect_max[146][2] = (mid_1[1183:1176] > top_0[1191:1184]) ? 1 : 0;
assign detect_max[146][3] = (mid_1[1183:1176] > top_1[1175:1168]) ? 1 : 0;
assign detect_max[146][4] = (mid_1[1183:1176] > top_1[1183:1176]) ? 1 : 0;
assign detect_max[146][5] = (mid_1[1183:1176] > top_1[1191:1184]) ? 1 : 0;
assign detect_max[146][6] = (mid_1[1183:1176] > top_2[1175:1168]) ? 1 : 0;
assign detect_max[146][7] = (mid_1[1183:1176] > top_2[1183:1176]) ? 1 : 0;
assign detect_max[146][8] = (mid_1[1183:1176] > top_2[1191:1184]) ? 1 : 0;
assign detect_max[146][9] = (mid_1[1183:1176] > mid_0[1175:1168]) ? 1 : 0;
assign detect_max[146][10] = (mid_1[1183:1176] > mid_0[1183:1176]) ? 1 : 0;
assign detect_max[146][11] = (mid_1[1183:1176] > mid_0[1191:1184]) ? 1 : 0;
assign detect_max[146][12] = (mid_1[1183:1176] > mid_1[1175:1168]) ? 1 : 0;
assign detect_max[146][13] = (mid_1[1183:1176] > mid_1[1191:1184]) ? 1 : 0;
assign detect_max[146][14] = (mid_1[1183:1176] > mid_2[1175:1168]) ? 1 : 0;
assign detect_max[146][15] = (mid_1[1183:1176] > mid_2[1183:1176]) ? 1 : 0;
assign detect_max[146][16] = (mid_1[1183:1176] > mid_2[1191:1184]) ? 1 : 0;
assign detect_max[146][17] = (mid_1[1183:1176] > btm_0[1175:1168]) ? 1 : 0;
assign detect_max[146][18] = (mid_1[1183:1176] > btm_0[1183:1176]) ? 1 : 0;
assign detect_max[146][19] = (mid_1[1183:1176] > btm_0[1191:1184]) ? 1 : 0;
assign detect_max[146][20] = (mid_1[1183:1176] > btm_1[1175:1168]) ? 1 : 0;
assign detect_max[146][21] = (mid_1[1183:1176] > btm_1[1183:1176]) ? 1 : 0;
assign detect_max[146][22] = (mid_1[1183:1176] > btm_1[1191:1184]) ? 1 : 0;
assign detect_max[146][23] = (mid_1[1183:1176] > btm_2[1175:1168]) ? 1 : 0;
assign detect_max[146][24] = (mid_1[1183:1176] > btm_2[1183:1176]) ? 1 : 0;
assign detect_max[146][25] = (mid_1[1183:1176] > btm_2[1191:1184]) ? 1 : 0;

assign detect_max[147][0] = (mid_1[1191:1184] > top_0[1183:1176]) ? 1 : 0;
assign detect_max[147][1] = (mid_1[1191:1184] > top_0[1191:1184]) ? 1 : 0;
assign detect_max[147][2] = (mid_1[1191:1184] > top_0[1199:1192]) ? 1 : 0;
assign detect_max[147][3] = (mid_1[1191:1184] > top_1[1183:1176]) ? 1 : 0;
assign detect_max[147][4] = (mid_1[1191:1184] > top_1[1191:1184]) ? 1 : 0;
assign detect_max[147][5] = (mid_1[1191:1184] > top_1[1199:1192]) ? 1 : 0;
assign detect_max[147][6] = (mid_1[1191:1184] > top_2[1183:1176]) ? 1 : 0;
assign detect_max[147][7] = (mid_1[1191:1184] > top_2[1191:1184]) ? 1 : 0;
assign detect_max[147][8] = (mid_1[1191:1184] > top_2[1199:1192]) ? 1 : 0;
assign detect_max[147][9] = (mid_1[1191:1184] > mid_0[1183:1176]) ? 1 : 0;
assign detect_max[147][10] = (mid_1[1191:1184] > mid_0[1191:1184]) ? 1 : 0;
assign detect_max[147][11] = (mid_1[1191:1184] > mid_0[1199:1192]) ? 1 : 0;
assign detect_max[147][12] = (mid_1[1191:1184] > mid_1[1183:1176]) ? 1 : 0;
assign detect_max[147][13] = (mid_1[1191:1184] > mid_1[1199:1192]) ? 1 : 0;
assign detect_max[147][14] = (mid_1[1191:1184] > mid_2[1183:1176]) ? 1 : 0;
assign detect_max[147][15] = (mid_1[1191:1184] > mid_2[1191:1184]) ? 1 : 0;
assign detect_max[147][16] = (mid_1[1191:1184] > mid_2[1199:1192]) ? 1 : 0;
assign detect_max[147][17] = (mid_1[1191:1184] > btm_0[1183:1176]) ? 1 : 0;
assign detect_max[147][18] = (mid_1[1191:1184] > btm_0[1191:1184]) ? 1 : 0;
assign detect_max[147][19] = (mid_1[1191:1184] > btm_0[1199:1192]) ? 1 : 0;
assign detect_max[147][20] = (mid_1[1191:1184] > btm_1[1183:1176]) ? 1 : 0;
assign detect_max[147][21] = (mid_1[1191:1184] > btm_1[1191:1184]) ? 1 : 0;
assign detect_max[147][22] = (mid_1[1191:1184] > btm_1[1199:1192]) ? 1 : 0;
assign detect_max[147][23] = (mid_1[1191:1184] > btm_2[1183:1176]) ? 1 : 0;
assign detect_max[147][24] = (mid_1[1191:1184] > btm_2[1191:1184]) ? 1 : 0;
assign detect_max[147][25] = (mid_1[1191:1184] > btm_2[1199:1192]) ? 1 : 0;

assign detect_max[148][0] = (mid_1[1199:1192] > top_0[1191:1184]) ? 1 : 0;
assign detect_max[148][1] = (mid_1[1199:1192] > top_0[1199:1192]) ? 1 : 0;
assign detect_max[148][2] = (mid_1[1199:1192] > top_0[1207:1200]) ? 1 : 0;
assign detect_max[148][3] = (mid_1[1199:1192] > top_1[1191:1184]) ? 1 : 0;
assign detect_max[148][4] = (mid_1[1199:1192] > top_1[1199:1192]) ? 1 : 0;
assign detect_max[148][5] = (mid_1[1199:1192] > top_1[1207:1200]) ? 1 : 0;
assign detect_max[148][6] = (mid_1[1199:1192] > top_2[1191:1184]) ? 1 : 0;
assign detect_max[148][7] = (mid_1[1199:1192] > top_2[1199:1192]) ? 1 : 0;
assign detect_max[148][8] = (mid_1[1199:1192] > top_2[1207:1200]) ? 1 : 0;
assign detect_max[148][9] = (mid_1[1199:1192] > mid_0[1191:1184]) ? 1 : 0;
assign detect_max[148][10] = (mid_1[1199:1192] > mid_0[1199:1192]) ? 1 : 0;
assign detect_max[148][11] = (mid_1[1199:1192] > mid_0[1207:1200]) ? 1 : 0;
assign detect_max[148][12] = (mid_1[1199:1192] > mid_1[1191:1184]) ? 1 : 0;
assign detect_max[148][13] = (mid_1[1199:1192] > mid_1[1207:1200]) ? 1 : 0;
assign detect_max[148][14] = (mid_1[1199:1192] > mid_2[1191:1184]) ? 1 : 0;
assign detect_max[148][15] = (mid_1[1199:1192] > mid_2[1199:1192]) ? 1 : 0;
assign detect_max[148][16] = (mid_1[1199:1192] > mid_2[1207:1200]) ? 1 : 0;
assign detect_max[148][17] = (mid_1[1199:1192] > btm_0[1191:1184]) ? 1 : 0;
assign detect_max[148][18] = (mid_1[1199:1192] > btm_0[1199:1192]) ? 1 : 0;
assign detect_max[148][19] = (mid_1[1199:1192] > btm_0[1207:1200]) ? 1 : 0;
assign detect_max[148][20] = (mid_1[1199:1192] > btm_1[1191:1184]) ? 1 : 0;
assign detect_max[148][21] = (mid_1[1199:1192] > btm_1[1199:1192]) ? 1 : 0;
assign detect_max[148][22] = (mid_1[1199:1192] > btm_1[1207:1200]) ? 1 : 0;
assign detect_max[148][23] = (mid_1[1199:1192] > btm_2[1191:1184]) ? 1 : 0;
assign detect_max[148][24] = (mid_1[1199:1192] > btm_2[1199:1192]) ? 1 : 0;
assign detect_max[148][25] = (mid_1[1199:1192] > btm_2[1207:1200]) ? 1 : 0;

assign detect_max[149][0] = (mid_1[1207:1200] > top_0[1199:1192]) ? 1 : 0;
assign detect_max[149][1] = (mid_1[1207:1200] > top_0[1207:1200]) ? 1 : 0;
assign detect_max[149][2] = (mid_1[1207:1200] > top_0[1215:1208]) ? 1 : 0;
assign detect_max[149][3] = (mid_1[1207:1200] > top_1[1199:1192]) ? 1 : 0;
assign detect_max[149][4] = (mid_1[1207:1200] > top_1[1207:1200]) ? 1 : 0;
assign detect_max[149][5] = (mid_1[1207:1200] > top_1[1215:1208]) ? 1 : 0;
assign detect_max[149][6] = (mid_1[1207:1200] > top_2[1199:1192]) ? 1 : 0;
assign detect_max[149][7] = (mid_1[1207:1200] > top_2[1207:1200]) ? 1 : 0;
assign detect_max[149][8] = (mid_1[1207:1200] > top_2[1215:1208]) ? 1 : 0;
assign detect_max[149][9] = (mid_1[1207:1200] > mid_0[1199:1192]) ? 1 : 0;
assign detect_max[149][10] = (mid_1[1207:1200] > mid_0[1207:1200]) ? 1 : 0;
assign detect_max[149][11] = (mid_1[1207:1200] > mid_0[1215:1208]) ? 1 : 0;
assign detect_max[149][12] = (mid_1[1207:1200] > mid_1[1199:1192]) ? 1 : 0;
assign detect_max[149][13] = (mid_1[1207:1200] > mid_1[1215:1208]) ? 1 : 0;
assign detect_max[149][14] = (mid_1[1207:1200] > mid_2[1199:1192]) ? 1 : 0;
assign detect_max[149][15] = (mid_1[1207:1200] > mid_2[1207:1200]) ? 1 : 0;
assign detect_max[149][16] = (mid_1[1207:1200] > mid_2[1215:1208]) ? 1 : 0;
assign detect_max[149][17] = (mid_1[1207:1200] > btm_0[1199:1192]) ? 1 : 0;
assign detect_max[149][18] = (mid_1[1207:1200] > btm_0[1207:1200]) ? 1 : 0;
assign detect_max[149][19] = (mid_1[1207:1200] > btm_0[1215:1208]) ? 1 : 0;
assign detect_max[149][20] = (mid_1[1207:1200] > btm_1[1199:1192]) ? 1 : 0;
assign detect_max[149][21] = (mid_1[1207:1200] > btm_1[1207:1200]) ? 1 : 0;
assign detect_max[149][22] = (mid_1[1207:1200] > btm_1[1215:1208]) ? 1 : 0;
assign detect_max[149][23] = (mid_1[1207:1200] > btm_2[1199:1192]) ? 1 : 0;
assign detect_max[149][24] = (mid_1[1207:1200] > btm_2[1207:1200]) ? 1 : 0;
assign detect_max[149][25] = (mid_1[1207:1200] > btm_2[1215:1208]) ? 1 : 0;

assign detect_max[150][0] = (mid_1[1215:1208] > top_0[1207:1200]) ? 1 : 0;
assign detect_max[150][1] = (mid_1[1215:1208] > top_0[1215:1208]) ? 1 : 0;
assign detect_max[150][2] = (mid_1[1215:1208] > top_0[1223:1216]) ? 1 : 0;
assign detect_max[150][3] = (mid_1[1215:1208] > top_1[1207:1200]) ? 1 : 0;
assign detect_max[150][4] = (mid_1[1215:1208] > top_1[1215:1208]) ? 1 : 0;
assign detect_max[150][5] = (mid_1[1215:1208] > top_1[1223:1216]) ? 1 : 0;
assign detect_max[150][6] = (mid_1[1215:1208] > top_2[1207:1200]) ? 1 : 0;
assign detect_max[150][7] = (mid_1[1215:1208] > top_2[1215:1208]) ? 1 : 0;
assign detect_max[150][8] = (mid_1[1215:1208] > top_2[1223:1216]) ? 1 : 0;
assign detect_max[150][9] = (mid_1[1215:1208] > mid_0[1207:1200]) ? 1 : 0;
assign detect_max[150][10] = (mid_1[1215:1208] > mid_0[1215:1208]) ? 1 : 0;
assign detect_max[150][11] = (mid_1[1215:1208] > mid_0[1223:1216]) ? 1 : 0;
assign detect_max[150][12] = (mid_1[1215:1208] > mid_1[1207:1200]) ? 1 : 0;
assign detect_max[150][13] = (mid_1[1215:1208] > mid_1[1223:1216]) ? 1 : 0;
assign detect_max[150][14] = (mid_1[1215:1208] > mid_2[1207:1200]) ? 1 : 0;
assign detect_max[150][15] = (mid_1[1215:1208] > mid_2[1215:1208]) ? 1 : 0;
assign detect_max[150][16] = (mid_1[1215:1208] > mid_2[1223:1216]) ? 1 : 0;
assign detect_max[150][17] = (mid_1[1215:1208] > btm_0[1207:1200]) ? 1 : 0;
assign detect_max[150][18] = (mid_1[1215:1208] > btm_0[1215:1208]) ? 1 : 0;
assign detect_max[150][19] = (mid_1[1215:1208] > btm_0[1223:1216]) ? 1 : 0;
assign detect_max[150][20] = (mid_1[1215:1208] > btm_1[1207:1200]) ? 1 : 0;
assign detect_max[150][21] = (mid_1[1215:1208] > btm_1[1215:1208]) ? 1 : 0;
assign detect_max[150][22] = (mid_1[1215:1208] > btm_1[1223:1216]) ? 1 : 0;
assign detect_max[150][23] = (mid_1[1215:1208] > btm_2[1207:1200]) ? 1 : 0;
assign detect_max[150][24] = (mid_1[1215:1208] > btm_2[1215:1208]) ? 1 : 0;
assign detect_max[150][25] = (mid_1[1215:1208] > btm_2[1223:1216]) ? 1 : 0;

assign detect_max[151][0] = (mid_1[1223:1216] > top_0[1215:1208]) ? 1 : 0;
assign detect_max[151][1] = (mid_1[1223:1216] > top_0[1223:1216]) ? 1 : 0;
assign detect_max[151][2] = (mid_1[1223:1216] > top_0[1231:1224]) ? 1 : 0;
assign detect_max[151][3] = (mid_1[1223:1216] > top_1[1215:1208]) ? 1 : 0;
assign detect_max[151][4] = (mid_1[1223:1216] > top_1[1223:1216]) ? 1 : 0;
assign detect_max[151][5] = (mid_1[1223:1216] > top_1[1231:1224]) ? 1 : 0;
assign detect_max[151][6] = (mid_1[1223:1216] > top_2[1215:1208]) ? 1 : 0;
assign detect_max[151][7] = (mid_1[1223:1216] > top_2[1223:1216]) ? 1 : 0;
assign detect_max[151][8] = (mid_1[1223:1216] > top_2[1231:1224]) ? 1 : 0;
assign detect_max[151][9] = (mid_1[1223:1216] > mid_0[1215:1208]) ? 1 : 0;
assign detect_max[151][10] = (mid_1[1223:1216] > mid_0[1223:1216]) ? 1 : 0;
assign detect_max[151][11] = (mid_1[1223:1216] > mid_0[1231:1224]) ? 1 : 0;
assign detect_max[151][12] = (mid_1[1223:1216] > mid_1[1215:1208]) ? 1 : 0;
assign detect_max[151][13] = (mid_1[1223:1216] > mid_1[1231:1224]) ? 1 : 0;
assign detect_max[151][14] = (mid_1[1223:1216] > mid_2[1215:1208]) ? 1 : 0;
assign detect_max[151][15] = (mid_1[1223:1216] > mid_2[1223:1216]) ? 1 : 0;
assign detect_max[151][16] = (mid_1[1223:1216] > mid_2[1231:1224]) ? 1 : 0;
assign detect_max[151][17] = (mid_1[1223:1216] > btm_0[1215:1208]) ? 1 : 0;
assign detect_max[151][18] = (mid_1[1223:1216] > btm_0[1223:1216]) ? 1 : 0;
assign detect_max[151][19] = (mid_1[1223:1216] > btm_0[1231:1224]) ? 1 : 0;
assign detect_max[151][20] = (mid_1[1223:1216] > btm_1[1215:1208]) ? 1 : 0;
assign detect_max[151][21] = (mid_1[1223:1216] > btm_1[1223:1216]) ? 1 : 0;
assign detect_max[151][22] = (mid_1[1223:1216] > btm_1[1231:1224]) ? 1 : 0;
assign detect_max[151][23] = (mid_1[1223:1216] > btm_2[1215:1208]) ? 1 : 0;
assign detect_max[151][24] = (mid_1[1223:1216] > btm_2[1223:1216]) ? 1 : 0;
assign detect_max[151][25] = (mid_1[1223:1216] > btm_2[1231:1224]) ? 1 : 0;

assign detect_max[152][0] = (mid_1[1231:1224] > top_0[1223:1216]) ? 1 : 0;
assign detect_max[152][1] = (mid_1[1231:1224] > top_0[1231:1224]) ? 1 : 0;
assign detect_max[152][2] = (mid_1[1231:1224] > top_0[1239:1232]) ? 1 : 0;
assign detect_max[152][3] = (mid_1[1231:1224] > top_1[1223:1216]) ? 1 : 0;
assign detect_max[152][4] = (mid_1[1231:1224] > top_1[1231:1224]) ? 1 : 0;
assign detect_max[152][5] = (mid_1[1231:1224] > top_1[1239:1232]) ? 1 : 0;
assign detect_max[152][6] = (mid_1[1231:1224] > top_2[1223:1216]) ? 1 : 0;
assign detect_max[152][7] = (mid_1[1231:1224] > top_2[1231:1224]) ? 1 : 0;
assign detect_max[152][8] = (mid_1[1231:1224] > top_2[1239:1232]) ? 1 : 0;
assign detect_max[152][9] = (mid_1[1231:1224] > mid_0[1223:1216]) ? 1 : 0;
assign detect_max[152][10] = (mid_1[1231:1224] > mid_0[1231:1224]) ? 1 : 0;
assign detect_max[152][11] = (mid_1[1231:1224] > mid_0[1239:1232]) ? 1 : 0;
assign detect_max[152][12] = (mid_1[1231:1224] > mid_1[1223:1216]) ? 1 : 0;
assign detect_max[152][13] = (mid_1[1231:1224] > mid_1[1239:1232]) ? 1 : 0;
assign detect_max[152][14] = (mid_1[1231:1224] > mid_2[1223:1216]) ? 1 : 0;
assign detect_max[152][15] = (mid_1[1231:1224] > mid_2[1231:1224]) ? 1 : 0;
assign detect_max[152][16] = (mid_1[1231:1224] > mid_2[1239:1232]) ? 1 : 0;
assign detect_max[152][17] = (mid_1[1231:1224] > btm_0[1223:1216]) ? 1 : 0;
assign detect_max[152][18] = (mid_1[1231:1224] > btm_0[1231:1224]) ? 1 : 0;
assign detect_max[152][19] = (mid_1[1231:1224] > btm_0[1239:1232]) ? 1 : 0;
assign detect_max[152][20] = (mid_1[1231:1224] > btm_1[1223:1216]) ? 1 : 0;
assign detect_max[152][21] = (mid_1[1231:1224] > btm_1[1231:1224]) ? 1 : 0;
assign detect_max[152][22] = (mid_1[1231:1224] > btm_1[1239:1232]) ? 1 : 0;
assign detect_max[152][23] = (mid_1[1231:1224] > btm_2[1223:1216]) ? 1 : 0;
assign detect_max[152][24] = (mid_1[1231:1224] > btm_2[1231:1224]) ? 1 : 0;
assign detect_max[152][25] = (mid_1[1231:1224] > btm_2[1239:1232]) ? 1 : 0;

assign detect_max[153][0] = (mid_1[1239:1232] > top_0[1231:1224]) ? 1 : 0;
assign detect_max[153][1] = (mid_1[1239:1232] > top_0[1239:1232]) ? 1 : 0;
assign detect_max[153][2] = (mid_1[1239:1232] > top_0[1247:1240]) ? 1 : 0;
assign detect_max[153][3] = (mid_1[1239:1232] > top_1[1231:1224]) ? 1 : 0;
assign detect_max[153][4] = (mid_1[1239:1232] > top_1[1239:1232]) ? 1 : 0;
assign detect_max[153][5] = (mid_1[1239:1232] > top_1[1247:1240]) ? 1 : 0;
assign detect_max[153][6] = (mid_1[1239:1232] > top_2[1231:1224]) ? 1 : 0;
assign detect_max[153][7] = (mid_1[1239:1232] > top_2[1239:1232]) ? 1 : 0;
assign detect_max[153][8] = (mid_1[1239:1232] > top_2[1247:1240]) ? 1 : 0;
assign detect_max[153][9] = (mid_1[1239:1232] > mid_0[1231:1224]) ? 1 : 0;
assign detect_max[153][10] = (mid_1[1239:1232] > mid_0[1239:1232]) ? 1 : 0;
assign detect_max[153][11] = (mid_1[1239:1232] > mid_0[1247:1240]) ? 1 : 0;
assign detect_max[153][12] = (mid_1[1239:1232] > mid_1[1231:1224]) ? 1 : 0;
assign detect_max[153][13] = (mid_1[1239:1232] > mid_1[1247:1240]) ? 1 : 0;
assign detect_max[153][14] = (mid_1[1239:1232] > mid_2[1231:1224]) ? 1 : 0;
assign detect_max[153][15] = (mid_1[1239:1232] > mid_2[1239:1232]) ? 1 : 0;
assign detect_max[153][16] = (mid_1[1239:1232] > mid_2[1247:1240]) ? 1 : 0;
assign detect_max[153][17] = (mid_1[1239:1232] > btm_0[1231:1224]) ? 1 : 0;
assign detect_max[153][18] = (mid_1[1239:1232] > btm_0[1239:1232]) ? 1 : 0;
assign detect_max[153][19] = (mid_1[1239:1232] > btm_0[1247:1240]) ? 1 : 0;
assign detect_max[153][20] = (mid_1[1239:1232] > btm_1[1231:1224]) ? 1 : 0;
assign detect_max[153][21] = (mid_1[1239:1232] > btm_1[1239:1232]) ? 1 : 0;
assign detect_max[153][22] = (mid_1[1239:1232] > btm_1[1247:1240]) ? 1 : 0;
assign detect_max[153][23] = (mid_1[1239:1232] > btm_2[1231:1224]) ? 1 : 0;
assign detect_max[153][24] = (mid_1[1239:1232] > btm_2[1239:1232]) ? 1 : 0;
assign detect_max[153][25] = (mid_1[1239:1232] > btm_2[1247:1240]) ? 1 : 0;

assign detect_max[154][0] = (mid_1[1247:1240] > top_0[1239:1232]) ? 1 : 0;
assign detect_max[154][1] = (mid_1[1247:1240] > top_0[1247:1240]) ? 1 : 0;
assign detect_max[154][2] = (mid_1[1247:1240] > top_0[1255:1248]) ? 1 : 0;
assign detect_max[154][3] = (mid_1[1247:1240] > top_1[1239:1232]) ? 1 : 0;
assign detect_max[154][4] = (mid_1[1247:1240] > top_1[1247:1240]) ? 1 : 0;
assign detect_max[154][5] = (mid_1[1247:1240] > top_1[1255:1248]) ? 1 : 0;
assign detect_max[154][6] = (mid_1[1247:1240] > top_2[1239:1232]) ? 1 : 0;
assign detect_max[154][7] = (mid_1[1247:1240] > top_2[1247:1240]) ? 1 : 0;
assign detect_max[154][8] = (mid_1[1247:1240] > top_2[1255:1248]) ? 1 : 0;
assign detect_max[154][9] = (mid_1[1247:1240] > mid_0[1239:1232]) ? 1 : 0;
assign detect_max[154][10] = (mid_1[1247:1240] > mid_0[1247:1240]) ? 1 : 0;
assign detect_max[154][11] = (mid_1[1247:1240] > mid_0[1255:1248]) ? 1 : 0;
assign detect_max[154][12] = (mid_1[1247:1240] > mid_1[1239:1232]) ? 1 : 0;
assign detect_max[154][13] = (mid_1[1247:1240] > mid_1[1255:1248]) ? 1 : 0;
assign detect_max[154][14] = (mid_1[1247:1240] > mid_2[1239:1232]) ? 1 : 0;
assign detect_max[154][15] = (mid_1[1247:1240] > mid_2[1247:1240]) ? 1 : 0;
assign detect_max[154][16] = (mid_1[1247:1240] > mid_2[1255:1248]) ? 1 : 0;
assign detect_max[154][17] = (mid_1[1247:1240] > btm_0[1239:1232]) ? 1 : 0;
assign detect_max[154][18] = (mid_1[1247:1240] > btm_0[1247:1240]) ? 1 : 0;
assign detect_max[154][19] = (mid_1[1247:1240] > btm_0[1255:1248]) ? 1 : 0;
assign detect_max[154][20] = (mid_1[1247:1240] > btm_1[1239:1232]) ? 1 : 0;
assign detect_max[154][21] = (mid_1[1247:1240] > btm_1[1247:1240]) ? 1 : 0;
assign detect_max[154][22] = (mid_1[1247:1240] > btm_1[1255:1248]) ? 1 : 0;
assign detect_max[154][23] = (mid_1[1247:1240] > btm_2[1239:1232]) ? 1 : 0;
assign detect_max[154][24] = (mid_1[1247:1240] > btm_2[1247:1240]) ? 1 : 0;
assign detect_max[154][25] = (mid_1[1247:1240] > btm_2[1255:1248]) ? 1 : 0;

assign detect_max[155][0] = (mid_1[1255:1248] > top_0[1247:1240]) ? 1 : 0;
assign detect_max[155][1] = (mid_1[1255:1248] > top_0[1255:1248]) ? 1 : 0;
assign detect_max[155][2] = (mid_1[1255:1248] > top_0[1263:1256]) ? 1 : 0;
assign detect_max[155][3] = (mid_1[1255:1248] > top_1[1247:1240]) ? 1 : 0;
assign detect_max[155][4] = (mid_1[1255:1248] > top_1[1255:1248]) ? 1 : 0;
assign detect_max[155][5] = (mid_1[1255:1248] > top_1[1263:1256]) ? 1 : 0;
assign detect_max[155][6] = (mid_1[1255:1248] > top_2[1247:1240]) ? 1 : 0;
assign detect_max[155][7] = (mid_1[1255:1248] > top_2[1255:1248]) ? 1 : 0;
assign detect_max[155][8] = (mid_1[1255:1248] > top_2[1263:1256]) ? 1 : 0;
assign detect_max[155][9] = (mid_1[1255:1248] > mid_0[1247:1240]) ? 1 : 0;
assign detect_max[155][10] = (mid_1[1255:1248] > mid_0[1255:1248]) ? 1 : 0;
assign detect_max[155][11] = (mid_1[1255:1248] > mid_0[1263:1256]) ? 1 : 0;
assign detect_max[155][12] = (mid_1[1255:1248] > mid_1[1247:1240]) ? 1 : 0;
assign detect_max[155][13] = (mid_1[1255:1248] > mid_1[1263:1256]) ? 1 : 0;
assign detect_max[155][14] = (mid_1[1255:1248] > mid_2[1247:1240]) ? 1 : 0;
assign detect_max[155][15] = (mid_1[1255:1248] > mid_2[1255:1248]) ? 1 : 0;
assign detect_max[155][16] = (mid_1[1255:1248] > mid_2[1263:1256]) ? 1 : 0;
assign detect_max[155][17] = (mid_1[1255:1248] > btm_0[1247:1240]) ? 1 : 0;
assign detect_max[155][18] = (mid_1[1255:1248] > btm_0[1255:1248]) ? 1 : 0;
assign detect_max[155][19] = (mid_1[1255:1248] > btm_0[1263:1256]) ? 1 : 0;
assign detect_max[155][20] = (mid_1[1255:1248] > btm_1[1247:1240]) ? 1 : 0;
assign detect_max[155][21] = (mid_1[1255:1248] > btm_1[1255:1248]) ? 1 : 0;
assign detect_max[155][22] = (mid_1[1255:1248] > btm_1[1263:1256]) ? 1 : 0;
assign detect_max[155][23] = (mid_1[1255:1248] > btm_2[1247:1240]) ? 1 : 0;
assign detect_max[155][24] = (mid_1[1255:1248] > btm_2[1255:1248]) ? 1 : 0;
assign detect_max[155][25] = (mid_1[1255:1248] > btm_2[1263:1256]) ? 1 : 0;

assign detect_max[156][0] = (mid_1[1263:1256] > top_0[1255:1248]) ? 1 : 0;
assign detect_max[156][1] = (mid_1[1263:1256] > top_0[1263:1256]) ? 1 : 0;
assign detect_max[156][2] = (mid_1[1263:1256] > top_0[1271:1264]) ? 1 : 0;
assign detect_max[156][3] = (mid_1[1263:1256] > top_1[1255:1248]) ? 1 : 0;
assign detect_max[156][4] = (mid_1[1263:1256] > top_1[1263:1256]) ? 1 : 0;
assign detect_max[156][5] = (mid_1[1263:1256] > top_1[1271:1264]) ? 1 : 0;
assign detect_max[156][6] = (mid_1[1263:1256] > top_2[1255:1248]) ? 1 : 0;
assign detect_max[156][7] = (mid_1[1263:1256] > top_2[1263:1256]) ? 1 : 0;
assign detect_max[156][8] = (mid_1[1263:1256] > top_2[1271:1264]) ? 1 : 0;
assign detect_max[156][9] = (mid_1[1263:1256] > mid_0[1255:1248]) ? 1 : 0;
assign detect_max[156][10] = (mid_1[1263:1256] > mid_0[1263:1256]) ? 1 : 0;
assign detect_max[156][11] = (mid_1[1263:1256] > mid_0[1271:1264]) ? 1 : 0;
assign detect_max[156][12] = (mid_1[1263:1256] > mid_1[1255:1248]) ? 1 : 0;
assign detect_max[156][13] = (mid_1[1263:1256] > mid_1[1271:1264]) ? 1 : 0;
assign detect_max[156][14] = (mid_1[1263:1256] > mid_2[1255:1248]) ? 1 : 0;
assign detect_max[156][15] = (mid_1[1263:1256] > mid_2[1263:1256]) ? 1 : 0;
assign detect_max[156][16] = (mid_1[1263:1256] > mid_2[1271:1264]) ? 1 : 0;
assign detect_max[156][17] = (mid_1[1263:1256] > btm_0[1255:1248]) ? 1 : 0;
assign detect_max[156][18] = (mid_1[1263:1256] > btm_0[1263:1256]) ? 1 : 0;
assign detect_max[156][19] = (mid_1[1263:1256] > btm_0[1271:1264]) ? 1 : 0;
assign detect_max[156][20] = (mid_1[1263:1256] > btm_1[1255:1248]) ? 1 : 0;
assign detect_max[156][21] = (mid_1[1263:1256] > btm_1[1263:1256]) ? 1 : 0;
assign detect_max[156][22] = (mid_1[1263:1256] > btm_1[1271:1264]) ? 1 : 0;
assign detect_max[156][23] = (mid_1[1263:1256] > btm_2[1255:1248]) ? 1 : 0;
assign detect_max[156][24] = (mid_1[1263:1256] > btm_2[1263:1256]) ? 1 : 0;
assign detect_max[156][25] = (mid_1[1263:1256] > btm_2[1271:1264]) ? 1 : 0;

assign detect_max[157][0] = (mid_1[1271:1264] > top_0[1263:1256]) ? 1 : 0;
assign detect_max[157][1] = (mid_1[1271:1264] > top_0[1271:1264]) ? 1 : 0;
assign detect_max[157][2] = (mid_1[1271:1264] > top_0[1279:1272]) ? 1 : 0;
assign detect_max[157][3] = (mid_1[1271:1264] > top_1[1263:1256]) ? 1 : 0;
assign detect_max[157][4] = (mid_1[1271:1264] > top_1[1271:1264]) ? 1 : 0;
assign detect_max[157][5] = (mid_1[1271:1264] > top_1[1279:1272]) ? 1 : 0;
assign detect_max[157][6] = (mid_1[1271:1264] > top_2[1263:1256]) ? 1 : 0;
assign detect_max[157][7] = (mid_1[1271:1264] > top_2[1271:1264]) ? 1 : 0;
assign detect_max[157][8] = (mid_1[1271:1264] > top_2[1279:1272]) ? 1 : 0;
assign detect_max[157][9] = (mid_1[1271:1264] > mid_0[1263:1256]) ? 1 : 0;
assign detect_max[157][10] = (mid_1[1271:1264] > mid_0[1271:1264]) ? 1 : 0;
assign detect_max[157][11] = (mid_1[1271:1264] > mid_0[1279:1272]) ? 1 : 0;
assign detect_max[157][12] = (mid_1[1271:1264] > mid_1[1263:1256]) ? 1 : 0;
assign detect_max[157][13] = (mid_1[1271:1264] > mid_1[1279:1272]) ? 1 : 0;
assign detect_max[157][14] = (mid_1[1271:1264] > mid_2[1263:1256]) ? 1 : 0;
assign detect_max[157][15] = (mid_1[1271:1264] > mid_2[1271:1264]) ? 1 : 0;
assign detect_max[157][16] = (mid_1[1271:1264] > mid_2[1279:1272]) ? 1 : 0;
assign detect_max[157][17] = (mid_1[1271:1264] > btm_0[1263:1256]) ? 1 : 0;
assign detect_max[157][18] = (mid_1[1271:1264] > btm_0[1271:1264]) ? 1 : 0;
assign detect_max[157][19] = (mid_1[1271:1264] > btm_0[1279:1272]) ? 1 : 0;
assign detect_max[157][20] = (mid_1[1271:1264] > btm_1[1263:1256]) ? 1 : 0;
assign detect_max[157][21] = (mid_1[1271:1264] > btm_1[1271:1264]) ? 1 : 0;
assign detect_max[157][22] = (mid_1[1271:1264] > btm_1[1279:1272]) ? 1 : 0;
assign detect_max[157][23] = (mid_1[1271:1264] > btm_2[1263:1256]) ? 1 : 0;
assign detect_max[157][24] = (mid_1[1271:1264] > btm_2[1271:1264]) ? 1 : 0;
assign detect_max[157][25] = (mid_1[1271:1264] > btm_2[1279:1272]) ? 1 : 0;

assign detect_max[158][0] = (mid_1[1279:1272] > top_0[1271:1264]) ? 1 : 0;
assign detect_max[158][1] = (mid_1[1279:1272] > top_0[1279:1272]) ? 1 : 0;
assign detect_max[158][2] = (mid_1[1279:1272] > top_0[1287:1280]) ? 1 : 0;
assign detect_max[158][3] = (mid_1[1279:1272] > top_1[1271:1264]) ? 1 : 0;
assign detect_max[158][4] = (mid_1[1279:1272] > top_1[1279:1272]) ? 1 : 0;
assign detect_max[158][5] = (mid_1[1279:1272] > top_1[1287:1280]) ? 1 : 0;
assign detect_max[158][6] = (mid_1[1279:1272] > top_2[1271:1264]) ? 1 : 0;
assign detect_max[158][7] = (mid_1[1279:1272] > top_2[1279:1272]) ? 1 : 0;
assign detect_max[158][8] = (mid_1[1279:1272] > top_2[1287:1280]) ? 1 : 0;
assign detect_max[158][9] = (mid_1[1279:1272] > mid_0[1271:1264]) ? 1 : 0;
assign detect_max[158][10] = (mid_1[1279:1272] > mid_0[1279:1272]) ? 1 : 0;
assign detect_max[158][11] = (mid_1[1279:1272] > mid_0[1287:1280]) ? 1 : 0;
assign detect_max[158][12] = (mid_1[1279:1272] > mid_1[1271:1264]) ? 1 : 0;
assign detect_max[158][13] = (mid_1[1279:1272] > mid_1[1287:1280]) ? 1 : 0;
assign detect_max[158][14] = (mid_1[1279:1272] > mid_2[1271:1264]) ? 1 : 0;
assign detect_max[158][15] = (mid_1[1279:1272] > mid_2[1279:1272]) ? 1 : 0;
assign detect_max[158][16] = (mid_1[1279:1272] > mid_2[1287:1280]) ? 1 : 0;
assign detect_max[158][17] = (mid_1[1279:1272] > btm_0[1271:1264]) ? 1 : 0;
assign detect_max[158][18] = (mid_1[1279:1272] > btm_0[1279:1272]) ? 1 : 0;
assign detect_max[158][19] = (mid_1[1279:1272] > btm_0[1287:1280]) ? 1 : 0;
assign detect_max[158][20] = (mid_1[1279:1272] > btm_1[1271:1264]) ? 1 : 0;
assign detect_max[158][21] = (mid_1[1279:1272] > btm_1[1279:1272]) ? 1 : 0;
assign detect_max[158][22] = (mid_1[1279:1272] > btm_1[1287:1280]) ? 1 : 0;
assign detect_max[158][23] = (mid_1[1279:1272] > btm_2[1271:1264]) ? 1 : 0;
assign detect_max[158][24] = (mid_1[1279:1272] > btm_2[1279:1272]) ? 1 : 0;
assign detect_max[158][25] = (mid_1[1279:1272] > btm_2[1287:1280]) ? 1 : 0;

assign detect_max[159][0] = (mid_1[1287:1280] > top_0[1279:1272]) ? 1 : 0;
assign detect_max[159][1] = (mid_1[1287:1280] > top_0[1287:1280]) ? 1 : 0;
assign detect_max[159][2] = (mid_1[1287:1280] > top_0[1295:1288]) ? 1 : 0;
assign detect_max[159][3] = (mid_1[1287:1280] > top_1[1279:1272]) ? 1 : 0;
assign detect_max[159][4] = (mid_1[1287:1280] > top_1[1287:1280]) ? 1 : 0;
assign detect_max[159][5] = (mid_1[1287:1280] > top_1[1295:1288]) ? 1 : 0;
assign detect_max[159][6] = (mid_1[1287:1280] > top_2[1279:1272]) ? 1 : 0;
assign detect_max[159][7] = (mid_1[1287:1280] > top_2[1287:1280]) ? 1 : 0;
assign detect_max[159][8] = (mid_1[1287:1280] > top_2[1295:1288]) ? 1 : 0;
assign detect_max[159][9] = (mid_1[1287:1280] > mid_0[1279:1272]) ? 1 : 0;
assign detect_max[159][10] = (mid_1[1287:1280] > mid_0[1287:1280]) ? 1 : 0;
assign detect_max[159][11] = (mid_1[1287:1280] > mid_0[1295:1288]) ? 1 : 0;
assign detect_max[159][12] = (mid_1[1287:1280] > mid_1[1279:1272]) ? 1 : 0;
assign detect_max[159][13] = (mid_1[1287:1280] > mid_1[1295:1288]) ? 1 : 0;
assign detect_max[159][14] = (mid_1[1287:1280] > mid_2[1279:1272]) ? 1 : 0;
assign detect_max[159][15] = (mid_1[1287:1280] > mid_2[1287:1280]) ? 1 : 0;
assign detect_max[159][16] = (mid_1[1287:1280] > mid_2[1295:1288]) ? 1 : 0;
assign detect_max[159][17] = (mid_1[1287:1280] > btm_0[1279:1272]) ? 1 : 0;
assign detect_max[159][18] = (mid_1[1287:1280] > btm_0[1287:1280]) ? 1 : 0;
assign detect_max[159][19] = (mid_1[1287:1280] > btm_0[1295:1288]) ? 1 : 0;
assign detect_max[159][20] = (mid_1[1287:1280] > btm_1[1279:1272]) ? 1 : 0;
assign detect_max[159][21] = (mid_1[1287:1280] > btm_1[1287:1280]) ? 1 : 0;
assign detect_max[159][22] = (mid_1[1287:1280] > btm_1[1295:1288]) ? 1 : 0;
assign detect_max[159][23] = (mid_1[1287:1280] > btm_2[1279:1272]) ? 1 : 0;
assign detect_max[159][24] = (mid_1[1287:1280] > btm_2[1287:1280]) ? 1 : 0;
assign detect_max[159][25] = (mid_1[1287:1280] > btm_2[1295:1288]) ? 1 : 0;

assign detect_max[160][0] = (mid_1[1295:1288] > top_0[1287:1280]) ? 1 : 0;
assign detect_max[160][1] = (mid_1[1295:1288] > top_0[1295:1288]) ? 1 : 0;
assign detect_max[160][2] = (mid_1[1295:1288] > top_0[1303:1296]) ? 1 : 0;
assign detect_max[160][3] = (mid_1[1295:1288] > top_1[1287:1280]) ? 1 : 0;
assign detect_max[160][4] = (mid_1[1295:1288] > top_1[1295:1288]) ? 1 : 0;
assign detect_max[160][5] = (mid_1[1295:1288] > top_1[1303:1296]) ? 1 : 0;
assign detect_max[160][6] = (mid_1[1295:1288] > top_2[1287:1280]) ? 1 : 0;
assign detect_max[160][7] = (mid_1[1295:1288] > top_2[1295:1288]) ? 1 : 0;
assign detect_max[160][8] = (mid_1[1295:1288] > top_2[1303:1296]) ? 1 : 0;
assign detect_max[160][9] = (mid_1[1295:1288] > mid_0[1287:1280]) ? 1 : 0;
assign detect_max[160][10] = (mid_1[1295:1288] > mid_0[1295:1288]) ? 1 : 0;
assign detect_max[160][11] = (mid_1[1295:1288] > mid_0[1303:1296]) ? 1 : 0;
assign detect_max[160][12] = (mid_1[1295:1288] > mid_1[1287:1280]) ? 1 : 0;
assign detect_max[160][13] = (mid_1[1295:1288] > mid_1[1303:1296]) ? 1 : 0;
assign detect_max[160][14] = (mid_1[1295:1288] > mid_2[1287:1280]) ? 1 : 0;
assign detect_max[160][15] = (mid_1[1295:1288] > mid_2[1295:1288]) ? 1 : 0;
assign detect_max[160][16] = (mid_1[1295:1288] > mid_2[1303:1296]) ? 1 : 0;
assign detect_max[160][17] = (mid_1[1295:1288] > btm_0[1287:1280]) ? 1 : 0;
assign detect_max[160][18] = (mid_1[1295:1288] > btm_0[1295:1288]) ? 1 : 0;
assign detect_max[160][19] = (mid_1[1295:1288] > btm_0[1303:1296]) ? 1 : 0;
assign detect_max[160][20] = (mid_1[1295:1288] > btm_1[1287:1280]) ? 1 : 0;
assign detect_max[160][21] = (mid_1[1295:1288] > btm_1[1295:1288]) ? 1 : 0;
assign detect_max[160][22] = (mid_1[1295:1288] > btm_1[1303:1296]) ? 1 : 0;
assign detect_max[160][23] = (mid_1[1295:1288] > btm_2[1287:1280]) ? 1 : 0;
assign detect_max[160][24] = (mid_1[1295:1288] > btm_2[1295:1288]) ? 1 : 0;
assign detect_max[160][25] = (mid_1[1295:1288] > btm_2[1303:1296]) ? 1 : 0;

assign detect_max[161][0] = (mid_1[1303:1296] > top_0[1295:1288]) ? 1 : 0;
assign detect_max[161][1] = (mid_1[1303:1296] > top_0[1303:1296]) ? 1 : 0;
assign detect_max[161][2] = (mid_1[1303:1296] > top_0[1311:1304]) ? 1 : 0;
assign detect_max[161][3] = (mid_1[1303:1296] > top_1[1295:1288]) ? 1 : 0;
assign detect_max[161][4] = (mid_1[1303:1296] > top_1[1303:1296]) ? 1 : 0;
assign detect_max[161][5] = (mid_1[1303:1296] > top_1[1311:1304]) ? 1 : 0;
assign detect_max[161][6] = (mid_1[1303:1296] > top_2[1295:1288]) ? 1 : 0;
assign detect_max[161][7] = (mid_1[1303:1296] > top_2[1303:1296]) ? 1 : 0;
assign detect_max[161][8] = (mid_1[1303:1296] > top_2[1311:1304]) ? 1 : 0;
assign detect_max[161][9] = (mid_1[1303:1296] > mid_0[1295:1288]) ? 1 : 0;
assign detect_max[161][10] = (mid_1[1303:1296] > mid_0[1303:1296]) ? 1 : 0;
assign detect_max[161][11] = (mid_1[1303:1296] > mid_0[1311:1304]) ? 1 : 0;
assign detect_max[161][12] = (mid_1[1303:1296] > mid_1[1295:1288]) ? 1 : 0;
assign detect_max[161][13] = (mid_1[1303:1296] > mid_1[1311:1304]) ? 1 : 0;
assign detect_max[161][14] = (mid_1[1303:1296] > mid_2[1295:1288]) ? 1 : 0;
assign detect_max[161][15] = (mid_1[1303:1296] > mid_2[1303:1296]) ? 1 : 0;
assign detect_max[161][16] = (mid_1[1303:1296] > mid_2[1311:1304]) ? 1 : 0;
assign detect_max[161][17] = (mid_1[1303:1296] > btm_0[1295:1288]) ? 1 : 0;
assign detect_max[161][18] = (mid_1[1303:1296] > btm_0[1303:1296]) ? 1 : 0;
assign detect_max[161][19] = (mid_1[1303:1296] > btm_0[1311:1304]) ? 1 : 0;
assign detect_max[161][20] = (mid_1[1303:1296] > btm_1[1295:1288]) ? 1 : 0;
assign detect_max[161][21] = (mid_1[1303:1296] > btm_1[1303:1296]) ? 1 : 0;
assign detect_max[161][22] = (mid_1[1303:1296] > btm_1[1311:1304]) ? 1 : 0;
assign detect_max[161][23] = (mid_1[1303:1296] > btm_2[1295:1288]) ? 1 : 0;
assign detect_max[161][24] = (mid_1[1303:1296] > btm_2[1303:1296]) ? 1 : 0;
assign detect_max[161][25] = (mid_1[1303:1296] > btm_2[1311:1304]) ? 1 : 0;

assign detect_max[162][0] = (mid_1[1311:1304] > top_0[1303:1296]) ? 1 : 0;
assign detect_max[162][1] = (mid_1[1311:1304] > top_0[1311:1304]) ? 1 : 0;
assign detect_max[162][2] = (mid_1[1311:1304] > top_0[1319:1312]) ? 1 : 0;
assign detect_max[162][3] = (mid_1[1311:1304] > top_1[1303:1296]) ? 1 : 0;
assign detect_max[162][4] = (mid_1[1311:1304] > top_1[1311:1304]) ? 1 : 0;
assign detect_max[162][5] = (mid_1[1311:1304] > top_1[1319:1312]) ? 1 : 0;
assign detect_max[162][6] = (mid_1[1311:1304] > top_2[1303:1296]) ? 1 : 0;
assign detect_max[162][7] = (mid_1[1311:1304] > top_2[1311:1304]) ? 1 : 0;
assign detect_max[162][8] = (mid_1[1311:1304] > top_2[1319:1312]) ? 1 : 0;
assign detect_max[162][9] = (mid_1[1311:1304] > mid_0[1303:1296]) ? 1 : 0;
assign detect_max[162][10] = (mid_1[1311:1304] > mid_0[1311:1304]) ? 1 : 0;
assign detect_max[162][11] = (mid_1[1311:1304] > mid_0[1319:1312]) ? 1 : 0;
assign detect_max[162][12] = (mid_1[1311:1304] > mid_1[1303:1296]) ? 1 : 0;
assign detect_max[162][13] = (mid_1[1311:1304] > mid_1[1319:1312]) ? 1 : 0;
assign detect_max[162][14] = (mid_1[1311:1304] > mid_2[1303:1296]) ? 1 : 0;
assign detect_max[162][15] = (mid_1[1311:1304] > mid_2[1311:1304]) ? 1 : 0;
assign detect_max[162][16] = (mid_1[1311:1304] > mid_2[1319:1312]) ? 1 : 0;
assign detect_max[162][17] = (mid_1[1311:1304] > btm_0[1303:1296]) ? 1 : 0;
assign detect_max[162][18] = (mid_1[1311:1304] > btm_0[1311:1304]) ? 1 : 0;
assign detect_max[162][19] = (mid_1[1311:1304] > btm_0[1319:1312]) ? 1 : 0;
assign detect_max[162][20] = (mid_1[1311:1304] > btm_1[1303:1296]) ? 1 : 0;
assign detect_max[162][21] = (mid_1[1311:1304] > btm_1[1311:1304]) ? 1 : 0;
assign detect_max[162][22] = (mid_1[1311:1304] > btm_1[1319:1312]) ? 1 : 0;
assign detect_max[162][23] = (mid_1[1311:1304] > btm_2[1303:1296]) ? 1 : 0;
assign detect_max[162][24] = (mid_1[1311:1304] > btm_2[1311:1304]) ? 1 : 0;
assign detect_max[162][25] = (mid_1[1311:1304] > btm_2[1319:1312]) ? 1 : 0;

assign detect_max[163][0] = (mid_1[1319:1312] > top_0[1311:1304]) ? 1 : 0;
assign detect_max[163][1] = (mid_1[1319:1312] > top_0[1319:1312]) ? 1 : 0;
assign detect_max[163][2] = (mid_1[1319:1312] > top_0[1327:1320]) ? 1 : 0;
assign detect_max[163][3] = (mid_1[1319:1312] > top_1[1311:1304]) ? 1 : 0;
assign detect_max[163][4] = (mid_1[1319:1312] > top_1[1319:1312]) ? 1 : 0;
assign detect_max[163][5] = (mid_1[1319:1312] > top_1[1327:1320]) ? 1 : 0;
assign detect_max[163][6] = (mid_1[1319:1312] > top_2[1311:1304]) ? 1 : 0;
assign detect_max[163][7] = (mid_1[1319:1312] > top_2[1319:1312]) ? 1 : 0;
assign detect_max[163][8] = (mid_1[1319:1312] > top_2[1327:1320]) ? 1 : 0;
assign detect_max[163][9] = (mid_1[1319:1312] > mid_0[1311:1304]) ? 1 : 0;
assign detect_max[163][10] = (mid_1[1319:1312] > mid_0[1319:1312]) ? 1 : 0;
assign detect_max[163][11] = (mid_1[1319:1312] > mid_0[1327:1320]) ? 1 : 0;
assign detect_max[163][12] = (mid_1[1319:1312] > mid_1[1311:1304]) ? 1 : 0;
assign detect_max[163][13] = (mid_1[1319:1312] > mid_1[1327:1320]) ? 1 : 0;
assign detect_max[163][14] = (mid_1[1319:1312] > mid_2[1311:1304]) ? 1 : 0;
assign detect_max[163][15] = (mid_1[1319:1312] > mid_2[1319:1312]) ? 1 : 0;
assign detect_max[163][16] = (mid_1[1319:1312] > mid_2[1327:1320]) ? 1 : 0;
assign detect_max[163][17] = (mid_1[1319:1312] > btm_0[1311:1304]) ? 1 : 0;
assign detect_max[163][18] = (mid_1[1319:1312] > btm_0[1319:1312]) ? 1 : 0;
assign detect_max[163][19] = (mid_1[1319:1312] > btm_0[1327:1320]) ? 1 : 0;
assign detect_max[163][20] = (mid_1[1319:1312] > btm_1[1311:1304]) ? 1 : 0;
assign detect_max[163][21] = (mid_1[1319:1312] > btm_1[1319:1312]) ? 1 : 0;
assign detect_max[163][22] = (mid_1[1319:1312] > btm_1[1327:1320]) ? 1 : 0;
assign detect_max[163][23] = (mid_1[1319:1312] > btm_2[1311:1304]) ? 1 : 0;
assign detect_max[163][24] = (mid_1[1319:1312] > btm_2[1319:1312]) ? 1 : 0;
assign detect_max[163][25] = (mid_1[1319:1312] > btm_2[1327:1320]) ? 1 : 0;

assign detect_max[164][0] = (mid_1[1327:1320] > top_0[1319:1312]) ? 1 : 0;
assign detect_max[164][1] = (mid_1[1327:1320] > top_0[1327:1320]) ? 1 : 0;
assign detect_max[164][2] = (mid_1[1327:1320] > top_0[1335:1328]) ? 1 : 0;
assign detect_max[164][3] = (mid_1[1327:1320] > top_1[1319:1312]) ? 1 : 0;
assign detect_max[164][4] = (mid_1[1327:1320] > top_1[1327:1320]) ? 1 : 0;
assign detect_max[164][5] = (mid_1[1327:1320] > top_1[1335:1328]) ? 1 : 0;
assign detect_max[164][6] = (mid_1[1327:1320] > top_2[1319:1312]) ? 1 : 0;
assign detect_max[164][7] = (mid_1[1327:1320] > top_2[1327:1320]) ? 1 : 0;
assign detect_max[164][8] = (mid_1[1327:1320] > top_2[1335:1328]) ? 1 : 0;
assign detect_max[164][9] = (mid_1[1327:1320] > mid_0[1319:1312]) ? 1 : 0;
assign detect_max[164][10] = (mid_1[1327:1320] > mid_0[1327:1320]) ? 1 : 0;
assign detect_max[164][11] = (mid_1[1327:1320] > mid_0[1335:1328]) ? 1 : 0;
assign detect_max[164][12] = (mid_1[1327:1320] > mid_1[1319:1312]) ? 1 : 0;
assign detect_max[164][13] = (mid_1[1327:1320] > mid_1[1335:1328]) ? 1 : 0;
assign detect_max[164][14] = (mid_1[1327:1320] > mid_2[1319:1312]) ? 1 : 0;
assign detect_max[164][15] = (mid_1[1327:1320] > mid_2[1327:1320]) ? 1 : 0;
assign detect_max[164][16] = (mid_1[1327:1320] > mid_2[1335:1328]) ? 1 : 0;
assign detect_max[164][17] = (mid_1[1327:1320] > btm_0[1319:1312]) ? 1 : 0;
assign detect_max[164][18] = (mid_1[1327:1320] > btm_0[1327:1320]) ? 1 : 0;
assign detect_max[164][19] = (mid_1[1327:1320] > btm_0[1335:1328]) ? 1 : 0;
assign detect_max[164][20] = (mid_1[1327:1320] > btm_1[1319:1312]) ? 1 : 0;
assign detect_max[164][21] = (mid_1[1327:1320] > btm_1[1327:1320]) ? 1 : 0;
assign detect_max[164][22] = (mid_1[1327:1320] > btm_1[1335:1328]) ? 1 : 0;
assign detect_max[164][23] = (mid_1[1327:1320] > btm_2[1319:1312]) ? 1 : 0;
assign detect_max[164][24] = (mid_1[1327:1320] > btm_2[1327:1320]) ? 1 : 0;
assign detect_max[164][25] = (mid_1[1327:1320] > btm_2[1335:1328]) ? 1 : 0;

assign detect_max[165][0] = (mid_1[1335:1328] > top_0[1327:1320]) ? 1 : 0;
assign detect_max[165][1] = (mid_1[1335:1328] > top_0[1335:1328]) ? 1 : 0;
assign detect_max[165][2] = (mid_1[1335:1328] > top_0[1343:1336]) ? 1 : 0;
assign detect_max[165][3] = (mid_1[1335:1328] > top_1[1327:1320]) ? 1 : 0;
assign detect_max[165][4] = (mid_1[1335:1328] > top_1[1335:1328]) ? 1 : 0;
assign detect_max[165][5] = (mid_1[1335:1328] > top_1[1343:1336]) ? 1 : 0;
assign detect_max[165][6] = (mid_1[1335:1328] > top_2[1327:1320]) ? 1 : 0;
assign detect_max[165][7] = (mid_1[1335:1328] > top_2[1335:1328]) ? 1 : 0;
assign detect_max[165][8] = (mid_1[1335:1328] > top_2[1343:1336]) ? 1 : 0;
assign detect_max[165][9] = (mid_1[1335:1328] > mid_0[1327:1320]) ? 1 : 0;
assign detect_max[165][10] = (mid_1[1335:1328] > mid_0[1335:1328]) ? 1 : 0;
assign detect_max[165][11] = (mid_1[1335:1328] > mid_0[1343:1336]) ? 1 : 0;
assign detect_max[165][12] = (mid_1[1335:1328] > mid_1[1327:1320]) ? 1 : 0;
assign detect_max[165][13] = (mid_1[1335:1328] > mid_1[1343:1336]) ? 1 : 0;
assign detect_max[165][14] = (mid_1[1335:1328] > mid_2[1327:1320]) ? 1 : 0;
assign detect_max[165][15] = (mid_1[1335:1328] > mid_2[1335:1328]) ? 1 : 0;
assign detect_max[165][16] = (mid_1[1335:1328] > mid_2[1343:1336]) ? 1 : 0;
assign detect_max[165][17] = (mid_1[1335:1328] > btm_0[1327:1320]) ? 1 : 0;
assign detect_max[165][18] = (mid_1[1335:1328] > btm_0[1335:1328]) ? 1 : 0;
assign detect_max[165][19] = (mid_1[1335:1328] > btm_0[1343:1336]) ? 1 : 0;
assign detect_max[165][20] = (mid_1[1335:1328] > btm_1[1327:1320]) ? 1 : 0;
assign detect_max[165][21] = (mid_1[1335:1328] > btm_1[1335:1328]) ? 1 : 0;
assign detect_max[165][22] = (mid_1[1335:1328] > btm_1[1343:1336]) ? 1 : 0;
assign detect_max[165][23] = (mid_1[1335:1328] > btm_2[1327:1320]) ? 1 : 0;
assign detect_max[165][24] = (mid_1[1335:1328] > btm_2[1335:1328]) ? 1 : 0;
assign detect_max[165][25] = (mid_1[1335:1328] > btm_2[1343:1336]) ? 1 : 0;

assign detect_max[166][0] = (mid_1[1343:1336] > top_0[1335:1328]) ? 1 : 0;
assign detect_max[166][1] = (mid_1[1343:1336] > top_0[1343:1336]) ? 1 : 0;
assign detect_max[166][2] = (mid_1[1343:1336] > top_0[1351:1344]) ? 1 : 0;
assign detect_max[166][3] = (mid_1[1343:1336] > top_1[1335:1328]) ? 1 : 0;
assign detect_max[166][4] = (mid_1[1343:1336] > top_1[1343:1336]) ? 1 : 0;
assign detect_max[166][5] = (mid_1[1343:1336] > top_1[1351:1344]) ? 1 : 0;
assign detect_max[166][6] = (mid_1[1343:1336] > top_2[1335:1328]) ? 1 : 0;
assign detect_max[166][7] = (mid_1[1343:1336] > top_2[1343:1336]) ? 1 : 0;
assign detect_max[166][8] = (mid_1[1343:1336] > top_2[1351:1344]) ? 1 : 0;
assign detect_max[166][9] = (mid_1[1343:1336] > mid_0[1335:1328]) ? 1 : 0;
assign detect_max[166][10] = (mid_1[1343:1336] > mid_0[1343:1336]) ? 1 : 0;
assign detect_max[166][11] = (mid_1[1343:1336] > mid_0[1351:1344]) ? 1 : 0;
assign detect_max[166][12] = (mid_1[1343:1336] > mid_1[1335:1328]) ? 1 : 0;
assign detect_max[166][13] = (mid_1[1343:1336] > mid_1[1351:1344]) ? 1 : 0;
assign detect_max[166][14] = (mid_1[1343:1336] > mid_2[1335:1328]) ? 1 : 0;
assign detect_max[166][15] = (mid_1[1343:1336] > mid_2[1343:1336]) ? 1 : 0;
assign detect_max[166][16] = (mid_1[1343:1336] > mid_2[1351:1344]) ? 1 : 0;
assign detect_max[166][17] = (mid_1[1343:1336] > btm_0[1335:1328]) ? 1 : 0;
assign detect_max[166][18] = (mid_1[1343:1336] > btm_0[1343:1336]) ? 1 : 0;
assign detect_max[166][19] = (mid_1[1343:1336] > btm_0[1351:1344]) ? 1 : 0;
assign detect_max[166][20] = (mid_1[1343:1336] > btm_1[1335:1328]) ? 1 : 0;
assign detect_max[166][21] = (mid_1[1343:1336] > btm_1[1343:1336]) ? 1 : 0;
assign detect_max[166][22] = (mid_1[1343:1336] > btm_1[1351:1344]) ? 1 : 0;
assign detect_max[166][23] = (mid_1[1343:1336] > btm_2[1335:1328]) ? 1 : 0;
assign detect_max[166][24] = (mid_1[1343:1336] > btm_2[1343:1336]) ? 1 : 0;
assign detect_max[166][25] = (mid_1[1343:1336] > btm_2[1351:1344]) ? 1 : 0;

assign detect_max[167][0] = (mid_1[1351:1344] > top_0[1343:1336]) ? 1 : 0;
assign detect_max[167][1] = (mid_1[1351:1344] > top_0[1351:1344]) ? 1 : 0;
assign detect_max[167][2] = (mid_1[1351:1344] > top_0[1359:1352]) ? 1 : 0;
assign detect_max[167][3] = (mid_1[1351:1344] > top_1[1343:1336]) ? 1 : 0;
assign detect_max[167][4] = (mid_1[1351:1344] > top_1[1351:1344]) ? 1 : 0;
assign detect_max[167][5] = (mid_1[1351:1344] > top_1[1359:1352]) ? 1 : 0;
assign detect_max[167][6] = (mid_1[1351:1344] > top_2[1343:1336]) ? 1 : 0;
assign detect_max[167][7] = (mid_1[1351:1344] > top_2[1351:1344]) ? 1 : 0;
assign detect_max[167][8] = (mid_1[1351:1344] > top_2[1359:1352]) ? 1 : 0;
assign detect_max[167][9] = (mid_1[1351:1344] > mid_0[1343:1336]) ? 1 : 0;
assign detect_max[167][10] = (mid_1[1351:1344] > mid_0[1351:1344]) ? 1 : 0;
assign detect_max[167][11] = (mid_1[1351:1344] > mid_0[1359:1352]) ? 1 : 0;
assign detect_max[167][12] = (mid_1[1351:1344] > mid_1[1343:1336]) ? 1 : 0;
assign detect_max[167][13] = (mid_1[1351:1344] > mid_1[1359:1352]) ? 1 : 0;
assign detect_max[167][14] = (mid_1[1351:1344] > mid_2[1343:1336]) ? 1 : 0;
assign detect_max[167][15] = (mid_1[1351:1344] > mid_2[1351:1344]) ? 1 : 0;
assign detect_max[167][16] = (mid_1[1351:1344] > mid_2[1359:1352]) ? 1 : 0;
assign detect_max[167][17] = (mid_1[1351:1344] > btm_0[1343:1336]) ? 1 : 0;
assign detect_max[167][18] = (mid_1[1351:1344] > btm_0[1351:1344]) ? 1 : 0;
assign detect_max[167][19] = (mid_1[1351:1344] > btm_0[1359:1352]) ? 1 : 0;
assign detect_max[167][20] = (mid_1[1351:1344] > btm_1[1343:1336]) ? 1 : 0;
assign detect_max[167][21] = (mid_1[1351:1344] > btm_1[1351:1344]) ? 1 : 0;
assign detect_max[167][22] = (mid_1[1351:1344] > btm_1[1359:1352]) ? 1 : 0;
assign detect_max[167][23] = (mid_1[1351:1344] > btm_2[1343:1336]) ? 1 : 0;
assign detect_max[167][24] = (mid_1[1351:1344] > btm_2[1351:1344]) ? 1 : 0;
assign detect_max[167][25] = (mid_1[1351:1344] > btm_2[1359:1352]) ? 1 : 0;

assign detect_max[168][0] = (mid_1[1359:1352] > top_0[1351:1344]) ? 1 : 0;
assign detect_max[168][1] = (mid_1[1359:1352] > top_0[1359:1352]) ? 1 : 0;
assign detect_max[168][2] = (mid_1[1359:1352] > top_0[1367:1360]) ? 1 : 0;
assign detect_max[168][3] = (mid_1[1359:1352] > top_1[1351:1344]) ? 1 : 0;
assign detect_max[168][4] = (mid_1[1359:1352] > top_1[1359:1352]) ? 1 : 0;
assign detect_max[168][5] = (mid_1[1359:1352] > top_1[1367:1360]) ? 1 : 0;
assign detect_max[168][6] = (mid_1[1359:1352] > top_2[1351:1344]) ? 1 : 0;
assign detect_max[168][7] = (mid_1[1359:1352] > top_2[1359:1352]) ? 1 : 0;
assign detect_max[168][8] = (mid_1[1359:1352] > top_2[1367:1360]) ? 1 : 0;
assign detect_max[168][9] = (mid_1[1359:1352] > mid_0[1351:1344]) ? 1 : 0;
assign detect_max[168][10] = (mid_1[1359:1352] > mid_0[1359:1352]) ? 1 : 0;
assign detect_max[168][11] = (mid_1[1359:1352] > mid_0[1367:1360]) ? 1 : 0;
assign detect_max[168][12] = (mid_1[1359:1352] > mid_1[1351:1344]) ? 1 : 0;
assign detect_max[168][13] = (mid_1[1359:1352] > mid_1[1367:1360]) ? 1 : 0;
assign detect_max[168][14] = (mid_1[1359:1352] > mid_2[1351:1344]) ? 1 : 0;
assign detect_max[168][15] = (mid_1[1359:1352] > mid_2[1359:1352]) ? 1 : 0;
assign detect_max[168][16] = (mid_1[1359:1352] > mid_2[1367:1360]) ? 1 : 0;
assign detect_max[168][17] = (mid_1[1359:1352] > btm_0[1351:1344]) ? 1 : 0;
assign detect_max[168][18] = (mid_1[1359:1352] > btm_0[1359:1352]) ? 1 : 0;
assign detect_max[168][19] = (mid_1[1359:1352] > btm_0[1367:1360]) ? 1 : 0;
assign detect_max[168][20] = (mid_1[1359:1352] > btm_1[1351:1344]) ? 1 : 0;
assign detect_max[168][21] = (mid_1[1359:1352] > btm_1[1359:1352]) ? 1 : 0;
assign detect_max[168][22] = (mid_1[1359:1352] > btm_1[1367:1360]) ? 1 : 0;
assign detect_max[168][23] = (mid_1[1359:1352] > btm_2[1351:1344]) ? 1 : 0;
assign detect_max[168][24] = (mid_1[1359:1352] > btm_2[1359:1352]) ? 1 : 0;
assign detect_max[168][25] = (mid_1[1359:1352] > btm_2[1367:1360]) ? 1 : 0;

assign detect_max[169][0] = (mid_1[1367:1360] > top_0[1359:1352]) ? 1 : 0;
assign detect_max[169][1] = (mid_1[1367:1360] > top_0[1367:1360]) ? 1 : 0;
assign detect_max[169][2] = (mid_1[1367:1360] > top_0[1375:1368]) ? 1 : 0;
assign detect_max[169][3] = (mid_1[1367:1360] > top_1[1359:1352]) ? 1 : 0;
assign detect_max[169][4] = (mid_1[1367:1360] > top_1[1367:1360]) ? 1 : 0;
assign detect_max[169][5] = (mid_1[1367:1360] > top_1[1375:1368]) ? 1 : 0;
assign detect_max[169][6] = (mid_1[1367:1360] > top_2[1359:1352]) ? 1 : 0;
assign detect_max[169][7] = (mid_1[1367:1360] > top_2[1367:1360]) ? 1 : 0;
assign detect_max[169][8] = (mid_1[1367:1360] > top_2[1375:1368]) ? 1 : 0;
assign detect_max[169][9] = (mid_1[1367:1360] > mid_0[1359:1352]) ? 1 : 0;
assign detect_max[169][10] = (mid_1[1367:1360] > mid_0[1367:1360]) ? 1 : 0;
assign detect_max[169][11] = (mid_1[1367:1360] > mid_0[1375:1368]) ? 1 : 0;
assign detect_max[169][12] = (mid_1[1367:1360] > mid_1[1359:1352]) ? 1 : 0;
assign detect_max[169][13] = (mid_1[1367:1360] > mid_1[1375:1368]) ? 1 : 0;
assign detect_max[169][14] = (mid_1[1367:1360] > mid_2[1359:1352]) ? 1 : 0;
assign detect_max[169][15] = (mid_1[1367:1360] > mid_2[1367:1360]) ? 1 : 0;
assign detect_max[169][16] = (mid_1[1367:1360] > mid_2[1375:1368]) ? 1 : 0;
assign detect_max[169][17] = (mid_1[1367:1360] > btm_0[1359:1352]) ? 1 : 0;
assign detect_max[169][18] = (mid_1[1367:1360] > btm_0[1367:1360]) ? 1 : 0;
assign detect_max[169][19] = (mid_1[1367:1360] > btm_0[1375:1368]) ? 1 : 0;
assign detect_max[169][20] = (mid_1[1367:1360] > btm_1[1359:1352]) ? 1 : 0;
assign detect_max[169][21] = (mid_1[1367:1360] > btm_1[1367:1360]) ? 1 : 0;
assign detect_max[169][22] = (mid_1[1367:1360] > btm_1[1375:1368]) ? 1 : 0;
assign detect_max[169][23] = (mid_1[1367:1360] > btm_2[1359:1352]) ? 1 : 0;
assign detect_max[169][24] = (mid_1[1367:1360] > btm_2[1367:1360]) ? 1 : 0;
assign detect_max[169][25] = (mid_1[1367:1360] > btm_2[1375:1368]) ? 1 : 0;

assign detect_max[170][0] = (mid_1[1375:1368] > top_0[1367:1360]) ? 1 : 0;
assign detect_max[170][1] = (mid_1[1375:1368] > top_0[1375:1368]) ? 1 : 0;
assign detect_max[170][2] = (mid_1[1375:1368] > top_0[1383:1376]) ? 1 : 0;
assign detect_max[170][3] = (mid_1[1375:1368] > top_1[1367:1360]) ? 1 : 0;
assign detect_max[170][4] = (mid_1[1375:1368] > top_1[1375:1368]) ? 1 : 0;
assign detect_max[170][5] = (mid_1[1375:1368] > top_1[1383:1376]) ? 1 : 0;
assign detect_max[170][6] = (mid_1[1375:1368] > top_2[1367:1360]) ? 1 : 0;
assign detect_max[170][7] = (mid_1[1375:1368] > top_2[1375:1368]) ? 1 : 0;
assign detect_max[170][8] = (mid_1[1375:1368] > top_2[1383:1376]) ? 1 : 0;
assign detect_max[170][9] = (mid_1[1375:1368] > mid_0[1367:1360]) ? 1 : 0;
assign detect_max[170][10] = (mid_1[1375:1368] > mid_0[1375:1368]) ? 1 : 0;
assign detect_max[170][11] = (mid_1[1375:1368] > mid_0[1383:1376]) ? 1 : 0;
assign detect_max[170][12] = (mid_1[1375:1368] > mid_1[1367:1360]) ? 1 : 0;
assign detect_max[170][13] = (mid_1[1375:1368] > mid_1[1383:1376]) ? 1 : 0;
assign detect_max[170][14] = (mid_1[1375:1368] > mid_2[1367:1360]) ? 1 : 0;
assign detect_max[170][15] = (mid_1[1375:1368] > mid_2[1375:1368]) ? 1 : 0;
assign detect_max[170][16] = (mid_1[1375:1368] > mid_2[1383:1376]) ? 1 : 0;
assign detect_max[170][17] = (mid_1[1375:1368] > btm_0[1367:1360]) ? 1 : 0;
assign detect_max[170][18] = (mid_1[1375:1368] > btm_0[1375:1368]) ? 1 : 0;
assign detect_max[170][19] = (mid_1[1375:1368] > btm_0[1383:1376]) ? 1 : 0;
assign detect_max[170][20] = (mid_1[1375:1368] > btm_1[1367:1360]) ? 1 : 0;
assign detect_max[170][21] = (mid_1[1375:1368] > btm_1[1375:1368]) ? 1 : 0;
assign detect_max[170][22] = (mid_1[1375:1368] > btm_1[1383:1376]) ? 1 : 0;
assign detect_max[170][23] = (mid_1[1375:1368] > btm_2[1367:1360]) ? 1 : 0;
assign detect_max[170][24] = (mid_1[1375:1368] > btm_2[1375:1368]) ? 1 : 0;
assign detect_max[170][25] = (mid_1[1375:1368] > btm_2[1383:1376]) ? 1 : 0;

assign detect_max[171][0] = (mid_1[1383:1376] > top_0[1375:1368]) ? 1 : 0;
assign detect_max[171][1] = (mid_1[1383:1376] > top_0[1383:1376]) ? 1 : 0;
assign detect_max[171][2] = (mid_1[1383:1376] > top_0[1391:1384]) ? 1 : 0;
assign detect_max[171][3] = (mid_1[1383:1376] > top_1[1375:1368]) ? 1 : 0;
assign detect_max[171][4] = (mid_1[1383:1376] > top_1[1383:1376]) ? 1 : 0;
assign detect_max[171][5] = (mid_1[1383:1376] > top_1[1391:1384]) ? 1 : 0;
assign detect_max[171][6] = (mid_1[1383:1376] > top_2[1375:1368]) ? 1 : 0;
assign detect_max[171][7] = (mid_1[1383:1376] > top_2[1383:1376]) ? 1 : 0;
assign detect_max[171][8] = (mid_1[1383:1376] > top_2[1391:1384]) ? 1 : 0;
assign detect_max[171][9] = (mid_1[1383:1376] > mid_0[1375:1368]) ? 1 : 0;
assign detect_max[171][10] = (mid_1[1383:1376] > mid_0[1383:1376]) ? 1 : 0;
assign detect_max[171][11] = (mid_1[1383:1376] > mid_0[1391:1384]) ? 1 : 0;
assign detect_max[171][12] = (mid_1[1383:1376] > mid_1[1375:1368]) ? 1 : 0;
assign detect_max[171][13] = (mid_1[1383:1376] > mid_1[1391:1384]) ? 1 : 0;
assign detect_max[171][14] = (mid_1[1383:1376] > mid_2[1375:1368]) ? 1 : 0;
assign detect_max[171][15] = (mid_1[1383:1376] > mid_2[1383:1376]) ? 1 : 0;
assign detect_max[171][16] = (mid_1[1383:1376] > mid_2[1391:1384]) ? 1 : 0;
assign detect_max[171][17] = (mid_1[1383:1376] > btm_0[1375:1368]) ? 1 : 0;
assign detect_max[171][18] = (mid_1[1383:1376] > btm_0[1383:1376]) ? 1 : 0;
assign detect_max[171][19] = (mid_1[1383:1376] > btm_0[1391:1384]) ? 1 : 0;
assign detect_max[171][20] = (mid_1[1383:1376] > btm_1[1375:1368]) ? 1 : 0;
assign detect_max[171][21] = (mid_1[1383:1376] > btm_1[1383:1376]) ? 1 : 0;
assign detect_max[171][22] = (mid_1[1383:1376] > btm_1[1391:1384]) ? 1 : 0;
assign detect_max[171][23] = (mid_1[1383:1376] > btm_2[1375:1368]) ? 1 : 0;
assign detect_max[171][24] = (mid_1[1383:1376] > btm_2[1383:1376]) ? 1 : 0;
assign detect_max[171][25] = (mid_1[1383:1376] > btm_2[1391:1384]) ? 1 : 0;

assign detect_max[172][0] = (mid_1[1391:1384] > top_0[1383:1376]) ? 1 : 0;
assign detect_max[172][1] = (mid_1[1391:1384] > top_0[1391:1384]) ? 1 : 0;
assign detect_max[172][2] = (mid_1[1391:1384] > top_0[1399:1392]) ? 1 : 0;
assign detect_max[172][3] = (mid_1[1391:1384] > top_1[1383:1376]) ? 1 : 0;
assign detect_max[172][4] = (mid_1[1391:1384] > top_1[1391:1384]) ? 1 : 0;
assign detect_max[172][5] = (mid_1[1391:1384] > top_1[1399:1392]) ? 1 : 0;
assign detect_max[172][6] = (mid_1[1391:1384] > top_2[1383:1376]) ? 1 : 0;
assign detect_max[172][7] = (mid_1[1391:1384] > top_2[1391:1384]) ? 1 : 0;
assign detect_max[172][8] = (mid_1[1391:1384] > top_2[1399:1392]) ? 1 : 0;
assign detect_max[172][9] = (mid_1[1391:1384] > mid_0[1383:1376]) ? 1 : 0;
assign detect_max[172][10] = (mid_1[1391:1384] > mid_0[1391:1384]) ? 1 : 0;
assign detect_max[172][11] = (mid_1[1391:1384] > mid_0[1399:1392]) ? 1 : 0;
assign detect_max[172][12] = (mid_1[1391:1384] > mid_1[1383:1376]) ? 1 : 0;
assign detect_max[172][13] = (mid_1[1391:1384] > mid_1[1399:1392]) ? 1 : 0;
assign detect_max[172][14] = (mid_1[1391:1384] > mid_2[1383:1376]) ? 1 : 0;
assign detect_max[172][15] = (mid_1[1391:1384] > mid_2[1391:1384]) ? 1 : 0;
assign detect_max[172][16] = (mid_1[1391:1384] > mid_2[1399:1392]) ? 1 : 0;
assign detect_max[172][17] = (mid_1[1391:1384] > btm_0[1383:1376]) ? 1 : 0;
assign detect_max[172][18] = (mid_1[1391:1384] > btm_0[1391:1384]) ? 1 : 0;
assign detect_max[172][19] = (mid_1[1391:1384] > btm_0[1399:1392]) ? 1 : 0;
assign detect_max[172][20] = (mid_1[1391:1384] > btm_1[1383:1376]) ? 1 : 0;
assign detect_max[172][21] = (mid_1[1391:1384] > btm_1[1391:1384]) ? 1 : 0;
assign detect_max[172][22] = (mid_1[1391:1384] > btm_1[1399:1392]) ? 1 : 0;
assign detect_max[172][23] = (mid_1[1391:1384] > btm_2[1383:1376]) ? 1 : 0;
assign detect_max[172][24] = (mid_1[1391:1384] > btm_2[1391:1384]) ? 1 : 0;
assign detect_max[172][25] = (mid_1[1391:1384] > btm_2[1399:1392]) ? 1 : 0;

assign detect_max[173][0] = (mid_1[1399:1392] > top_0[1391:1384]) ? 1 : 0;
assign detect_max[173][1] = (mid_1[1399:1392] > top_0[1399:1392]) ? 1 : 0;
assign detect_max[173][2] = (mid_1[1399:1392] > top_0[1407:1400]) ? 1 : 0;
assign detect_max[173][3] = (mid_1[1399:1392] > top_1[1391:1384]) ? 1 : 0;
assign detect_max[173][4] = (mid_1[1399:1392] > top_1[1399:1392]) ? 1 : 0;
assign detect_max[173][5] = (mid_1[1399:1392] > top_1[1407:1400]) ? 1 : 0;
assign detect_max[173][6] = (mid_1[1399:1392] > top_2[1391:1384]) ? 1 : 0;
assign detect_max[173][7] = (mid_1[1399:1392] > top_2[1399:1392]) ? 1 : 0;
assign detect_max[173][8] = (mid_1[1399:1392] > top_2[1407:1400]) ? 1 : 0;
assign detect_max[173][9] = (mid_1[1399:1392] > mid_0[1391:1384]) ? 1 : 0;
assign detect_max[173][10] = (mid_1[1399:1392] > mid_0[1399:1392]) ? 1 : 0;
assign detect_max[173][11] = (mid_1[1399:1392] > mid_0[1407:1400]) ? 1 : 0;
assign detect_max[173][12] = (mid_1[1399:1392] > mid_1[1391:1384]) ? 1 : 0;
assign detect_max[173][13] = (mid_1[1399:1392] > mid_1[1407:1400]) ? 1 : 0;
assign detect_max[173][14] = (mid_1[1399:1392] > mid_2[1391:1384]) ? 1 : 0;
assign detect_max[173][15] = (mid_1[1399:1392] > mid_2[1399:1392]) ? 1 : 0;
assign detect_max[173][16] = (mid_1[1399:1392] > mid_2[1407:1400]) ? 1 : 0;
assign detect_max[173][17] = (mid_1[1399:1392] > btm_0[1391:1384]) ? 1 : 0;
assign detect_max[173][18] = (mid_1[1399:1392] > btm_0[1399:1392]) ? 1 : 0;
assign detect_max[173][19] = (mid_1[1399:1392] > btm_0[1407:1400]) ? 1 : 0;
assign detect_max[173][20] = (mid_1[1399:1392] > btm_1[1391:1384]) ? 1 : 0;
assign detect_max[173][21] = (mid_1[1399:1392] > btm_1[1399:1392]) ? 1 : 0;
assign detect_max[173][22] = (mid_1[1399:1392] > btm_1[1407:1400]) ? 1 : 0;
assign detect_max[173][23] = (mid_1[1399:1392] > btm_2[1391:1384]) ? 1 : 0;
assign detect_max[173][24] = (mid_1[1399:1392] > btm_2[1399:1392]) ? 1 : 0;
assign detect_max[173][25] = (mid_1[1399:1392] > btm_2[1407:1400]) ? 1 : 0;

assign detect_max[174][0] = (mid_1[1407:1400] > top_0[1399:1392]) ? 1 : 0;
assign detect_max[174][1] = (mid_1[1407:1400] > top_0[1407:1400]) ? 1 : 0;
assign detect_max[174][2] = (mid_1[1407:1400] > top_0[1415:1408]) ? 1 : 0;
assign detect_max[174][3] = (mid_1[1407:1400] > top_1[1399:1392]) ? 1 : 0;
assign detect_max[174][4] = (mid_1[1407:1400] > top_1[1407:1400]) ? 1 : 0;
assign detect_max[174][5] = (mid_1[1407:1400] > top_1[1415:1408]) ? 1 : 0;
assign detect_max[174][6] = (mid_1[1407:1400] > top_2[1399:1392]) ? 1 : 0;
assign detect_max[174][7] = (mid_1[1407:1400] > top_2[1407:1400]) ? 1 : 0;
assign detect_max[174][8] = (mid_1[1407:1400] > top_2[1415:1408]) ? 1 : 0;
assign detect_max[174][9] = (mid_1[1407:1400] > mid_0[1399:1392]) ? 1 : 0;
assign detect_max[174][10] = (mid_1[1407:1400] > mid_0[1407:1400]) ? 1 : 0;
assign detect_max[174][11] = (mid_1[1407:1400] > mid_0[1415:1408]) ? 1 : 0;
assign detect_max[174][12] = (mid_1[1407:1400] > mid_1[1399:1392]) ? 1 : 0;
assign detect_max[174][13] = (mid_1[1407:1400] > mid_1[1415:1408]) ? 1 : 0;
assign detect_max[174][14] = (mid_1[1407:1400] > mid_2[1399:1392]) ? 1 : 0;
assign detect_max[174][15] = (mid_1[1407:1400] > mid_2[1407:1400]) ? 1 : 0;
assign detect_max[174][16] = (mid_1[1407:1400] > mid_2[1415:1408]) ? 1 : 0;
assign detect_max[174][17] = (mid_1[1407:1400] > btm_0[1399:1392]) ? 1 : 0;
assign detect_max[174][18] = (mid_1[1407:1400] > btm_0[1407:1400]) ? 1 : 0;
assign detect_max[174][19] = (mid_1[1407:1400] > btm_0[1415:1408]) ? 1 : 0;
assign detect_max[174][20] = (mid_1[1407:1400] > btm_1[1399:1392]) ? 1 : 0;
assign detect_max[174][21] = (mid_1[1407:1400] > btm_1[1407:1400]) ? 1 : 0;
assign detect_max[174][22] = (mid_1[1407:1400] > btm_1[1415:1408]) ? 1 : 0;
assign detect_max[174][23] = (mid_1[1407:1400] > btm_2[1399:1392]) ? 1 : 0;
assign detect_max[174][24] = (mid_1[1407:1400] > btm_2[1407:1400]) ? 1 : 0;
assign detect_max[174][25] = (mid_1[1407:1400] > btm_2[1415:1408]) ? 1 : 0;

assign detect_max[175][0] = (mid_1[1415:1408] > top_0[1407:1400]) ? 1 : 0;
assign detect_max[175][1] = (mid_1[1415:1408] > top_0[1415:1408]) ? 1 : 0;
assign detect_max[175][2] = (mid_1[1415:1408] > top_0[1423:1416]) ? 1 : 0;
assign detect_max[175][3] = (mid_1[1415:1408] > top_1[1407:1400]) ? 1 : 0;
assign detect_max[175][4] = (mid_1[1415:1408] > top_1[1415:1408]) ? 1 : 0;
assign detect_max[175][5] = (mid_1[1415:1408] > top_1[1423:1416]) ? 1 : 0;
assign detect_max[175][6] = (mid_1[1415:1408] > top_2[1407:1400]) ? 1 : 0;
assign detect_max[175][7] = (mid_1[1415:1408] > top_2[1415:1408]) ? 1 : 0;
assign detect_max[175][8] = (mid_1[1415:1408] > top_2[1423:1416]) ? 1 : 0;
assign detect_max[175][9] = (mid_1[1415:1408] > mid_0[1407:1400]) ? 1 : 0;
assign detect_max[175][10] = (mid_1[1415:1408] > mid_0[1415:1408]) ? 1 : 0;
assign detect_max[175][11] = (mid_1[1415:1408] > mid_0[1423:1416]) ? 1 : 0;
assign detect_max[175][12] = (mid_1[1415:1408] > mid_1[1407:1400]) ? 1 : 0;
assign detect_max[175][13] = (mid_1[1415:1408] > mid_1[1423:1416]) ? 1 : 0;
assign detect_max[175][14] = (mid_1[1415:1408] > mid_2[1407:1400]) ? 1 : 0;
assign detect_max[175][15] = (mid_1[1415:1408] > mid_2[1415:1408]) ? 1 : 0;
assign detect_max[175][16] = (mid_1[1415:1408] > mid_2[1423:1416]) ? 1 : 0;
assign detect_max[175][17] = (mid_1[1415:1408] > btm_0[1407:1400]) ? 1 : 0;
assign detect_max[175][18] = (mid_1[1415:1408] > btm_0[1415:1408]) ? 1 : 0;
assign detect_max[175][19] = (mid_1[1415:1408] > btm_0[1423:1416]) ? 1 : 0;
assign detect_max[175][20] = (mid_1[1415:1408] > btm_1[1407:1400]) ? 1 : 0;
assign detect_max[175][21] = (mid_1[1415:1408] > btm_1[1415:1408]) ? 1 : 0;
assign detect_max[175][22] = (mid_1[1415:1408] > btm_1[1423:1416]) ? 1 : 0;
assign detect_max[175][23] = (mid_1[1415:1408] > btm_2[1407:1400]) ? 1 : 0;
assign detect_max[175][24] = (mid_1[1415:1408] > btm_2[1415:1408]) ? 1 : 0;
assign detect_max[175][25] = (mid_1[1415:1408] > btm_2[1423:1416]) ? 1 : 0;

assign detect_max[176][0] = (mid_1[1423:1416] > top_0[1415:1408]) ? 1 : 0;
assign detect_max[176][1] = (mid_1[1423:1416] > top_0[1423:1416]) ? 1 : 0;
assign detect_max[176][2] = (mid_1[1423:1416] > top_0[1431:1424]) ? 1 : 0;
assign detect_max[176][3] = (mid_1[1423:1416] > top_1[1415:1408]) ? 1 : 0;
assign detect_max[176][4] = (mid_1[1423:1416] > top_1[1423:1416]) ? 1 : 0;
assign detect_max[176][5] = (mid_1[1423:1416] > top_1[1431:1424]) ? 1 : 0;
assign detect_max[176][6] = (mid_1[1423:1416] > top_2[1415:1408]) ? 1 : 0;
assign detect_max[176][7] = (mid_1[1423:1416] > top_2[1423:1416]) ? 1 : 0;
assign detect_max[176][8] = (mid_1[1423:1416] > top_2[1431:1424]) ? 1 : 0;
assign detect_max[176][9] = (mid_1[1423:1416] > mid_0[1415:1408]) ? 1 : 0;
assign detect_max[176][10] = (mid_1[1423:1416] > mid_0[1423:1416]) ? 1 : 0;
assign detect_max[176][11] = (mid_1[1423:1416] > mid_0[1431:1424]) ? 1 : 0;
assign detect_max[176][12] = (mid_1[1423:1416] > mid_1[1415:1408]) ? 1 : 0;
assign detect_max[176][13] = (mid_1[1423:1416] > mid_1[1431:1424]) ? 1 : 0;
assign detect_max[176][14] = (mid_1[1423:1416] > mid_2[1415:1408]) ? 1 : 0;
assign detect_max[176][15] = (mid_1[1423:1416] > mid_2[1423:1416]) ? 1 : 0;
assign detect_max[176][16] = (mid_1[1423:1416] > mid_2[1431:1424]) ? 1 : 0;
assign detect_max[176][17] = (mid_1[1423:1416] > btm_0[1415:1408]) ? 1 : 0;
assign detect_max[176][18] = (mid_1[1423:1416] > btm_0[1423:1416]) ? 1 : 0;
assign detect_max[176][19] = (mid_1[1423:1416] > btm_0[1431:1424]) ? 1 : 0;
assign detect_max[176][20] = (mid_1[1423:1416] > btm_1[1415:1408]) ? 1 : 0;
assign detect_max[176][21] = (mid_1[1423:1416] > btm_1[1423:1416]) ? 1 : 0;
assign detect_max[176][22] = (mid_1[1423:1416] > btm_1[1431:1424]) ? 1 : 0;
assign detect_max[176][23] = (mid_1[1423:1416] > btm_2[1415:1408]) ? 1 : 0;
assign detect_max[176][24] = (mid_1[1423:1416] > btm_2[1423:1416]) ? 1 : 0;
assign detect_max[176][25] = (mid_1[1423:1416] > btm_2[1431:1424]) ? 1 : 0;

assign detect_max[177][0] = (mid_1[1431:1424] > top_0[1423:1416]) ? 1 : 0;
assign detect_max[177][1] = (mid_1[1431:1424] > top_0[1431:1424]) ? 1 : 0;
assign detect_max[177][2] = (mid_1[1431:1424] > top_0[1439:1432]) ? 1 : 0;
assign detect_max[177][3] = (mid_1[1431:1424] > top_1[1423:1416]) ? 1 : 0;
assign detect_max[177][4] = (mid_1[1431:1424] > top_1[1431:1424]) ? 1 : 0;
assign detect_max[177][5] = (mid_1[1431:1424] > top_1[1439:1432]) ? 1 : 0;
assign detect_max[177][6] = (mid_1[1431:1424] > top_2[1423:1416]) ? 1 : 0;
assign detect_max[177][7] = (mid_1[1431:1424] > top_2[1431:1424]) ? 1 : 0;
assign detect_max[177][8] = (mid_1[1431:1424] > top_2[1439:1432]) ? 1 : 0;
assign detect_max[177][9] = (mid_1[1431:1424] > mid_0[1423:1416]) ? 1 : 0;
assign detect_max[177][10] = (mid_1[1431:1424] > mid_0[1431:1424]) ? 1 : 0;
assign detect_max[177][11] = (mid_1[1431:1424] > mid_0[1439:1432]) ? 1 : 0;
assign detect_max[177][12] = (mid_1[1431:1424] > mid_1[1423:1416]) ? 1 : 0;
assign detect_max[177][13] = (mid_1[1431:1424] > mid_1[1439:1432]) ? 1 : 0;
assign detect_max[177][14] = (mid_1[1431:1424] > mid_2[1423:1416]) ? 1 : 0;
assign detect_max[177][15] = (mid_1[1431:1424] > mid_2[1431:1424]) ? 1 : 0;
assign detect_max[177][16] = (mid_1[1431:1424] > mid_2[1439:1432]) ? 1 : 0;
assign detect_max[177][17] = (mid_1[1431:1424] > btm_0[1423:1416]) ? 1 : 0;
assign detect_max[177][18] = (mid_1[1431:1424] > btm_0[1431:1424]) ? 1 : 0;
assign detect_max[177][19] = (mid_1[1431:1424] > btm_0[1439:1432]) ? 1 : 0;
assign detect_max[177][20] = (mid_1[1431:1424] > btm_1[1423:1416]) ? 1 : 0;
assign detect_max[177][21] = (mid_1[1431:1424] > btm_1[1431:1424]) ? 1 : 0;
assign detect_max[177][22] = (mid_1[1431:1424] > btm_1[1439:1432]) ? 1 : 0;
assign detect_max[177][23] = (mid_1[1431:1424] > btm_2[1423:1416]) ? 1 : 0;
assign detect_max[177][24] = (mid_1[1431:1424] > btm_2[1431:1424]) ? 1 : 0;
assign detect_max[177][25] = (mid_1[1431:1424] > btm_2[1439:1432]) ? 1 : 0;

assign detect_max[178][0] = (mid_1[1439:1432] > top_0[1431:1424]) ? 1 : 0;
assign detect_max[178][1] = (mid_1[1439:1432] > top_0[1439:1432]) ? 1 : 0;
assign detect_max[178][2] = (mid_1[1439:1432] > top_0[1447:1440]) ? 1 : 0;
assign detect_max[178][3] = (mid_1[1439:1432] > top_1[1431:1424]) ? 1 : 0;
assign detect_max[178][4] = (mid_1[1439:1432] > top_1[1439:1432]) ? 1 : 0;
assign detect_max[178][5] = (mid_1[1439:1432] > top_1[1447:1440]) ? 1 : 0;
assign detect_max[178][6] = (mid_1[1439:1432] > top_2[1431:1424]) ? 1 : 0;
assign detect_max[178][7] = (mid_1[1439:1432] > top_2[1439:1432]) ? 1 : 0;
assign detect_max[178][8] = (mid_1[1439:1432] > top_2[1447:1440]) ? 1 : 0;
assign detect_max[178][9] = (mid_1[1439:1432] > mid_0[1431:1424]) ? 1 : 0;
assign detect_max[178][10] = (mid_1[1439:1432] > mid_0[1439:1432]) ? 1 : 0;
assign detect_max[178][11] = (mid_1[1439:1432] > mid_0[1447:1440]) ? 1 : 0;
assign detect_max[178][12] = (mid_1[1439:1432] > mid_1[1431:1424]) ? 1 : 0;
assign detect_max[178][13] = (mid_1[1439:1432] > mid_1[1447:1440]) ? 1 : 0;
assign detect_max[178][14] = (mid_1[1439:1432] > mid_2[1431:1424]) ? 1 : 0;
assign detect_max[178][15] = (mid_1[1439:1432] > mid_2[1439:1432]) ? 1 : 0;
assign detect_max[178][16] = (mid_1[1439:1432] > mid_2[1447:1440]) ? 1 : 0;
assign detect_max[178][17] = (mid_1[1439:1432] > btm_0[1431:1424]) ? 1 : 0;
assign detect_max[178][18] = (mid_1[1439:1432] > btm_0[1439:1432]) ? 1 : 0;
assign detect_max[178][19] = (mid_1[1439:1432] > btm_0[1447:1440]) ? 1 : 0;
assign detect_max[178][20] = (mid_1[1439:1432] > btm_1[1431:1424]) ? 1 : 0;
assign detect_max[178][21] = (mid_1[1439:1432] > btm_1[1439:1432]) ? 1 : 0;
assign detect_max[178][22] = (mid_1[1439:1432] > btm_1[1447:1440]) ? 1 : 0;
assign detect_max[178][23] = (mid_1[1439:1432] > btm_2[1431:1424]) ? 1 : 0;
assign detect_max[178][24] = (mid_1[1439:1432] > btm_2[1439:1432]) ? 1 : 0;
assign detect_max[178][25] = (mid_1[1439:1432] > btm_2[1447:1440]) ? 1 : 0;

assign detect_max[179][0] = (mid_1[1447:1440] > top_0[1439:1432]) ? 1 : 0;
assign detect_max[179][1] = (mid_1[1447:1440] > top_0[1447:1440]) ? 1 : 0;
assign detect_max[179][2] = (mid_1[1447:1440] > top_0[1455:1448]) ? 1 : 0;
assign detect_max[179][3] = (mid_1[1447:1440] > top_1[1439:1432]) ? 1 : 0;
assign detect_max[179][4] = (mid_1[1447:1440] > top_1[1447:1440]) ? 1 : 0;
assign detect_max[179][5] = (mid_1[1447:1440] > top_1[1455:1448]) ? 1 : 0;
assign detect_max[179][6] = (mid_1[1447:1440] > top_2[1439:1432]) ? 1 : 0;
assign detect_max[179][7] = (mid_1[1447:1440] > top_2[1447:1440]) ? 1 : 0;
assign detect_max[179][8] = (mid_1[1447:1440] > top_2[1455:1448]) ? 1 : 0;
assign detect_max[179][9] = (mid_1[1447:1440] > mid_0[1439:1432]) ? 1 : 0;
assign detect_max[179][10] = (mid_1[1447:1440] > mid_0[1447:1440]) ? 1 : 0;
assign detect_max[179][11] = (mid_1[1447:1440] > mid_0[1455:1448]) ? 1 : 0;
assign detect_max[179][12] = (mid_1[1447:1440] > mid_1[1439:1432]) ? 1 : 0;
assign detect_max[179][13] = (mid_1[1447:1440] > mid_1[1455:1448]) ? 1 : 0;
assign detect_max[179][14] = (mid_1[1447:1440] > mid_2[1439:1432]) ? 1 : 0;
assign detect_max[179][15] = (mid_1[1447:1440] > mid_2[1447:1440]) ? 1 : 0;
assign detect_max[179][16] = (mid_1[1447:1440] > mid_2[1455:1448]) ? 1 : 0;
assign detect_max[179][17] = (mid_1[1447:1440] > btm_0[1439:1432]) ? 1 : 0;
assign detect_max[179][18] = (mid_1[1447:1440] > btm_0[1447:1440]) ? 1 : 0;
assign detect_max[179][19] = (mid_1[1447:1440] > btm_0[1455:1448]) ? 1 : 0;
assign detect_max[179][20] = (mid_1[1447:1440] > btm_1[1439:1432]) ? 1 : 0;
assign detect_max[179][21] = (mid_1[1447:1440] > btm_1[1447:1440]) ? 1 : 0;
assign detect_max[179][22] = (mid_1[1447:1440] > btm_1[1455:1448]) ? 1 : 0;
assign detect_max[179][23] = (mid_1[1447:1440] > btm_2[1439:1432]) ? 1 : 0;
assign detect_max[179][24] = (mid_1[1447:1440] > btm_2[1447:1440]) ? 1 : 0;
assign detect_max[179][25] = (mid_1[1447:1440] > btm_2[1455:1448]) ? 1 : 0;

assign detect_max[180][0] = (mid_1[1455:1448] > top_0[1447:1440]) ? 1 : 0;
assign detect_max[180][1] = (mid_1[1455:1448] > top_0[1455:1448]) ? 1 : 0;
assign detect_max[180][2] = (mid_1[1455:1448] > top_0[1463:1456]) ? 1 : 0;
assign detect_max[180][3] = (mid_1[1455:1448] > top_1[1447:1440]) ? 1 : 0;
assign detect_max[180][4] = (mid_1[1455:1448] > top_1[1455:1448]) ? 1 : 0;
assign detect_max[180][5] = (mid_1[1455:1448] > top_1[1463:1456]) ? 1 : 0;
assign detect_max[180][6] = (mid_1[1455:1448] > top_2[1447:1440]) ? 1 : 0;
assign detect_max[180][7] = (mid_1[1455:1448] > top_2[1455:1448]) ? 1 : 0;
assign detect_max[180][8] = (mid_1[1455:1448] > top_2[1463:1456]) ? 1 : 0;
assign detect_max[180][9] = (mid_1[1455:1448] > mid_0[1447:1440]) ? 1 : 0;
assign detect_max[180][10] = (mid_1[1455:1448] > mid_0[1455:1448]) ? 1 : 0;
assign detect_max[180][11] = (mid_1[1455:1448] > mid_0[1463:1456]) ? 1 : 0;
assign detect_max[180][12] = (mid_1[1455:1448] > mid_1[1447:1440]) ? 1 : 0;
assign detect_max[180][13] = (mid_1[1455:1448] > mid_1[1463:1456]) ? 1 : 0;
assign detect_max[180][14] = (mid_1[1455:1448] > mid_2[1447:1440]) ? 1 : 0;
assign detect_max[180][15] = (mid_1[1455:1448] > mid_2[1455:1448]) ? 1 : 0;
assign detect_max[180][16] = (mid_1[1455:1448] > mid_2[1463:1456]) ? 1 : 0;
assign detect_max[180][17] = (mid_1[1455:1448] > btm_0[1447:1440]) ? 1 : 0;
assign detect_max[180][18] = (mid_1[1455:1448] > btm_0[1455:1448]) ? 1 : 0;
assign detect_max[180][19] = (mid_1[1455:1448] > btm_0[1463:1456]) ? 1 : 0;
assign detect_max[180][20] = (mid_1[1455:1448] > btm_1[1447:1440]) ? 1 : 0;
assign detect_max[180][21] = (mid_1[1455:1448] > btm_1[1455:1448]) ? 1 : 0;
assign detect_max[180][22] = (mid_1[1455:1448] > btm_1[1463:1456]) ? 1 : 0;
assign detect_max[180][23] = (mid_1[1455:1448] > btm_2[1447:1440]) ? 1 : 0;
assign detect_max[180][24] = (mid_1[1455:1448] > btm_2[1455:1448]) ? 1 : 0;
assign detect_max[180][25] = (mid_1[1455:1448] > btm_2[1463:1456]) ? 1 : 0;

assign detect_max[181][0] = (mid_1[1463:1456] > top_0[1455:1448]) ? 1 : 0;
assign detect_max[181][1] = (mid_1[1463:1456] > top_0[1463:1456]) ? 1 : 0;
assign detect_max[181][2] = (mid_1[1463:1456] > top_0[1471:1464]) ? 1 : 0;
assign detect_max[181][3] = (mid_1[1463:1456] > top_1[1455:1448]) ? 1 : 0;
assign detect_max[181][4] = (mid_1[1463:1456] > top_1[1463:1456]) ? 1 : 0;
assign detect_max[181][5] = (mid_1[1463:1456] > top_1[1471:1464]) ? 1 : 0;
assign detect_max[181][6] = (mid_1[1463:1456] > top_2[1455:1448]) ? 1 : 0;
assign detect_max[181][7] = (mid_1[1463:1456] > top_2[1463:1456]) ? 1 : 0;
assign detect_max[181][8] = (mid_1[1463:1456] > top_2[1471:1464]) ? 1 : 0;
assign detect_max[181][9] = (mid_1[1463:1456] > mid_0[1455:1448]) ? 1 : 0;
assign detect_max[181][10] = (mid_1[1463:1456] > mid_0[1463:1456]) ? 1 : 0;
assign detect_max[181][11] = (mid_1[1463:1456] > mid_0[1471:1464]) ? 1 : 0;
assign detect_max[181][12] = (mid_1[1463:1456] > mid_1[1455:1448]) ? 1 : 0;
assign detect_max[181][13] = (mid_1[1463:1456] > mid_1[1471:1464]) ? 1 : 0;
assign detect_max[181][14] = (mid_1[1463:1456] > mid_2[1455:1448]) ? 1 : 0;
assign detect_max[181][15] = (mid_1[1463:1456] > mid_2[1463:1456]) ? 1 : 0;
assign detect_max[181][16] = (mid_1[1463:1456] > mid_2[1471:1464]) ? 1 : 0;
assign detect_max[181][17] = (mid_1[1463:1456] > btm_0[1455:1448]) ? 1 : 0;
assign detect_max[181][18] = (mid_1[1463:1456] > btm_0[1463:1456]) ? 1 : 0;
assign detect_max[181][19] = (mid_1[1463:1456] > btm_0[1471:1464]) ? 1 : 0;
assign detect_max[181][20] = (mid_1[1463:1456] > btm_1[1455:1448]) ? 1 : 0;
assign detect_max[181][21] = (mid_1[1463:1456] > btm_1[1463:1456]) ? 1 : 0;
assign detect_max[181][22] = (mid_1[1463:1456] > btm_1[1471:1464]) ? 1 : 0;
assign detect_max[181][23] = (mid_1[1463:1456] > btm_2[1455:1448]) ? 1 : 0;
assign detect_max[181][24] = (mid_1[1463:1456] > btm_2[1463:1456]) ? 1 : 0;
assign detect_max[181][25] = (mid_1[1463:1456] > btm_2[1471:1464]) ? 1 : 0;

assign detect_max[182][0] = (mid_1[1471:1464] > top_0[1463:1456]) ? 1 : 0;
assign detect_max[182][1] = (mid_1[1471:1464] > top_0[1471:1464]) ? 1 : 0;
assign detect_max[182][2] = (mid_1[1471:1464] > top_0[1479:1472]) ? 1 : 0;
assign detect_max[182][3] = (mid_1[1471:1464] > top_1[1463:1456]) ? 1 : 0;
assign detect_max[182][4] = (mid_1[1471:1464] > top_1[1471:1464]) ? 1 : 0;
assign detect_max[182][5] = (mid_1[1471:1464] > top_1[1479:1472]) ? 1 : 0;
assign detect_max[182][6] = (mid_1[1471:1464] > top_2[1463:1456]) ? 1 : 0;
assign detect_max[182][7] = (mid_1[1471:1464] > top_2[1471:1464]) ? 1 : 0;
assign detect_max[182][8] = (mid_1[1471:1464] > top_2[1479:1472]) ? 1 : 0;
assign detect_max[182][9] = (mid_1[1471:1464] > mid_0[1463:1456]) ? 1 : 0;
assign detect_max[182][10] = (mid_1[1471:1464] > mid_0[1471:1464]) ? 1 : 0;
assign detect_max[182][11] = (mid_1[1471:1464] > mid_0[1479:1472]) ? 1 : 0;
assign detect_max[182][12] = (mid_1[1471:1464] > mid_1[1463:1456]) ? 1 : 0;
assign detect_max[182][13] = (mid_1[1471:1464] > mid_1[1479:1472]) ? 1 : 0;
assign detect_max[182][14] = (mid_1[1471:1464] > mid_2[1463:1456]) ? 1 : 0;
assign detect_max[182][15] = (mid_1[1471:1464] > mid_2[1471:1464]) ? 1 : 0;
assign detect_max[182][16] = (mid_1[1471:1464] > mid_2[1479:1472]) ? 1 : 0;
assign detect_max[182][17] = (mid_1[1471:1464] > btm_0[1463:1456]) ? 1 : 0;
assign detect_max[182][18] = (mid_1[1471:1464] > btm_0[1471:1464]) ? 1 : 0;
assign detect_max[182][19] = (mid_1[1471:1464] > btm_0[1479:1472]) ? 1 : 0;
assign detect_max[182][20] = (mid_1[1471:1464] > btm_1[1463:1456]) ? 1 : 0;
assign detect_max[182][21] = (mid_1[1471:1464] > btm_1[1471:1464]) ? 1 : 0;
assign detect_max[182][22] = (mid_1[1471:1464] > btm_1[1479:1472]) ? 1 : 0;
assign detect_max[182][23] = (mid_1[1471:1464] > btm_2[1463:1456]) ? 1 : 0;
assign detect_max[182][24] = (mid_1[1471:1464] > btm_2[1471:1464]) ? 1 : 0;
assign detect_max[182][25] = (mid_1[1471:1464] > btm_2[1479:1472]) ? 1 : 0;

assign detect_max[183][0] = (mid_1[1479:1472] > top_0[1471:1464]) ? 1 : 0;
assign detect_max[183][1] = (mid_1[1479:1472] > top_0[1479:1472]) ? 1 : 0;
assign detect_max[183][2] = (mid_1[1479:1472] > top_0[1487:1480]) ? 1 : 0;
assign detect_max[183][3] = (mid_1[1479:1472] > top_1[1471:1464]) ? 1 : 0;
assign detect_max[183][4] = (mid_1[1479:1472] > top_1[1479:1472]) ? 1 : 0;
assign detect_max[183][5] = (mid_1[1479:1472] > top_1[1487:1480]) ? 1 : 0;
assign detect_max[183][6] = (mid_1[1479:1472] > top_2[1471:1464]) ? 1 : 0;
assign detect_max[183][7] = (mid_1[1479:1472] > top_2[1479:1472]) ? 1 : 0;
assign detect_max[183][8] = (mid_1[1479:1472] > top_2[1487:1480]) ? 1 : 0;
assign detect_max[183][9] = (mid_1[1479:1472] > mid_0[1471:1464]) ? 1 : 0;
assign detect_max[183][10] = (mid_1[1479:1472] > mid_0[1479:1472]) ? 1 : 0;
assign detect_max[183][11] = (mid_1[1479:1472] > mid_0[1487:1480]) ? 1 : 0;
assign detect_max[183][12] = (mid_1[1479:1472] > mid_1[1471:1464]) ? 1 : 0;
assign detect_max[183][13] = (mid_1[1479:1472] > mid_1[1487:1480]) ? 1 : 0;
assign detect_max[183][14] = (mid_1[1479:1472] > mid_2[1471:1464]) ? 1 : 0;
assign detect_max[183][15] = (mid_1[1479:1472] > mid_2[1479:1472]) ? 1 : 0;
assign detect_max[183][16] = (mid_1[1479:1472] > mid_2[1487:1480]) ? 1 : 0;
assign detect_max[183][17] = (mid_1[1479:1472] > btm_0[1471:1464]) ? 1 : 0;
assign detect_max[183][18] = (mid_1[1479:1472] > btm_0[1479:1472]) ? 1 : 0;
assign detect_max[183][19] = (mid_1[1479:1472] > btm_0[1487:1480]) ? 1 : 0;
assign detect_max[183][20] = (mid_1[1479:1472] > btm_1[1471:1464]) ? 1 : 0;
assign detect_max[183][21] = (mid_1[1479:1472] > btm_1[1479:1472]) ? 1 : 0;
assign detect_max[183][22] = (mid_1[1479:1472] > btm_1[1487:1480]) ? 1 : 0;
assign detect_max[183][23] = (mid_1[1479:1472] > btm_2[1471:1464]) ? 1 : 0;
assign detect_max[183][24] = (mid_1[1479:1472] > btm_2[1479:1472]) ? 1 : 0;
assign detect_max[183][25] = (mid_1[1479:1472] > btm_2[1487:1480]) ? 1 : 0;

assign detect_max[184][0] = (mid_1[1487:1480] > top_0[1479:1472]) ? 1 : 0;
assign detect_max[184][1] = (mid_1[1487:1480] > top_0[1487:1480]) ? 1 : 0;
assign detect_max[184][2] = (mid_1[1487:1480] > top_0[1495:1488]) ? 1 : 0;
assign detect_max[184][3] = (mid_1[1487:1480] > top_1[1479:1472]) ? 1 : 0;
assign detect_max[184][4] = (mid_1[1487:1480] > top_1[1487:1480]) ? 1 : 0;
assign detect_max[184][5] = (mid_1[1487:1480] > top_1[1495:1488]) ? 1 : 0;
assign detect_max[184][6] = (mid_1[1487:1480] > top_2[1479:1472]) ? 1 : 0;
assign detect_max[184][7] = (mid_1[1487:1480] > top_2[1487:1480]) ? 1 : 0;
assign detect_max[184][8] = (mid_1[1487:1480] > top_2[1495:1488]) ? 1 : 0;
assign detect_max[184][9] = (mid_1[1487:1480] > mid_0[1479:1472]) ? 1 : 0;
assign detect_max[184][10] = (mid_1[1487:1480] > mid_0[1487:1480]) ? 1 : 0;
assign detect_max[184][11] = (mid_1[1487:1480] > mid_0[1495:1488]) ? 1 : 0;
assign detect_max[184][12] = (mid_1[1487:1480] > mid_1[1479:1472]) ? 1 : 0;
assign detect_max[184][13] = (mid_1[1487:1480] > mid_1[1495:1488]) ? 1 : 0;
assign detect_max[184][14] = (mid_1[1487:1480] > mid_2[1479:1472]) ? 1 : 0;
assign detect_max[184][15] = (mid_1[1487:1480] > mid_2[1487:1480]) ? 1 : 0;
assign detect_max[184][16] = (mid_1[1487:1480] > mid_2[1495:1488]) ? 1 : 0;
assign detect_max[184][17] = (mid_1[1487:1480] > btm_0[1479:1472]) ? 1 : 0;
assign detect_max[184][18] = (mid_1[1487:1480] > btm_0[1487:1480]) ? 1 : 0;
assign detect_max[184][19] = (mid_1[1487:1480] > btm_0[1495:1488]) ? 1 : 0;
assign detect_max[184][20] = (mid_1[1487:1480] > btm_1[1479:1472]) ? 1 : 0;
assign detect_max[184][21] = (mid_1[1487:1480] > btm_1[1487:1480]) ? 1 : 0;
assign detect_max[184][22] = (mid_1[1487:1480] > btm_1[1495:1488]) ? 1 : 0;
assign detect_max[184][23] = (mid_1[1487:1480] > btm_2[1479:1472]) ? 1 : 0;
assign detect_max[184][24] = (mid_1[1487:1480] > btm_2[1487:1480]) ? 1 : 0;
assign detect_max[184][25] = (mid_1[1487:1480] > btm_2[1495:1488]) ? 1 : 0;

assign detect_max[185][0] = (mid_1[1495:1488] > top_0[1487:1480]) ? 1 : 0;
assign detect_max[185][1] = (mid_1[1495:1488] > top_0[1495:1488]) ? 1 : 0;
assign detect_max[185][2] = (mid_1[1495:1488] > top_0[1503:1496]) ? 1 : 0;
assign detect_max[185][3] = (mid_1[1495:1488] > top_1[1487:1480]) ? 1 : 0;
assign detect_max[185][4] = (mid_1[1495:1488] > top_1[1495:1488]) ? 1 : 0;
assign detect_max[185][5] = (mid_1[1495:1488] > top_1[1503:1496]) ? 1 : 0;
assign detect_max[185][6] = (mid_1[1495:1488] > top_2[1487:1480]) ? 1 : 0;
assign detect_max[185][7] = (mid_1[1495:1488] > top_2[1495:1488]) ? 1 : 0;
assign detect_max[185][8] = (mid_1[1495:1488] > top_2[1503:1496]) ? 1 : 0;
assign detect_max[185][9] = (mid_1[1495:1488] > mid_0[1487:1480]) ? 1 : 0;
assign detect_max[185][10] = (mid_1[1495:1488] > mid_0[1495:1488]) ? 1 : 0;
assign detect_max[185][11] = (mid_1[1495:1488] > mid_0[1503:1496]) ? 1 : 0;
assign detect_max[185][12] = (mid_1[1495:1488] > mid_1[1487:1480]) ? 1 : 0;
assign detect_max[185][13] = (mid_1[1495:1488] > mid_1[1503:1496]) ? 1 : 0;
assign detect_max[185][14] = (mid_1[1495:1488] > mid_2[1487:1480]) ? 1 : 0;
assign detect_max[185][15] = (mid_1[1495:1488] > mid_2[1495:1488]) ? 1 : 0;
assign detect_max[185][16] = (mid_1[1495:1488] > mid_2[1503:1496]) ? 1 : 0;
assign detect_max[185][17] = (mid_1[1495:1488] > btm_0[1487:1480]) ? 1 : 0;
assign detect_max[185][18] = (mid_1[1495:1488] > btm_0[1495:1488]) ? 1 : 0;
assign detect_max[185][19] = (mid_1[1495:1488] > btm_0[1503:1496]) ? 1 : 0;
assign detect_max[185][20] = (mid_1[1495:1488] > btm_1[1487:1480]) ? 1 : 0;
assign detect_max[185][21] = (mid_1[1495:1488] > btm_1[1495:1488]) ? 1 : 0;
assign detect_max[185][22] = (mid_1[1495:1488] > btm_1[1503:1496]) ? 1 : 0;
assign detect_max[185][23] = (mid_1[1495:1488] > btm_2[1487:1480]) ? 1 : 0;
assign detect_max[185][24] = (mid_1[1495:1488] > btm_2[1495:1488]) ? 1 : 0;
assign detect_max[185][25] = (mid_1[1495:1488] > btm_2[1503:1496]) ? 1 : 0;

assign detect_max[186][0] = (mid_1[1503:1496] > top_0[1495:1488]) ? 1 : 0;
assign detect_max[186][1] = (mid_1[1503:1496] > top_0[1503:1496]) ? 1 : 0;
assign detect_max[186][2] = (mid_1[1503:1496] > top_0[1511:1504]) ? 1 : 0;
assign detect_max[186][3] = (mid_1[1503:1496] > top_1[1495:1488]) ? 1 : 0;
assign detect_max[186][4] = (mid_1[1503:1496] > top_1[1503:1496]) ? 1 : 0;
assign detect_max[186][5] = (mid_1[1503:1496] > top_1[1511:1504]) ? 1 : 0;
assign detect_max[186][6] = (mid_1[1503:1496] > top_2[1495:1488]) ? 1 : 0;
assign detect_max[186][7] = (mid_1[1503:1496] > top_2[1503:1496]) ? 1 : 0;
assign detect_max[186][8] = (mid_1[1503:1496] > top_2[1511:1504]) ? 1 : 0;
assign detect_max[186][9] = (mid_1[1503:1496] > mid_0[1495:1488]) ? 1 : 0;
assign detect_max[186][10] = (mid_1[1503:1496] > mid_0[1503:1496]) ? 1 : 0;
assign detect_max[186][11] = (mid_1[1503:1496] > mid_0[1511:1504]) ? 1 : 0;
assign detect_max[186][12] = (mid_1[1503:1496] > mid_1[1495:1488]) ? 1 : 0;
assign detect_max[186][13] = (mid_1[1503:1496] > mid_1[1511:1504]) ? 1 : 0;
assign detect_max[186][14] = (mid_1[1503:1496] > mid_2[1495:1488]) ? 1 : 0;
assign detect_max[186][15] = (mid_1[1503:1496] > mid_2[1503:1496]) ? 1 : 0;
assign detect_max[186][16] = (mid_1[1503:1496] > mid_2[1511:1504]) ? 1 : 0;
assign detect_max[186][17] = (mid_1[1503:1496] > btm_0[1495:1488]) ? 1 : 0;
assign detect_max[186][18] = (mid_1[1503:1496] > btm_0[1503:1496]) ? 1 : 0;
assign detect_max[186][19] = (mid_1[1503:1496] > btm_0[1511:1504]) ? 1 : 0;
assign detect_max[186][20] = (mid_1[1503:1496] > btm_1[1495:1488]) ? 1 : 0;
assign detect_max[186][21] = (mid_1[1503:1496] > btm_1[1503:1496]) ? 1 : 0;
assign detect_max[186][22] = (mid_1[1503:1496] > btm_1[1511:1504]) ? 1 : 0;
assign detect_max[186][23] = (mid_1[1503:1496] > btm_2[1495:1488]) ? 1 : 0;
assign detect_max[186][24] = (mid_1[1503:1496] > btm_2[1503:1496]) ? 1 : 0;
assign detect_max[186][25] = (mid_1[1503:1496] > btm_2[1511:1504]) ? 1 : 0;

assign detect_max[187][0] = (mid_1[1511:1504] > top_0[1503:1496]) ? 1 : 0;
assign detect_max[187][1] = (mid_1[1511:1504] > top_0[1511:1504]) ? 1 : 0;
assign detect_max[187][2] = (mid_1[1511:1504] > top_0[1519:1512]) ? 1 : 0;
assign detect_max[187][3] = (mid_1[1511:1504] > top_1[1503:1496]) ? 1 : 0;
assign detect_max[187][4] = (mid_1[1511:1504] > top_1[1511:1504]) ? 1 : 0;
assign detect_max[187][5] = (mid_1[1511:1504] > top_1[1519:1512]) ? 1 : 0;
assign detect_max[187][6] = (mid_1[1511:1504] > top_2[1503:1496]) ? 1 : 0;
assign detect_max[187][7] = (mid_1[1511:1504] > top_2[1511:1504]) ? 1 : 0;
assign detect_max[187][8] = (mid_1[1511:1504] > top_2[1519:1512]) ? 1 : 0;
assign detect_max[187][9] = (mid_1[1511:1504] > mid_0[1503:1496]) ? 1 : 0;
assign detect_max[187][10] = (mid_1[1511:1504] > mid_0[1511:1504]) ? 1 : 0;
assign detect_max[187][11] = (mid_1[1511:1504] > mid_0[1519:1512]) ? 1 : 0;
assign detect_max[187][12] = (mid_1[1511:1504] > mid_1[1503:1496]) ? 1 : 0;
assign detect_max[187][13] = (mid_1[1511:1504] > mid_1[1519:1512]) ? 1 : 0;
assign detect_max[187][14] = (mid_1[1511:1504] > mid_2[1503:1496]) ? 1 : 0;
assign detect_max[187][15] = (mid_1[1511:1504] > mid_2[1511:1504]) ? 1 : 0;
assign detect_max[187][16] = (mid_1[1511:1504] > mid_2[1519:1512]) ? 1 : 0;
assign detect_max[187][17] = (mid_1[1511:1504] > btm_0[1503:1496]) ? 1 : 0;
assign detect_max[187][18] = (mid_1[1511:1504] > btm_0[1511:1504]) ? 1 : 0;
assign detect_max[187][19] = (mid_1[1511:1504] > btm_0[1519:1512]) ? 1 : 0;
assign detect_max[187][20] = (mid_1[1511:1504] > btm_1[1503:1496]) ? 1 : 0;
assign detect_max[187][21] = (mid_1[1511:1504] > btm_1[1511:1504]) ? 1 : 0;
assign detect_max[187][22] = (mid_1[1511:1504] > btm_1[1519:1512]) ? 1 : 0;
assign detect_max[187][23] = (mid_1[1511:1504] > btm_2[1503:1496]) ? 1 : 0;
assign detect_max[187][24] = (mid_1[1511:1504] > btm_2[1511:1504]) ? 1 : 0;
assign detect_max[187][25] = (mid_1[1511:1504] > btm_2[1519:1512]) ? 1 : 0;

assign detect_max[188][0] = (mid_1[1519:1512] > top_0[1511:1504]) ? 1 : 0;
assign detect_max[188][1] = (mid_1[1519:1512] > top_0[1519:1512]) ? 1 : 0;
assign detect_max[188][2] = (mid_1[1519:1512] > top_0[1527:1520]) ? 1 : 0;
assign detect_max[188][3] = (mid_1[1519:1512] > top_1[1511:1504]) ? 1 : 0;
assign detect_max[188][4] = (mid_1[1519:1512] > top_1[1519:1512]) ? 1 : 0;
assign detect_max[188][5] = (mid_1[1519:1512] > top_1[1527:1520]) ? 1 : 0;
assign detect_max[188][6] = (mid_1[1519:1512] > top_2[1511:1504]) ? 1 : 0;
assign detect_max[188][7] = (mid_1[1519:1512] > top_2[1519:1512]) ? 1 : 0;
assign detect_max[188][8] = (mid_1[1519:1512] > top_2[1527:1520]) ? 1 : 0;
assign detect_max[188][9] = (mid_1[1519:1512] > mid_0[1511:1504]) ? 1 : 0;
assign detect_max[188][10] = (mid_1[1519:1512] > mid_0[1519:1512]) ? 1 : 0;
assign detect_max[188][11] = (mid_1[1519:1512] > mid_0[1527:1520]) ? 1 : 0;
assign detect_max[188][12] = (mid_1[1519:1512] > mid_1[1511:1504]) ? 1 : 0;
assign detect_max[188][13] = (mid_1[1519:1512] > mid_1[1527:1520]) ? 1 : 0;
assign detect_max[188][14] = (mid_1[1519:1512] > mid_2[1511:1504]) ? 1 : 0;
assign detect_max[188][15] = (mid_1[1519:1512] > mid_2[1519:1512]) ? 1 : 0;
assign detect_max[188][16] = (mid_1[1519:1512] > mid_2[1527:1520]) ? 1 : 0;
assign detect_max[188][17] = (mid_1[1519:1512] > btm_0[1511:1504]) ? 1 : 0;
assign detect_max[188][18] = (mid_1[1519:1512] > btm_0[1519:1512]) ? 1 : 0;
assign detect_max[188][19] = (mid_1[1519:1512] > btm_0[1527:1520]) ? 1 : 0;
assign detect_max[188][20] = (mid_1[1519:1512] > btm_1[1511:1504]) ? 1 : 0;
assign detect_max[188][21] = (mid_1[1519:1512] > btm_1[1519:1512]) ? 1 : 0;
assign detect_max[188][22] = (mid_1[1519:1512] > btm_1[1527:1520]) ? 1 : 0;
assign detect_max[188][23] = (mid_1[1519:1512] > btm_2[1511:1504]) ? 1 : 0;
assign detect_max[188][24] = (mid_1[1519:1512] > btm_2[1519:1512]) ? 1 : 0;
assign detect_max[188][25] = (mid_1[1519:1512] > btm_2[1527:1520]) ? 1 : 0;

assign detect_max[189][0] = (mid_1[1527:1520] > top_0[1519:1512]) ? 1 : 0;
assign detect_max[189][1] = (mid_1[1527:1520] > top_0[1527:1520]) ? 1 : 0;
assign detect_max[189][2] = (mid_1[1527:1520] > top_0[1535:1528]) ? 1 : 0;
assign detect_max[189][3] = (mid_1[1527:1520] > top_1[1519:1512]) ? 1 : 0;
assign detect_max[189][4] = (mid_1[1527:1520] > top_1[1527:1520]) ? 1 : 0;
assign detect_max[189][5] = (mid_1[1527:1520] > top_1[1535:1528]) ? 1 : 0;
assign detect_max[189][6] = (mid_1[1527:1520] > top_2[1519:1512]) ? 1 : 0;
assign detect_max[189][7] = (mid_1[1527:1520] > top_2[1527:1520]) ? 1 : 0;
assign detect_max[189][8] = (mid_1[1527:1520] > top_2[1535:1528]) ? 1 : 0;
assign detect_max[189][9] = (mid_1[1527:1520] > mid_0[1519:1512]) ? 1 : 0;
assign detect_max[189][10] = (mid_1[1527:1520] > mid_0[1527:1520]) ? 1 : 0;
assign detect_max[189][11] = (mid_1[1527:1520] > mid_0[1535:1528]) ? 1 : 0;
assign detect_max[189][12] = (mid_1[1527:1520] > mid_1[1519:1512]) ? 1 : 0;
assign detect_max[189][13] = (mid_1[1527:1520] > mid_1[1535:1528]) ? 1 : 0;
assign detect_max[189][14] = (mid_1[1527:1520] > mid_2[1519:1512]) ? 1 : 0;
assign detect_max[189][15] = (mid_1[1527:1520] > mid_2[1527:1520]) ? 1 : 0;
assign detect_max[189][16] = (mid_1[1527:1520] > mid_2[1535:1528]) ? 1 : 0;
assign detect_max[189][17] = (mid_1[1527:1520] > btm_0[1519:1512]) ? 1 : 0;
assign detect_max[189][18] = (mid_1[1527:1520] > btm_0[1527:1520]) ? 1 : 0;
assign detect_max[189][19] = (mid_1[1527:1520] > btm_0[1535:1528]) ? 1 : 0;
assign detect_max[189][20] = (mid_1[1527:1520] > btm_1[1519:1512]) ? 1 : 0;
assign detect_max[189][21] = (mid_1[1527:1520] > btm_1[1527:1520]) ? 1 : 0;
assign detect_max[189][22] = (mid_1[1527:1520] > btm_1[1535:1528]) ? 1 : 0;
assign detect_max[189][23] = (mid_1[1527:1520] > btm_2[1519:1512]) ? 1 : 0;
assign detect_max[189][24] = (mid_1[1527:1520] > btm_2[1527:1520]) ? 1 : 0;
assign detect_max[189][25] = (mid_1[1527:1520] > btm_2[1535:1528]) ? 1 : 0;

assign detect_max[190][0] = (mid_1[1535:1528] > top_0[1527:1520]) ? 1 : 0;
assign detect_max[190][1] = (mid_1[1535:1528] > top_0[1535:1528]) ? 1 : 0;
assign detect_max[190][2] = (mid_1[1535:1528] > top_0[1543:1536]) ? 1 : 0;
assign detect_max[190][3] = (mid_1[1535:1528] > top_1[1527:1520]) ? 1 : 0;
assign detect_max[190][4] = (mid_1[1535:1528] > top_1[1535:1528]) ? 1 : 0;
assign detect_max[190][5] = (mid_1[1535:1528] > top_1[1543:1536]) ? 1 : 0;
assign detect_max[190][6] = (mid_1[1535:1528] > top_2[1527:1520]) ? 1 : 0;
assign detect_max[190][7] = (mid_1[1535:1528] > top_2[1535:1528]) ? 1 : 0;
assign detect_max[190][8] = (mid_1[1535:1528] > top_2[1543:1536]) ? 1 : 0;
assign detect_max[190][9] = (mid_1[1535:1528] > mid_0[1527:1520]) ? 1 : 0;
assign detect_max[190][10] = (mid_1[1535:1528] > mid_0[1535:1528]) ? 1 : 0;
assign detect_max[190][11] = (mid_1[1535:1528] > mid_0[1543:1536]) ? 1 : 0;
assign detect_max[190][12] = (mid_1[1535:1528] > mid_1[1527:1520]) ? 1 : 0;
assign detect_max[190][13] = (mid_1[1535:1528] > mid_1[1543:1536]) ? 1 : 0;
assign detect_max[190][14] = (mid_1[1535:1528] > mid_2[1527:1520]) ? 1 : 0;
assign detect_max[190][15] = (mid_1[1535:1528] > mid_2[1535:1528]) ? 1 : 0;
assign detect_max[190][16] = (mid_1[1535:1528] > mid_2[1543:1536]) ? 1 : 0;
assign detect_max[190][17] = (mid_1[1535:1528] > btm_0[1527:1520]) ? 1 : 0;
assign detect_max[190][18] = (mid_1[1535:1528] > btm_0[1535:1528]) ? 1 : 0;
assign detect_max[190][19] = (mid_1[1535:1528] > btm_0[1543:1536]) ? 1 : 0;
assign detect_max[190][20] = (mid_1[1535:1528] > btm_1[1527:1520]) ? 1 : 0;
assign detect_max[190][21] = (mid_1[1535:1528] > btm_1[1535:1528]) ? 1 : 0;
assign detect_max[190][22] = (mid_1[1535:1528] > btm_1[1543:1536]) ? 1 : 0;
assign detect_max[190][23] = (mid_1[1535:1528] > btm_2[1527:1520]) ? 1 : 0;
assign detect_max[190][24] = (mid_1[1535:1528] > btm_2[1535:1528]) ? 1 : 0;
assign detect_max[190][25] = (mid_1[1535:1528] > btm_2[1543:1536]) ? 1 : 0;

assign detect_max[191][0] = (mid_1[1543:1536] > top_0[1535:1528]) ? 1 : 0;
assign detect_max[191][1] = (mid_1[1543:1536] > top_0[1543:1536]) ? 1 : 0;
assign detect_max[191][2] = (mid_1[1543:1536] > top_0[1551:1544]) ? 1 : 0;
assign detect_max[191][3] = (mid_1[1543:1536] > top_1[1535:1528]) ? 1 : 0;
assign detect_max[191][4] = (mid_1[1543:1536] > top_1[1543:1536]) ? 1 : 0;
assign detect_max[191][5] = (mid_1[1543:1536] > top_1[1551:1544]) ? 1 : 0;
assign detect_max[191][6] = (mid_1[1543:1536] > top_2[1535:1528]) ? 1 : 0;
assign detect_max[191][7] = (mid_1[1543:1536] > top_2[1543:1536]) ? 1 : 0;
assign detect_max[191][8] = (mid_1[1543:1536] > top_2[1551:1544]) ? 1 : 0;
assign detect_max[191][9] = (mid_1[1543:1536] > mid_0[1535:1528]) ? 1 : 0;
assign detect_max[191][10] = (mid_1[1543:1536] > mid_0[1543:1536]) ? 1 : 0;
assign detect_max[191][11] = (mid_1[1543:1536] > mid_0[1551:1544]) ? 1 : 0;
assign detect_max[191][12] = (mid_1[1543:1536] > mid_1[1535:1528]) ? 1 : 0;
assign detect_max[191][13] = (mid_1[1543:1536] > mid_1[1551:1544]) ? 1 : 0;
assign detect_max[191][14] = (mid_1[1543:1536] > mid_2[1535:1528]) ? 1 : 0;
assign detect_max[191][15] = (mid_1[1543:1536] > mid_2[1543:1536]) ? 1 : 0;
assign detect_max[191][16] = (mid_1[1543:1536] > mid_2[1551:1544]) ? 1 : 0;
assign detect_max[191][17] = (mid_1[1543:1536] > btm_0[1535:1528]) ? 1 : 0;
assign detect_max[191][18] = (mid_1[1543:1536] > btm_0[1543:1536]) ? 1 : 0;
assign detect_max[191][19] = (mid_1[1543:1536] > btm_0[1551:1544]) ? 1 : 0;
assign detect_max[191][20] = (mid_1[1543:1536] > btm_1[1535:1528]) ? 1 : 0;
assign detect_max[191][21] = (mid_1[1543:1536] > btm_1[1543:1536]) ? 1 : 0;
assign detect_max[191][22] = (mid_1[1543:1536] > btm_1[1551:1544]) ? 1 : 0;
assign detect_max[191][23] = (mid_1[1543:1536] > btm_2[1535:1528]) ? 1 : 0;
assign detect_max[191][24] = (mid_1[1543:1536] > btm_2[1543:1536]) ? 1 : 0;
assign detect_max[191][25] = (mid_1[1543:1536] > btm_2[1551:1544]) ? 1 : 0;

assign detect_max[192][0] = (mid_1[1551:1544] > top_0[1543:1536]) ? 1 : 0;
assign detect_max[192][1] = (mid_1[1551:1544] > top_0[1551:1544]) ? 1 : 0;
assign detect_max[192][2] = (mid_1[1551:1544] > top_0[1559:1552]) ? 1 : 0;
assign detect_max[192][3] = (mid_1[1551:1544] > top_1[1543:1536]) ? 1 : 0;
assign detect_max[192][4] = (mid_1[1551:1544] > top_1[1551:1544]) ? 1 : 0;
assign detect_max[192][5] = (mid_1[1551:1544] > top_1[1559:1552]) ? 1 : 0;
assign detect_max[192][6] = (mid_1[1551:1544] > top_2[1543:1536]) ? 1 : 0;
assign detect_max[192][7] = (mid_1[1551:1544] > top_2[1551:1544]) ? 1 : 0;
assign detect_max[192][8] = (mid_1[1551:1544] > top_2[1559:1552]) ? 1 : 0;
assign detect_max[192][9] = (mid_1[1551:1544] > mid_0[1543:1536]) ? 1 : 0;
assign detect_max[192][10] = (mid_1[1551:1544] > mid_0[1551:1544]) ? 1 : 0;
assign detect_max[192][11] = (mid_1[1551:1544] > mid_0[1559:1552]) ? 1 : 0;
assign detect_max[192][12] = (mid_1[1551:1544] > mid_1[1543:1536]) ? 1 : 0;
assign detect_max[192][13] = (mid_1[1551:1544] > mid_1[1559:1552]) ? 1 : 0;
assign detect_max[192][14] = (mid_1[1551:1544] > mid_2[1543:1536]) ? 1 : 0;
assign detect_max[192][15] = (mid_1[1551:1544] > mid_2[1551:1544]) ? 1 : 0;
assign detect_max[192][16] = (mid_1[1551:1544] > mid_2[1559:1552]) ? 1 : 0;
assign detect_max[192][17] = (mid_1[1551:1544] > btm_0[1543:1536]) ? 1 : 0;
assign detect_max[192][18] = (mid_1[1551:1544] > btm_0[1551:1544]) ? 1 : 0;
assign detect_max[192][19] = (mid_1[1551:1544] > btm_0[1559:1552]) ? 1 : 0;
assign detect_max[192][20] = (mid_1[1551:1544] > btm_1[1543:1536]) ? 1 : 0;
assign detect_max[192][21] = (mid_1[1551:1544] > btm_1[1551:1544]) ? 1 : 0;
assign detect_max[192][22] = (mid_1[1551:1544] > btm_1[1559:1552]) ? 1 : 0;
assign detect_max[192][23] = (mid_1[1551:1544] > btm_2[1543:1536]) ? 1 : 0;
assign detect_max[192][24] = (mid_1[1551:1544] > btm_2[1551:1544]) ? 1 : 0;
assign detect_max[192][25] = (mid_1[1551:1544] > btm_2[1559:1552]) ? 1 : 0;

assign detect_max[193][0] = (mid_1[1559:1552] > top_0[1551:1544]) ? 1 : 0;
assign detect_max[193][1] = (mid_1[1559:1552] > top_0[1559:1552]) ? 1 : 0;
assign detect_max[193][2] = (mid_1[1559:1552] > top_0[1567:1560]) ? 1 : 0;
assign detect_max[193][3] = (mid_1[1559:1552] > top_1[1551:1544]) ? 1 : 0;
assign detect_max[193][4] = (mid_1[1559:1552] > top_1[1559:1552]) ? 1 : 0;
assign detect_max[193][5] = (mid_1[1559:1552] > top_1[1567:1560]) ? 1 : 0;
assign detect_max[193][6] = (mid_1[1559:1552] > top_2[1551:1544]) ? 1 : 0;
assign detect_max[193][7] = (mid_1[1559:1552] > top_2[1559:1552]) ? 1 : 0;
assign detect_max[193][8] = (mid_1[1559:1552] > top_2[1567:1560]) ? 1 : 0;
assign detect_max[193][9] = (mid_1[1559:1552] > mid_0[1551:1544]) ? 1 : 0;
assign detect_max[193][10] = (mid_1[1559:1552] > mid_0[1559:1552]) ? 1 : 0;
assign detect_max[193][11] = (mid_1[1559:1552] > mid_0[1567:1560]) ? 1 : 0;
assign detect_max[193][12] = (mid_1[1559:1552] > mid_1[1551:1544]) ? 1 : 0;
assign detect_max[193][13] = (mid_1[1559:1552] > mid_1[1567:1560]) ? 1 : 0;
assign detect_max[193][14] = (mid_1[1559:1552] > mid_2[1551:1544]) ? 1 : 0;
assign detect_max[193][15] = (mid_1[1559:1552] > mid_2[1559:1552]) ? 1 : 0;
assign detect_max[193][16] = (mid_1[1559:1552] > mid_2[1567:1560]) ? 1 : 0;
assign detect_max[193][17] = (mid_1[1559:1552] > btm_0[1551:1544]) ? 1 : 0;
assign detect_max[193][18] = (mid_1[1559:1552] > btm_0[1559:1552]) ? 1 : 0;
assign detect_max[193][19] = (mid_1[1559:1552] > btm_0[1567:1560]) ? 1 : 0;
assign detect_max[193][20] = (mid_1[1559:1552] > btm_1[1551:1544]) ? 1 : 0;
assign detect_max[193][21] = (mid_1[1559:1552] > btm_1[1559:1552]) ? 1 : 0;
assign detect_max[193][22] = (mid_1[1559:1552] > btm_1[1567:1560]) ? 1 : 0;
assign detect_max[193][23] = (mid_1[1559:1552] > btm_2[1551:1544]) ? 1 : 0;
assign detect_max[193][24] = (mid_1[1559:1552] > btm_2[1559:1552]) ? 1 : 0;
assign detect_max[193][25] = (mid_1[1559:1552] > btm_2[1567:1560]) ? 1 : 0;

assign detect_max[194][0] = (mid_1[1567:1560] > top_0[1559:1552]) ? 1 : 0;
assign detect_max[194][1] = (mid_1[1567:1560] > top_0[1567:1560]) ? 1 : 0;
assign detect_max[194][2] = (mid_1[1567:1560] > top_0[1575:1568]) ? 1 : 0;
assign detect_max[194][3] = (mid_1[1567:1560] > top_1[1559:1552]) ? 1 : 0;
assign detect_max[194][4] = (mid_1[1567:1560] > top_1[1567:1560]) ? 1 : 0;
assign detect_max[194][5] = (mid_1[1567:1560] > top_1[1575:1568]) ? 1 : 0;
assign detect_max[194][6] = (mid_1[1567:1560] > top_2[1559:1552]) ? 1 : 0;
assign detect_max[194][7] = (mid_1[1567:1560] > top_2[1567:1560]) ? 1 : 0;
assign detect_max[194][8] = (mid_1[1567:1560] > top_2[1575:1568]) ? 1 : 0;
assign detect_max[194][9] = (mid_1[1567:1560] > mid_0[1559:1552]) ? 1 : 0;
assign detect_max[194][10] = (mid_1[1567:1560] > mid_0[1567:1560]) ? 1 : 0;
assign detect_max[194][11] = (mid_1[1567:1560] > mid_0[1575:1568]) ? 1 : 0;
assign detect_max[194][12] = (mid_1[1567:1560] > mid_1[1559:1552]) ? 1 : 0;
assign detect_max[194][13] = (mid_1[1567:1560] > mid_1[1575:1568]) ? 1 : 0;
assign detect_max[194][14] = (mid_1[1567:1560] > mid_2[1559:1552]) ? 1 : 0;
assign detect_max[194][15] = (mid_1[1567:1560] > mid_2[1567:1560]) ? 1 : 0;
assign detect_max[194][16] = (mid_1[1567:1560] > mid_2[1575:1568]) ? 1 : 0;
assign detect_max[194][17] = (mid_1[1567:1560] > btm_0[1559:1552]) ? 1 : 0;
assign detect_max[194][18] = (mid_1[1567:1560] > btm_0[1567:1560]) ? 1 : 0;
assign detect_max[194][19] = (mid_1[1567:1560] > btm_0[1575:1568]) ? 1 : 0;
assign detect_max[194][20] = (mid_1[1567:1560] > btm_1[1559:1552]) ? 1 : 0;
assign detect_max[194][21] = (mid_1[1567:1560] > btm_1[1567:1560]) ? 1 : 0;
assign detect_max[194][22] = (mid_1[1567:1560] > btm_1[1575:1568]) ? 1 : 0;
assign detect_max[194][23] = (mid_1[1567:1560] > btm_2[1559:1552]) ? 1 : 0;
assign detect_max[194][24] = (mid_1[1567:1560] > btm_2[1567:1560]) ? 1 : 0;
assign detect_max[194][25] = (mid_1[1567:1560] > btm_2[1575:1568]) ? 1 : 0;

assign detect_max[195][0] = (mid_1[1575:1568] > top_0[1567:1560]) ? 1 : 0;
assign detect_max[195][1] = (mid_1[1575:1568] > top_0[1575:1568]) ? 1 : 0;
assign detect_max[195][2] = (mid_1[1575:1568] > top_0[1583:1576]) ? 1 : 0;
assign detect_max[195][3] = (mid_1[1575:1568] > top_1[1567:1560]) ? 1 : 0;
assign detect_max[195][4] = (mid_1[1575:1568] > top_1[1575:1568]) ? 1 : 0;
assign detect_max[195][5] = (mid_1[1575:1568] > top_1[1583:1576]) ? 1 : 0;
assign detect_max[195][6] = (mid_1[1575:1568] > top_2[1567:1560]) ? 1 : 0;
assign detect_max[195][7] = (mid_1[1575:1568] > top_2[1575:1568]) ? 1 : 0;
assign detect_max[195][8] = (mid_1[1575:1568] > top_2[1583:1576]) ? 1 : 0;
assign detect_max[195][9] = (mid_1[1575:1568] > mid_0[1567:1560]) ? 1 : 0;
assign detect_max[195][10] = (mid_1[1575:1568] > mid_0[1575:1568]) ? 1 : 0;
assign detect_max[195][11] = (mid_1[1575:1568] > mid_0[1583:1576]) ? 1 : 0;
assign detect_max[195][12] = (mid_1[1575:1568] > mid_1[1567:1560]) ? 1 : 0;
assign detect_max[195][13] = (mid_1[1575:1568] > mid_1[1583:1576]) ? 1 : 0;
assign detect_max[195][14] = (mid_1[1575:1568] > mid_2[1567:1560]) ? 1 : 0;
assign detect_max[195][15] = (mid_1[1575:1568] > mid_2[1575:1568]) ? 1 : 0;
assign detect_max[195][16] = (mid_1[1575:1568] > mid_2[1583:1576]) ? 1 : 0;
assign detect_max[195][17] = (mid_1[1575:1568] > btm_0[1567:1560]) ? 1 : 0;
assign detect_max[195][18] = (mid_1[1575:1568] > btm_0[1575:1568]) ? 1 : 0;
assign detect_max[195][19] = (mid_1[1575:1568] > btm_0[1583:1576]) ? 1 : 0;
assign detect_max[195][20] = (mid_1[1575:1568] > btm_1[1567:1560]) ? 1 : 0;
assign detect_max[195][21] = (mid_1[1575:1568] > btm_1[1575:1568]) ? 1 : 0;
assign detect_max[195][22] = (mid_1[1575:1568] > btm_1[1583:1576]) ? 1 : 0;
assign detect_max[195][23] = (mid_1[1575:1568] > btm_2[1567:1560]) ? 1 : 0;
assign detect_max[195][24] = (mid_1[1575:1568] > btm_2[1575:1568]) ? 1 : 0;
assign detect_max[195][25] = (mid_1[1575:1568] > btm_2[1583:1576]) ? 1 : 0;

assign detect_max[196][0] = (mid_1[1583:1576] > top_0[1575:1568]) ? 1 : 0;
assign detect_max[196][1] = (mid_1[1583:1576] > top_0[1583:1576]) ? 1 : 0;
assign detect_max[196][2] = (mid_1[1583:1576] > top_0[1591:1584]) ? 1 : 0;
assign detect_max[196][3] = (mid_1[1583:1576] > top_1[1575:1568]) ? 1 : 0;
assign detect_max[196][4] = (mid_1[1583:1576] > top_1[1583:1576]) ? 1 : 0;
assign detect_max[196][5] = (mid_1[1583:1576] > top_1[1591:1584]) ? 1 : 0;
assign detect_max[196][6] = (mid_1[1583:1576] > top_2[1575:1568]) ? 1 : 0;
assign detect_max[196][7] = (mid_1[1583:1576] > top_2[1583:1576]) ? 1 : 0;
assign detect_max[196][8] = (mid_1[1583:1576] > top_2[1591:1584]) ? 1 : 0;
assign detect_max[196][9] = (mid_1[1583:1576] > mid_0[1575:1568]) ? 1 : 0;
assign detect_max[196][10] = (mid_1[1583:1576] > mid_0[1583:1576]) ? 1 : 0;
assign detect_max[196][11] = (mid_1[1583:1576] > mid_0[1591:1584]) ? 1 : 0;
assign detect_max[196][12] = (mid_1[1583:1576] > mid_1[1575:1568]) ? 1 : 0;
assign detect_max[196][13] = (mid_1[1583:1576] > mid_1[1591:1584]) ? 1 : 0;
assign detect_max[196][14] = (mid_1[1583:1576] > mid_2[1575:1568]) ? 1 : 0;
assign detect_max[196][15] = (mid_1[1583:1576] > mid_2[1583:1576]) ? 1 : 0;
assign detect_max[196][16] = (mid_1[1583:1576] > mid_2[1591:1584]) ? 1 : 0;
assign detect_max[196][17] = (mid_1[1583:1576] > btm_0[1575:1568]) ? 1 : 0;
assign detect_max[196][18] = (mid_1[1583:1576] > btm_0[1583:1576]) ? 1 : 0;
assign detect_max[196][19] = (mid_1[1583:1576] > btm_0[1591:1584]) ? 1 : 0;
assign detect_max[196][20] = (mid_1[1583:1576] > btm_1[1575:1568]) ? 1 : 0;
assign detect_max[196][21] = (mid_1[1583:1576] > btm_1[1583:1576]) ? 1 : 0;
assign detect_max[196][22] = (mid_1[1583:1576] > btm_1[1591:1584]) ? 1 : 0;
assign detect_max[196][23] = (mid_1[1583:1576] > btm_2[1575:1568]) ? 1 : 0;
assign detect_max[196][24] = (mid_1[1583:1576] > btm_2[1583:1576]) ? 1 : 0;
assign detect_max[196][25] = (mid_1[1583:1576] > btm_2[1591:1584]) ? 1 : 0;

assign detect_max[197][0] = (mid_1[1591:1584] > top_0[1583:1576]) ? 1 : 0;
assign detect_max[197][1] = (mid_1[1591:1584] > top_0[1591:1584]) ? 1 : 0;
assign detect_max[197][2] = (mid_1[1591:1584] > top_0[1599:1592]) ? 1 : 0;
assign detect_max[197][3] = (mid_1[1591:1584] > top_1[1583:1576]) ? 1 : 0;
assign detect_max[197][4] = (mid_1[1591:1584] > top_1[1591:1584]) ? 1 : 0;
assign detect_max[197][5] = (mid_1[1591:1584] > top_1[1599:1592]) ? 1 : 0;
assign detect_max[197][6] = (mid_1[1591:1584] > top_2[1583:1576]) ? 1 : 0;
assign detect_max[197][7] = (mid_1[1591:1584] > top_2[1591:1584]) ? 1 : 0;
assign detect_max[197][8] = (mid_1[1591:1584] > top_2[1599:1592]) ? 1 : 0;
assign detect_max[197][9] = (mid_1[1591:1584] > mid_0[1583:1576]) ? 1 : 0;
assign detect_max[197][10] = (mid_1[1591:1584] > mid_0[1591:1584]) ? 1 : 0;
assign detect_max[197][11] = (mid_1[1591:1584] > mid_0[1599:1592]) ? 1 : 0;
assign detect_max[197][12] = (mid_1[1591:1584] > mid_1[1583:1576]) ? 1 : 0;
assign detect_max[197][13] = (mid_1[1591:1584] > mid_1[1599:1592]) ? 1 : 0;
assign detect_max[197][14] = (mid_1[1591:1584] > mid_2[1583:1576]) ? 1 : 0;
assign detect_max[197][15] = (mid_1[1591:1584] > mid_2[1591:1584]) ? 1 : 0;
assign detect_max[197][16] = (mid_1[1591:1584] > mid_2[1599:1592]) ? 1 : 0;
assign detect_max[197][17] = (mid_1[1591:1584] > btm_0[1583:1576]) ? 1 : 0;
assign detect_max[197][18] = (mid_1[1591:1584] > btm_0[1591:1584]) ? 1 : 0;
assign detect_max[197][19] = (mid_1[1591:1584] > btm_0[1599:1592]) ? 1 : 0;
assign detect_max[197][20] = (mid_1[1591:1584] > btm_1[1583:1576]) ? 1 : 0;
assign detect_max[197][21] = (mid_1[1591:1584] > btm_1[1591:1584]) ? 1 : 0;
assign detect_max[197][22] = (mid_1[1591:1584] > btm_1[1599:1592]) ? 1 : 0;
assign detect_max[197][23] = (mid_1[1591:1584] > btm_2[1583:1576]) ? 1 : 0;
assign detect_max[197][24] = (mid_1[1591:1584] > btm_2[1591:1584]) ? 1 : 0;
assign detect_max[197][25] = (mid_1[1591:1584] > btm_2[1599:1592]) ? 1 : 0;

assign detect_max[198][0] = (mid_1[1599:1592] > top_0[1591:1584]) ? 1 : 0;
assign detect_max[198][1] = (mid_1[1599:1592] > top_0[1599:1592]) ? 1 : 0;
assign detect_max[198][2] = (mid_1[1599:1592] > top_0[1607:1600]) ? 1 : 0;
assign detect_max[198][3] = (mid_1[1599:1592] > top_1[1591:1584]) ? 1 : 0;
assign detect_max[198][4] = (mid_1[1599:1592] > top_1[1599:1592]) ? 1 : 0;
assign detect_max[198][5] = (mid_1[1599:1592] > top_1[1607:1600]) ? 1 : 0;
assign detect_max[198][6] = (mid_1[1599:1592] > top_2[1591:1584]) ? 1 : 0;
assign detect_max[198][7] = (mid_1[1599:1592] > top_2[1599:1592]) ? 1 : 0;
assign detect_max[198][8] = (mid_1[1599:1592] > top_2[1607:1600]) ? 1 : 0;
assign detect_max[198][9] = (mid_1[1599:1592] > mid_0[1591:1584]) ? 1 : 0;
assign detect_max[198][10] = (mid_1[1599:1592] > mid_0[1599:1592]) ? 1 : 0;
assign detect_max[198][11] = (mid_1[1599:1592] > mid_0[1607:1600]) ? 1 : 0;
assign detect_max[198][12] = (mid_1[1599:1592] > mid_1[1591:1584]) ? 1 : 0;
assign detect_max[198][13] = (mid_1[1599:1592] > mid_1[1607:1600]) ? 1 : 0;
assign detect_max[198][14] = (mid_1[1599:1592] > mid_2[1591:1584]) ? 1 : 0;
assign detect_max[198][15] = (mid_1[1599:1592] > mid_2[1599:1592]) ? 1 : 0;
assign detect_max[198][16] = (mid_1[1599:1592] > mid_2[1607:1600]) ? 1 : 0;
assign detect_max[198][17] = (mid_1[1599:1592] > btm_0[1591:1584]) ? 1 : 0;
assign detect_max[198][18] = (mid_1[1599:1592] > btm_0[1599:1592]) ? 1 : 0;
assign detect_max[198][19] = (mid_1[1599:1592] > btm_0[1607:1600]) ? 1 : 0;
assign detect_max[198][20] = (mid_1[1599:1592] > btm_1[1591:1584]) ? 1 : 0;
assign detect_max[198][21] = (mid_1[1599:1592] > btm_1[1599:1592]) ? 1 : 0;
assign detect_max[198][22] = (mid_1[1599:1592] > btm_1[1607:1600]) ? 1 : 0;
assign detect_max[198][23] = (mid_1[1599:1592] > btm_2[1591:1584]) ? 1 : 0;
assign detect_max[198][24] = (mid_1[1599:1592] > btm_2[1599:1592]) ? 1 : 0;
assign detect_max[198][25] = (mid_1[1599:1592] > btm_2[1607:1600]) ? 1 : 0;

assign detect_max[199][0] = (mid_1[1607:1600] > top_0[1599:1592]) ? 1 : 0;
assign detect_max[199][1] = (mid_1[1607:1600] > top_0[1607:1600]) ? 1 : 0;
assign detect_max[199][2] = (mid_1[1607:1600] > top_0[1615:1608]) ? 1 : 0;
assign detect_max[199][3] = (mid_1[1607:1600] > top_1[1599:1592]) ? 1 : 0;
assign detect_max[199][4] = (mid_1[1607:1600] > top_1[1607:1600]) ? 1 : 0;
assign detect_max[199][5] = (mid_1[1607:1600] > top_1[1615:1608]) ? 1 : 0;
assign detect_max[199][6] = (mid_1[1607:1600] > top_2[1599:1592]) ? 1 : 0;
assign detect_max[199][7] = (mid_1[1607:1600] > top_2[1607:1600]) ? 1 : 0;
assign detect_max[199][8] = (mid_1[1607:1600] > top_2[1615:1608]) ? 1 : 0;
assign detect_max[199][9] = (mid_1[1607:1600] > mid_0[1599:1592]) ? 1 : 0;
assign detect_max[199][10] = (mid_1[1607:1600] > mid_0[1607:1600]) ? 1 : 0;
assign detect_max[199][11] = (mid_1[1607:1600] > mid_0[1615:1608]) ? 1 : 0;
assign detect_max[199][12] = (mid_1[1607:1600] > mid_1[1599:1592]) ? 1 : 0;
assign detect_max[199][13] = (mid_1[1607:1600] > mid_1[1615:1608]) ? 1 : 0;
assign detect_max[199][14] = (mid_1[1607:1600] > mid_2[1599:1592]) ? 1 : 0;
assign detect_max[199][15] = (mid_1[1607:1600] > mid_2[1607:1600]) ? 1 : 0;
assign detect_max[199][16] = (mid_1[1607:1600] > mid_2[1615:1608]) ? 1 : 0;
assign detect_max[199][17] = (mid_1[1607:1600] > btm_0[1599:1592]) ? 1 : 0;
assign detect_max[199][18] = (mid_1[1607:1600] > btm_0[1607:1600]) ? 1 : 0;
assign detect_max[199][19] = (mid_1[1607:1600] > btm_0[1615:1608]) ? 1 : 0;
assign detect_max[199][20] = (mid_1[1607:1600] > btm_1[1599:1592]) ? 1 : 0;
assign detect_max[199][21] = (mid_1[1607:1600] > btm_1[1607:1600]) ? 1 : 0;
assign detect_max[199][22] = (mid_1[1607:1600] > btm_1[1615:1608]) ? 1 : 0;
assign detect_max[199][23] = (mid_1[1607:1600] > btm_2[1599:1592]) ? 1 : 0;
assign detect_max[199][24] = (mid_1[1607:1600] > btm_2[1607:1600]) ? 1 : 0;
assign detect_max[199][25] = (mid_1[1607:1600] > btm_2[1615:1608]) ? 1 : 0;

assign detect_max[200][0] = (mid_1[1615:1608] > top_0[1607:1600]) ? 1 : 0;
assign detect_max[200][1] = (mid_1[1615:1608] > top_0[1615:1608]) ? 1 : 0;
assign detect_max[200][2] = (mid_1[1615:1608] > top_0[1623:1616]) ? 1 : 0;
assign detect_max[200][3] = (mid_1[1615:1608] > top_1[1607:1600]) ? 1 : 0;
assign detect_max[200][4] = (mid_1[1615:1608] > top_1[1615:1608]) ? 1 : 0;
assign detect_max[200][5] = (mid_1[1615:1608] > top_1[1623:1616]) ? 1 : 0;
assign detect_max[200][6] = (mid_1[1615:1608] > top_2[1607:1600]) ? 1 : 0;
assign detect_max[200][7] = (mid_1[1615:1608] > top_2[1615:1608]) ? 1 : 0;
assign detect_max[200][8] = (mid_1[1615:1608] > top_2[1623:1616]) ? 1 : 0;
assign detect_max[200][9] = (mid_1[1615:1608] > mid_0[1607:1600]) ? 1 : 0;
assign detect_max[200][10] = (mid_1[1615:1608] > mid_0[1615:1608]) ? 1 : 0;
assign detect_max[200][11] = (mid_1[1615:1608] > mid_0[1623:1616]) ? 1 : 0;
assign detect_max[200][12] = (mid_1[1615:1608] > mid_1[1607:1600]) ? 1 : 0;
assign detect_max[200][13] = (mid_1[1615:1608] > mid_1[1623:1616]) ? 1 : 0;
assign detect_max[200][14] = (mid_1[1615:1608] > mid_2[1607:1600]) ? 1 : 0;
assign detect_max[200][15] = (mid_1[1615:1608] > mid_2[1615:1608]) ? 1 : 0;
assign detect_max[200][16] = (mid_1[1615:1608] > mid_2[1623:1616]) ? 1 : 0;
assign detect_max[200][17] = (mid_1[1615:1608] > btm_0[1607:1600]) ? 1 : 0;
assign detect_max[200][18] = (mid_1[1615:1608] > btm_0[1615:1608]) ? 1 : 0;
assign detect_max[200][19] = (mid_1[1615:1608] > btm_0[1623:1616]) ? 1 : 0;
assign detect_max[200][20] = (mid_1[1615:1608] > btm_1[1607:1600]) ? 1 : 0;
assign detect_max[200][21] = (mid_1[1615:1608] > btm_1[1615:1608]) ? 1 : 0;
assign detect_max[200][22] = (mid_1[1615:1608] > btm_1[1623:1616]) ? 1 : 0;
assign detect_max[200][23] = (mid_1[1615:1608] > btm_2[1607:1600]) ? 1 : 0;
assign detect_max[200][24] = (mid_1[1615:1608] > btm_2[1615:1608]) ? 1 : 0;
assign detect_max[200][25] = (mid_1[1615:1608] > btm_2[1623:1616]) ? 1 : 0;

assign detect_max[201][0] = (mid_1[1623:1616] > top_0[1615:1608]) ? 1 : 0;
assign detect_max[201][1] = (mid_1[1623:1616] > top_0[1623:1616]) ? 1 : 0;
assign detect_max[201][2] = (mid_1[1623:1616] > top_0[1631:1624]) ? 1 : 0;
assign detect_max[201][3] = (mid_1[1623:1616] > top_1[1615:1608]) ? 1 : 0;
assign detect_max[201][4] = (mid_1[1623:1616] > top_1[1623:1616]) ? 1 : 0;
assign detect_max[201][5] = (mid_1[1623:1616] > top_1[1631:1624]) ? 1 : 0;
assign detect_max[201][6] = (mid_1[1623:1616] > top_2[1615:1608]) ? 1 : 0;
assign detect_max[201][7] = (mid_1[1623:1616] > top_2[1623:1616]) ? 1 : 0;
assign detect_max[201][8] = (mid_1[1623:1616] > top_2[1631:1624]) ? 1 : 0;
assign detect_max[201][9] = (mid_1[1623:1616] > mid_0[1615:1608]) ? 1 : 0;
assign detect_max[201][10] = (mid_1[1623:1616] > mid_0[1623:1616]) ? 1 : 0;
assign detect_max[201][11] = (mid_1[1623:1616] > mid_0[1631:1624]) ? 1 : 0;
assign detect_max[201][12] = (mid_1[1623:1616] > mid_1[1615:1608]) ? 1 : 0;
assign detect_max[201][13] = (mid_1[1623:1616] > mid_1[1631:1624]) ? 1 : 0;
assign detect_max[201][14] = (mid_1[1623:1616] > mid_2[1615:1608]) ? 1 : 0;
assign detect_max[201][15] = (mid_1[1623:1616] > mid_2[1623:1616]) ? 1 : 0;
assign detect_max[201][16] = (mid_1[1623:1616] > mid_2[1631:1624]) ? 1 : 0;
assign detect_max[201][17] = (mid_1[1623:1616] > btm_0[1615:1608]) ? 1 : 0;
assign detect_max[201][18] = (mid_1[1623:1616] > btm_0[1623:1616]) ? 1 : 0;
assign detect_max[201][19] = (mid_1[1623:1616] > btm_0[1631:1624]) ? 1 : 0;
assign detect_max[201][20] = (mid_1[1623:1616] > btm_1[1615:1608]) ? 1 : 0;
assign detect_max[201][21] = (mid_1[1623:1616] > btm_1[1623:1616]) ? 1 : 0;
assign detect_max[201][22] = (mid_1[1623:1616] > btm_1[1631:1624]) ? 1 : 0;
assign detect_max[201][23] = (mid_1[1623:1616] > btm_2[1615:1608]) ? 1 : 0;
assign detect_max[201][24] = (mid_1[1623:1616] > btm_2[1623:1616]) ? 1 : 0;
assign detect_max[201][25] = (mid_1[1623:1616] > btm_2[1631:1624]) ? 1 : 0;

assign detect_max[202][0] = (mid_1[1631:1624] > top_0[1623:1616]) ? 1 : 0;
assign detect_max[202][1] = (mid_1[1631:1624] > top_0[1631:1624]) ? 1 : 0;
assign detect_max[202][2] = (mid_1[1631:1624] > top_0[1639:1632]) ? 1 : 0;
assign detect_max[202][3] = (mid_1[1631:1624] > top_1[1623:1616]) ? 1 : 0;
assign detect_max[202][4] = (mid_1[1631:1624] > top_1[1631:1624]) ? 1 : 0;
assign detect_max[202][5] = (mid_1[1631:1624] > top_1[1639:1632]) ? 1 : 0;
assign detect_max[202][6] = (mid_1[1631:1624] > top_2[1623:1616]) ? 1 : 0;
assign detect_max[202][7] = (mid_1[1631:1624] > top_2[1631:1624]) ? 1 : 0;
assign detect_max[202][8] = (mid_1[1631:1624] > top_2[1639:1632]) ? 1 : 0;
assign detect_max[202][9] = (mid_1[1631:1624] > mid_0[1623:1616]) ? 1 : 0;
assign detect_max[202][10] = (mid_1[1631:1624] > mid_0[1631:1624]) ? 1 : 0;
assign detect_max[202][11] = (mid_1[1631:1624] > mid_0[1639:1632]) ? 1 : 0;
assign detect_max[202][12] = (mid_1[1631:1624] > mid_1[1623:1616]) ? 1 : 0;
assign detect_max[202][13] = (mid_1[1631:1624] > mid_1[1639:1632]) ? 1 : 0;
assign detect_max[202][14] = (mid_1[1631:1624] > mid_2[1623:1616]) ? 1 : 0;
assign detect_max[202][15] = (mid_1[1631:1624] > mid_2[1631:1624]) ? 1 : 0;
assign detect_max[202][16] = (mid_1[1631:1624] > mid_2[1639:1632]) ? 1 : 0;
assign detect_max[202][17] = (mid_1[1631:1624] > btm_0[1623:1616]) ? 1 : 0;
assign detect_max[202][18] = (mid_1[1631:1624] > btm_0[1631:1624]) ? 1 : 0;
assign detect_max[202][19] = (mid_1[1631:1624] > btm_0[1639:1632]) ? 1 : 0;
assign detect_max[202][20] = (mid_1[1631:1624] > btm_1[1623:1616]) ? 1 : 0;
assign detect_max[202][21] = (mid_1[1631:1624] > btm_1[1631:1624]) ? 1 : 0;
assign detect_max[202][22] = (mid_1[1631:1624] > btm_1[1639:1632]) ? 1 : 0;
assign detect_max[202][23] = (mid_1[1631:1624] > btm_2[1623:1616]) ? 1 : 0;
assign detect_max[202][24] = (mid_1[1631:1624] > btm_2[1631:1624]) ? 1 : 0;
assign detect_max[202][25] = (mid_1[1631:1624] > btm_2[1639:1632]) ? 1 : 0;

assign detect_max[203][0] = (mid_1[1639:1632] > top_0[1631:1624]) ? 1 : 0;
assign detect_max[203][1] = (mid_1[1639:1632] > top_0[1639:1632]) ? 1 : 0;
assign detect_max[203][2] = (mid_1[1639:1632] > top_0[1647:1640]) ? 1 : 0;
assign detect_max[203][3] = (mid_1[1639:1632] > top_1[1631:1624]) ? 1 : 0;
assign detect_max[203][4] = (mid_1[1639:1632] > top_1[1639:1632]) ? 1 : 0;
assign detect_max[203][5] = (mid_1[1639:1632] > top_1[1647:1640]) ? 1 : 0;
assign detect_max[203][6] = (mid_1[1639:1632] > top_2[1631:1624]) ? 1 : 0;
assign detect_max[203][7] = (mid_1[1639:1632] > top_2[1639:1632]) ? 1 : 0;
assign detect_max[203][8] = (mid_1[1639:1632] > top_2[1647:1640]) ? 1 : 0;
assign detect_max[203][9] = (mid_1[1639:1632] > mid_0[1631:1624]) ? 1 : 0;
assign detect_max[203][10] = (mid_1[1639:1632] > mid_0[1639:1632]) ? 1 : 0;
assign detect_max[203][11] = (mid_1[1639:1632] > mid_0[1647:1640]) ? 1 : 0;
assign detect_max[203][12] = (mid_1[1639:1632] > mid_1[1631:1624]) ? 1 : 0;
assign detect_max[203][13] = (mid_1[1639:1632] > mid_1[1647:1640]) ? 1 : 0;
assign detect_max[203][14] = (mid_1[1639:1632] > mid_2[1631:1624]) ? 1 : 0;
assign detect_max[203][15] = (mid_1[1639:1632] > mid_2[1639:1632]) ? 1 : 0;
assign detect_max[203][16] = (mid_1[1639:1632] > mid_2[1647:1640]) ? 1 : 0;
assign detect_max[203][17] = (mid_1[1639:1632] > btm_0[1631:1624]) ? 1 : 0;
assign detect_max[203][18] = (mid_1[1639:1632] > btm_0[1639:1632]) ? 1 : 0;
assign detect_max[203][19] = (mid_1[1639:1632] > btm_0[1647:1640]) ? 1 : 0;
assign detect_max[203][20] = (mid_1[1639:1632] > btm_1[1631:1624]) ? 1 : 0;
assign detect_max[203][21] = (mid_1[1639:1632] > btm_1[1639:1632]) ? 1 : 0;
assign detect_max[203][22] = (mid_1[1639:1632] > btm_1[1647:1640]) ? 1 : 0;
assign detect_max[203][23] = (mid_1[1639:1632] > btm_2[1631:1624]) ? 1 : 0;
assign detect_max[203][24] = (mid_1[1639:1632] > btm_2[1639:1632]) ? 1 : 0;
assign detect_max[203][25] = (mid_1[1639:1632] > btm_2[1647:1640]) ? 1 : 0;

assign detect_max[204][0] = (mid_1[1647:1640] > top_0[1639:1632]) ? 1 : 0;
assign detect_max[204][1] = (mid_1[1647:1640] > top_0[1647:1640]) ? 1 : 0;
assign detect_max[204][2] = (mid_1[1647:1640] > top_0[1655:1648]) ? 1 : 0;
assign detect_max[204][3] = (mid_1[1647:1640] > top_1[1639:1632]) ? 1 : 0;
assign detect_max[204][4] = (mid_1[1647:1640] > top_1[1647:1640]) ? 1 : 0;
assign detect_max[204][5] = (mid_1[1647:1640] > top_1[1655:1648]) ? 1 : 0;
assign detect_max[204][6] = (mid_1[1647:1640] > top_2[1639:1632]) ? 1 : 0;
assign detect_max[204][7] = (mid_1[1647:1640] > top_2[1647:1640]) ? 1 : 0;
assign detect_max[204][8] = (mid_1[1647:1640] > top_2[1655:1648]) ? 1 : 0;
assign detect_max[204][9] = (mid_1[1647:1640] > mid_0[1639:1632]) ? 1 : 0;
assign detect_max[204][10] = (mid_1[1647:1640] > mid_0[1647:1640]) ? 1 : 0;
assign detect_max[204][11] = (mid_1[1647:1640] > mid_0[1655:1648]) ? 1 : 0;
assign detect_max[204][12] = (mid_1[1647:1640] > mid_1[1639:1632]) ? 1 : 0;
assign detect_max[204][13] = (mid_1[1647:1640] > mid_1[1655:1648]) ? 1 : 0;
assign detect_max[204][14] = (mid_1[1647:1640] > mid_2[1639:1632]) ? 1 : 0;
assign detect_max[204][15] = (mid_1[1647:1640] > mid_2[1647:1640]) ? 1 : 0;
assign detect_max[204][16] = (mid_1[1647:1640] > mid_2[1655:1648]) ? 1 : 0;
assign detect_max[204][17] = (mid_1[1647:1640] > btm_0[1639:1632]) ? 1 : 0;
assign detect_max[204][18] = (mid_1[1647:1640] > btm_0[1647:1640]) ? 1 : 0;
assign detect_max[204][19] = (mid_1[1647:1640] > btm_0[1655:1648]) ? 1 : 0;
assign detect_max[204][20] = (mid_1[1647:1640] > btm_1[1639:1632]) ? 1 : 0;
assign detect_max[204][21] = (mid_1[1647:1640] > btm_1[1647:1640]) ? 1 : 0;
assign detect_max[204][22] = (mid_1[1647:1640] > btm_1[1655:1648]) ? 1 : 0;
assign detect_max[204][23] = (mid_1[1647:1640] > btm_2[1639:1632]) ? 1 : 0;
assign detect_max[204][24] = (mid_1[1647:1640] > btm_2[1647:1640]) ? 1 : 0;
assign detect_max[204][25] = (mid_1[1647:1640] > btm_2[1655:1648]) ? 1 : 0;

assign detect_max[205][0] = (mid_1[1655:1648] > top_0[1647:1640]) ? 1 : 0;
assign detect_max[205][1] = (mid_1[1655:1648] > top_0[1655:1648]) ? 1 : 0;
assign detect_max[205][2] = (mid_1[1655:1648] > top_0[1663:1656]) ? 1 : 0;
assign detect_max[205][3] = (mid_1[1655:1648] > top_1[1647:1640]) ? 1 : 0;
assign detect_max[205][4] = (mid_1[1655:1648] > top_1[1655:1648]) ? 1 : 0;
assign detect_max[205][5] = (mid_1[1655:1648] > top_1[1663:1656]) ? 1 : 0;
assign detect_max[205][6] = (mid_1[1655:1648] > top_2[1647:1640]) ? 1 : 0;
assign detect_max[205][7] = (mid_1[1655:1648] > top_2[1655:1648]) ? 1 : 0;
assign detect_max[205][8] = (mid_1[1655:1648] > top_2[1663:1656]) ? 1 : 0;
assign detect_max[205][9] = (mid_1[1655:1648] > mid_0[1647:1640]) ? 1 : 0;
assign detect_max[205][10] = (mid_1[1655:1648] > mid_0[1655:1648]) ? 1 : 0;
assign detect_max[205][11] = (mid_1[1655:1648] > mid_0[1663:1656]) ? 1 : 0;
assign detect_max[205][12] = (mid_1[1655:1648] > mid_1[1647:1640]) ? 1 : 0;
assign detect_max[205][13] = (mid_1[1655:1648] > mid_1[1663:1656]) ? 1 : 0;
assign detect_max[205][14] = (mid_1[1655:1648] > mid_2[1647:1640]) ? 1 : 0;
assign detect_max[205][15] = (mid_1[1655:1648] > mid_2[1655:1648]) ? 1 : 0;
assign detect_max[205][16] = (mid_1[1655:1648] > mid_2[1663:1656]) ? 1 : 0;
assign detect_max[205][17] = (mid_1[1655:1648] > btm_0[1647:1640]) ? 1 : 0;
assign detect_max[205][18] = (mid_1[1655:1648] > btm_0[1655:1648]) ? 1 : 0;
assign detect_max[205][19] = (mid_1[1655:1648] > btm_0[1663:1656]) ? 1 : 0;
assign detect_max[205][20] = (mid_1[1655:1648] > btm_1[1647:1640]) ? 1 : 0;
assign detect_max[205][21] = (mid_1[1655:1648] > btm_1[1655:1648]) ? 1 : 0;
assign detect_max[205][22] = (mid_1[1655:1648] > btm_1[1663:1656]) ? 1 : 0;
assign detect_max[205][23] = (mid_1[1655:1648] > btm_2[1647:1640]) ? 1 : 0;
assign detect_max[205][24] = (mid_1[1655:1648] > btm_2[1655:1648]) ? 1 : 0;
assign detect_max[205][25] = (mid_1[1655:1648] > btm_2[1663:1656]) ? 1 : 0;

assign detect_max[206][0] = (mid_1[1663:1656] > top_0[1655:1648]) ? 1 : 0;
assign detect_max[206][1] = (mid_1[1663:1656] > top_0[1663:1656]) ? 1 : 0;
assign detect_max[206][2] = (mid_1[1663:1656] > top_0[1671:1664]) ? 1 : 0;
assign detect_max[206][3] = (mid_1[1663:1656] > top_1[1655:1648]) ? 1 : 0;
assign detect_max[206][4] = (mid_1[1663:1656] > top_1[1663:1656]) ? 1 : 0;
assign detect_max[206][5] = (mid_1[1663:1656] > top_1[1671:1664]) ? 1 : 0;
assign detect_max[206][6] = (mid_1[1663:1656] > top_2[1655:1648]) ? 1 : 0;
assign detect_max[206][7] = (mid_1[1663:1656] > top_2[1663:1656]) ? 1 : 0;
assign detect_max[206][8] = (mid_1[1663:1656] > top_2[1671:1664]) ? 1 : 0;
assign detect_max[206][9] = (mid_1[1663:1656] > mid_0[1655:1648]) ? 1 : 0;
assign detect_max[206][10] = (mid_1[1663:1656] > mid_0[1663:1656]) ? 1 : 0;
assign detect_max[206][11] = (mid_1[1663:1656] > mid_0[1671:1664]) ? 1 : 0;
assign detect_max[206][12] = (mid_1[1663:1656] > mid_1[1655:1648]) ? 1 : 0;
assign detect_max[206][13] = (mid_1[1663:1656] > mid_1[1671:1664]) ? 1 : 0;
assign detect_max[206][14] = (mid_1[1663:1656] > mid_2[1655:1648]) ? 1 : 0;
assign detect_max[206][15] = (mid_1[1663:1656] > mid_2[1663:1656]) ? 1 : 0;
assign detect_max[206][16] = (mid_1[1663:1656] > mid_2[1671:1664]) ? 1 : 0;
assign detect_max[206][17] = (mid_1[1663:1656] > btm_0[1655:1648]) ? 1 : 0;
assign detect_max[206][18] = (mid_1[1663:1656] > btm_0[1663:1656]) ? 1 : 0;
assign detect_max[206][19] = (mid_1[1663:1656] > btm_0[1671:1664]) ? 1 : 0;
assign detect_max[206][20] = (mid_1[1663:1656] > btm_1[1655:1648]) ? 1 : 0;
assign detect_max[206][21] = (mid_1[1663:1656] > btm_1[1663:1656]) ? 1 : 0;
assign detect_max[206][22] = (mid_1[1663:1656] > btm_1[1671:1664]) ? 1 : 0;
assign detect_max[206][23] = (mid_1[1663:1656] > btm_2[1655:1648]) ? 1 : 0;
assign detect_max[206][24] = (mid_1[1663:1656] > btm_2[1663:1656]) ? 1 : 0;
assign detect_max[206][25] = (mid_1[1663:1656] > btm_2[1671:1664]) ? 1 : 0;

assign detect_max[207][0] = (mid_1[1671:1664] > top_0[1663:1656]) ? 1 : 0;
assign detect_max[207][1] = (mid_1[1671:1664] > top_0[1671:1664]) ? 1 : 0;
assign detect_max[207][2] = (mid_1[1671:1664] > top_0[1679:1672]) ? 1 : 0;
assign detect_max[207][3] = (mid_1[1671:1664] > top_1[1663:1656]) ? 1 : 0;
assign detect_max[207][4] = (mid_1[1671:1664] > top_1[1671:1664]) ? 1 : 0;
assign detect_max[207][5] = (mid_1[1671:1664] > top_1[1679:1672]) ? 1 : 0;
assign detect_max[207][6] = (mid_1[1671:1664] > top_2[1663:1656]) ? 1 : 0;
assign detect_max[207][7] = (mid_1[1671:1664] > top_2[1671:1664]) ? 1 : 0;
assign detect_max[207][8] = (mid_1[1671:1664] > top_2[1679:1672]) ? 1 : 0;
assign detect_max[207][9] = (mid_1[1671:1664] > mid_0[1663:1656]) ? 1 : 0;
assign detect_max[207][10] = (mid_1[1671:1664] > mid_0[1671:1664]) ? 1 : 0;
assign detect_max[207][11] = (mid_1[1671:1664] > mid_0[1679:1672]) ? 1 : 0;
assign detect_max[207][12] = (mid_1[1671:1664] > mid_1[1663:1656]) ? 1 : 0;
assign detect_max[207][13] = (mid_1[1671:1664] > mid_1[1679:1672]) ? 1 : 0;
assign detect_max[207][14] = (mid_1[1671:1664] > mid_2[1663:1656]) ? 1 : 0;
assign detect_max[207][15] = (mid_1[1671:1664] > mid_2[1671:1664]) ? 1 : 0;
assign detect_max[207][16] = (mid_1[1671:1664] > mid_2[1679:1672]) ? 1 : 0;
assign detect_max[207][17] = (mid_1[1671:1664] > btm_0[1663:1656]) ? 1 : 0;
assign detect_max[207][18] = (mid_1[1671:1664] > btm_0[1671:1664]) ? 1 : 0;
assign detect_max[207][19] = (mid_1[1671:1664] > btm_0[1679:1672]) ? 1 : 0;
assign detect_max[207][20] = (mid_1[1671:1664] > btm_1[1663:1656]) ? 1 : 0;
assign detect_max[207][21] = (mid_1[1671:1664] > btm_1[1671:1664]) ? 1 : 0;
assign detect_max[207][22] = (mid_1[1671:1664] > btm_1[1679:1672]) ? 1 : 0;
assign detect_max[207][23] = (mid_1[1671:1664] > btm_2[1663:1656]) ? 1 : 0;
assign detect_max[207][24] = (mid_1[1671:1664] > btm_2[1671:1664]) ? 1 : 0;
assign detect_max[207][25] = (mid_1[1671:1664] > btm_2[1679:1672]) ? 1 : 0;

assign detect_max[208][0] = (mid_1[1679:1672] > top_0[1671:1664]) ? 1 : 0;
assign detect_max[208][1] = (mid_1[1679:1672] > top_0[1679:1672]) ? 1 : 0;
assign detect_max[208][2] = (mid_1[1679:1672] > top_0[1687:1680]) ? 1 : 0;
assign detect_max[208][3] = (mid_1[1679:1672] > top_1[1671:1664]) ? 1 : 0;
assign detect_max[208][4] = (mid_1[1679:1672] > top_1[1679:1672]) ? 1 : 0;
assign detect_max[208][5] = (mid_1[1679:1672] > top_1[1687:1680]) ? 1 : 0;
assign detect_max[208][6] = (mid_1[1679:1672] > top_2[1671:1664]) ? 1 : 0;
assign detect_max[208][7] = (mid_1[1679:1672] > top_2[1679:1672]) ? 1 : 0;
assign detect_max[208][8] = (mid_1[1679:1672] > top_2[1687:1680]) ? 1 : 0;
assign detect_max[208][9] = (mid_1[1679:1672] > mid_0[1671:1664]) ? 1 : 0;
assign detect_max[208][10] = (mid_1[1679:1672] > mid_0[1679:1672]) ? 1 : 0;
assign detect_max[208][11] = (mid_1[1679:1672] > mid_0[1687:1680]) ? 1 : 0;
assign detect_max[208][12] = (mid_1[1679:1672] > mid_1[1671:1664]) ? 1 : 0;
assign detect_max[208][13] = (mid_1[1679:1672] > mid_1[1687:1680]) ? 1 : 0;
assign detect_max[208][14] = (mid_1[1679:1672] > mid_2[1671:1664]) ? 1 : 0;
assign detect_max[208][15] = (mid_1[1679:1672] > mid_2[1679:1672]) ? 1 : 0;
assign detect_max[208][16] = (mid_1[1679:1672] > mid_2[1687:1680]) ? 1 : 0;
assign detect_max[208][17] = (mid_1[1679:1672] > btm_0[1671:1664]) ? 1 : 0;
assign detect_max[208][18] = (mid_1[1679:1672] > btm_0[1679:1672]) ? 1 : 0;
assign detect_max[208][19] = (mid_1[1679:1672] > btm_0[1687:1680]) ? 1 : 0;
assign detect_max[208][20] = (mid_1[1679:1672] > btm_1[1671:1664]) ? 1 : 0;
assign detect_max[208][21] = (mid_1[1679:1672] > btm_1[1679:1672]) ? 1 : 0;
assign detect_max[208][22] = (mid_1[1679:1672] > btm_1[1687:1680]) ? 1 : 0;
assign detect_max[208][23] = (mid_1[1679:1672] > btm_2[1671:1664]) ? 1 : 0;
assign detect_max[208][24] = (mid_1[1679:1672] > btm_2[1679:1672]) ? 1 : 0;
assign detect_max[208][25] = (mid_1[1679:1672] > btm_2[1687:1680]) ? 1 : 0;

assign detect_max[209][0] = (mid_1[1687:1680] > top_0[1679:1672]) ? 1 : 0;
assign detect_max[209][1] = (mid_1[1687:1680] > top_0[1687:1680]) ? 1 : 0;
assign detect_max[209][2] = (mid_1[1687:1680] > top_0[1695:1688]) ? 1 : 0;
assign detect_max[209][3] = (mid_1[1687:1680] > top_1[1679:1672]) ? 1 : 0;
assign detect_max[209][4] = (mid_1[1687:1680] > top_1[1687:1680]) ? 1 : 0;
assign detect_max[209][5] = (mid_1[1687:1680] > top_1[1695:1688]) ? 1 : 0;
assign detect_max[209][6] = (mid_1[1687:1680] > top_2[1679:1672]) ? 1 : 0;
assign detect_max[209][7] = (mid_1[1687:1680] > top_2[1687:1680]) ? 1 : 0;
assign detect_max[209][8] = (mid_1[1687:1680] > top_2[1695:1688]) ? 1 : 0;
assign detect_max[209][9] = (mid_1[1687:1680] > mid_0[1679:1672]) ? 1 : 0;
assign detect_max[209][10] = (mid_1[1687:1680] > mid_0[1687:1680]) ? 1 : 0;
assign detect_max[209][11] = (mid_1[1687:1680] > mid_0[1695:1688]) ? 1 : 0;
assign detect_max[209][12] = (mid_1[1687:1680] > mid_1[1679:1672]) ? 1 : 0;
assign detect_max[209][13] = (mid_1[1687:1680] > mid_1[1695:1688]) ? 1 : 0;
assign detect_max[209][14] = (mid_1[1687:1680] > mid_2[1679:1672]) ? 1 : 0;
assign detect_max[209][15] = (mid_1[1687:1680] > mid_2[1687:1680]) ? 1 : 0;
assign detect_max[209][16] = (mid_1[1687:1680] > mid_2[1695:1688]) ? 1 : 0;
assign detect_max[209][17] = (mid_1[1687:1680] > btm_0[1679:1672]) ? 1 : 0;
assign detect_max[209][18] = (mid_1[1687:1680] > btm_0[1687:1680]) ? 1 : 0;
assign detect_max[209][19] = (mid_1[1687:1680] > btm_0[1695:1688]) ? 1 : 0;
assign detect_max[209][20] = (mid_1[1687:1680] > btm_1[1679:1672]) ? 1 : 0;
assign detect_max[209][21] = (mid_1[1687:1680] > btm_1[1687:1680]) ? 1 : 0;
assign detect_max[209][22] = (mid_1[1687:1680] > btm_1[1695:1688]) ? 1 : 0;
assign detect_max[209][23] = (mid_1[1687:1680] > btm_2[1679:1672]) ? 1 : 0;
assign detect_max[209][24] = (mid_1[1687:1680] > btm_2[1687:1680]) ? 1 : 0;
assign detect_max[209][25] = (mid_1[1687:1680] > btm_2[1695:1688]) ? 1 : 0;

assign detect_max[210][0] = (mid_1[1695:1688] > top_0[1687:1680]) ? 1 : 0;
assign detect_max[210][1] = (mid_1[1695:1688] > top_0[1695:1688]) ? 1 : 0;
assign detect_max[210][2] = (mid_1[1695:1688] > top_0[1703:1696]) ? 1 : 0;
assign detect_max[210][3] = (mid_1[1695:1688] > top_1[1687:1680]) ? 1 : 0;
assign detect_max[210][4] = (mid_1[1695:1688] > top_1[1695:1688]) ? 1 : 0;
assign detect_max[210][5] = (mid_1[1695:1688] > top_1[1703:1696]) ? 1 : 0;
assign detect_max[210][6] = (mid_1[1695:1688] > top_2[1687:1680]) ? 1 : 0;
assign detect_max[210][7] = (mid_1[1695:1688] > top_2[1695:1688]) ? 1 : 0;
assign detect_max[210][8] = (mid_1[1695:1688] > top_2[1703:1696]) ? 1 : 0;
assign detect_max[210][9] = (mid_1[1695:1688] > mid_0[1687:1680]) ? 1 : 0;
assign detect_max[210][10] = (mid_1[1695:1688] > mid_0[1695:1688]) ? 1 : 0;
assign detect_max[210][11] = (mid_1[1695:1688] > mid_0[1703:1696]) ? 1 : 0;
assign detect_max[210][12] = (mid_1[1695:1688] > mid_1[1687:1680]) ? 1 : 0;
assign detect_max[210][13] = (mid_1[1695:1688] > mid_1[1703:1696]) ? 1 : 0;
assign detect_max[210][14] = (mid_1[1695:1688] > mid_2[1687:1680]) ? 1 : 0;
assign detect_max[210][15] = (mid_1[1695:1688] > mid_2[1695:1688]) ? 1 : 0;
assign detect_max[210][16] = (mid_1[1695:1688] > mid_2[1703:1696]) ? 1 : 0;
assign detect_max[210][17] = (mid_1[1695:1688] > btm_0[1687:1680]) ? 1 : 0;
assign detect_max[210][18] = (mid_1[1695:1688] > btm_0[1695:1688]) ? 1 : 0;
assign detect_max[210][19] = (mid_1[1695:1688] > btm_0[1703:1696]) ? 1 : 0;
assign detect_max[210][20] = (mid_1[1695:1688] > btm_1[1687:1680]) ? 1 : 0;
assign detect_max[210][21] = (mid_1[1695:1688] > btm_1[1695:1688]) ? 1 : 0;
assign detect_max[210][22] = (mid_1[1695:1688] > btm_1[1703:1696]) ? 1 : 0;
assign detect_max[210][23] = (mid_1[1695:1688] > btm_2[1687:1680]) ? 1 : 0;
assign detect_max[210][24] = (mid_1[1695:1688] > btm_2[1695:1688]) ? 1 : 0;
assign detect_max[210][25] = (mid_1[1695:1688] > btm_2[1703:1696]) ? 1 : 0;

assign detect_max[211][0] = (mid_1[1703:1696] > top_0[1695:1688]) ? 1 : 0;
assign detect_max[211][1] = (mid_1[1703:1696] > top_0[1703:1696]) ? 1 : 0;
assign detect_max[211][2] = (mid_1[1703:1696] > top_0[1711:1704]) ? 1 : 0;
assign detect_max[211][3] = (mid_1[1703:1696] > top_1[1695:1688]) ? 1 : 0;
assign detect_max[211][4] = (mid_1[1703:1696] > top_1[1703:1696]) ? 1 : 0;
assign detect_max[211][5] = (mid_1[1703:1696] > top_1[1711:1704]) ? 1 : 0;
assign detect_max[211][6] = (mid_1[1703:1696] > top_2[1695:1688]) ? 1 : 0;
assign detect_max[211][7] = (mid_1[1703:1696] > top_2[1703:1696]) ? 1 : 0;
assign detect_max[211][8] = (mid_1[1703:1696] > top_2[1711:1704]) ? 1 : 0;
assign detect_max[211][9] = (mid_1[1703:1696] > mid_0[1695:1688]) ? 1 : 0;
assign detect_max[211][10] = (mid_1[1703:1696] > mid_0[1703:1696]) ? 1 : 0;
assign detect_max[211][11] = (mid_1[1703:1696] > mid_0[1711:1704]) ? 1 : 0;
assign detect_max[211][12] = (mid_1[1703:1696] > mid_1[1695:1688]) ? 1 : 0;
assign detect_max[211][13] = (mid_1[1703:1696] > mid_1[1711:1704]) ? 1 : 0;
assign detect_max[211][14] = (mid_1[1703:1696] > mid_2[1695:1688]) ? 1 : 0;
assign detect_max[211][15] = (mid_1[1703:1696] > mid_2[1703:1696]) ? 1 : 0;
assign detect_max[211][16] = (mid_1[1703:1696] > mid_2[1711:1704]) ? 1 : 0;
assign detect_max[211][17] = (mid_1[1703:1696] > btm_0[1695:1688]) ? 1 : 0;
assign detect_max[211][18] = (mid_1[1703:1696] > btm_0[1703:1696]) ? 1 : 0;
assign detect_max[211][19] = (mid_1[1703:1696] > btm_0[1711:1704]) ? 1 : 0;
assign detect_max[211][20] = (mid_1[1703:1696] > btm_1[1695:1688]) ? 1 : 0;
assign detect_max[211][21] = (mid_1[1703:1696] > btm_1[1703:1696]) ? 1 : 0;
assign detect_max[211][22] = (mid_1[1703:1696] > btm_1[1711:1704]) ? 1 : 0;
assign detect_max[211][23] = (mid_1[1703:1696] > btm_2[1695:1688]) ? 1 : 0;
assign detect_max[211][24] = (mid_1[1703:1696] > btm_2[1703:1696]) ? 1 : 0;
assign detect_max[211][25] = (mid_1[1703:1696] > btm_2[1711:1704]) ? 1 : 0;

assign detect_max[212][0] = (mid_1[1711:1704] > top_0[1703:1696]) ? 1 : 0;
assign detect_max[212][1] = (mid_1[1711:1704] > top_0[1711:1704]) ? 1 : 0;
assign detect_max[212][2] = (mid_1[1711:1704] > top_0[1719:1712]) ? 1 : 0;
assign detect_max[212][3] = (mid_1[1711:1704] > top_1[1703:1696]) ? 1 : 0;
assign detect_max[212][4] = (mid_1[1711:1704] > top_1[1711:1704]) ? 1 : 0;
assign detect_max[212][5] = (mid_1[1711:1704] > top_1[1719:1712]) ? 1 : 0;
assign detect_max[212][6] = (mid_1[1711:1704] > top_2[1703:1696]) ? 1 : 0;
assign detect_max[212][7] = (mid_1[1711:1704] > top_2[1711:1704]) ? 1 : 0;
assign detect_max[212][8] = (mid_1[1711:1704] > top_2[1719:1712]) ? 1 : 0;
assign detect_max[212][9] = (mid_1[1711:1704] > mid_0[1703:1696]) ? 1 : 0;
assign detect_max[212][10] = (mid_1[1711:1704] > mid_0[1711:1704]) ? 1 : 0;
assign detect_max[212][11] = (mid_1[1711:1704] > mid_0[1719:1712]) ? 1 : 0;
assign detect_max[212][12] = (mid_1[1711:1704] > mid_1[1703:1696]) ? 1 : 0;
assign detect_max[212][13] = (mid_1[1711:1704] > mid_1[1719:1712]) ? 1 : 0;
assign detect_max[212][14] = (mid_1[1711:1704] > mid_2[1703:1696]) ? 1 : 0;
assign detect_max[212][15] = (mid_1[1711:1704] > mid_2[1711:1704]) ? 1 : 0;
assign detect_max[212][16] = (mid_1[1711:1704] > mid_2[1719:1712]) ? 1 : 0;
assign detect_max[212][17] = (mid_1[1711:1704] > btm_0[1703:1696]) ? 1 : 0;
assign detect_max[212][18] = (mid_1[1711:1704] > btm_0[1711:1704]) ? 1 : 0;
assign detect_max[212][19] = (mid_1[1711:1704] > btm_0[1719:1712]) ? 1 : 0;
assign detect_max[212][20] = (mid_1[1711:1704] > btm_1[1703:1696]) ? 1 : 0;
assign detect_max[212][21] = (mid_1[1711:1704] > btm_1[1711:1704]) ? 1 : 0;
assign detect_max[212][22] = (mid_1[1711:1704] > btm_1[1719:1712]) ? 1 : 0;
assign detect_max[212][23] = (mid_1[1711:1704] > btm_2[1703:1696]) ? 1 : 0;
assign detect_max[212][24] = (mid_1[1711:1704] > btm_2[1711:1704]) ? 1 : 0;
assign detect_max[212][25] = (mid_1[1711:1704] > btm_2[1719:1712]) ? 1 : 0;

assign detect_max[213][0] = (mid_1[1719:1712] > top_0[1711:1704]) ? 1 : 0;
assign detect_max[213][1] = (mid_1[1719:1712] > top_0[1719:1712]) ? 1 : 0;
assign detect_max[213][2] = (mid_1[1719:1712] > top_0[1727:1720]) ? 1 : 0;
assign detect_max[213][3] = (mid_1[1719:1712] > top_1[1711:1704]) ? 1 : 0;
assign detect_max[213][4] = (mid_1[1719:1712] > top_1[1719:1712]) ? 1 : 0;
assign detect_max[213][5] = (mid_1[1719:1712] > top_1[1727:1720]) ? 1 : 0;
assign detect_max[213][6] = (mid_1[1719:1712] > top_2[1711:1704]) ? 1 : 0;
assign detect_max[213][7] = (mid_1[1719:1712] > top_2[1719:1712]) ? 1 : 0;
assign detect_max[213][8] = (mid_1[1719:1712] > top_2[1727:1720]) ? 1 : 0;
assign detect_max[213][9] = (mid_1[1719:1712] > mid_0[1711:1704]) ? 1 : 0;
assign detect_max[213][10] = (mid_1[1719:1712] > mid_0[1719:1712]) ? 1 : 0;
assign detect_max[213][11] = (mid_1[1719:1712] > mid_0[1727:1720]) ? 1 : 0;
assign detect_max[213][12] = (mid_1[1719:1712] > mid_1[1711:1704]) ? 1 : 0;
assign detect_max[213][13] = (mid_1[1719:1712] > mid_1[1727:1720]) ? 1 : 0;
assign detect_max[213][14] = (mid_1[1719:1712] > mid_2[1711:1704]) ? 1 : 0;
assign detect_max[213][15] = (mid_1[1719:1712] > mid_2[1719:1712]) ? 1 : 0;
assign detect_max[213][16] = (mid_1[1719:1712] > mid_2[1727:1720]) ? 1 : 0;
assign detect_max[213][17] = (mid_1[1719:1712] > btm_0[1711:1704]) ? 1 : 0;
assign detect_max[213][18] = (mid_1[1719:1712] > btm_0[1719:1712]) ? 1 : 0;
assign detect_max[213][19] = (mid_1[1719:1712] > btm_0[1727:1720]) ? 1 : 0;
assign detect_max[213][20] = (mid_1[1719:1712] > btm_1[1711:1704]) ? 1 : 0;
assign detect_max[213][21] = (mid_1[1719:1712] > btm_1[1719:1712]) ? 1 : 0;
assign detect_max[213][22] = (mid_1[1719:1712] > btm_1[1727:1720]) ? 1 : 0;
assign detect_max[213][23] = (mid_1[1719:1712] > btm_2[1711:1704]) ? 1 : 0;
assign detect_max[213][24] = (mid_1[1719:1712] > btm_2[1719:1712]) ? 1 : 0;
assign detect_max[213][25] = (mid_1[1719:1712] > btm_2[1727:1720]) ? 1 : 0;

assign detect_max[214][0] = (mid_1[1727:1720] > top_0[1719:1712]) ? 1 : 0;
assign detect_max[214][1] = (mid_1[1727:1720] > top_0[1727:1720]) ? 1 : 0;
assign detect_max[214][2] = (mid_1[1727:1720] > top_0[1735:1728]) ? 1 : 0;
assign detect_max[214][3] = (mid_1[1727:1720] > top_1[1719:1712]) ? 1 : 0;
assign detect_max[214][4] = (mid_1[1727:1720] > top_1[1727:1720]) ? 1 : 0;
assign detect_max[214][5] = (mid_1[1727:1720] > top_1[1735:1728]) ? 1 : 0;
assign detect_max[214][6] = (mid_1[1727:1720] > top_2[1719:1712]) ? 1 : 0;
assign detect_max[214][7] = (mid_1[1727:1720] > top_2[1727:1720]) ? 1 : 0;
assign detect_max[214][8] = (mid_1[1727:1720] > top_2[1735:1728]) ? 1 : 0;
assign detect_max[214][9] = (mid_1[1727:1720] > mid_0[1719:1712]) ? 1 : 0;
assign detect_max[214][10] = (mid_1[1727:1720] > mid_0[1727:1720]) ? 1 : 0;
assign detect_max[214][11] = (mid_1[1727:1720] > mid_0[1735:1728]) ? 1 : 0;
assign detect_max[214][12] = (mid_1[1727:1720] > mid_1[1719:1712]) ? 1 : 0;
assign detect_max[214][13] = (mid_1[1727:1720] > mid_1[1735:1728]) ? 1 : 0;
assign detect_max[214][14] = (mid_1[1727:1720] > mid_2[1719:1712]) ? 1 : 0;
assign detect_max[214][15] = (mid_1[1727:1720] > mid_2[1727:1720]) ? 1 : 0;
assign detect_max[214][16] = (mid_1[1727:1720] > mid_2[1735:1728]) ? 1 : 0;
assign detect_max[214][17] = (mid_1[1727:1720] > btm_0[1719:1712]) ? 1 : 0;
assign detect_max[214][18] = (mid_1[1727:1720] > btm_0[1727:1720]) ? 1 : 0;
assign detect_max[214][19] = (mid_1[1727:1720] > btm_0[1735:1728]) ? 1 : 0;
assign detect_max[214][20] = (mid_1[1727:1720] > btm_1[1719:1712]) ? 1 : 0;
assign detect_max[214][21] = (mid_1[1727:1720] > btm_1[1727:1720]) ? 1 : 0;
assign detect_max[214][22] = (mid_1[1727:1720] > btm_1[1735:1728]) ? 1 : 0;
assign detect_max[214][23] = (mid_1[1727:1720] > btm_2[1719:1712]) ? 1 : 0;
assign detect_max[214][24] = (mid_1[1727:1720] > btm_2[1727:1720]) ? 1 : 0;
assign detect_max[214][25] = (mid_1[1727:1720] > btm_2[1735:1728]) ? 1 : 0;

assign detect_max[215][0] = (mid_1[1735:1728] > top_0[1727:1720]) ? 1 : 0;
assign detect_max[215][1] = (mid_1[1735:1728] > top_0[1735:1728]) ? 1 : 0;
assign detect_max[215][2] = (mid_1[1735:1728] > top_0[1743:1736]) ? 1 : 0;
assign detect_max[215][3] = (mid_1[1735:1728] > top_1[1727:1720]) ? 1 : 0;
assign detect_max[215][4] = (mid_1[1735:1728] > top_1[1735:1728]) ? 1 : 0;
assign detect_max[215][5] = (mid_1[1735:1728] > top_1[1743:1736]) ? 1 : 0;
assign detect_max[215][6] = (mid_1[1735:1728] > top_2[1727:1720]) ? 1 : 0;
assign detect_max[215][7] = (mid_1[1735:1728] > top_2[1735:1728]) ? 1 : 0;
assign detect_max[215][8] = (mid_1[1735:1728] > top_2[1743:1736]) ? 1 : 0;
assign detect_max[215][9] = (mid_1[1735:1728] > mid_0[1727:1720]) ? 1 : 0;
assign detect_max[215][10] = (mid_1[1735:1728] > mid_0[1735:1728]) ? 1 : 0;
assign detect_max[215][11] = (mid_1[1735:1728] > mid_0[1743:1736]) ? 1 : 0;
assign detect_max[215][12] = (mid_1[1735:1728] > mid_1[1727:1720]) ? 1 : 0;
assign detect_max[215][13] = (mid_1[1735:1728] > mid_1[1743:1736]) ? 1 : 0;
assign detect_max[215][14] = (mid_1[1735:1728] > mid_2[1727:1720]) ? 1 : 0;
assign detect_max[215][15] = (mid_1[1735:1728] > mid_2[1735:1728]) ? 1 : 0;
assign detect_max[215][16] = (mid_1[1735:1728] > mid_2[1743:1736]) ? 1 : 0;
assign detect_max[215][17] = (mid_1[1735:1728] > btm_0[1727:1720]) ? 1 : 0;
assign detect_max[215][18] = (mid_1[1735:1728] > btm_0[1735:1728]) ? 1 : 0;
assign detect_max[215][19] = (mid_1[1735:1728] > btm_0[1743:1736]) ? 1 : 0;
assign detect_max[215][20] = (mid_1[1735:1728] > btm_1[1727:1720]) ? 1 : 0;
assign detect_max[215][21] = (mid_1[1735:1728] > btm_1[1735:1728]) ? 1 : 0;
assign detect_max[215][22] = (mid_1[1735:1728] > btm_1[1743:1736]) ? 1 : 0;
assign detect_max[215][23] = (mid_1[1735:1728] > btm_2[1727:1720]) ? 1 : 0;
assign detect_max[215][24] = (mid_1[1735:1728] > btm_2[1735:1728]) ? 1 : 0;
assign detect_max[215][25] = (mid_1[1735:1728] > btm_2[1743:1736]) ? 1 : 0;

assign detect_max[216][0] = (mid_1[1743:1736] > top_0[1735:1728]) ? 1 : 0;
assign detect_max[216][1] = (mid_1[1743:1736] > top_0[1743:1736]) ? 1 : 0;
assign detect_max[216][2] = (mid_1[1743:1736] > top_0[1751:1744]) ? 1 : 0;
assign detect_max[216][3] = (mid_1[1743:1736] > top_1[1735:1728]) ? 1 : 0;
assign detect_max[216][4] = (mid_1[1743:1736] > top_1[1743:1736]) ? 1 : 0;
assign detect_max[216][5] = (mid_1[1743:1736] > top_1[1751:1744]) ? 1 : 0;
assign detect_max[216][6] = (mid_1[1743:1736] > top_2[1735:1728]) ? 1 : 0;
assign detect_max[216][7] = (mid_1[1743:1736] > top_2[1743:1736]) ? 1 : 0;
assign detect_max[216][8] = (mid_1[1743:1736] > top_2[1751:1744]) ? 1 : 0;
assign detect_max[216][9] = (mid_1[1743:1736] > mid_0[1735:1728]) ? 1 : 0;
assign detect_max[216][10] = (mid_1[1743:1736] > mid_0[1743:1736]) ? 1 : 0;
assign detect_max[216][11] = (mid_1[1743:1736] > mid_0[1751:1744]) ? 1 : 0;
assign detect_max[216][12] = (mid_1[1743:1736] > mid_1[1735:1728]) ? 1 : 0;
assign detect_max[216][13] = (mid_1[1743:1736] > mid_1[1751:1744]) ? 1 : 0;
assign detect_max[216][14] = (mid_1[1743:1736] > mid_2[1735:1728]) ? 1 : 0;
assign detect_max[216][15] = (mid_1[1743:1736] > mid_2[1743:1736]) ? 1 : 0;
assign detect_max[216][16] = (mid_1[1743:1736] > mid_2[1751:1744]) ? 1 : 0;
assign detect_max[216][17] = (mid_1[1743:1736] > btm_0[1735:1728]) ? 1 : 0;
assign detect_max[216][18] = (mid_1[1743:1736] > btm_0[1743:1736]) ? 1 : 0;
assign detect_max[216][19] = (mid_1[1743:1736] > btm_0[1751:1744]) ? 1 : 0;
assign detect_max[216][20] = (mid_1[1743:1736] > btm_1[1735:1728]) ? 1 : 0;
assign detect_max[216][21] = (mid_1[1743:1736] > btm_1[1743:1736]) ? 1 : 0;
assign detect_max[216][22] = (mid_1[1743:1736] > btm_1[1751:1744]) ? 1 : 0;
assign detect_max[216][23] = (mid_1[1743:1736] > btm_2[1735:1728]) ? 1 : 0;
assign detect_max[216][24] = (mid_1[1743:1736] > btm_2[1743:1736]) ? 1 : 0;
assign detect_max[216][25] = (mid_1[1743:1736] > btm_2[1751:1744]) ? 1 : 0;

assign detect_max[217][0] = (mid_1[1751:1744] > top_0[1743:1736]) ? 1 : 0;
assign detect_max[217][1] = (mid_1[1751:1744] > top_0[1751:1744]) ? 1 : 0;
assign detect_max[217][2] = (mid_1[1751:1744] > top_0[1759:1752]) ? 1 : 0;
assign detect_max[217][3] = (mid_1[1751:1744] > top_1[1743:1736]) ? 1 : 0;
assign detect_max[217][4] = (mid_1[1751:1744] > top_1[1751:1744]) ? 1 : 0;
assign detect_max[217][5] = (mid_1[1751:1744] > top_1[1759:1752]) ? 1 : 0;
assign detect_max[217][6] = (mid_1[1751:1744] > top_2[1743:1736]) ? 1 : 0;
assign detect_max[217][7] = (mid_1[1751:1744] > top_2[1751:1744]) ? 1 : 0;
assign detect_max[217][8] = (mid_1[1751:1744] > top_2[1759:1752]) ? 1 : 0;
assign detect_max[217][9] = (mid_1[1751:1744] > mid_0[1743:1736]) ? 1 : 0;
assign detect_max[217][10] = (mid_1[1751:1744] > mid_0[1751:1744]) ? 1 : 0;
assign detect_max[217][11] = (mid_1[1751:1744] > mid_0[1759:1752]) ? 1 : 0;
assign detect_max[217][12] = (mid_1[1751:1744] > mid_1[1743:1736]) ? 1 : 0;
assign detect_max[217][13] = (mid_1[1751:1744] > mid_1[1759:1752]) ? 1 : 0;
assign detect_max[217][14] = (mid_1[1751:1744] > mid_2[1743:1736]) ? 1 : 0;
assign detect_max[217][15] = (mid_1[1751:1744] > mid_2[1751:1744]) ? 1 : 0;
assign detect_max[217][16] = (mid_1[1751:1744] > mid_2[1759:1752]) ? 1 : 0;
assign detect_max[217][17] = (mid_1[1751:1744] > btm_0[1743:1736]) ? 1 : 0;
assign detect_max[217][18] = (mid_1[1751:1744] > btm_0[1751:1744]) ? 1 : 0;
assign detect_max[217][19] = (mid_1[1751:1744] > btm_0[1759:1752]) ? 1 : 0;
assign detect_max[217][20] = (mid_1[1751:1744] > btm_1[1743:1736]) ? 1 : 0;
assign detect_max[217][21] = (mid_1[1751:1744] > btm_1[1751:1744]) ? 1 : 0;
assign detect_max[217][22] = (mid_1[1751:1744] > btm_1[1759:1752]) ? 1 : 0;
assign detect_max[217][23] = (mid_1[1751:1744] > btm_2[1743:1736]) ? 1 : 0;
assign detect_max[217][24] = (mid_1[1751:1744] > btm_2[1751:1744]) ? 1 : 0;
assign detect_max[217][25] = (mid_1[1751:1744] > btm_2[1759:1752]) ? 1 : 0;

assign detect_max[218][0] = (mid_1[1759:1752] > top_0[1751:1744]) ? 1 : 0;
assign detect_max[218][1] = (mid_1[1759:1752] > top_0[1759:1752]) ? 1 : 0;
assign detect_max[218][2] = (mid_1[1759:1752] > top_0[1767:1760]) ? 1 : 0;
assign detect_max[218][3] = (mid_1[1759:1752] > top_1[1751:1744]) ? 1 : 0;
assign detect_max[218][4] = (mid_1[1759:1752] > top_1[1759:1752]) ? 1 : 0;
assign detect_max[218][5] = (mid_1[1759:1752] > top_1[1767:1760]) ? 1 : 0;
assign detect_max[218][6] = (mid_1[1759:1752] > top_2[1751:1744]) ? 1 : 0;
assign detect_max[218][7] = (mid_1[1759:1752] > top_2[1759:1752]) ? 1 : 0;
assign detect_max[218][8] = (mid_1[1759:1752] > top_2[1767:1760]) ? 1 : 0;
assign detect_max[218][9] = (mid_1[1759:1752] > mid_0[1751:1744]) ? 1 : 0;
assign detect_max[218][10] = (mid_1[1759:1752] > mid_0[1759:1752]) ? 1 : 0;
assign detect_max[218][11] = (mid_1[1759:1752] > mid_0[1767:1760]) ? 1 : 0;
assign detect_max[218][12] = (mid_1[1759:1752] > mid_1[1751:1744]) ? 1 : 0;
assign detect_max[218][13] = (mid_1[1759:1752] > mid_1[1767:1760]) ? 1 : 0;
assign detect_max[218][14] = (mid_1[1759:1752] > mid_2[1751:1744]) ? 1 : 0;
assign detect_max[218][15] = (mid_1[1759:1752] > mid_2[1759:1752]) ? 1 : 0;
assign detect_max[218][16] = (mid_1[1759:1752] > mid_2[1767:1760]) ? 1 : 0;
assign detect_max[218][17] = (mid_1[1759:1752] > btm_0[1751:1744]) ? 1 : 0;
assign detect_max[218][18] = (mid_1[1759:1752] > btm_0[1759:1752]) ? 1 : 0;
assign detect_max[218][19] = (mid_1[1759:1752] > btm_0[1767:1760]) ? 1 : 0;
assign detect_max[218][20] = (mid_1[1759:1752] > btm_1[1751:1744]) ? 1 : 0;
assign detect_max[218][21] = (mid_1[1759:1752] > btm_1[1759:1752]) ? 1 : 0;
assign detect_max[218][22] = (mid_1[1759:1752] > btm_1[1767:1760]) ? 1 : 0;
assign detect_max[218][23] = (mid_1[1759:1752] > btm_2[1751:1744]) ? 1 : 0;
assign detect_max[218][24] = (mid_1[1759:1752] > btm_2[1759:1752]) ? 1 : 0;
assign detect_max[218][25] = (mid_1[1759:1752] > btm_2[1767:1760]) ? 1 : 0;

assign detect_max[219][0] = (mid_1[1767:1760] > top_0[1759:1752]) ? 1 : 0;
assign detect_max[219][1] = (mid_1[1767:1760] > top_0[1767:1760]) ? 1 : 0;
assign detect_max[219][2] = (mid_1[1767:1760] > top_0[1775:1768]) ? 1 : 0;
assign detect_max[219][3] = (mid_1[1767:1760] > top_1[1759:1752]) ? 1 : 0;
assign detect_max[219][4] = (mid_1[1767:1760] > top_1[1767:1760]) ? 1 : 0;
assign detect_max[219][5] = (mid_1[1767:1760] > top_1[1775:1768]) ? 1 : 0;
assign detect_max[219][6] = (mid_1[1767:1760] > top_2[1759:1752]) ? 1 : 0;
assign detect_max[219][7] = (mid_1[1767:1760] > top_2[1767:1760]) ? 1 : 0;
assign detect_max[219][8] = (mid_1[1767:1760] > top_2[1775:1768]) ? 1 : 0;
assign detect_max[219][9] = (mid_1[1767:1760] > mid_0[1759:1752]) ? 1 : 0;
assign detect_max[219][10] = (mid_1[1767:1760] > mid_0[1767:1760]) ? 1 : 0;
assign detect_max[219][11] = (mid_1[1767:1760] > mid_0[1775:1768]) ? 1 : 0;
assign detect_max[219][12] = (mid_1[1767:1760] > mid_1[1759:1752]) ? 1 : 0;
assign detect_max[219][13] = (mid_1[1767:1760] > mid_1[1775:1768]) ? 1 : 0;
assign detect_max[219][14] = (mid_1[1767:1760] > mid_2[1759:1752]) ? 1 : 0;
assign detect_max[219][15] = (mid_1[1767:1760] > mid_2[1767:1760]) ? 1 : 0;
assign detect_max[219][16] = (mid_1[1767:1760] > mid_2[1775:1768]) ? 1 : 0;
assign detect_max[219][17] = (mid_1[1767:1760] > btm_0[1759:1752]) ? 1 : 0;
assign detect_max[219][18] = (mid_1[1767:1760] > btm_0[1767:1760]) ? 1 : 0;
assign detect_max[219][19] = (mid_1[1767:1760] > btm_0[1775:1768]) ? 1 : 0;
assign detect_max[219][20] = (mid_1[1767:1760] > btm_1[1759:1752]) ? 1 : 0;
assign detect_max[219][21] = (mid_1[1767:1760] > btm_1[1767:1760]) ? 1 : 0;
assign detect_max[219][22] = (mid_1[1767:1760] > btm_1[1775:1768]) ? 1 : 0;
assign detect_max[219][23] = (mid_1[1767:1760] > btm_2[1759:1752]) ? 1 : 0;
assign detect_max[219][24] = (mid_1[1767:1760] > btm_2[1767:1760]) ? 1 : 0;
assign detect_max[219][25] = (mid_1[1767:1760] > btm_2[1775:1768]) ? 1 : 0;

assign detect_max[220][0] = (mid_1[1775:1768] > top_0[1767:1760]) ? 1 : 0;
assign detect_max[220][1] = (mid_1[1775:1768] > top_0[1775:1768]) ? 1 : 0;
assign detect_max[220][2] = (mid_1[1775:1768] > top_0[1783:1776]) ? 1 : 0;
assign detect_max[220][3] = (mid_1[1775:1768] > top_1[1767:1760]) ? 1 : 0;
assign detect_max[220][4] = (mid_1[1775:1768] > top_1[1775:1768]) ? 1 : 0;
assign detect_max[220][5] = (mid_1[1775:1768] > top_1[1783:1776]) ? 1 : 0;
assign detect_max[220][6] = (mid_1[1775:1768] > top_2[1767:1760]) ? 1 : 0;
assign detect_max[220][7] = (mid_1[1775:1768] > top_2[1775:1768]) ? 1 : 0;
assign detect_max[220][8] = (mid_1[1775:1768] > top_2[1783:1776]) ? 1 : 0;
assign detect_max[220][9] = (mid_1[1775:1768] > mid_0[1767:1760]) ? 1 : 0;
assign detect_max[220][10] = (mid_1[1775:1768] > mid_0[1775:1768]) ? 1 : 0;
assign detect_max[220][11] = (mid_1[1775:1768] > mid_0[1783:1776]) ? 1 : 0;
assign detect_max[220][12] = (mid_1[1775:1768] > mid_1[1767:1760]) ? 1 : 0;
assign detect_max[220][13] = (mid_1[1775:1768] > mid_1[1783:1776]) ? 1 : 0;
assign detect_max[220][14] = (mid_1[1775:1768] > mid_2[1767:1760]) ? 1 : 0;
assign detect_max[220][15] = (mid_1[1775:1768] > mid_2[1775:1768]) ? 1 : 0;
assign detect_max[220][16] = (mid_1[1775:1768] > mid_2[1783:1776]) ? 1 : 0;
assign detect_max[220][17] = (mid_1[1775:1768] > btm_0[1767:1760]) ? 1 : 0;
assign detect_max[220][18] = (mid_1[1775:1768] > btm_0[1775:1768]) ? 1 : 0;
assign detect_max[220][19] = (mid_1[1775:1768] > btm_0[1783:1776]) ? 1 : 0;
assign detect_max[220][20] = (mid_1[1775:1768] > btm_1[1767:1760]) ? 1 : 0;
assign detect_max[220][21] = (mid_1[1775:1768] > btm_1[1775:1768]) ? 1 : 0;
assign detect_max[220][22] = (mid_1[1775:1768] > btm_1[1783:1776]) ? 1 : 0;
assign detect_max[220][23] = (mid_1[1775:1768] > btm_2[1767:1760]) ? 1 : 0;
assign detect_max[220][24] = (mid_1[1775:1768] > btm_2[1775:1768]) ? 1 : 0;
assign detect_max[220][25] = (mid_1[1775:1768] > btm_2[1783:1776]) ? 1 : 0;

assign detect_max[221][0] = (mid_1[1783:1776] > top_0[1775:1768]) ? 1 : 0;
assign detect_max[221][1] = (mid_1[1783:1776] > top_0[1783:1776]) ? 1 : 0;
assign detect_max[221][2] = (mid_1[1783:1776] > top_0[1791:1784]) ? 1 : 0;
assign detect_max[221][3] = (mid_1[1783:1776] > top_1[1775:1768]) ? 1 : 0;
assign detect_max[221][4] = (mid_1[1783:1776] > top_1[1783:1776]) ? 1 : 0;
assign detect_max[221][5] = (mid_1[1783:1776] > top_1[1791:1784]) ? 1 : 0;
assign detect_max[221][6] = (mid_1[1783:1776] > top_2[1775:1768]) ? 1 : 0;
assign detect_max[221][7] = (mid_1[1783:1776] > top_2[1783:1776]) ? 1 : 0;
assign detect_max[221][8] = (mid_1[1783:1776] > top_2[1791:1784]) ? 1 : 0;
assign detect_max[221][9] = (mid_1[1783:1776] > mid_0[1775:1768]) ? 1 : 0;
assign detect_max[221][10] = (mid_1[1783:1776] > mid_0[1783:1776]) ? 1 : 0;
assign detect_max[221][11] = (mid_1[1783:1776] > mid_0[1791:1784]) ? 1 : 0;
assign detect_max[221][12] = (mid_1[1783:1776] > mid_1[1775:1768]) ? 1 : 0;
assign detect_max[221][13] = (mid_1[1783:1776] > mid_1[1791:1784]) ? 1 : 0;
assign detect_max[221][14] = (mid_1[1783:1776] > mid_2[1775:1768]) ? 1 : 0;
assign detect_max[221][15] = (mid_1[1783:1776] > mid_2[1783:1776]) ? 1 : 0;
assign detect_max[221][16] = (mid_1[1783:1776] > mid_2[1791:1784]) ? 1 : 0;
assign detect_max[221][17] = (mid_1[1783:1776] > btm_0[1775:1768]) ? 1 : 0;
assign detect_max[221][18] = (mid_1[1783:1776] > btm_0[1783:1776]) ? 1 : 0;
assign detect_max[221][19] = (mid_1[1783:1776] > btm_0[1791:1784]) ? 1 : 0;
assign detect_max[221][20] = (mid_1[1783:1776] > btm_1[1775:1768]) ? 1 : 0;
assign detect_max[221][21] = (mid_1[1783:1776] > btm_1[1783:1776]) ? 1 : 0;
assign detect_max[221][22] = (mid_1[1783:1776] > btm_1[1791:1784]) ? 1 : 0;
assign detect_max[221][23] = (mid_1[1783:1776] > btm_2[1775:1768]) ? 1 : 0;
assign detect_max[221][24] = (mid_1[1783:1776] > btm_2[1783:1776]) ? 1 : 0;
assign detect_max[221][25] = (mid_1[1783:1776] > btm_2[1791:1784]) ? 1 : 0;

assign detect_max[222][0] = (mid_1[1791:1784] > top_0[1783:1776]) ? 1 : 0;
assign detect_max[222][1] = (mid_1[1791:1784] > top_0[1791:1784]) ? 1 : 0;
assign detect_max[222][2] = (mid_1[1791:1784] > top_0[1799:1792]) ? 1 : 0;
assign detect_max[222][3] = (mid_1[1791:1784] > top_1[1783:1776]) ? 1 : 0;
assign detect_max[222][4] = (mid_1[1791:1784] > top_1[1791:1784]) ? 1 : 0;
assign detect_max[222][5] = (mid_1[1791:1784] > top_1[1799:1792]) ? 1 : 0;
assign detect_max[222][6] = (mid_1[1791:1784] > top_2[1783:1776]) ? 1 : 0;
assign detect_max[222][7] = (mid_1[1791:1784] > top_2[1791:1784]) ? 1 : 0;
assign detect_max[222][8] = (mid_1[1791:1784] > top_2[1799:1792]) ? 1 : 0;
assign detect_max[222][9] = (mid_1[1791:1784] > mid_0[1783:1776]) ? 1 : 0;
assign detect_max[222][10] = (mid_1[1791:1784] > mid_0[1791:1784]) ? 1 : 0;
assign detect_max[222][11] = (mid_1[1791:1784] > mid_0[1799:1792]) ? 1 : 0;
assign detect_max[222][12] = (mid_1[1791:1784] > mid_1[1783:1776]) ? 1 : 0;
assign detect_max[222][13] = (mid_1[1791:1784] > mid_1[1799:1792]) ? 1 : 0;
assign detect_max[222][14] = (mid_1[1791:1784] > mid_2[1783:1776]) ? 1 : 0;
assign detect_max[222][15] = (mid_1[1791:1784] > mid_2[1791:1784]) ? 1 : 0;
assign detect_max[222][16] = (mid_1[1791:1784] > mid_2[1799:1792]) ? 1 : 0;
assign detect_max[222][17] = (mid_1[1791:1784] > btm_0[1783:1776]) ? 1 : 0;
assign detect_max[222][18] = (mid_1[1791:1784] > btm_0[1791:1784]) ? 1 : 0;
assign detect_max[222][19] = (mid_1[1791:1784] > btm_0[1799:1792]) ? 1 : 0;
assign detect_max[222][20] = (mid_1[1791:1784] > btm_1[1783:1776]) ? 1 : 0;
assign detect_max[222][21] = (mid_1[1791:1784] > btm_1[1791:1784]) ? 1 : 0;
assign detect_max[222][22] = (mid_1[1791:1784] > btm_1[1799:1792]) ? 1 : 0;
assign detect_max[222][23] = (mid_1[1791:1784] > btm_2[1783:1776]) ? 1 : 0;
assign detect_max[222][24] = (mid_1[1791:1784] > btm_2[1791:1784]) ? 1 : 0;
assign detect_max[222][25] = (mid_1[1791:1784] > btm_2[1799:1792]) ? 1 : 0;

assign detect_max[223][0] = (mid_1[1799:1792] > top_0[1791:1784]) ? 1 : 0;
assign detect_max[223][1] = (mid_1[1799:1792] > top_0[1799:1792]) ? 1 : 0;
assign detect_max[223][2] = (mid_1[1799:1792] > top_0[1807:1800]) ? 1 : 0;
assign detect_max[223][3] = (mid_1[1799:1792] > top_1[1791:1784]) ? 1 : 0;
assign detect_max[223][4] = (mid_1[1799:1792] > top_1[1799:1792]) ? 1 : 0;
assign detect_max[223][5] = (mid_1[1799:1792] > top_1[1807:1800]) ? 1 : 0;
assign detect_max[223][6] = (mid_1[1799:1792] > top_2[1791:1784]) ? 1 : 0;
assign detect_max[223][7] = (mid_1[1799:1792] > top_2[1799:1792]) ? 1 : 0;
assign detect_max[223][8] = (mid_1[1799:1792] > top_2[1807:1800]) ? 1 : 0;
assign detect_max[223][9] = (mid_1[1799:1792] > mid_0[1791:1784]) ? 1 : 0;
assign detect_max[223][10] = (mid_1[1799:1792] > mid_0[1799:1792]) ? 1 : 0;
assign detect_max[223][11] = (mid_1[1799:1792] > mid_0[1807:1800]) ? 1 : 0;
assign detect_max[223][12] = (mid_1[1799:1792] > mid_1[1791:1784]) ? 1 : 0;
assign detect_max[223][13] = (mid_1[1799:1792] > mid_1[1807:1800]) ? 1 : 0;
assign detect_max[223][14] = (mid_1[1799:1792] > mid_2[1791:1784]) ? 1 : 0;
assign detect_max[223][15] = (mid_1[1799:1792] > mid_2[1799:1792]) ? 1 : 0;
assign detect_max[223][16] = (mid_1[1799:1792] > mid_2[1807:1800]) ? 1 : 0;
assign detect_max[223][17] = (mid_1[1799:1792] > btm_0[1791:1784]) ? 1 : 0;
assign detect_max[223][18] = (mid_1[1799:1792] > btm_0[1799:1792]) ? 1 : 0;
assign detect_max[223][19] = (mid_1[1799:1792] > btm_0[1807:1800]) ? 1 : 0;
assign detect_max[223][20] = (mid_1[1799:1792] > btm_1[1791:1784]) ? 1 : 0;
assign detect_max[223][21] = (mid_1[1799:1792] > btm_1[1799:1792]) ? 1 : 0;
assign detect_max[223][22] = (mid_1[1799:1792] > btm_1[1807:1800]) ? 1 : 0;
assign detect_max[223][23] = (mid_1[1799:1792] > btm_2[1791:1784]) ? 1 : 0;
assign detect_max[223][24] = (mid_1[1799:1792] > btm_2[1799:1792]) ? 1 : 0;
assign detect_max[223][25] = (mid_1[1799:1792] > btm_2[1807:1800]) ? 1 : 0;

assign detect_max[224][0] = (mid_1[1807:1800] > top_0[1799:1792]) ? 1 : 0;
assign detect_max[224][1] = (mid_1[1807:1800] > top_0[1807:1800]) ? 1 : 0;
assign detect_max[224][2] = (mid_1[1807:1800] > top_0[1815:1808]) ? 1 : 0;
assign detect_max[224][3] = (mid_1[1807:1800] > top_1[1799:1792]) ? 1 : 0;
assign detect_max[224][4] = (mid_1[1807:1800] > top_1[1807:1800]) ? 1 : 0;
assign detect_max[224][5] = (mid_1[1807:1800] > top_1[1815:1808]) ? 1 : 0;
assign detect_max[224][6] = (mid_1[1807:1800] > top_2[1799:1792]) ? 1 : 0;
assign detect_max[224][7] = (mid_1[1807:1800] > top_2[1807:1800]) ? 1 : 0;
assign detect_max[224][8] = (mid_1[1807:1800] > top_2[1815:1808]) ? 1 : 0;
assign detect_max[224][9] = (mid_1[1807:1800] > mid_0[1799:1792]) ? 1 : 0;
assign detect_max[224][10] = (mid_1[1807:1800] > mid_0[1807:1800]) ? 1 : 0;
assign detect_max[224][11] = (mid_1[1807:1800] > mid_0[1815:1808]) ? 1 : 0;
assign detect_max[224][12] = (mid_1[1807:1800] > mid_1[1799:1792]) ? 1 : 0;
assign detect_max[224][13] = (mid_1[1807:1800] > mid_1[1815:1808]) ? 1 : 0;
assign detect_max[224][14] = (mid_1[1807:1800] > mid_2[1799:1792]) ? 1 : 0;
assign detect_max[224][15] = (mid_1[1807:1800] > mid_2[1807:1800]) ? 1 : 0;
assign detect_max[224][16] = (mid_1[1807:1800] > mid_2[1815:1808]) ? 1 : 0;
assign detect_max[224][17] = (mid_1[1807:1800] > btm_0[1799:1792]) ? 1 : 0;
assign detect_max[224][18] = (mid_1[1807:1800] > btm_0[1807:1800]) ? 1 : 0;
assign detect_max[224][19] = (mid_1[1807:1800] > btm_0[1815:1808]) ? 1 : 0;
assign detect_max[224][20] = (mid_1[1807:1800] > btm_1[1799:1792]) ? 1 : 0;
assign detect_max[224][21] = (mid_1[1807:1800] > btm_1[1807:1800]) ? 1 : 0;
assign detect_max[224][22] = (mid_1[1807:1800] > btm_1[1815:1808]) ? 1 : 0;
assign detect_max[224][23] = (mid_1[1807:1800] > btm_2[1799:1792]) ? 1 : 0;
assign detect_max[224][24] = (mid_1[1807:1800] > btm_2[1807:1800]) ? 1 : 0;
assign detect_max[224][25] = (mid_1[1807:1800] > btm_2[1815:1808]) ? 1 : 0;

assign detect_max[225][0] = (mid_1[1815:1808] > top_0[1807:1800]) ? 1 : 0;
assign detect_max[225][1] = (mid_1[1815:1808] > top_0[1815:1808]) ? 1 : 0;
assign detect_max[225][2] = (mid_1[1815:1808] > top_0[1823:1816]) ? 1 : 0;
assign detect_max[225][3] = (mid_1[1815:1808] > top_1[1807:1800]) ? 1 : 0;
assign detect_max[225][4] = (mid_1[1815:1808] > top_1[1815:1808]) ? 1 : 0;
assign detect_max[225][5] = (mid_1[1815:1808] > top_1[1823:1816]) ? 1 : 0;
assign detect_max[225][6] = (mid_1[1815:1808] > top_2[1807:1800]) ? 1 : 0;
assign detect_max[225][7] = (mid_1[1815:1808] > top_2[1815:1808]) ? 1 : 0;
assign detect_max[225][8] = (mid_1[1815:1808] > top_2[1823:1816]) ? 1 : 0;
assign detect_max[225][9] = (mid_1[1815:1808] > mid_0[1807:1800]) ? 1 : 0;
assign detect_max[225][10] = (mid_1[1815:1808] > mid_0[1815:1808]) ? 1 : 0;
assign detect_max[225][11] = (mid_1[1815:1808] > mid_0[1823:1816]) ? 1 : 0;
assign detect_max[225][12] = (mid_1[1815:1808] > mid_1[1807:1800]) ? 1 : 0;
assign detect_max[225][13] = (mid_1[1815:1808] > mid_1[1823:1816]) ? 1 : 0;
assign detect_max[225][14] = (mid_1[1815:1808] > mid_2[1807:1800]) ? 1 : 0;
assign detect_max[225][15] = (mid_1[1815:1808] > mid_2[1815:1808]) ? 1 : 0;
assign detect_max[225][16] = (mid_1[1815:1808] > mid_2[1823:1816]) ? 1 : 0;
assign detect_max[225][17] = (mid_1[1815:1808] > btm_0[1807:1800]) ? 1 : 0;
assign detect_max[225][18] = (mid_1[1815:1808] > btm_0[1815:1808]) ? 1 : 0;
assign detect_max[225][19] = (mid_1[1815:1808] > btm_0[1823:1816]) ? 1 : 0;
assign detect_max[225][20] = (mid_1[1815:1808] > btm_1[1807:1800]) ? 1 : 0;
assign detect_max[225][21] = (mid_1[1815:1808] > btm_1[1815:1808]) ? 1 : 0;
assign detect_max[225][22] = (mid_1[1815:1808] > btm_1[1823:1816]) ? 1 : 0;
assign detect_max[225][23] = (mid_1[1815:1808] > btm_2[1807:1800]) ? 1 : 0;
assign detect_max[225][24] = (mid_1[1815:1808] > btm_2[1815:1808]) ? 1 : 0;
assign detect_max[225][25] = (mid_1[1815:1808] > btm_2[1823:1816]) ? 1 : 0;

assign detect_max[226][0] = (mid_1[1823:1816] > top_0[1815:1808]) ? 1 : 0;
assign detect_max[226][1] = (mid_1[1823:1816] > top_0[1823:1816]) ? 1 : 0;
assign detect_max[226][2] = (mid_1[1823:1816] > top_0[1831:1824]) ? 1 : 0;
assign detect_max[226][3] = (mid_1[1823:1816] > top_1[1815:1808]) ? 1 : 0;
assign detect_max[226][4] = (mid_1[1823:1816] > top_1[1823:1816]) ? 1 : 0;
assign detect_max[226][5] = (mid_1[1823:1816] > top_1[1831:1824]) ? 1 : 0;
assign detect_max[226][6] = (mid_1[1823:1816] > top_2[1815:1808]) ? 1 : 0;
assign detect_max[226][7] = (mid_1[1823:1816] > top_2[1823:1816]) ? 1 : 0;
assign detect_max[226][8] = (mid_1[1823:1816] > top_2[1831:1824]) ? 1 : 0;
assign detect_max[226][9] = (mid_1[1823:1816] > mid_0[1815:1808]) ? 1 : 0;
assign detect_max[226][10] = (mid_1[1823:1816] > mid_0[1823:1816]) ? 1 : 0;
assign detect_max[226][11] = (mid_1[1823:1816] > mid_0[1831:1824]) ? 1 : 0;
assign detect_max[226][12] = (mid_1[1823:1816] > mid_1[1815:1808]) ? 1 : 0;
assign detect_max[226][13] = (mid_1[1823:1816] > mid_1[1831:1824]) ? 1 : 0;
assign detect_max[226][14] = (mid_1[1823:1816] > mid_2[1815:1808]) ? 1 : 0;
assign detect_max[226][15] = (mid_1[1823:1816] > mid_2[1823:1816]) ? 1 : 0;
assign detect_max[226][16] = (mid_1[1823:1816] > mid_2[1831:1824]) ? 1 : 0;
assign detect_max[226][17] = (mid_1[1823:1816] > btm_0[1815:1808]) ? 1 : 0;
assign detect_max[226][18] = (mid_1[1823:1816] > btm_0[1823:1816]) ? 1 : 0;
assign detect_max[226][19] = (mid_1[1823:1816] > btm_0[1831:1824]) ? 1 : 0;
assign detect_max[226][20] = (mid_1[1823:1816] > btm_1[1815:1808]) ? 1 : 0;
assign detect_max[226][21] = (mid_1[1823:1816] > btm_1[1823:1816]) ? 1 : 0;
assign detect_max[226][22] = (mid_1[1823:1816] > btm_1[1831:1824]) ? 1 : 0;
assign detect_max[226][23] = (mid_1[1823:1816] > btm_2[1815:1808]) ? 1 : 0;
assign detect_max[226][24] = (mid_1[1823:1816] > btm_2[1823:1816]) ? 1 : 0;
assign detect_max[226][25] = (mid_1[1823:1816] > btm_2[1831:1824]) ? 1 : 0;

assign detect_max[227][0] = (mid_1[1831:1824] > top_0[1823:1816]) ? 1 : 0;
assign detect_max[227][1] = (mid_1[1831:1824] > top_0[1831:1824]) ? 1 : 0;
assign detect_max[227][2] = (mid_1[1831:1824] > top_0[1839:1832]) ? 1 : 0;
assign detect_max[227][3] = (mid_1[1831:1824] > top_1[1823:1816]) ? 1 : 0;
assign detect_max[227][4] = (mid_1[1831:1824] > top_1[1831:1824]) ? 1 : 0;
assign detect_max[227][5] = (mid_1[1831:1824] > top_1[1839:1832]) ? 1 : 0;
assign detect_max[227][6] = (mid_1[1831:1824] > top_2[1823:1816]) ? 1 : 0;
assign detect_max[227][7] = (mid_1[1831:1824] > top_2[1831:1824]) ? 1 : 0;
assign detect_max[227][8] = (mid_1[1831:1824] > top_2[1839:1832]) ? 1 : 0;
assign detect_max[227][9] = (mid_1[1831:1824] > mid_0[1823:1816]) ? 1 : 0;
assign detect_max[227][10] = (mid_1[1831:1824] > mid_0[1831:1824]) ? 1 : 0;
assign detect_max[227][11] = (mid_1[1831:1824] > mid_0[1839:1832]) ? 1 : 0;
assign detect_max[227][12] = (mid_1[1831:1824] > mid_1[1823:1816]) ? 1 : 0;
assign detect_max[227][13] = (mid_1[1831:1824] > mid_1[1839:1832]) ? 1 : 0;
assign detect_max[227][14] = (mid_1[1831:1824] > mid_2[1823:1816]) ? 1 : 0;
assign detect_max[227][15] = (mid_1[1831:1824] > mid_2[1831:1824]) ? 1 : 0;
assign detect_max[227][16] = (mid_1[1831:1824] > mid_2[1839:1832]) ? 1 : 0;
assign detect_max[227][17] = (mid_1[1831:1824] > btm_0[1823:1816]) ? 1 : 0;
assign detect_max[227][18] = (mid_1[1831:1824] > btm_0[1831:1824]) ? 1 : 0;
assign detect_max[227][19] = (mid_1[1831:1824] > btm_0[1839:1832]) ? 1 : 0;
assign detect_max[227][20] = (mid_1[1831:1824] > btm_1[1823:1816]) ? 1 : 0;
assign detect_max[227][21] = (mid_1[1831:1824] > btm_1[1831:1824]) ? 1 : 0;
assign detect_max[227][22] = (mid_1[1831:1824] > btm_1[1839:1832]) ? 1 : 0;
assign detect_max[227][23] = (mid_1[1831:1824] > btm_2[1823:1816]) ? 1 : 0;
assign detect_max[227][24] = (mid_1[1831:1824] > btm_2[1831:1824]) ? 1 : 0;
assign detect_max[227][25] = (mid_1[1831:1824] > btm_2[1839:1832]) ? 1 : 0;

assign detect_max[228][0] = (mid_1[1839:1832] > top_0[1831:1824]) ? 1 : 0;
assign detect_max[228][1] = (mid_1[1839:1832] > top_0[1839:1832]) ? 1 : 0;
assign detect_max[228][2] = (mid_1[1839:1832] > top_0[1847:1840]) ? 1 : 0;
assign detect_max[228][3] = (mid_1[1839:1832] > top_1[1831:1824]) ? 1 : 0;
assign detect_max[228][4] = (mid_1[1839:1832] > top_1[1839:1832]) ? 1 : 0;
assign detect_max[228][5] = (mid_1[1839:1832] > top_1[1847:1840]) ? 1 : 0;
assign detect_max[228][6] = (mid_1[1839:1832] > top_2[1831:1824]) ? 1 : 0;
assign detect_max[228][7] = (mid_1[1839:1832] > top_2[1839:1832]) ? 1 : 0;
assign detect_max[228][8] = (mid_1[1839:1832] > top_2[1847:1840]) ? 1 : 0;
assign detect_max[228][9] = (mid_1[1839:1832] > mid_0[1831:1824]) ? 1 : 0;
assign detect_max[228][10] = (mid_1[1839:1832] > mid_0[1839:1832]) ? 1 : 0;
assign detect_max[228][11] = (mid_1[1839:1832] > mid_0[1847:1840]) ? 1 : 0;
assign detect_max[228][12] = (mid_1[1839:1832] > mid_1[1831:1824]) ? 1 : 0;
assign detect_max[228][13] = (mid_1[1839:1832] > mid_1[1847:1840]) ? 1 : 0;
assign detect_max[228][14] = (mid_1[1839:1832] > mid_2[1831:1824]) ? 1 : 0;
assign detect_max[228][15] = (mid_1[1839:1832] > mid_2[1839:1832]) ? 1 : 0;
assign detect_max[228][16] = (mid_1[1839:1832] > mid_2[1847:1840]) ? 1 : 0;
assign detect_max[228][17] = (mid_1[1839:1832] > btm_0[1831:1824]) ? 1 : 0;
assign detect_max[228][18] = (mid_1[1839:1832] > btm_0[1839:1832]) ? 1 : 0;
assign detect_max[228][19] = (mid_1[1839:1832] > btm_0[1847:1840]) ? 1 : 0;
assign detect_max[228][20] = (mid_1[1839:1832] > btm_1[1831:1824]) ? 1 : 0;
assign detect_max[228][21] = (mid_1[1839:1832] > btm_1[1839:1832]) ? 1 : 0;
assign detect_max[228][22] = (mid_1[1839:1832] > btm_1[1847:1840]) ? 1 : 0;
assign detect_max[228][23] = (mid_1[1839:1832] > btm_2[1831:1824]) ? 1 : 0;
assign detect_max[228][24] = (mid_1[1839:1832] > btm_2[1839:1832]) ? 1 : 0;
assign detect_max[228][25] = (mid_1[1839:1832] > btm_2[1847:1840]) ? 1 : 0;

assign detect_max[229][0] = (mid_1[1847:1840] > top_0[1839:1832]) ? 1 : 0;
assign detect_max[229][1] = (mid_1[1847:1840] > top_0[1847:1840]) ? 1 : 0;
assign detect_max[229][2] = (mid_1[1847:1840] > top_0[1855:1848]) ? 1 : 0;
assign detect_max[229][3] = (mid_1[1847:1840] > top_1[1839:1832]) ? 1 : 0;
assign detect_max[229][4] = (mid_1[1847:1840] > top_1[1847:1840]) ? 1 : 0;
assign detect_max[229][5] = (mid_1[1847:1840] > top_1[1855:1848]) ? 1 : 0;
assign detect_max[229][6] = (mid_1[1847:1840] > top_2[1839:1832]) ? 1 : 0;
assign detect_max[229][7] = (mid_1[1847:1840] > top_2[1847:1840]) ? 1 : 0;
assign detect_max[229][8] = (mid_1[1847:1840] > top_2[1855:1848]) ? 1 : 0;
assign detect_max[229][9] = (mid_1[1847:1840] > mid_0[1839:1832]) ? 1 : 0;
assign detect_max[229][10] = (mid_1[1847:1840] > mid_0[1847:1840]) ? 1 : 0;
assign detect_max[229][11] = (mid_1[1847:1840] > mid_0[1855:1848]) ? 1 : 0;
assign detect_max[229][12] = (mid_1[1847:1840] > mid_1[1839:1832]) ? 1 : 0;
assign detect_max[229][13] = (mid_1[1847:1840] > mid_1[1855:1848]) ? 1 : 0;
assign detect_max[229][14] = (mid_1[1847:1840] > mid_2[1839:1832]) ? 1 : 0;
assign detect_max[229][15] = (mid_1[1847:1840] > mid_2[1847:1840]) ? 1 : 0;
assign detect_max[229][16] = (mid_1[1847:1840] > mid_2[1855:1848]) ? 1 : 0;
assign detect_max[229][17] = (mid_1[1847:1840] > btm_0[1839:1832]) ? 1 : 0;
assign detect_max[229][18] = (mid_1[1847:1840] > btm_0[1847:1840]) ? 1 : 0;
assign detect_max[229][19] = (mid_1[1847:1840] > btm_0[1855:1848]) ? 1 : 0;
assign detect_max[229][20] = (mid_1[1847:1840] > btm_1[1839:1832]) ? 1 : 0;
assign detect_max[229][21] = (mid_1[1847:1840] > btm_1[1847:1840]) ? 1 : 0;
assign detect_max[229][22] = (mid_1[1847:1840] > btm_1[1855:1848]) ? 1 : 0;
assign detect_max[229][23] = (mid_1[1847:1840] > btm_2[1839:1832]) ? 1 : 0;
assign detect_max[229][24] = (mid_1[1847:1840] > btm_2[1847:1840]) ? 1 : 0;
assign detect_max[229][25] = (mid_1[1847:1840] > btm_2[1855:1848]) ? 1 : 0;

assign detect_max[230][0] = (mid_1[1855:1848] > top_0[1847:1840]) ? 1 : 0;
assign detect_max[230][1] = (mid_1[1855:1848] > top_0[1855:1848]) ? 1 : 0;
assign detect_max[230][2] = (mid_1[1855:1848] > top_0[1863:1856]) ? 1 : 0;
assign detect_max[230][3] = (mid_1[1855:1848] > top_1[1847:1840]) ? 1 : 0;
assign detect_max[230][4] = (mid_1[1855:1848] > top_1[1855:1848]) ? 1 : 0;
assign detect_max[230][5] = (mid_1[1855:1848] > top_1[1863:1856]) ? 1 : 0;
assign detect_max[230][6] = (mid_1[1855:1848] > top_2[1847:1840]) ? 1 : 0;
assign detect_max[230][7] = (mid_1[1855:1848] > top_2[1855:1848]) ? 1 : 0;
assign detect_max[230][8] = (mid_1[1855:1848] > top_2[1863:1856]) ? 1 : 0;
assign detect_max[230][9] = (mid_1[1855:1848] > mid_0[1847:1840]) ? 1 : 0;
assign detect_max[230][10] = (mid_1[1855:1848] > mid_0[1855:1848]) ? 1 : 0;
assign detect_max[230][11] = (mid_1[1855:1848] > mid_0[1863:1856]) ? 1 : 0;
assign detect_max[230][12] = (mid_1[1855:1848] > mid_1[1847:1840]) ? 1 : 0;
assign detect_max[230][13] = (mid_1[1855:1848] > mid_1[1863:1856]) ? 1 : 0;
assign detect_max[230][14] = (mid_1[1855:1848] > mid_2[1847:1840]) ? 1 : 0;
assign detect_max[230][15] = (mid_1[1855:1848] > mid_2[1855:1848]) ? 1 : 0;
assign detect_max[230][16] = (mid_1[1855:1848] > mid_2[1863:1856]) ? 1 : 0;
assign detect_max[230][17] = (mid_1[1855:1848] > btm_0[1847:1840]) ? 1 : 0;
assign detect_max[230][18] = (mid_1[1855:1848] > btm_0[1855:1848]) ? 1 : 0;
assign detect_max[230][19] = (mid_1[1855:1848] > btm_0[1863:1856]) ? 1 : 0;
assign detect_max[230][20] = (mid_1[1855:1848] > btm_1[1847:1840]) ? 1 : 0;
assign detect_max[230][21] = (mid_1[1855:1848] > btm_1[1855:1848]) ? 1 : 0;
assign detect_max[230][22] = (mid_1[1855:1848] > btm_1[1863:1856]) ? 1 : 0;
assign detect_max[230][23] = (mid_1[1855:1848] > btm_2[1847:1840]) ? 1 : 0;
assign detect_max[230][24] = (mid_1[1855:1848] > btm_2[1855:1848]) ? 1 : 0;
assign detect_max[230][25] = (mid_1[1855:1848] > btm_2[1863:1856]) ? 1 : 0;

assign detect_max[231][0] = (mid_1[1863:1856] > top_0[1855:1848]) ? 1 : 0;
assign detect_max[231][1] = (mid_1[1863:1856] > top_0[1863:1856]) ? 1 : 0;
assign detect_max[231][2] = (mid_1[1863:1856] > top_0[1871:1864]) ? 1 : 0;
assign detect_max[231][3] = (mid_1[1863:1856] > top_1[1855:1848]) ? 1 : 0;
assign detect_max[231][4] = (mid_1[1863:1856] > top_1[1863:1856]) ? 1 : 0;
assign detect_max[231][5] = (mid_1[1863:1856] > top_1[1871:1864]) ? 1 : 0;
assign detect_max[231][6] = (mid_1[1863:1856] > top_2[1855:1848]) ? 1 : 0;
assign detect_max[231][7] = (mid_1[1863:1856] > top_2[1863:1856]) ? 1 : 0;
assign detect_max[231][8] = (mid_1[1863:1856] > top_2[1871:1864]) ? 1 : 0;
assign detect_max[231][9] = (mid_1[1863:1856] > mid_0[1855:1848]) ? 1 : 0;
assign detect_max[231][10] = (mid_1[1863:1856] > mid_0[1863:1856]) ? 1 : 0;
assign detect_max[231][11] = (mid_1[1863:1856] > mid_0[1871:1864]) ? 1 : 0;
assign detect_max[231][12] = (mid_1[1863:1856] > mid_1[1855:1848]) ? 1 : 0;
assign detect_max[231][13] = (mid_1[1863:1856] > mid_1[1871:1864]) ? 1 : 0;
assign detect_max[231][14] = (mid_1[1863:1856] > mid_2[1855:1848]) ? 1 : 0;
assign detect_max[231][15] = (mid_1[1863:1856] > mid_2[1863:1856]) ? 1 : 0;
assign detect_max[231][16] = (mid_1[1863:1856] > mid_2[1871:1864]) ? 1 : 0;
assign detect_max[231][17] = (mid_1[1863:1856] > btm_0[1855:1848]) ? 1 : 0;
assign detect_max[231][18] = (mid_1[1863:1856] > btm_0[1863:1856]) ? 1 : 0;
assign detect_max[231][19] = (mid_1[1863:1856] > btm_0[1871:1864]) ? 1 : 0;
assign detect_max[231][20] = (mid_1[1863:1856] > btm_1[1855:1848]) ? 1 : 0;
assign detect_max[231][21] = (mid_1[1863:1856] > btm_1[1863:1856]) ? 1 : 0;
assign detect_max[231][22] = (mid_1[1863:1856] > btm_1[1871:1864]) ? 1 : 0;
assign detect_max[231][23] = (mid_1[1863:1856] > btm_2[1855:1848]) ? 1 : 0;
assign detect_max[231][24] = (mid_1[1863:1856] > btm_2[1863:1856]) ? 1 : 0;
assign detect_max[231][25] = (mid_1[1863:1856] > btm_2[1871:1864]) ? 1 : 0;

assign detect_max[232][0] = (mid_1[1871:1864] > top_0[1863:1856]) ? 1 : 0;
assign detect_max[232][1] = (mid_1[1871:1864] > top_0[1871:1864]) ? 1 : 0;
assign detect_max[232][2] = (mid_1[1871:1864] > top_0[1879:1872]) ? 1 : 0;
assign detect_max[232][3] = (mid_1[1871:1864] > top_1[1863:1856]) ? 1 : 0;
assign detect_max[232][4] = (mid_1[1871:1864] > top_1[1871:1864]) ? 1 : 0;
assign detect_max[232][5] = (mid_1[1871:1864] > top_1[1879:1872]) ? 1 : 0;
assign detect_max[232][6] = (mid_1[1871:1864] > top_2[1863:1856]) ? 1 : 0;
assign detect_max[232][7] = (mid_1[1871:1864] > top_2[1871:1864]) ? 1 : 0;
assign detect_max[232][8] = (mid_1[1871:1864] > top_2[1879:1872]) ? 1 : 0;
assign detect_max[232][9] = (mid_1[1871:1864] > mid_0[1863:1856]) ? 1 : 0;
assign detect_max[232][10] = (mid_1[1871:1864] > mid_0[1871:1864]) ? 1 : 0;
assign detect_max[232][11] = (mid_1[1871:1864] > mid_0[1879:1872]) ? 1 : 0;
assign detect_max[232][12] = (mid_1[1871:1864] > mid_1[1863:1856]) ? 1 : 0;
assign detect_max[232][13] = (mid_1[1871:1864] > mid_1[1879:1872]) ? 1 : 0;
assign detect_max[232][14] = (mid_1[1871:1864] > mid_2[1863:1856]) ? 1 : 0;
assign detect_max[232][15] = (mid_1[1871:1864] > mid_2[1871:1864]) ? 1 : 0;
assign detect_max[232][16] = (mid_1[1871:1864] > mid_2[1879:1872]) ? 1 : 0;
assign detect_max[232][17] = (mid_1[1871:1864] > btm_0[1863:1856]) ? 1 : 0;
assign detect_max[232][18] = (mid_1[1871:1864] > btm_0[1871:1864]) ? 1 : 0;
assign detect_max[232][19] = (mid_1[1871:1864] > btm_0[1879:1872]) ? 1 : 0;
assign detect_max[232][20] = (mid_1[1871:1864] > btm_1[1863:1856]) ? 1 : 0;
assign detect_max[232][21] = (mid_1[1871:1864] > btm_1[1871:1864]) ? 1 : 0;
assign detect_max[232][22] = (mid_1[1871:1864] > btm_1[1879:1872]) ? 1 : 0;
assign detect_max[232][23] = (mid_1[1871:1864] > btm_2[1863:1856]) ? 1 : 0;
assign detect_max[232][24] = (mid_1[1871:1864] > btm_2[1871:1864]) ? 1 : 0;
assign detect_max[232][25] = (mid_1[1871:1864] > btm_2[1879:1872]) ? 1 : 0;

assign detect_max[233][0] = (mid_1[1879:1872] > top_0[1871:1864]) ? 1 : 0;
assign detect_max[233][1] = (mid_1[1879:1872] > top_0[1879:1872]) ? 1 : 0;
assign detect_max[233][2] = (mid_1[1879:1872] > top_0[1887:1880]) ? 1 : 0;
assign detect_max[233][3] = (mid_1[1879:1872] > top_1[1871:1864]) ? 1 : 0;
assign detect_max[233][4] = (mid_1[1879:1872] > top_1[1879:1872]) ? 1 : 0;
assign detect_max[233][5] = (mid_1[1879:1872] > top_1[1887:1880]) ? 1 : 0;
assign detect_max[233][6] = (mid_1[1879:1872] > top_2[1871:1864]) ? 1 : 0;
assign detect_max[233][7] = (mid_1[1879:1872] > top_2[1879:1872]) ? 1 : 0;
assign detect_max[233][8] = (mid_1[1879:1872] > top_2[1887:1880]) ? 1 : 0;
assign detect_max[233][9] = (mid_1[1879:1872] > mid_0[1871:1864]) ? 1 : 0;
assign detect_max[233][10] = (mid_1[1879:1872] > mid_0[1879:1872]) ? 1 : 0;
assign detect_max[233][11] = (mid_1[1879:1872] > mid_0[1887:1880]) ? 1 : 0;
assign detect_max[233][12] = (mid_1[1879:1872] > mid_1[1871:1864]) ? 1 : 0;
assign detect_max[233][13] = (mid_1[1879:1872] > mid_1[1887:1880]) ? 1 : 0;
assign detect_max[233][14] = (mid_1[1879:1872] > mid_2[1871:1864]) ? 1 : 0;
assign detect_max[233][15] = (mid_1[1879:1872] > mid_2[1879:1872]) ? 1 : 0;
assign detect_max[233][16] = (mid_1[1879:1872] > mid_2[1887:1880]) ? 1 : 0;
assign detect_max[233][17] = (mid_1[1879:1872] > btm_0[1871:1864]) ? 1 : 0;
assign detect_max[233][18] = (mid_1[1879:1872] > btm_0[1879:1872]) ? 1 : 0;
assign detect_max[233][19] = (mid_1[1879:1872] > btm_0[1887:1880]) ? 1 : 0;
assign detect_max[233][20] = (mid_1[1879:1872] > btm_1[1871:1864]) ? 1 : 0;
assign detect_max[233][21] = (mid_1[1879:1872] > btm_1[1879:1872]) ? 1 : 0;
assign detect_max[233][22] = (mid_1[1879:1872] > btm_1[1887:1880]) ? 1 : 0;
assign detect_max[233][23] = (mid_1[1879:1872] > btm_2[1871:1864]) ? 1 : 0;
assign detect_max[233][24] = (mid_1[1879:1872] > btm_2[1879:1872]) ? 1 : 0;
assign detect_max[233][25] = (mid_1[1879:1872] > btm_2[1887:1880]) ? 1 : 0;

assign detect_max[234][0] = (mid_1[1887:1880] > top_0[1879:1872]) ? 1 : 0;
assign detect_max[234][1] = (mid_1[1887:1880] > top_0[1887:1880]) ? 1 : 0;
assign detect_max[234][2] = (mid_1[1887:1880] > top_0[1895:1888]) ? 1 : 0;
assign detect_max[234][3] = (mid_1[1887:1880] > top_1[1879:1872]) ? 1 : 0;
assign detect_max[234][4] = (mid_1[1887:1880] > top_1[1887:1880]) ? 1 : 0;
assign detect_max[234][5] = (mid_1[1887:1880] > top_1[1895:1888]) ? 1 : 0;
assign detect_max[234][6] = (mid_1[1887:1880] > top_2[1879:1872]) ? 1 : 0;
assign detect_max[234][7] = (mid_1[1887:1880] > top_2[1887:1880]) ? 1 : 0;
assign detect_max[234][8] = (mid_1[1887:1880] > top_2[1895:1888]) ? 1 : 0;
assign detect_max[234][9] = (mid_1[1887:1880] > mid_0[1879:1872]) ? 1 : 0;
assign detect_max[234][10] = (mid_1[1887:1880] > mid_0[1887:1880]) ? 1 : 0;
assign detect_max[234][11] = (mid_1[1887:1880] > mid_0[1895:1888]) ? 1 : 0;
assign detect_max[234][12] = (mid_1[1887:1880] > mid_1[1879:1872]) ? 1 : 0;
assign detect_max[234][13] = (mid_1[1887:1880] > mid_1[1895:1888]) ? 1 : 0;
assign detect_max[234][14] = (mid_1[1887:1880] > mid_2[1879:1872]) ? 1 : 0;
assign detect_max[234][15] = (mid_1[1887:1880] > mid_2[1887:1880]) ? 1 : 0;
assign detect_max[234][16] = (mid_1[1887:1880] > mid_2[1895:1888]) ? 1 : 0;
assign detect_max[234][17] = (mid_1[1887:1880] > btm_0[1879:1872]) ? 1 : 0;
assign detect_max[234][18] = (mid_1[1887:1880] > btm_0[1887:1880]) ? 1 : 0;
assign detect_max[234][19] = (mid_1[1887:1880] > btm_0[1895:1888]) ? 1 : 0;
assign detect_max[234][20] = (mid_1[1887:1880] > btm_1[1879:1872]) ? 1 : 0;
assign detect_max[234][21] = (mid_1[1887:1880] > btm_1[1887:1880]) ? 1 : 0;
assign detect_max[234][22] = (mid_1[1887:1880] > btm_1[1895:1888]) ? 1 : 0;
assign detect_max[234][23] = (mid_1[1887:1880] > btm_2[1879:1872]) ? 1 : 0;
assign detect_max[234][24] = (mid_1[1887:1880] > btm_2[1887:1880]) ? 1 : 0;
assign detect_max[234][25] = (mid_1[1887:1880] > btm_2[1895:1888]) ? 1 : 0;

assign detect_max[235][0] = (mid_1[1895:1888] > top_0[1887:1880]) ? 1 : 0;
assign detect_max[235][1] = (mid_1[1895:1888] > top_0[1895:1888]) ? 1 : 0;
assign detect_max[235][2] = (mid_1[1895:1888] > top_0[1903:1896]) ? 1 : 0;
assign detect_max[235][3] = (mid_1[1895:1888] > top_1[1887:1880]) ? 1 : 0;
assign detect_max[235][4] = (mid_1[1895:1888] > top_1[1895:1888]) ? 1 : 0;
assign detect_max[235][5] = (mid_1[1895:1888] > top_1[1903:1896]) ? 1 : 0;
assign detect_max[235][6] = (mid_1[1895:1888] > top_2[1887:1880]) ? 1 : 0;
assign detect_max[235][7] = (mid_1[1895:1888] > top_2[1895:1888]) ? 1 : 0;
assign detect_max[235][8] = (mid_1[1895:1888] > top_2[1903:1896]) ? 1 : 0;
assign detect_max[235][9] = (mid_1[1895:1888] > mid_0[1887:1880]) ? 1 : 0;
assign detect_max[235][10] = (mid_1[1895:1888] > mid_0[1895:1888]) ? 1 : 0;
assign detect_max[235][11] = (mid_1[1895:1888] > mid_0[1903:1896]) ? 1 : 0;
assign detect_max[235][12] = (mid_1[1895:1888] > mid_1[1887:1880]) ? 1 : 0;
assign detect_max[235][13] = (mid_1[1895:1888] > mid_1[1903:1896]) ? 1 : 0;
assign detect_max[235][14] = (mid_1[1895:1888] > mid_2[1887:1880]) ? 1 : 0;
assign detect_max[235][15] = (mid_1[1895:1888] > mid_2[1895:1888]) ? 1 : 0;
assign detect_max[235][16] = (mid_1[1895:1888] > mid_2[1903:1896]) ? 1 : 0;
assign detect_max[235][17] = (mid_1[1895:1888] > btm_0[1887:1880]) ? 1 : 0;
assign detect_max[235][18] = (mid_1[1895:1888] > btm_0[1895:1888]) ? 1 : 0;
assign detect_max[235][19] = (mid_1[1895:1888] > btm_0[1903:1896]) ? 1 : 0;
assign detect_max[235][20] = (mid_1[1895:1888] > btm_1[1887:1880]) ? 1 : 0;
assign detect_max[235][21] = (mid_1[1895:1888] > btm_1[1895:1888]) ? 1 : 0;
assign detect_max[235][22] = (mid_1[1895:1888] > btm_1[1903:1896]) ? 1 : 0;
assign detect_max[235][23] = (mid_1[1895:1888] > btm_2[1887:1880]) ? 1 : 0;
assign detect_max[235][24] = (mid_1[1895:1888] > btm_2[1895:1888]) ? 1 : 0;
assign detect_max[235][25] = (mid_1[1895:1888] > btm_2[1903:1896]) ? 1 : 0;

assign detect_max[236][0] = (mid_1[1903:1896] > top_0[1895:1888]) ? 1 : 0;
assign detect_max[236][1] = (mid_1[1903:1896] > top_0[1903:1896]) ? 1 : 0;
assign detect_max[236][2] = (mid_1[1903:1896] > top_0[1911:1904]) ? 1 : 0;
assign detect_max[236][3] = (mid_1[1903:1896] > top_1[1895:1888]) ? 1 : 0;
assign detect_max[236][4] = (mid_1[1903:1896] > top_1[1903:1896]) ? 1 : 0;
assign detect_max[236][5] = (mid_1[1903:1896] > top_1[1911:1904]) ? 1 : 0;
assign detect_max[236][6] = (mid_1[1903:1896] > top_2[1895:1888]) ? 1 : 0;
assign detect_max[236][7] = (mid_1[1903:1896] > top_2[1903:1896]) ? 1 : 0;
assign detect_max[236][8] = (mid_1[1903:1896] > top_2[1911:1904]) ? 1 : 0;
assign detect_max[236][9] = (mid_1[1903:1896] > mid_0[1895:1888]) ? 1 : 0;
assign detect_max[236][10] = (mid_1[1903:1896] > mid_0[1903:1896]) ? 1 : 0;
assign detect_max[236][11] = (mid_1[1903:1896] > mid_0[1911:1904]) ? 1 : 0;
assign detect_max[236][12] = (mid_1[1903:1896] > mid_1[1895:1888]) ? 1 : 0;
assign detect_max[236][13] = (mid_1[1903:1896] > mid_1[1911:1904]) ? 1 : 0;
assign detect_max[236][14] = (mid_1[1903:1896] > mid_2[1895:1888]) ? 1 : 0;
assign detect_max[236][15] = (mid_1[1903:1896] > mid_2[1903:1896]) ? 1 : 0;
assign detect_max[236][16] = (mid_1[1903:1896] > mid_2[1911:1904]) ? 1 : 0;
assign detect_max[236][17] = (mid_1[1903:1896] > btm_0[1895:1888]) ? 1 : 0;
assign detect_max[236][18] = (mid_1[1903:1896] > btm_0[1903:1896]) ? 1 : 0;
assign detect_max[236][19] = (mid_1[1903:1896] > btm_0[1911:1904]) ? 1 : 0;
assign detect_max[236][20] = (mid_1[1903:1896] > btm_1[1895:1888]) ? 1 : 0;
assign detect_max[236][21] = (mid_1[1903:1896] > btm_1[1903:1896]) ? 1 : 0;
assign detect_max[236][22] = (mid_1[1903:1896] > btm_1[1911:1904]) ? 1 : 0;
assign detect_max[236][23] = (mid_1[1903:1896] > btm_2[1895:1888]) ? 1 : 0;
assign detect_max[236][24] = (mid_1[1903:1896] > btm_2[1903:1896]) ? 1 : 0;
assign detect_max[236][25] = (mid_1[1903:1896] > btm_2[1911:1904]) ? 1 : 0;

assign detect_max[237][0] = (mid_1[1911:1904] > top_0[1903:1896]) ? 1 : 0;
assign detect_max[237][1] = (mid_1[1911:1904] > top_0[1911:1904]) ? 1 : 0;
assign detect_max[237][2] = (mid_1[1911:1904] > top_0[1919:1912]) ? 1 : 0;
assign detect_max[237][3] = (mid_1[1911:1904] > top_1[1903:1896]) ? 1 : 0;
assign detect_max[237][4] = (mid_1[1911:1904] > top_1[1911:1904]) ? 1 : 0;
assign detect_max[237][5] = (mid_1[1911:1904] > top_1[1919:1912]) ? 1 : 0;
assign detect_max[237][6] = (mid_1[1911:1904] > top_2[1903:1896]) ? 1 : 0;
assign detect_max[237][7] = (mid_1[1911:1904] > top_2[1911:1904]) ? 1 : 0;
assign detect_max[237][8] = (mid_1[1911:1904] > top_2[1919:1912]) ? 1 : 0;
assign detect_max[237][9] = (mid_1[1911:1904] > mid_0[1903:1896]) ? 1 : 0;
assign detect_max[237][10] = (mid_1[1911:1904] > mid_0[1911:1904]) ? 1 : 0;
assign detect_max[237][11] = (mid_1[1911:1904] > mid_0[1919:1912]) ? 1 : 0;
assign detect_max[237][12] = (mid_1[1911:1904] > mid_1[1903:1896]) ? 1 : 0;
assign detect_max[237][13] = (mid_1[1911:1904] > mid_1[1919:1912]) ? 1 : 0;
assign detect_max[237][14] = (mid_1[1911:1904] > mid_2[1903:1896]) ? 1 : 0;
assign detect_max[237][15] = (mid_1[1911:1904] > mid_2[1911:1904]) ? 1 : 0;
assign detect_max[237][16] = (mid_1[1911:1904] > mid_2[1919:1912]) ? 1 : 0;
assign detect_max[237][17] = (mid_1[1911:1904] > btm_0[1903:1896]) ? 1 : 0;
assign detect_max[237][18] = (mid_1[1911:1904] > btm_0[1911:1904]) ? 1 : 0;
assign detect_max[237][19] = (mid_1[1911:1904] > btm_0[1919:1912]) ? 1 : 0;
assign detect_max[237][20] = (mid_1[1911:1904] > btm_1[1903:1896]) ? 1 : 0;
assign detect_max[237][21] = (mid_1[1911:1904] > btm_1[1911:1904]) ? 1 : 0;
assign detect_max[237][22] = (mid_1[1911:1904] > btm_1[1919:1912]) ? 1 : 0;
assign detect_max[237][23] = (mid_1[1911:1904] > btm_2[1903:1896]) ? 1 : 0;
assign detect_max[237][24] = (mid_1[1911:1904] > btm_2[1911:1904]) ? 1 : 0;
assign detect_max[237][25] = (mid_1[1911:1904] > btm_2[1919:1912]) ? 1 : 0;

assign detect_max[238][0] = (mid_1[1919:1912] > top_0[1911:1904]) ? 1 : 0;
assign detect_max[238][1] = (mid_1[1919:1912] > top_0[1919:1912]) ? 1 : 0;
assign detect_max[238][2] = (mid_1[1919:1912] > top_0[1927:1920]) ? 1 : 0;
assign detect_max[238][3] = (mid_1[1919:1912] > top_1[1911:1904]) ? 1 : 0;
assign detect_max[238][4] = (mid_1[1919:1912] > top_1[1919:1912]) ? 1 : 0;
assign detect_max[238][5] = (mid_1[1919:1912] > top_1[1927:1920]) ? 1 : 0;
assign detect_max[238][6] = (mid_1[1919:1912] > top_2[1911:1904]) ? 1 : 0;
assign detect_max[238][7] = (mid_1[1919:1912] > top_2[1919:1912]) ? 1 : 0;
assign detect_max[238][8] = (mid_1[1919:1912] > top_2[1927:1920]) ? 1 : 0;
assign detect_max[238][9] = (mid_1[1919:1912] > mid_0[1911:1904]) ? 1 : 0;
assign detect_max[238][10] = (mid_1[1919:1912] > mid_0[1919:1912]) ? 1 : 0;
assign detect_max[238][11] = (mid_1[1919:1912] > mid_0[1927:1920]) ? 1 : 0;
assign detect_max[238][12] = (mid_1[1919:1912] > mid_1[1911:1904]) ? 1 : 0;
assign detect_max[238][13] = (mid_1[1919:1912] > mid_1[1927:1920]) ? 1 : 0;
assign detect_max[238][14] = (mid_1[1919:1912] > mid_2[1911:1904]) ? 1 : 0;
assign detect_max[238][15] = (mid_1[1919:1912] > mid_2[1919:1912]) ? 1 : 0;
assign detect_max[238][16] = (mid_1[1919:1912] > mid_2[1927:1920]) ? 1 : 0;
assign detect_max[238][17] = (mid_1[1919:1912] > btm_0[1911:1904]) ? 1 : 0;
assign detect_max[238][18] = (mid_1[1919:1912] > btm_0[1919:1912]) ? 1 : 0;
assign detect_max[238][19] = (mid_1[1919:1912] > btm_0[1927:1920]) ? 1 : 0;
assign detect_max[238][20] = (mid_1[1919:1912] > btm_1[1911:1904]) ? 1 : 0;
assign detect_max[238][21] = (mid_1[1919:1912] > btm_1[1919:1912]) ? 1 : 0;
assign detect_max[238][22] = (mid_1[1919:1912] > btm_1[1927:1920]) ? 1 : 0;
assign detect_max[238][23] = (mid_1[1919:1912] > btm_2[1911:1904]) ? 1 : 0;
assign detect_max[238][24] = (mid_1[1919:1912] > btm_2[1919:1912]) ? 1 : 0;
assign detect_max[238][25] = (mid_1[1919:1912] > btm_2[1927:1920]) ? 1 : 0;

assign detect_max[239][0] = (mid_1[1927:1920] > top_0[1919:1912]) ? 1 : 0;
assign detect_max[239][1] = (mid_1[1927:1920] > top_0[1927:1920]) ? 1 : 0;
assign detect_max[239][2] = (mid_1[1927:1920] > top_0[1935:1928]) ? 1 : 0;
assign detect_max[239][3] = (mid_1[1927:1920] > top_1[1919:1912]) ? 1 : 0;
assign detect_max[239][4] = (mid_1[1927:1920] > top_1[1927:1920]) ? 1 : 0;
assign detect_max[239][5] = (mid_1[1927:1920] > top_1[1935:1928]) ? 1 : 0;
assign detect_max[239][6] = (mid_1[1927:1920] > top_2[1919:1912]) ? 1 : 0;
assign detect_max[239][7] = (mid_1[1927:1920] > top_2[1927:1920]) ? 1 : 0;
assign detect_max[239][8] = (mid_1[1927:1920] > top_2[1935:1928]) ? 1 : 0;
assign detect_max[239][9] = (mid_1[1927:1920] > mid_0[1919:1912]) ? 1 : 0;
assign detect_max[239][10] = (mid_1[1927:1920] > mid_0[1927:1920]) ? 1 : 0;
assign detect_max[239][11] = (mid_1[1927:1920] > mid_0[1935:1928]) ? 1 : 0;
assign detect_max[239][12] = (mid_1[1927:1920] > mid_1[1919:1912]) ? 1 : 0;
assign detect_max[239][13] = (mid_1[1927:1920] > mid_1[1935:1928]) ? 1 : 0;
assign detect_max[239][14] = (mid_1[1927:1920] > mid_2[1919:1912]) ? 1 : 0;
assign detect_max[239][15] = (mid_1[1927:1920] > mid_2[1927:1920]) ? 1 : 0;
assign detect_max[239][16] = (mid_1[1927:1920] > mid_2[1935:1928]) ? 1 : 0;
assign detect_max[239][17] = (mid_1[1927:1920] > btm_0[1919:1912]) ? 1 : 0;
assign detect_max[239][18] = (mid_1[1927:1920] > btm_0[1927:1920]) ? 1 : 0;
assign detect_max[239][19] = (mid_1[1927:1920] > btm_0[1935:1928]) ? 1 : 0;
assign detect_max[239][20] = (mid_1[1927:1920] > btm_1[1919:1912]) ? 1 : 0;
assign detect_max[239][21] = (mid_1[1927:1920] > btm_1[1927:1920]) ? 1 : 0;
assign detect_max[239][22] = (mid_1[1927:1920] > btm_1[1935:1928]) ? 1 : 0;
assign detect_max[239][23] = (mid_1[1927:1920] > btm_2[1919:1912]) ? 1 : 0;
assign detect_max[239][24] = (mid_1[1927:1920] > btm_2[1927:1920]) ? 1 : 0;
assign detect_max[239][25] = (mid_1[1927:1920] > btm_2[1935:1928]) ? 1 : 0;

assign detect_max[240][0] = (mid_1[1935:1928] > top_0[1927:1920]) ? 1 : 0;
assign detect_max[240][1] = (mid_1[1935:1928] > top_0[1935:1928]) ? 1 : 0;
assign detect_max[240][2] = (mid_1[1935:1928] > top_0[1943:1936]) ? 1 : 0;
assign detect_max[240][3] = (mid_1[1935:1928] > top_1[1927:1920]) ? 1 : 0;
assign detect_max[240][4] = (mid_1[1935:1928] > top_1[1935:1928]) ? 1 : 0;
assign detect_max[240][5] = (mid_1[1935:1928] > top_1[1943:1936]) ? 1 : 0;
assign detect_max[240][6] = (mid_1[1935:1928] > top_2[1927:1920]) ? 1 : 0;
assign detect_max[240][7] = (mid_1[1935:1928] > top_2[1935:1928]) ? 1 : 0;
assign detect_max[240][8] = (mid_1[1935:1928] > top_2[1943:1936]) ? 1 : 0;
assign detect_max[240][9] = (mid_1[1935:1928] > mid_0[1927:1920]) ? 1 : 0;
assign detect_max[240][10] = (mid_1[1935:1928] > mid_0[1935:1928]) ? 1 : 0;
assign detect_max[240][11] = (mid_1[1935:1928] > mid_0[1943:1936]) ? 1 : 0;
assign detect_max[240][12] = (mid_1[1935:1928] > mid_1[1927:1920]) ? 1 : 0;
assign detect_max[240][13] = (mid_1[1935:1928] > mid_1[1943:1936]) ? 1 : 0;
assign detect_max[240][14] = (mid_1[1935:1928] > mid_2[1927:1920]) ? 1 : 0;
assign detect_max[240][15] = (mid_1[1935:1928] > mid_2[1935:1928]) ? 1 : 0;
assign detect_max[240][16] = (mid_1[1935:1928] > mid_2[1943:1936]) ? 1 : 0;
assign detect_max[240][17] = (mid_1[1935:1928] > btm_0[1927:1920]) ? 1 : 0;
assign detect_max[240][18] = (mid_1[1935:1928] > btm_0[1935:1928]) ? 1 : 0;
assign detect_max[240][19] = (mid_1[1935:1928] > btm_0[1943:1936]) ? 1 : 0;
assign detect_max[240][20] = (mid_1[1935:1928] > btm_1[1927:1920]) ? 1 : 0;
assign detect_max[240][21] = (mid_1[1935:1928] > btm_1[1935:1928]) ? 1 : 0;
assign detect_max[240][22] = (mid_1[1935:1928] > btm_1[1943:1936]) ? 1 : 0;
assign detect_max[240][23] = (mid_1[1935:1928] > btm_2[1927:1920]) ? 1 : 0;
assign detect_max[240][24] = (mid_1[1935:1928] > btm_2[1935:1928]) ? 1 : 0;
assign detect_max[240][25] = (mid_1[1935:1928] > btm_2[1943:1936]) ? 1 : 0;

assign detect_max[241][0] = (mid_1[1943:1936] > top_0[1935:1928]) ? 1 : 0;
assign detect_max[241][1] = (mid_1[1943:1936] > top_0[1943:1936]) ? 1 : 0;
assign detect_max[241][2] = (mid_1[1943:1936] > top_0[1951:1944]) ? 1 : 0;
assign detect_max[241][3] = (mid_1[1943:1936] > top_1[1935:1928]) ? 1 : 0;
assign detect_max[241][4] = (mid_1[1943:1936] > top_1[1943:1936]) ? 1 : 0;
assign detect_max[241][5] = (mid_1[1943:1936] > top_1[1951:1944]) ? 1 : 0;
assign detect_max[241][6] = (mid_1[1943:1936] > top_2[1935:1928]) ? 1 : 0;
assign detect_max[241][7] = (mid_1[1943:1936] > top_2[1943:1936]) ? 1 : 0;
assign detect_max[241][8] = (mid_1[1943:1936] > top_2[1951:1944]) ? 1 : 0;
assign detect_max[241][9] = (mid_1[1943:1936] > mid_0[1935:1928]) ? 1 : 0;
assign detect_max[241][10] = (mid_1[1943:1936] > mid_0[1943:1936]) ? 1 : 0;
assign detect_max[241][11] = (mid_1[1943:1936] > mid_0[1951:1944]) ? 1 : 0;
assign detect_max[241][12] = (mid_1[1943:1936] > mid_1[1935:1928]) ? 1 : 0;
assign detect_max[241][13] = (mid_1[1943:1936] > mid_1[1951:1944]) ? 1 : 0;
assign detect_max[241][14] = (mid_1[1943:1936] > mid_2[1935:1928]) ? 1 : 0;
assign detect_max[241][15] = (mid_1[1943:1936] > mid_2[1943:1936]) ? 1 : 0;
assign detect_max[241][16] = (mid_1[1943:1936] > mid_2[1951:1944]) ? 1 : 0;
assign detect_max[241][17] = (mid_1[1943:1936] > btm_0[1935:1928]) ? 1 : 0;
assign detect_max[241][18] = (mid_1[1943:1936] > btm_0[1943:1936]) ? 1 : 0;
assign detect_max[241][19] = (mid_1[1943:1936] > btm_0[1951:1944]) ? 1 : 0;
assign detect_max[241][20] = (mid_1[1943:1936] > btm_1[1935:1928]) ? 1 : 0;
assign detect_max[241][21] = (mid_1[1943:1936] > btm_1[1943:1936]) ? 1 : 0;
assign detect_max[241][22] = (mid_1[1943:1936] > btm_1[1951:1944]) ? 1 : 0;
assign detect_max[241][23] = (mid_1[1943:1936] > btm_2[1935:1928]) ? 1 : 0;
assign detect_max[241][24] = (mid_1[1943:1936] > btm_2[1943:1936]) ? 1 : 0;
assign detect_max[241][25] = (mid_1[1943:1936] > btm_2[1951:1944]) ? 1 : 0;

assign detect_max[242][0] = (mid_1[1951:1944] > top_0[1943:1936]) ? 1 : 0;
assign detect_max[242][1] = (mid_1[1951:1944] > top_0[1951:1944]) ? 1 : 0;
assign detect_max[242][2] = (mid_1[1951:1944] > top_0[1959:1952]) ? 1 : 0;
assign detect_max[242][3] = (mid_1[1951:1944] > top_1[1943:1936]) ? 1 : 0;
assign detect_max[242][4] = (mid_1[1951:1944] > top_1[1951:1944]) ? 1 : 0;
assign detect_max[242][5] = (mid_1[1951:1944] > top_1[1959:1952]) ? 1 : 0;
assign detect_max[242][6] = (mid_1[1951:1944] > top_2[1943:1936]) ? 1 : 0;
assign detect_max[242][7] = (mid_1[1951:1944] > top_2[1951:1944]) ? 1 : 0;
assign detect_max[242][8] = (mid_1[1951:1944] > top_2[1959:1952]) ? 1 : 0;
assign detect_max[242][9] = (mid_1[1951:1944] > mid_0[1943:1936]) ? 1 : 0;
assign detect_max[242][10] = (mid_1[1951:1944] > mid_0[1951:1944]) ? 1 : 0;
assign detect_max[242][11] = (mid_1[1951:1944] > mid_0[1959:1952]) ? 1 : 0;
assign detect_max[242][12] = (mid_1[1951:1944] > mid_1[1943:1936]) ? 1 : 0;
assign detect_max[242][13] = (mid_1[1951:1944] > mid_1[1959:1952]) ? 1 : 0;
assign detect_max[242][14] = (mid_1[1951:1944] > mid_2[1943:1936]) ? 1 : 0;
assign detect_max[242][15] = (mid_1[1951:1944] > mid_2[1951:1944]) ? 1 : 0;
assign detect_max[242][16] = (mid_1[1951:1944] > mid_2[1959:1952]) ? 1 : 0;
assign detect_max[242][17] = (mid_1[1951:1944] > btm_0[1943:1936]) ? 1 : 0;
assign detect_max[242][18] = (mid_1[1951:1944] > btm_0[1951:1944]) ? 1 : 0;
assign detect_max[242][19] = (mid_1[1951:1944] > btm_0[1959:1952]) ? 1 : 0;
assign detect_max[242][20] = (mid_1[1951:1944] > btm_1[1943:1936]) ? 1 : 0;
assign detect_max[242][21] = (mid_1[1951:1944] > btm_1[1951:1944]) ? 1 : 0;
assign detect_max[242][22] = (mid_1[1951:1944] > btm_1[1959:1952]) ? 1 : 0;
assign detect_max[242][23] = (mid_1[1951:1944] > btm_2[1943:1936]) ? 1 : 0;
assign detect_max[242][24] = (mid_1[1951:1944] > btm_2[1951:1944]) ? 1 : 0;
assign detect_max[242][25] = (mid_1[1951:1944] > btm_2[1959:1952]) ? 1 : 0;

assign detect_max[243][0] = (mid_1[1959:1952] > top_0[1951:1944]) ? 1 : 0;
assign detect_max[243][1] = (mid_1[1959:1952] > top_0[1959:1952]) ? 1 : 0;
assign detect_max[243][2] = (mid_1[1959:1952] > top_0[1967:1960]) ? 1 : 0;
assign detect_max[243][3] = (mid_1[1959:1952] > top_1[1951:1944]) ? 1 : 0;
assign detect_max[243][4] = (mid_1[1959:1952] > top_1[1959:1952]) ? 1 : 0;
assign detect_max[243][5] = (mid_1[1959:1952] > top_1[1967:1960]) ? 1 : 0;
assign detect_max[243][6] = (mid_1[1959:1952] > top_2[1951:1944]) ? 1 : 0;
assign detect_max[243][7] = (mid_1[1959:1952] > top_2[1959:1952]) ? 1 : 0;
assign detect_max[243][8] = (mid_1[1959:1952] > top_2[1967:1960]) ? 1 : 0;
assign detect_max[243][9] = (mid_1[1959:1952] > mid_0[1951:1944]) ? 1 : 0;
assign detect_max[243][10] = (mid_1[1959:1952] > mid_0[1959:1952]) ? 1 : 0;
assign detect_max[243][11] = (mid_1[1959:1952] > mid_0[1967:1960]) ? 1 : 0;
assign detect_max[243][12] = (mid_1[1959:1952] > mid_1[1951:1944]) ? 1 : 0;
assign detect_max[243][13] = (mid_1[1959:1952] > mid_1[1967:1960]) ? 1 : 0;
assign detect_max[243][14] = (mid_1[1959:1952] > mid_2[1951:1944]) ? 1 : 0;
assign detect_max[243][15] = (mid_1[1959:1952] > mid_2[1959:1952]) ? 1 : 0;
assign detect_max[243][16] = (mid_1[1959:1952] > mid_2[1967:1960]) ? 1 : 0;
assign detect_max[243][17] = (mid_1[1959:1952] > btm_0[1951:1944]) ? 1 : 0;
assign detect_max[243][18] = (mid_1[1959:1952] > btm_0[1959:1952]) ? 1 : 0;
assign detect_max[243][19] = (mid_1[1959:1952] > btm_0[1967:1960]) ? 1 : 0;
assign detect_max[243][20] = (mid_1[1959:1952] > btm_1[1951:1944]) ? 1 : 0;
assign detect_max[243][21] = (mid_1[1959:1952] > btm_1[1959:1952]) ? 1 : 0;
assign detect_max[243][22] = (mid_1[1959:1952] > btm_1[1967:1960]) ? 1 : 0;
assign detect_max[243][23] = (mid_1[1959:1952] > btm_2[1951:1944]) ? 1 : 0;
assign detect_max[243][24] = (mid_1[1959:1952] > btm_2[1959:1952]) ? 1 : 0;
assign detect_max[243][25] = (mid_1[1959:1952] > btm_2[1967:1960]) ? 1 : 0;

assign detect_max[244][0] = (mid_1[1967:1960] > top_0[1959:1952]) ? 1 : 0;
assign detect_max[244][1] = (mid_1[1967:1960] > top_0[1967:1960]) ? 1 : 0;
assign detect_max[244][2] = (mid_1[1967:1960] > top_0[1975:1968]) ? 1 : 0;
assign detect_max[244][3] = (mid_1[1967:1960] > top_1[1959:1952]) ? 1 : 0;
assign detect_max[244][4] = (mid_1[1967:1960] > top_1[1967:1960]) ? 1 : 0;
assign detect_max[244][5] = (mid_1[1967:1960] > top_1[1975:1968]) ? 1 : 0;
assign detect_max[244][6] = (mid_1[1967:1960] > top_2[1959:1952]) ? 1 : 0;
assign detect_max[244][7] = (mid_1[1967:1960] > top_2[1967:1960]) ? 1 : 0;
assign detect_max[244][8] = (mid_1[1967:1960] > top_2[1975:1968]) ? 1 : 0;
assign detect_max[244][9] = (mid_1[1967:1960] > mid_0[1959:1952]) ? 1 : 0;
assign detect_max[244][10] = (mid_1[1967:1960] > mid_0[1967:1960]) ? 1 : 0;
assign detect_max[244][11] = (mid_1[1967:1960] > mid_0[1975:1968]) ? 1 : 0;
assign detect_max[244][12] = (mid_1[1967:1960] > mid_1[1959:1952]) ? 1 : 0;
assign detect_max[244][13] = (mid_1[1967:1960] > mid_1[1975:1968]) ? 1 : 0;
assign detect_max[244][14] = (mid_1[1967:1960] > mid_2[1959:1952]) ? 1 : 0;
assign detect_max[244][15] = (mid_1[1967:1960] > mid_2[1967:1960]) ? 1 : 0;
assign detect_max[244][16] = (mid_1[1967:1960] > mid_2[1975:1968]) ? 1 : 0;
assign detect_max[244][17] = (mid_1[1967:1960] > btm_0[1959:1952]) ? 1 : 0;
assign detect_max[244][18] = (mid_1[1967:1960] > btm_0[1967:1960]) ? 1 : 0;
assign detect_max[244][19] = (mid_1[1967:1960] > btm_0[1975:1968]) ? 1 : 0;
assign detect_max[244][20] = (mid_1[1967:1960] > btm_1[1959:1952]) ? 1 : 0;
assign detect_max[244][21] = (mid_1[1967:1960] > btm_1[1967:1960]) ? 1 : 0;
assign detect_max[244][22] = (mid_1[1967:1960] > btm_1[1975:1968]) ? 1 : 0;
assign detect_max[244][23] = (mid_1[1967:1960] > btm_2[1959:1952]) ? 1 : 0;
assign detect_max[244][24] = (mid_1[1967:1960] > btm_2[1967:1960]) ? 1 : 0;
assign detect_max[244][25] = (mid_1[1967:1960] > btm_2[1975:1968]) ? 1 : 0;

assign detect_max[245][0] = (mid_1[1975:1968] > top_0[1967:1960]) ? 1 : 0;
assign detect_max[245][1] = (mid_1[1975:1968] > top_0[1975:1968]) ? 1 : 0;
assign detect_max[245][2] = (mid_1[1975:1968] > top_0[1983:1976]) ? 1 : 0;
assign detect_max[245][3] = (mid_1[1975:1968] > top_1[1967:1960]) ? 1 : 0;
assign detect_max[245][4] = (mid_1[1975:1968] > top_1[1975:1968]) ? 1 : 0;
assign detect_max[245][5] = (mid_1[1975:1968] > top_1[1983:1976]) ? 1 : 0;
assign detect_max[245][6] = (mid_1[1975:1968] > top_2[1967:1960]) ? 1 : 0;
assign detect_max[245][7] = (mid_1[1975:1968] > top_2[1975:1968]) ? 1 : 0;
assign detect_max[245][8] = (mid_1[1975:1968] > top_2[1983:1976]) ? 1 : 0;
assign detect_max[245][9] = (mid_1[1975:1968] > mid_0[1967:1960]) ? 1 : 0;
assign detect_max[245][10] = (mid_1[1975:1968] > mid_0[1975:1968]) ? 1 : 0;
assign detect_max[245][11] = (mid_1[1975:1968] > mid_0[1983:1976]) ? 1 : 0;
assign detect_max[245][12] = (mid_1[1975:1968] > mid_1[1967:1960]) ? 1 : 0;
assign detect_max[245][13] = (mid_1[1975:1968] > mid_1[1983:1976]) ? 1 : 0;
assign detect_max[245][14] = (mid_1[1975:1968] > mid_2[1967:1960]) ? 1 : 0;
assign detect_max[245][15] = (mid_1[1975:1968] > mid_2[1975:1968]) ? 1 : 0;
assign detect_max[245][16] = (mid_1[1975:1968] > mid_2[1983:1976]) ? 1 : 0;
assign detect_max[245][17] = (mid_1[1975:1968] > btm_0[1967:1960]) ? 1 : 0;
assign detect_max[245][18] = (mid_1[1975:1968] > btm_0[1975:1968]) ? 1 : 0;
assign detect_max[245][19] = (mid_1[1975:1968] > btm_0[1983:1976]) ? 1 : 0;
assign detect_max[245][20] = (mid_1[1975:1968] > btm_1[1967:1960]) ? 1 : 0;
assign detect_max[245][21] = (mid_1[1975:1968] > btm_1[1975:1968]) ? 1 : 0;
assign detect_max[245][22] = (mid_1[1975:1968] > btm_1[1983:1976]) ? 1 : 0;
assign detect_max[245][23] = (mid_1[1975:1968] > btm_2[1967:1960]) ? 1 : 0;
assign detect_max[245][24] = (mid_1[1975:1968] > btm_2[1975:1968]) ? 1 : 0;
assign detect_max[245][25] = (mid_1[1975:1968] > btm_2[1983:1976]) ? 1 : 0;

assign detect_max[246][0] = (mid_1[1983:1976] > top_0[1975:1968]) ? 1 : 0;
assign detect_max[246][1] = (mid_1[1983:1976] > top_0[1983:1976]) ? 1 : 0;
assign detect_max[246][2] = (mid_1[1983:1976] > top_0[1991:1984]) ? 1 : 0;
assign detect_max[246][3] = (mid_1[1983:1976] > top_1[1975:1968]) ? 1 : 0;
assign detect_max[246][4] = (mid_1[1983:1976] > top_1[1983:1976]) ? 1 : 0;
assign detect_max[246][5] = (mid_1[1983:1976] > top_1[1991:1984]) ? 1 : 0;
assign detect_max[246][6] = (mid_1[1983:1976] > top_2[1975:1968]) ? 1 : 0;
assign detect_max[246][7] = (mid_1[1983:1976] > top_2[1983:1976]) ? 1 : 0;
assign detect_max[246][8] = (mid_1[1983:1976] > top_2[1991:1984]) ? 1 : 0;
assign detect_max[246][9] = (mid_1[1983:1976] > mid_0[1975:1968]) ? 1 : 0;
assign detect_max[246][10] = (mid_1[1983:1976] > mid_0[1983:1976]) ? 1 : 0;
assign detect_max[246][11] = (mid_1[1983:1976] > mid_0[1991:1984]) ? 1 : 0;
assign detect_max[246][12] = (mid_1[1983:1976] > mid_1[1975:1968]) ? 1 : 0;
assign detect_max[246][13] = (mid_1[1983:1976] > mid_1[1991:1984]) ? 1 : 0;
assign detect_max[246][14] = (mid_1[1983:1976] > mid_2[1975:1968]) ? 1 : 0;
assign detect_max[246][15] = (mid_1[1983:1976] > mid_2[1983:1976]) ? 1 : 0;
assign detect_max[246][16] = (mid_1[1983:1976] > mid_2[1991:1984]) ? 1 : 0;
assign detect_max[246][17] = (mid_1[1983:1976] > btm_0[1975:1968]) ? 1 : 0;
assign detect_max[246][18] = (mid_1[1983:1976] > btm_0[1983:1976]) ? 1 : 0;
assign detect_max[246][19] = (mid_1[1983:1976] > btm_0[1991:1984]) ? 1 : 0;
assign detect_max[246][20] = (mid_1[1983:1976] > btm_1[1975:1968]) ? 1 : 0;
assign detect_max[246][21] = (mid_1[1983:1976] > btm_1[1983:1976]) ? 1 : 0;
assign detect_max[246][22] = (mid_1[1983:1976] > btm_1[1991:1984]) ? 1 : 0;
assign detect_max[246][23] = (mid_1[1983:1976] > btm_2[1975:1968]) ? 1 : 0;
assign detect_max[246][24] = (mid_1[1983:1976] > btm_2[1983:1976]) ? 1 : 0;
assign detect_max[246][25] = (mid_1[1983:1976] > btm_2[1991:1984]) ? 1 : 0;

assign detect_max[247][0] = (mid_1[1991:1984] > top_0[1983:1976]) ? 1 : 0;
assign detect_max[247][1] = (mid_1[1991:1984] > top_0[1991:1984]) ? 1 : 0;
assign detect_max[247][2] = (mid_1[1991:1984] > top_0[1999:1992]) ? 1 : 0;
assign detect_max[247][3] = (mid_1[1991:1984] > top_1[1983:1976]) ? 1 : 0;
assign detect_max[247][4] = (mid_1[1991:1984] > top_1[1991:1984]) ? 1 : 0;
assign detect_max[247][5] = (mid_1[1991:1984] > top_1[1999:1992]) ? 1 : 0;
assign detect_max[247][6] = (mid_1[1991:1984] > top_2[1983:1976]) ? 1 : 0;
assign detect_max[247][7] = (mid_1[1991:1984] > top_2[1991:1984]) ? 1 : 0;
assign detect_max[247][8] = (mid_1[1991:1984] > top_2[1999:1992]) ? 1 : 0;
assign detect_max[247][9] = (mid_1[1991:1984] > mid_0[1983:1976]) ? 1 : 0;
assign detect_max[247][10] = (mid_1[1991:1984] > mid_0[1991:1984]) ? 1 : 0;
assign detect_max[247][11] = (mid_1[1991:1984] > mid_0[1999:1992]) ? 1 : 0;
assign detect_max[247][12] = (mid_1[1991:1984] > mid_1[1983:1976]) ? 1 : 0;
assign detect_max[247][13] = (mid_1[1991:1984] > mid_1[1999:1992]) ? 1 : 0;
assign detect_max[247][14] = (mid_1[1991:1984] > mid_2[1983:1976]) ? 1 : 0;
assign detect_max[247][15] = (mid_1[1991:1984] > mid_2[1991:1984]) ? 1 : 0;
assign detect_max[247][16] = (mid_1[1991:1984] > mid_2[1999:1992]) ? 1 : 0;
assign detect_max[247][17] = (mid_1[1991:1984] > btm_0[1983:1976]) ? 1 : 0;
assign detect_max[247][18] = (mid_1[1991:1984] > btm_0[1991:1984]) ? 1 : 0;
assign detect_max[247][19] = (mid_1[1991:1984] > btm_0[1999:1992]) ? 1 : 0;
assign detect_max[247][20] = (mid_1[1991:1984] > btm_1[1983:1976]) ? 1 : 0;
assign detect_max[247][21] = (mid_1[1991:1984] > btm_1[1991:1984]) ? 1 : 0;
assign detect_max[247][22] = (mid_1[1991:1984] > btm_1[1999:1992]) ? 1 : 0;
assign detect_max[247][23] = (mid_1[1991:1984] > btm_2[1983:1976]) ? 1 : 0;
assign detect_max[247][24] = (mid_1[1991:1984] > btm_2[1991:1984]) ? 1 : 0;
assign detect_max[247][25] = (mid_1[1991:1984] > btm_2[1999:1992]) ? 1 : 0;

assign detect_max[248][0] = (mid_1[1999:1992] > top_0[1991:1984]) ? 1 : 0;
assign detect_max[248][1] = (mid_1[1999:1992] > top_0[1999:1992]) ? 1 : 0;
assign detect_max[248][2] = (mid_1[1999:1992] > top_0[2007:2000]) ? 1 : 0;
assign detect_max[248][3] = (mid_1[1999:1992] > top_1[1991:1984]) ? 1 : 0;
assign detect_max[248][4] = (mid_1[1999:1992] > top_1[1999:1992]) ? 1 : 0;
assign detect_max[248][5] = (mid_1[1999:1992] > top_1[2007:2000]) ? 1 : 0;
assign detect_max[248][6] = (mid_1[1999:1992] > top_2[1991:1984]) ? 1 : 0;
assign detect_max[248][7] = (mid_1[1999:1992] > top_2[1999:1992]) ? 1 : 0;
assign detect_max[248][8] = (mid_1[1999:1992] > top_2[2007:2000]) ? 1 : 0;
assign detect_max[248][9] = (mid_1[1999:1992] > mid_0[1991:1984]) ? 1 : 0;
assign detect_max[248][10] = (mid_1[1999:1992] > mid_0[1999:1992]) ? 1 : 0;
assign detect_max[248][11] = (mid_1[1999:1992] > mid_0[2007:2000]) ? 1 : 0;
assign detect_max[248][12] = (mid_1[1999:1992] > mid_1[1991:1984]) ? 1 : 0;
assign detect_max[248][13] = (mid_1[1999:1992] > mid_1[2007:2000]) ? 1 : 0;
assign detect_max[248][14] = (mid_1[1999:1992] > mid_2[1991:1984]) ? 1 : 0;
assign detect_max[248][15] = (mid_1[1999:1992] > mid_2[1999:1992]) ? 1 : 0;
assign detect_max[248][16] = (mid_1[1999:1992] > mid_2[2007:2000]) ? 1 : 0;
assign detect_max[248][17] = (mid_1[1999:1992] > btm_0[1991:1984]) ? 1 : 0;
assign detect_max[248][18] = (mid_1[1999:1992] > btm_0[1999:1992]) ? 1 : 0;
assign detect_max[248][19] = (mid_1[1999:1992] > btm_0[2007:2000]) ? 1 : 0;
assign detect_max[248][20] = (mid_1[1999:1992] > btm_1[1991:1984]) ? 1 : 0;
assign detect_max[248][21] = (mid_1[1999:1992] > btm_1[1999:1992]) ? 1 : 0;
assign detect_max[248][22] = (mid_1[1999:1992] > btm_1[2007:2000]) ? 1 : 0;
assign detect_max[248][23] = (mid_1[1999:1992] > btm_2[1991:1984]) ? 1 : 0;
assign detect_max[248][24] = (mid_1[1999:1992] > btm_2[1999:1992]) ? 1 : 0;
assign detect_max[248][25] = (mid_1[1999:1992] > btm_2[2007:2000]) ? 1 : 0;

assign detect_max[249][0] = (mid_1[2007:2000] > top_0[1999:1992]) ? 1 : 0;
assign detect_max[249][1] = (mid_1[2007:2000] > top_0[2007:2000]) ? 1 : 0;
assign detect_max[249][2] = (mid_1[2007:2000] > top_0[2015:2008]) ? 1 : 0;
assign detect_max[249][3] = (mid_1[2007:2000] > top_1[1999:1992]) ? 1 : 0;
assign detect_max[249][4] = (mid_1[2007:2000] > top_1[2007:2000]) ? 1 : 0;
assign detect_max[249][5] = (mid_1[2007:2000] > top_1[2015:2008]) ? 1 : 0;
assign detect_max[249][6] = (mid_1[2007:2000] > top_2[1999:1992]) ? 1 : 0;
assign detect_max[249][7] = (mid_1[2007:2000] > top_2[2007:2000]) ? 1 : 0;
assign detect_max[249][8] = (mid_1[2007:2000] > top_2[2015:2008]) ? 1 : 0;
assign detect_max[249][9] = (mid_1[2007:2000] > mid_0[1999:1992]) ? 1 : 0;
assign detect_max[249][10] = (mid_1[2007:2000] > mid_0[2007:2000]) ? 1 : 0;
assign detect_max[249][11] = (mid_1[2007:2000] > mid_0[2015:2008]) ? 1 : 0;
assign detect_max[249][12] = (mid_1[2007:2000] > mid_1[1999:1992]) ? 1 : 0;
assign detect_max[249][13] = (mid_1[2007:2000] > mid_1[2015:2008]) ? 1 : 0;
assign detect_max[249][14] = (mid_1[2007:2000] > mid_2[1999:1992]) ? 1 : 0;
assign detect_max[249][15] = (mid_1[2007:2000] > mid_2[2007:2000]) ? 1 : 0;
assign detect_max[249][16] = (mid_1[2007:2000] > mid_2[2015:2008]) ? 1 : 0;
assign detect_max[249][17] = (mid_1[2007:2000] > btm_0[1999:1992]) ? 1 : 0;
assign detect_max[249][18] = (mid_1[2007:2000] > btm_0[2007:2000]) ? 1 : 0;
assign detect_max[249][19] = (mid_1[2007:2000] > btm_0[2015:2008]) ? 1 : 0;
assign detect_max[249][20] = (mid_1[2007:2000] > btm_1[1999:1992]) ? 1 : 0;
assign detect_max[249][21] = (mid_1[2007:2000] > btm_1[2007:2000]) ? 1 : 0;
assign detect_max[249][22] = (mid_1[2007:2000] > btm_1[2015:2008]) ? 1 : 0;
assign detect_max[249][23] = (mid_1[2007:2000] > btm_2[1999:1992]) ? 1 : 0;
assign detect_max[249][24] = (mid_1[2007:2000] > btm_2[2007:2000]) ? 1 : 0;
assign detect_max[249][25] = (mid_1[2007:2000] > btm_2[2015:2008]) ? 1 : 0;

assign detect_max[250][0] = (mid_1[2015:2008] > top_0[2007:2000]) ? 1 : 0;
assign detect_max[250][1] = (mid_1[2015:2008] > top_0[2015:2008]) ? 1 : 0;
assign detect_max[250][2] = (mid_1[2015:2008] > top_0[2023:2016]) ? 1 : 0;
assign detect_max[250][3] = (mid_1[2015:2008] > top_1[2007:2000]) ? 1 : 0;
assign detect_max[250][4] = (mid_1[2015:2008] > top_1[2015:2008]) ? 1 : 0;
assign detect_max[250][5] = (mid_1[2015:2008] > top_1[2023:2016]) ? 1 : 0;
assign detect_max[250][6] = (mid_1[2015:2008] > top_2[2007:2000]) ? 1 : 0;
assign detect_max[250][7] = (mid_1[2015:2008] > top_2[2015:2008]) ? 1 : 0;
assign detect_max[250][8] = (mid_1[2015:2008] > top_2[2023:2016]) ? 1 : 0;
assign detect_max[250][9] = (mid_1[2015:2008] > mid_0[2007:2000]) ? 1 : 0;
assign detect_max[250][10] = (mid_1[2015:2008] > mid_0[2015:2008]) ? 1 : 0;
assign detect_max[250][11] = (mid_1[2015:2008] > mid_0[2023:2016]) ? 1 : 0;
assign detect_max[250][12] = (mid_1[2015:2008] > mid_1[2007:2000]) ? 1 : 0;
assign detect_max[250][13] = (mid_1[2015:2008] > mid_1[2023:2016]) ? 1 : 0;
assign detect_max[250][14] = (mid_1[2015:2008] > mid_2[2007:2000]) ? 1 : 0;
assign detect_max[250][15] = (mid_1[2015:2008] > mid_2[2015:2008]) ? 1 : 0;
assign detect_max[250][16] = (mid_1[2015:2008] > mid_2[2023:2016]) ? 1 : 0;
assign detect_max[250][17] = (mid_1[2015:2008] > btm_0[2007:2000]) ? 1 : 0;
assign detect_max[250][18] = (mid_1[2015:2008] > btm_0[2015:2008]) ? 1 : 0;
assign detect_max[250][19] = (mid_1[2015:2008] > btm_0[2023:2016]) ? 1 : 0;
assign detect_max[250][20] = (mid_1[2015:2008] > btm_1[2007:2000]) ? 1 : 0;
assign detect_max[250][21] = (mid_1[2015:2008] > btm_1[2015:2008]) ? 1 : 0;
assign detect_max[250][22] = (mid_1[2015:2008] > btm_1[2023:2016]) ? 1 : 0;
assign detect_max[250][23] = (mid_1[2015:2008] > btm_2[2007:2000]) ? 1 : 0;
assign detect_max[250][24] = (mid_1[2015:2008] > btm_2[2015:2008]) ? 1 : 0;
assign detect_max[250][25] = (mid_1[2015:2008] > btm_2[2023:2016]) ? 1 : 0;

assign detect_max[251][0] = (mid_1[2023:2016] > top_0[2015:2008]) ? 1 : 0;
assign detect_max[251][1] = (mid_1[2023:2016] > top_0[2023:2016]) ? 1 : 0;
assign detect_max[251][2] = (mid_1[2023:2016] > top_0[2031:2024]) ? 1 : 0;
assign detect_max[251][3] = (mid_1[2023:2016] > top_1[2015:2008]) ? 1 : 0;
assign detect_max[251][4] = (mid_1[2023:2016] > top_1[2023:2016]) ? 1 : 0;
assign detect_max[251][5] = (mid_1[2023:2016] > top_1[2031:2024]) ? 1 : 0;
assign detect_max[251][6] = (mid_1[2023:2016] > top_2[2015:2008]) ? 1 : 0;
assign detect_max[251][7] = (mid_1[2023:2016] > top_2[2023:2016]) ? 1 : 0;
assign detect_max[251][8] = (mid_1[2023:2016] > top_2[2031:2024]) ? 1 : 0;
assign detect_max[251][9] = (mid_1[2023:2016] > mid_0[2015:2008]) ? 1 : 0;
assign detect_max[251][10] = (mid_1[2023:2016] > mid_0[2023:2016]) ? 1 : 0;
assign detect_max[251][11] = (mid_1[2023:2016] > mid_0[2031:2024]) ? 1 : 0;
assign detect_max[251][12] = (mid_1[2023:2016] > mid_1[2015:2008]) ? 1 : 0;
assign detect_max[251][13] = (mid_1[2023:2016] > mid_1[2031:2024]) ? 1 : 0;
assign detect_max[251][14] = (mid_1[2023:2016] > mid_2[2015:2008]) ? 1 : 0;
assign detect_max[251][15] = (mid_1[2023:2016] > mid_2[2023:2016]) ? 1 : 0;
assign detect_max[251][16] = (mid_1[2023:2016] > mid_2[2031:2024]) ? 1 : 0;
assign detect_max[251][17] = (mid_1[2023:2016] > btm_0[2015:2008]) ? 1 : 0;
assign detect_max[251][18] = (mid_1[2023:2016] > btm_0[2023:2016]) ? 1 : 0;
assign detect_max[251][19] = (mid_1[2023:2016] > btm_0[2031:2024]) ? 1 : 0;
assign detect_max[251][20] = (mid_1[2023:2016] > btm_1[2015:2008]) ? 1 : 0;
assign detect_max[251][21] = (mid_1[2023:2016] > btm_1[2023:2016]) ? 1 : 0;
assign detect_max[251][22] = (mid_1[2023:2016] > btm_1[2031:2024]) ? 1 : 0;
assign detect_max[251][23] = (mid_1[2023:2016] > btm_2[2015:2008]) ? 1 : 0;
assign detect_max[251][24] = (mid_1[2023:2016] > btm_2[2023:2016]) ? 1 : 0;
assign detect_max[251][25] = (mid_1[2023:2016] > btm_2[2031:2024]) ? 1 : 0;

assign detect_max[252][0] = (mid_1[2031:2024] > top_0[2023:2016]) ? 1 : 0;
assign detect_max[252][1] = (mid_1[2031:2024] > top_0[2031:2024]) ? 1 : 0;
assign detect_max[252][2] = (mid_1[2031:2024] > top_0[2039:2032]) ? 1 : 0;
assign detect_max[252][3] = (mid_1[2031:2024] > top_1[2023:2016]) ? 1 : 0;
assign detect_max[252][4] = (mid_1[2031:2024] > top_1[2031:2024]) ? 1 : 0;
assign detect_max[252][5] = (mid_1[2031:2024] > top_1[2039:2032]) ? 1 : 0;
assign detect_max[252][6] = (mid_1[2031:2024] > top_2[2023:2016]) ? 1 : 0;
assign detect_max[252][7] = (mid_1[2031:2024] > top_2[2031:2024]) ? 1 : 0;
assign detect_max[252][8] = (mid_1[2031:2024] > top_2[2039:2032]) ? 1 : 0;
assign detect_max[252][9] = (mid_1[2031:2024] > mid_0[2023:2016]) ? 1 : 0;
assign detect_max[252][10] = (mid_1[2031:2024] > mid_0[2031:2024]) ? 1 : 0;
assign detect_max[252][11] = (mid_1[2031:2024] > mid_0[2039:2032]) ? 1 : 0;
assign detect_max[252][12] = (mid_1[2031:2024] > mid_1[2023:2016]) ? 1 : 0;
assign detect_max[252][13] = (mid_1[2031:2024] > mid_1[2039:2032]) ? 1 : 0;
assign detect_max[252][14] = (mid_1[2031:2024] > mid_2[2023:2016]) ? 1 : 0;
assign detect_max[252][15] = (mid_1[2031:2024] > mid_2[2031:2024]) ? 1 : 0;
assign detect_max[252][16] = (mid_1[2031:2024] > mid_2[2039:2032]) ? 1 : 0;
assign detect_max[252][17] = (mid_1[2031:2024] > btm_0[2023:2016]) ? 1 : 0;
assign detect_max[252][18] = (mid_1[2031:2024] > btm_0[2031:2024]) ? 1 : 0;
assign detect_max[252][19] = (mid_1[2031:2024] > btm_0[2039:2032]) ? 1 : 0;
assign detect_max[252][20] = (mid_1[2031:2024] > btm_1[2023:2016]) ? 1 : 0;
assign detect_max[252][21] = (mid_1[2031:2024] > btm_1[2031:2024]) ? 1 : 0;
assign detect_max[252][22] = (mid_1[2031:2024] > btm_1[2039:2032]) ? 1 : 0;
assign detect_max[252][23] = (mid_1[2031:2024] > btm_2[2023:2016]) ? 1 : 0;
assign detect_max[252][24] = (mid_1[2031:2024] > btm_2[2031:2024]) ? 1 : 0;
assign detect_max[252][25] = (mid_1[2031:2024] > btm_2[2039:2032]) ? 1 : 0;

assign detect_max[253][0] = (mid_1[2039:2032] > top_0[2031:2024]) ? 1 : 0;
assign detect_max[253][1] = (mid_1[2039:2032] > top_0[2039:2032]) ? 1 : 0;
assign detect_max[253][2] = (mid_1[2039:2032] > top_0[2047:2040]) ? 1 : 0;
assign detect_max[253][3] = (mid_1[2039:2032] > top_1[2031:2024]) ? 1 : 0;
assign detect_max[253][4] = (mid_1[2039:2032] > top_1[2039:2032]) ? 1 : 0;
assign detect_max[253][5] = (mid_1[2039:2032] > top_1[2047:2040]) ? 1 : 0;
assign detect_max[253][6] = (mid_1[2039:2032] > top_2[2031:2024]) ? 1 : 0;
assign detect_max[253][7] = (mid_1[2039:2032] > top_2[2039:2032]) ? 1 : 0;
assign detect_max[253][8] = (mid_1[2039:2032] > top_2[2047:2040]) ? 1 : 0;
assign detect_max[253][9] = (mid_1[2039:2032] > mid_0[2031:2024]) ? 1 : 0;
assign detect_max[253][10] = (mid_1[2039:2032] > mid_0[2039:2032]) ? 1 : 0;
assign detect_max[253][11] = (mid_1[2039:2032] > mid_0[2047:2040]) ? 1 : 0;
assign detect_max[253][12] = (mid_1[2039:2032] > mid_1[2031:2024]) ? 1 : 0;
assign detect_max[253][13] = (mid_1[2039:2032] > mid_1[2047:2040]) ? 1 : 0;
assign detect_max[253][14] = (mid_1[2039:2032] > mid_2[2031:2024]) ? 1 : 0;
assign detect_max[253][15] = (mid_1[2039:2032] > mid_2[2039:2032]) ? 1 : 0;
assign detect_max[253][16] = (mid_1[2039:2032] > mid_2[2047:2040]) ? 1 : 0;
assign detect_max[253][17] = (mid_1[2039:2032] > btm_0[2031:2024]) ? 1 : 0;
assign detect_max[253][18] = (mid_1[2039:2032] > btm_0[2039:2032]) ? 1 : 0;
assign detect_max[253][19] = (mid_1[2039:2032] > btm_0[2047:2040]) ? 1 : 0;
assign detect_max[253][20] = (mid_1[2039:2032] > btm_1[2031:2024]) ? 1 : 0;
assign detect_max[253][21] = (mid_1[2039:2032] > btm_1[2039:2032]) ? 1 : 0;
assign detect_max[253][22] = (mid_1[2039:2032] > btm_1[2047:2040]) ? 1 : 0;
assign detect_max[253][23] = (mid_1[2039:2032] > btm_2[2031:2024]) ? 1 : 0;
assign detect_max[253][24] = (mid_1[2039:2032] > btm_2[2039:2032]) ? 1 : 0;
assign detect_max[253][25] = (mid_1[2039:2032] > btm_2[2047:2040]) ? 1 : 0;

assign detect_max[254][0] = (mid_1[2047:2040] > top_0[2039:2032]) ? 1 : 0;
assign detect_max[254][1] = (mid_1[2047:2040] > top_0[2047:2040]) ? 1 : 0;
assign detect_max[254][2] = (mid_1[2047:2040] > top_0[2055:2048]) ? 1 : 0;
assign detect_max[254][3] = (mid_1[2047:2040] > top_1[2039:2032]) ? 1 : 0;
assign detect_max[254][4] = (mid_1[2047:2040] > top_1[2047:2040]) ? 1 : 0;
assign detect_max[254][5] = (mid_1[2047:2040] > top_1[2055:2048]) ? 1 : 0;
assign detect_max[254][6] = (mid_1[2047:2040] > top_2[2039:2032]) ? 1 : 0;
assign detect_max[254][7] = (mid_1[2047:2040] > top_2[2047:2040]) ? 1 : 0;
assign detect_max[254][8] = (mid_1[2047:2040] > top_2[2055:2048]) ? 1 : 0;
assign detect_max[254][9] = (mid_1[2047:2040] > mid_0[2039:2032]) ? 1 : 0;
assign detect_max[254][10] = (mid_1[2047:2040] > mid_0[2047:2040]) ? 1 : 0;
assign detect_max[254][11] = (mid_1[2047:2040] > mid_0[2055:2048]) ? 1 : 0;
assign detect_max[254][12] = (mid_1[2047:2040] > mid_1[2039:2032]) ? 1 : 0;
assign detect_max[254][13] = (mid_1[2047:2040] > mid_1[2055:2048]) ? 1 : 0;
assign detect_max[254][14] = (mid_1[2047:2040] > mid_2[2039:2032]) ? 1 : 0;
assign detect_max[254][15] = (mid_1[2047:2040] > mid_2[2047:2040]) ? 1 : 0;
assign detect_max[254][16] = (mid_1[2047:2040] > mid_2[2055:2048]) ? 1 : 0;
assign detect_max[254][17] = (mid_1[2047:2040] > btm_0[2039:2032]) ? 1 : 0;
assign detect_max[254][18] = (mid_1[2047:2040] > btm_0[2047:2040]) ? 1 : 0;
assign detect_max[254][19] = (mid_1[2047:2040] > btm_0[2055:2048]) ? 1 : 0;
assign detect_max[254][20] = (mid_1[2047:2040] > btm_1[2039:2032]) ? 1 : 0;
assign detect_max[254][21] = (mid_1[2047:2040] > btm_1[2047:2040]) ? 1 : 0;
assign detect_max[254][22] = (mid_1[2047:2040] > btm_1[2055:2048]) ? 1 : 0;
assign detect_max[254][23] = (mid_1[2047:2040] > btm_2[2039:2032]) ? 1 : 0;
assign detect_max[254][24] = (mid_1[2047:2040] > btm_2[2047:2040]) ? 1 : 0;
assign detect_max[254][25] = (mid_1[2047:2040] > btm_2[2055:2048]) ? 1 : 0;

assign detect_max[255][0] = (mid_1[2055:2048] > top_0[2047:2040]) ? 1 : 0;
assign detect_max[255][1] = (mid_1[2055:2048] > top_0[2055:2048]) ? 1 : 0;
assign detect_max[255][2] = (mid_1[2055:2048] > top_0[2063:2056]) ? 1 : 0;
assign detect_max[255][3] = (mid_1[2055:2048] > top_1[2047:2040]) ? 1 : 0;
assign detect_max[255][4] = (mid_1[2055:2048] > top_1[2055:2048]) ? 1 : 0;
assign detect_max[255][5] = (mid_1[2055:2048] > top_1[2063:2056]) ? 1 : 0;
assign detect_max[255][6] = (mid_1[2055:2048] > top_2[2047:2040]) ? 1 : 0;
assign detect_max[255][7] = (mid_1[2055:2048] > top_2[2055:2048]) ? 1 : 0;
assign detect_max[255][8] = (mid_1[2055:2048] > top_2[2063:2056]) ? 1 : 0;
assign detect_max[255][9] = (mid_1[2055:2048] > mid_0[2047:2040]) ? 1 : 0;
assign detect_max[255][10] = (mid_1[2055:2048] > mid_0[2055:2048]) ? 1 : 0;
assign detect_max[255][11] = (mid_1[2055:2048] > mid_0[2063:2056]) ? 1 : 0;
assign detect_max[255][12] = (mid_1[2055:2048] > mid_1[2047:2040]) ? 1 : 0;
assign detect_max[255][13] = (mid_1[2055:2048] > mid_1[2063:2056]) ? 1 : 0;
assign detect_max[255][14] = (mid_1[2055:2048] > mid_2[2047:2040]) ? 1 : 0;
assign detect_max[255][15] = (mid_1[2055:2048] > mid_2[2055:2048]) ? 1 : 0;
assign detect_max[255][16] = (mid_1[2055:2048] > mid_2[2063:2056]) ? 1 : 0;
assign detect_max[255][17] = (mid_1[2055:2048] > btm_0[2047:2040]) ? 1 : 0;
assign detect_max[255][18] = (mid_1[2055:2048] > btm_0[2055:2048]) ? 1 : 0;
assign detect_max[255][19] = (mid_1[2055:2048] > btm_0[2063:2056]) ? 1 : 0;
assign detect_max[255][20] = (mid_1[2055:2048] > btm_1[2047:2040]) ? 1 : 0;
assign detect_max[255][21] = (mid_1[2055:2048] > btm_1[2055:2048]) ? 1 : 0;
assign detect_max[255][22] = (mid_1[2055:2048] > btm_1[2063:2056]) ? 1 : 0;
assign detect_max[255][23] = (mid_1[2055:2048] > btm_2[2047:2040]) ? 1 : 0;
assign detect_max[255][24] = (mid_1[2055:2048] > btm_2[2055:2048]) ? 1 : 0;
assign detect_max[255][25] = (mid_1[2055:2048] > btm_2[2063:2056]) ? 1 : 0;

assign detect_max[256][0] = (mid_1[2063:2056] > top_0[2055:2048]) ? 1 : 0;
assign detect_max[256][1] = (mid_1[2063:2056] > top_0[2063:2056]) ? 1 : 0;
assign detect_max[256][2] = (mid_1[2063:2056] > top_0[2071:2064]) ? 1 : 0;
assign detect_max[256][3] = (mid_1[2063:2056] > top_1[2055:2048]) ? 1 : 0;
assign detect_max[256][4] = (mid_1[2063:2056] > top_1[2063:2056]) ? 1 : 0;
assign detect_max[256][5] = (mid_1[2063:2056] > top_1[2071:2064]) ? 1 : 0;
assign detect_max[256][6] = (mid_1[2063:2056] > top_2[2055:2048]) ? 1 : 0;
assign detect_max[256][7] = (mid_1[2063:2056] > top_2[2063:2056]) ? 1 : 0;
assign detect_max[256][8] = (mid_1[2063:2056] > top_2[2071:2064]) ? 1 : 0;
assign detect_max[256][9] = (mid_1[2063:2056] > mid_0[2055:2048]) ? 1 : 0;
assign detect_max[256][10] = (mid_1[2063:2056] > mid_0[2063:2056]) ? 1 : 0;
assign detect_max[256][11] = (mid_1[2063:2056] > mid_0[2071:2064]) ? 1 : 0;
assign detect_max[256][12] = (mid_1[2063:2056] > mid_1[2055:2048]) ? 1 : 0;
assign detect_max[256][13] = (mid_1[2063:2056] > mid_1[2071:2064]) ? 1 : 0;
assign detect_max[256][14] = (mid_1[2063:2056] > mid_2[2055:2048]) ? 1 : 0;
assign detect_max[256][15] = (mid_1[2063:2056] > mid_2[2063:2056]) ? 1 : 0;
assign detect_max[256][16] = (mid_1[2063:2056] > mid_2[2071:2064]) ? 1 : 0;
assign detect_max[256][17] = (mid_1[2063:2056] > btm_0[2055:2048]) ? 1 : 0;
assign detect_max[256][18] = (mid_1[2063:2056] > btm_0[2063:2056]) ? 1 : 0;
assign detect_max[256][19] = (mid_1[2063:2056] > btm_0[2071:2064]) ? 1 : 0;
assign detect_max[256][20] = (mid_1[2063:2056] > btm_1[2055:2048]) ? 1 : 0;
assign detect_max[256][21] = (mid_1[2063:2056] > btm_1[2063:2056]) ? 1 : 0;
assign detect_max[256][22] = (mid_1[2063:2056] > btm_1[2071:2064]) ? 1 : 0;
assign detect_max[256][23] = (mid_1[2063:2056] > btm_2[2055:2048]) ? 1 : 0;
assign detect_max[256][24] = (mid_1[2063:2056] > btm_2[2063:2056]) ? 1 : 0;
assign detect_max[256][25] = (mid_1[2063:2056] > btm_2[2071:2064]) ? 1 : 0;

assign detect_max[257][0] = (mid_1[2071:2064] > top_0[2063:2056]) ? 1 : 0;
assign detect_max[257][1] = (mid_1[2071:2064] > top_0[2071:2064]) ? 1 : 0;
assign detect_max[257][2] = (mid_1[2071:2064] > top_0[2079:2072]) ? 1 : 0;
assign detect_max[257][3] = (mid_1[2071:2064] > top_1[2063:2056]) ? 1 : 0;
assign detect_max[257][4] = (mid_1[2071:2064] > top_1[2071:2064]) ? 1 : 0;
assign detect_max[257][5] = (mid_1[2071:2064] > top_1[2079:2072]) ? 1 : 0;
assign detect_max[257][6] = (mid_1[2071:2064] > top_2[2063:2056]) ? 1 : 0;
assign detect_max[257][7] = (mid_1[2071:2064] > top_2[2071:2064]) ? 1 : 0;
assign detect_max[257][8] = (mid_1[2071:2064] > top_2[2079:2072]) ? 1 : 0;
assign detect_max[257][9] = (mid_1[2071:2064] > mid_0[2063:2056]) ? 1 : 0;
assign detect_max[257][10] = (mid_1[2071:2064] > mid_0[2071:2064]) ? 1 : 0;
assign detect_max[257][11] = (mid_1[2071:2064] > mid_0[2079:2072]) ? 1 : 0;
assign detect_max[257][12] = (mid_1[2071:2064] > mid_1[2063:2056]) ? 1 : 0;
assign detect_max[257][13] = (mid_1[2071:2064] > mid_1[2079:2072]) ? 1 : 0;
assign detect_max[257][14] = (mid_1[2071:2064] > mid_2[2063:2056]) ? 1 : 0;
assign detect_max[257][15] = (mid_1[2071:2064] > mid_2[2071:2064]) ? 1 : 0;
assign detect_max[257][16] = (mid_1[2071:2064] > mid_2[2079:2072]) ? 1 : 0;
assign detect_max[257][17] = (mid_1[2071:2064] > btm_0[2063:2056]) ? 1 : 0;
assign detect_max[257][18] = (mid_1[2071:2064] > btm_0[2071:2064]) ? 1 : 0;
assign detect_max[257][19] = (mid_1[2071:2064] > btm_0[2079:2072]) ? 1 : 0;
assign detect_max[257][20] = (mid_1[2071:2064] > btm_1[2063:2056]) ? 1 : 0;
assign detect_max[257][21] = (mid_1[2071:2064] > btm_1[2071:2064]) ? 1 : 0;
assign detect_max[257][22] = (mid_1[2071:2064] > btm_1[2079:2072]) ? 1 : 0;
assign detect_max[257][23] = (mid_1[2071:2064] > btm_2[2063:2056]) ? 1 : 0;
assign detect_max[257][24] = (mid_1[2071:2064] > btm_2[2071:2064]) ? 1 : 0;
assign detect_max[257][25] = (mid_1[2071:2064] > btm_2[2079:2072]) ? 1 : 0;

assign detect_max[258][0] = (mid_1[2079:2072] > top_0[2071:2064]) ? 1 : 0;
assign detect_max[258][1] = (mid_1[2079:2072] > top_0[2079:2072]) ? 1 : 0;
assign detect_max[258][2] = (mid_1[2079:2072] > top_0[2087:2080]) ? 1 : 0;
assign detect_max[258][3] = (mid_1[2079:2072] > top_1[2071:2064]) ? 1 : 0;
assign detect_max[258][4] = (mid_1[2079:2072] > top_1[2079:2072]) ? 1 : 0;
assign detect_max[258][5] = (mid_1[2079:2072] > top_1[2087:2080]) ? 1 : 0;
assign detect_max[258][6] = (mid_1[2079:2072] > top_2[2071:2064]) ? 1 : 0;
assign detect_max[258][7] = (mid_1[2079:2072] > top_2[2079:2072]) ? 1 : 0;
assign detect_max[258][8] = (mid_1[2079:2072] > top_2[2087:2080]) ? 1 : 0;
assign detect_max[258][9] = (mid_1[2079:2072] > mid_0[2071:2064]) ? 1 : 0;
assign detect_max[258][10] = (mid_1[2079:2072] > mid_0[2079:2072]) ? 1 : 0;
assign detect_max[258][11] = (mid_1[2079:2072] > mid_0[2087:2080]) ? 1 : 0;
assign detect_max[258][12] = (mid_1[2079:2072] > mid_1[2071:2064]) ? 1 : 0;
assign detect_max[258][13] = (mid_1[2079:2072] > mid_1[2087:2080]) ? 1 : 0;
assign detect_max[258][14] = (mid_1[2079:2072] > mid_2[2071:2064]) ? 1 : 0;
assign detect_max[258][15] = (mid_1[2079:2072] > mid_2[2079:2072]) ? 1 : 0;
assign detect_max[258][16] = (mid_1[2079:2072] > mid_2[2087:2080]) ? 1 : 0;
assign detect_max[258][17] = (mid_1[2079:2072] > btm_0[2071:2064]) ? 1 : 0;
assign detect_max[258][18] = (mid_1[2079:2072] > btm_0[2079:2072]) ? 1 : 0;
assign detect_max[258][19] = (mid_1[2079:2072] > btm_0[2087:2080]) ? 1 : 0;
assign detect_max[258][20] = (mid_1[2079:2072] > btm_1[2071:2064]) ? 1 : 0;
assign detect_max[258][21] = (mid_1[2079:2072] > btm_1[2079:2072]) ? 1 : 0;
assign detect_max[258][22] = (mid_1[2079:2072] > btm_1[2087:2080]) ? 1 : 0;
assign detect_max[258][23] = (mid_1[2079:2072] > btm_2[2071:2064]) ? 1 : 0;
assign detect_max[258][24] = (mid_1[2079:2072] > btm_2[2079:2072]) ? 1 : 0;
assign detect_max[258][25] = (mid_1[2079:2072] > btm_2[2087:2080]) ? 1 : 0;

assign detect_max[259][0] = (mid_1[2087:2080] > top_0[2079:2072]) ? 1 : 0;
assign detect_max[259][1] = (mid_1[2087:2080] > top_0[2087:2080]) ? 1 : 0;
assign detect_max[259][2] = (mid_1[2087:2080] > top_0[2095:2088]) ? 1 : 0;
assign detect_max[259][3] = (mid_1[2087:2080] > top_1[2079:2072]) ? 1 : 0;
assign detect_max[259][4] = (mid_1[2087:2080] > top_1[2087:2080]) ? 1 : 0;
assign detect_max[259][5] = (mid_1[2087:2080] > top_1[2095:2088]) ? 1 : 0;
assign detect_max[259][6] = (mid_1[2087:2080] > top_2[2079:2072]) ? 1 : 0;
assign detect_max[259][7] = (mid_1[2087:2080] > top_2[2087:2080]) ? 1 : 0;
assign detect_max[259][8] = (mid_1[2087:2080] > top_2[2095:2088]) ? 1 : 0;
assign detect_max[259][9] = (mid_1[2087:2080] > mid_0[2079:2072]) ? 1 : 0;
assign detect_max[259][10] = (mid_1[2087:2080] > mid_0[2087:2080]) ? 1 : 0;
assign detect_max[259][11] = (mid_1[2087:2080] > mid_0[2095:2088]) ? 1 : 0;
assign detect_max[259][12] = (mid_1[2087:2080] > mid_1[2079:2072]) ? 1 : 0;
assign detect_max[259][13] = (mid_1[2087:2080] > mid_1[2095:2088]) ? 1 : 0;
assign detect_max[259][14] = (mid_1[2087:2080] > mid_2[2079:2072]) ? 1 : 0;
assign detect_max[259][15] = (mid_1[2087:2080] > mid_2[2087:2080]) ? 1 : 0;
assign detect_max[259][16] = (mid_1[2087:2080] > mid_2[2095:2088]) ? 1 : 0;
assign detect_max[259][17] = (mid_1[2087:2080] > btm_0[2079:2072]) ? 1 : 0;
assign detect_max[259][18] = (mid_1[2087:2080] > btm_0[2087:2080]) ? 1 : 0;
assign detect_max[259][19] = (mid_1[2087:2080] > btm_0[2095:2088]) ? 1 : 0;
assign detect_max[259][20] = (mid_1[2087:2080] > btm_1[2079:2072]) ? 1 : 0;
assign detect_max[259][21] = (mid_1[2087:2080] > btm_1[2087:2080]) ? 1 : 0;
assign detect_max[259][22] = (mid_1[2087:2080] > btm_1[2095:2088]) ? 1 : 0;
assign detect_max[259][23] = (mid_1[2087:2080] > btm_2[2079:2072]) ? 1 : 0;
assign detect_max[259][24] = (mid_1[2087:2080] > btm_2[2087:2080]) ? 1 : 0;
assign detect_max[259][25] = (mid_1[2087:2080] > btm_2[2095:2088]) ? 1 : 0;

assign detect_max[260][0] = (mid_1[2095:2088] > top_0[2087:2080]) ? 1 : 0;
assign detect_max[260][1] = (mid_1[2095:2088] > top_0[2095:2088]) ? 1 : 0;
assign detect_max[260][2] = (mid_1[2095:2088] > top_0[2103:2096]) ? 1 : 0;
assign detect_max[260][3] = (mid_1[2095:2088] > top_1[2087:2080]) ? 1 : 0;
assign detect_max[260][4] = (mid_1[2095:2088] > top_1[2095:2088]) ? 1 : 0;
assign detect_max[260][5] = (mid_1[2095:2088] > top_1[2103:2096]) ? 1 : 0;
assign detect_max[260][6] = (mid_1[2095:2088] > top_2[2087:2080]) ? 1 : 0;
assign detect_max[260][7] = (mid_1[2095:2088] > top_2[2095:2088]) ? 1 : 0;
assign detect_max[260][8] = (mid_1[2095:2088] > top_2[2103:2096]) ? 1 : 0;
assign detect_max[260][9] = (mid_1[2095:2088] > mid_0[2087:2080]) ? 1 : 0;
assign detect_max[260][10] = (mid_1[2095:2088] > mid_0[2095:2088]) ? 1 : 0;
assign detect_max[260][11] = (mid_1[2095:2088] > mid_0[2103:2096]) ? 1 : 0;
assign detect_max[260][12] = (mid_1[2095:2088] > mid_1[2087:2080]) ? 1 : 0;
assign detect_max[260][13] = (mid_1[2095:2088] > mid_1[2103:2096]) ? 1 : 0;
assign detect_max[260][14] = (mid_1[2095:2088] > mid_2[2087:2080]) ? 1 : 0;
assign detect_max[260][15] = (mid_1[2095:2088] > mid_2[2095:2088]) ? 1 : 0;
assign detect_max[260][16] = (mid_1[2095:2088] > mid_2[2103:2096]) ? 1 : 0;
assign detect_max[260][17] = (mid_1[2095:2088] > btm_0[2087:2080]) ? 1 : 0;
assign detect_max[260][18] = (mid_1[2095:2088] > btm_0[2095:2088]) ? 1 : 0;
assign detect_max[260][19] = (mid_1[2095:2088] > btm_0[2103:2096]) ? 1 : 0;
assign detect_max[260][20] = (mid_1[2095:2088] > btm_1[2087:2080]) ? 1 : 0;
assign detect_max[260][21] = (mid_1[2095:2088] > btm_1[2095:2088]) ? 1 : 0;
assign detect_max[260][22] = (mid_1[2095:2088] > btm_1[2103:2096]) ? 1 : 0;
assign detect_max[260][23] = (mid_1[2095:2088] > btm_2[2087:2080]) ? 1 : 0;
assign detect_max[260][24] = (mid_1[2095:2088] > btm_2[2095:2088]) ? 1 : 0;
assign detect_max[260][25] = (mid_1[2095:2088] > btm_2[2103:2096]) ? 1 : 0;

assign detect_max[261][0] = (mid_1[2103:2096] > top_0[2095:2088]) ? 1 : 0;
assign detect_max[261][1] = (mid_1[2103:2096] > top_0[2103:2096]) ? 1 : 0;
assign detect_max[261][2] = (mid_1[2103:2096] > top_0[2111:2104]) ? 1 : 0;
assign detect_max[261][3] = (mid_1[2103:2096] > top_1[2095:2088]) ? 1 : 0;
assign detect_max[261][4] = (mid_1[2103:2096] > top_1[2103:2096]) ? 1 : 0;
assign detect_max[261][5] = (mid_1[2103:2096] > top_1[2111:2104]) ? 1 : 0;
assign detect_max[261][6] = (mid_1[2103:2096] > top_2[2095:2088]) ? 1 : 0;
assign detect_max[261][7] = (mid_1[2103:2096] > top_2[2103:2096]) ? 1 : 0;
assign detect_max[261][8] = (mid_1[2103:2096] > top_2[2111:2104]) ? 1 : 0;
assign detect_max[261][9] = (mid_1[2103:2096] > mid_0[2095:2088]) ? 1 : 0;
assign detect_max[261][10] = (mid_1[2103:2096] > mid_0[2103:2096]) ? 1 : 0;
assign detect_max[261][11] = (mid_1[2103:2096] > mid_0[2111:2104]) ? 1 : 0;
assign detect_max[261][12] = (mid_1[2103:2096] > mid_1[2095:2088]) ? 1 : 0;
assign detect_max[261][13] = (mid_1[2103:2096] > mid_1[2111:2104]) ? 1 : 0;
assign detect_max[261][14] = (mid_1[2103:2096] > mid_2[2095:2088]) ? 1 : 0;
assign detect_max[261][15] = (mid_1[2103:2096] > mid_2[2103:2096]) ? 1 : 0;
assign detect_max[261][16] = (mid_1[2103:2096] > mid_2[2111:2104]) ? 1 : 0;
assign detect_max[261][17] = (mid_1[2103:2096] > btm_0[2095:2088]) ? 1 : 0;
assign detect_max[261][18] = (mid_1[2103:2096] > btm_0[2103:2096]) ? 1 : 0;
assign detect_max[261][19] = (mid_1[2103:2096] > btm_0[2111:2104]) ? 1 : 0;
assign detect_max[261][20] = (mid_1[2103:2096] > btm_1[2095:2088]) ? 1 : 0;
assign detect_max[261][21] = (mid_1[2103:2096] > btm_1[2103:2096]) ? 1 : 0;
assign detect_max[261][22] = (mid_1[2103:2096] > btm_1[2111:2104]) ? 1 : 0;
assign detect_max[261][23] = (mid_1[2103:2096] > btm_2[2095:2088]) ? 1 : 0;
assign detect_max[261][24] = (mid_1[2103:2096] > btm_2[2103:2096]) ? 1 : 0;
assign detect_max[261][25] = (mid_1[2103:2096] > btm_2[2111:2104]) ? 1 : 0;

assign detect_max[262][0] = (mid_1[2111:2104] > top_0[2103:2096]) ? 1 : 0;
assign detect_max[262][1] = (mid_1[2111:2104] > top_0[2111:2104]) ? 1 : 0;
assign detect_max[262][2] = (mid_1[2111:2104] > top_0[2119:2112]) ? 1 : 0;
assign detect_max[262][3] = (mid_1[2111:2104] > top_1[2103:2096]) ? 1 : 0;
assign detect_max[262][4] = (mid_1[2111:2104] > top_1[2111:2104]) ? 1 : 0;
assign detect_max[262][5] = (mid_1[2111:2104] > top_1[2119:2112]) ? 1 : 0;
assign detect_max[262][6] = (mid_1[2111:2104] > top_2[2103:2096]) ? 1 : 0;
assign detect_max[262][7] = (mid_1[2111:2104] > top_2[2111:2104]) ? 1 : 0;
assign detect_max[262][8] = (mid_1[2111:2104] > top_2[2119:2112]) ? 1 : 0;
assign detect_max[262][9] = (mid_1[2111:2104] > mid_0[2103:2096]) ? 1 : 0;
assign detect_max[262][10] = (mid_1[2111:2104] > mid_0[2111:2104]) ? 1 : 0;
assign detect_max[262][11] = (mid_1[2111:2104] > mid_0[2119:2112]) ? 1 : 0;
assign detect_max[262][12] = (mid_1[2111:2104] > mid_1[2103:2096]) ? 1 : 0;
assign detect_max[262][13] = (mid_1[2111:2104] > mid_1[2119:2112]) ? 1 : 0;
assign detect_max[262][14] = (mid_1[2111:2104] > mid_2[2103:2096]) ? 1 : 0;
assign detect_max[262][15] = (mid_1[2111:2104] > mid_2[2111:2104]) ? 1 : 0;
assign detect_max[262][16] = (mid_1[2111:2104] > mid_2[2119:2112]) ? 1 : 0;
assign detect_max[262][17] = (mid_1[2111:2104] > btm_0[2103:2096]) ? 1 : 0;
assign detect_max[262][18] = (mid_1[2111:2104] > btm_0[2111:2104]) ? 1 : 0;
assign detect_max[262][19] = (mid_1[2111:2104] > btm_0[2119:2112]) ? 1 : 0;
assign detect_max[262][20] = (mid_1[2111:2104] > btm_1[2103:2096]) ? 1 : 0;
assign detect_max[262][21] = (mid_1[2111:2104] > btm_1[2111:2104]) ? 1 : 0;
assign detect_max[262][22] = (mid_1[2111:2104] > btm_1[2119:2112]) ? 1 : 0;
assign detect_max[262][23] = (mid_1[2111:2104] > btm_2[2103:2096]) ? 1 : 0;
assign detect_max[262][24] = (mid_1[2111:2104] > btm_2[2111:2104]) ? 1 : 0;
assign detect_max[262][25] = (mid_1[2111:2104] > btm_2[2119:2112]) ? 1 : 0;

assign detect_max[263][0] = (mid_1[2119:2112] > top_0[2111:2104]) ? 1 : 0;
assign detect_max[263][1] = (mid_1[2119:2112] > top_0[2119:2112]) ? 1 : 0;
assign detect_max[263][2] = (mid_1[2119:2112] > top_0[2127:2120]) ? 1 : 0;
assign detect_max[263][3] = (mid_1[2119:2112] > top_1[2111:2104]) ? 1 : 0;
assign detect_max[263][4] = (mid_1[2119:2112] > top_1[2119:2112]) ? 1 : 0;
assign detect_max[263][5] = (mid_1[2119:2112] > top_1[2127:2120]) ? 1 : 0;
assign detect_max[263][6] = (mid_1[2119:2112] > top_2[2111:2104]) ? 1 : 0;
assign detect_max[263][7] = (mid_1[2119:2112] > top_2[2119:2112]) ? 1 : 0;
assign detect_max[263][8] = (mid_1[2119:2112] > top_2[2127:2120]) ? 1 : 0;
assign detect_max[263][9] = (mid_1[2119:2112] > mid_0[2111:2104]) ? 1 : 0;
assign detect_max[263][10] = (mid_1[2119:2112] > mid_0[2119:2112]) ? 1 : 0;
assign detect_max[263][11] = (mid_1[2119:2112] > mid_0[2127:2120]) ? 1 : 0;
assign detect_max[263][12] = (mid_1[2119:2112] > mid_1[2111:2104]) ? 1 : 0;
assign detect_max[263][13] = (mid_1[2119:2112] > mid_1[2127:2120]) ? 1 : 0;
assign detect_max[263][14] = (mid_1[2119:2112] > mid_2[2111:2104]) ? 1 : 0;
assign detect_max[263][15] = (mid_1[2119:2112] > mid_2[2119:2112]) ? 1 : 0;
assign detect_max[263][16] = (mid_1[2119:2112] > mid_2[2127:2120]) ? 1 : 0;
assign detect_max[263][17] = (mid_1[2119:2112] > btm_0[2111:2104]) ? 1 : 0;
assign detect_max[263][18] = (mid_1[2119:2112] > btm_0[2119:2112]) ? 1 : 0;
assign detect_max[263][19] = (mid_1[2119:2112] > btm_0[2127:2120]) ? 1 : 0;
assign detect_max[263][20] = (mid_1[2119:2112] > btm_1[2111:2104]) ? 1 : 0;
assign detect_max[263][21] = (mid_1[2119:2112] > btm_1[2119:2112]) ? 1 : 0;
assign detect_max[263][22] = (mid_1[2119:2112] > btm_1[2127:2120]) ? 1 : 0;
assign detect_max[263][23] = (mid_1[2119:2112] > btm_2[2111:2104]) ? 1 : 0;
assign detect_max[263][24] = (mid_1[2119:2112] > btm_2[2119:2112]) ? 1 : 0;
assign detect_max[263][25] = (mid_1[2119:2112] > btm_2[2127:2120]) ? 1 : 0;

assign detect_max[264][0] = (mid_1[2127:2120] > top_0[2119:2112]) ? 1 : 0;
assign detect_max[264][1] = (mid_1[2127:2120] > top_0[2127:2120]) ? 1 : 0;
assign detect_max[264][2] = (mid_1[2127:2120] > top_0[2135:2128]) ? 1 : 0;
assign detect_max[264][3] = (mid_1[2127:2120] > top_1[2119:2112]) ? 1 : 0;
assign detect_max[264][4] = (mid_1[2127:2120] > top_1[2127:2120]) ? 1 : 0;
assign detect_max[264][5] = (mid_1[2127:2120] > top_1[2135:2128]) ? 1 : 0;
assign detect_max[264][6] = (mid_1[2127:2120] > top_2[2119:2112]) ? 1 : 0;
assign detect_max[264][7] = (mid_1[2127:2120] > top_2[2127:2120]) ? 1 : 0;
assign detect_max[264][8] = (mid_1[2127:2120] > top_2[2135:2128]) ? 1 : 0;
assign detect_max[264][9] = (mid_1[2127:2120] > mid_0[2119:2112]) ? 1 : 0;
assign detect_max[264][10] = (mid_1[2127:2120] > mid_0[2127:2120]) ? 1 : 0;
assign detect_max[264][11] = (mid_1[2127:2120] > mid_0[2135:2128]) ? 1 : 0;
assign detect_max[264][12] = (mid_1[2127:2120] > mid_1[2119:2112]) ? 1 : 0;
assign detect_max[264][13] = (mid_1[2127:2120] > mid_1[2135:2128]) ? 1 : 0;
assign detect_max[264][14] = (mid_1[2127:2120] > mid_2[2119:2112]) ? 1 : 0;
assign detect_max[264][15] = (mid_1[2127:2120] > mid_2[2127:2120]) ? 1 : 0;
assign detect_max[264][16] = (mid_1[2127:2120] > mid_2[2135:2128]) ? 1 : 0;
assign detect_max[264][17] = (mid_1[2127:2120] > btm_0[2119:2112]) ? 1 : 0;
assign detect_max[264][18] = (mid_1[2127:2120] > btm_0[2127:2120]) ? 1 : 0;
assign detect_max[264][19] = (mid_1[2127:2120] > btm_0[2135:2128]) ? 1 : 0;
assign detect_max[264][20] = (mid_1[2127:2120] > btm_1[2119:2112]) ? 1 : 0;
assign detect_max[264][21] = (mid_1[2127:2120] > btm_1[2127:2120]) ? 1 : 0;
assign detect_max[264][22] = (mid_1[2127:2120] > btm_1[2135:2128]) ? 1 : 0;
assign detect_max[264][23] = (mid_1[2127:2120] > btm_2[2119:2112]) ? 1 : 0;
assign detect_max[264][24] = (mid_1[2127:2120] > btm_2[2127:2120]) ? 1 : 0;
assign detect_max[264][25] = (mid_1[2127:2120] > btm_2[2135:2128]) ? 1 : 0;

assign detect_max[265][0] = (mid_1[2135:2128] > top_0[2127:2120]) ? 1 : 0;
assign detect_max[265][1] = (mid_1[2135:2128] > top_0[2135:2128]) ? 1 : 0;
assign detect_max[265][2] = (mid_1[2135:2128] > top_0[2143:2136]) ? 1 : 0;
assign detect_max[265][3] = (mid_1[2135:2128] > top_1[2127:2120]) ? 1 : 0;
assign detect_max[265][4] = (mid_1[2135:2128] > top_1[2135:2128]) ? 1 : 0;
assign detect_max[265][5] = (mid_1[2135:2128] > top_1[2143:2136]) ? 1 : 0;
assign detect_max[265][6] = (mid_1[2135:2128] > top_2[2127:2120]) ? 1 : 0;
assign detect_max[265][7] = (mid_1[2135:2128] > top_2[2135:2128]) ? 1 : 0;
assign detect_max[265][8] = (mid_1[2135:2128] > top_2[2143:2136]) ? 1 : 0;
assign detect_max[265][9] = (mid_1[2135:2128] > mid_0[2127:2120]) ? 1 : 0;
assign detect_max[265][10] = (mid_1[2135:2128] > mid_0[2135:2128]) ? 1 : 0;
assign detect_max[265][11] = (mid_1[2135:2128] > mid_0[2143:2136]) ? 1 : 0;
assign detect_max[265][12] = (mid_1[2135:2128] > mid_1[2127:2120]) ? 1 : 0;
assign detect_max[265][13] = (mid_1[2135:2128] > mid_1[2143:2136]) ? 1 : 0;
assign detect_max[265][14] = (mid_1[2135:2128] > mid_2[2127:2120]) ? 1 : 0;
assign detect_max[265][15] = (mid_1[2135:2128] > mid_2[2135:2128]) ? 1 : 0;
assign detect_max[265][16] = (mid_1[2135:2128] > mid_2[2143:2136]) ? 1 : 0;
assign detect_max[265][17] = (mid_1[2135:2128] > btm_0[2127:2120]) ? 1 : 0;
assign detect_max[265][18] = (mid_1[2135:2128] > btm_0[2135:2128]) ? 1 : 0;
assign detect_max[265][19] = (mid_1[2135:2128] > btm_0[2143:2136]) ? 1 : 0;
assign detect_max[265][20] = (mid_1[2135:2128] > btm_1[2127:2120]) ? 1 : 0;
assign detect_max[265][21] = (mid_1[2135:2128] > btm_1[2135:2128]) ? 1 : 0;
assign detect_max[265][22] = (mid_1[2135:2128] > btm_1[2143:2136]) ? 1 : 0;
assign detect_max[265][23] = (mid_1[2135:2128] > btm_2[2127:2120]) ? 1 : 0;
assign detect_max[265][24] = (mid_1[2135:2128] > btm_2[2135:2128]) ? 1 : 0;
assign detect_max[265][25] = (mid_1[2135:2128] > btm_2[2143:2136]) ? 1 : 0;

assign detect_max[266][0] = (mid_1[2143:2136] > top_0[2135:2128]) ? 1 : 0;
assign detect_max[266][1] = (mid_1[2143:2136] > top_0[2143:2136]) ? 1 : 0;
assign detect_max[266][2] = (mid_1[2143:2136] > top_0[2151:2144]) ? 1 : 0;
assign detect_max[266][3] = (mid_1[2143:2136] > top_1[2135:2128]) ? 1 : 0;
assign detect_max[266][4] = (mid_1[2143:2136] > top_1[2143:2136]) ? 1 : 0;
assign detect_max[266][5] = (mid_1[2143:2136] > top_1[2151:2144]) ? 1 : 0;
assign detect_max[266][6] = (mid_1[2143:2136] > top_2[2135:2128]) ? 1 : 0;
assign detect_max[266][7] = (mid_1[2143:2136] > top_2[2143:2136]) ? 1 : 0;
assign detect_max[266][8] = (mid_1[2143:2136] > top_2[2151:2144]) ? 1 : 0;
assign detect_max[266][9] = (mid_1[2143:2136] > mid_0[2135:2128]) ? 1 : 0;
assign detect_max[266][10] = (mid_1[2143:2136] > mid_0[2143:2136]) ? 1 : 0;
assign detect_max[266][11] = (mid_1[2143:2136] > mid_0[2151:2144]) ? 1 : 0;
assign detect_max[266][12] = (mid_1[2143:2136] > mid_1[2135:2128]) ? 1 : 0;
assign detect_max[266][13] = (mid_1[2143:2136] > mid_1[2151:2144]) ? 1 : 0;
assign detect_max[266][14] = (mid_1[2143:2136] > mid_2[2135:2128]) ? 1 : 0;
assign detect_max[266][15] = (mid_1[2143:2136] > mid_2[2143:2136]) ? 1 : 0;
assign detect_max[266][16] = (mid_1[2143:2136] > mid_2[2151:2144]) ? 1 : 0;
assign detect_max[266][17] = (mid_1[2143:2136] > btm_0[2135:2128]) ? 1 : 0;
assign detect_max[266][18] = (mid_1[2143:2136] > btm_0[2143:2136]) ? 1 : 0;
assign detect_max[266][19] = (mid_1[2143:2136] > btm_0[2151:2144]) ? 1 : 0;
assign detect_max[266][20] = (mid_1[2143:2136] > btm_1[2135:2128]) ? 1 : 0;
assign detect_max[266][21] = (mid_1[2143:2136] > btm_1[2143:2136]) ? 1 : 0;
assign detect_max[266][22] = (mid_1[2143:2136] > btm_1[2151:2144]) ? 1 : 0;
assign detect_max[266][23] = (mid_1[2143:2136] > btm_2[2135:2128]) ? 1 : 0;
assign detect_max[266][24] = (mid_1[2143:2136] > btm_2[2143:2136]) ? 1 : 0;
assign detect_max[266][25] = (mid_1[2143:2136] > btm_2[2151:2144]) ? 1 : 0;

assign detect_max[267][0] = (mid_1[2151:2144] > top_0[2143:2136]) ? 1 : 0;
assign detect_max[267][1] = (mid_1[2151:2144] > top_0[2151:2144]) ? 1 : 0;
assign detect_max[267][2] = (mid_1[2151:2144] > top_0[2159:2152]) ? 1 : 0;
assign detect_max[267][3] = (mid_1[2151:2144] > top_1[2143:2136]) ? 1 : 0;
assign detect_max[267][4] = (mid_1[2151:2144] > top_1[2151:2144]) ? 1 : 0;
assign detect_max[267][5] = (mid_1[2151:2144] > top_1[2159:2152]) ? 1 : 0;
assign detect_max[267][6] = (mid_1[2151:2144] > top_2[2143:2136]) ? 1 : 0;
assign detect_max[267][7] = (mid_1[2151:2144] > top_2[2151:2144]) ? 1 : 0;
assign detect_max[267][8] = (mid_1[2151:2144] > top_2[2159:2152]) ? 1 : 0;
assign detect_max[267][9] = (mid_1[2151:2144] > mid_0[2143:2136]) ? 1 : 0;
assign detect_max[267][10] = (mid_1[2151:2144] > mid_0[2151:2144]) ? 1 : 0;
assign detect_max[267][11] = (mid_1[2151:2144] > mid_0[2159:2152]) ? 1 : 0;
assign detect_max[267][12] = (mid_1[2151:2144] > mid_1[2143:2136]) ? 1 : 0;
assign detect_max[267][13] = (mid_1[2151:2144] > mid_1[2159:2152]) ? 1 : 0;
assign detect_max[267][14] = (mid_1[2151:2144] > mid_2[2143:2136]) ? 1 : 0;
assign detect_max[267][15] = (mid_1[2151:2144] > mid_2[2151:2144]) ? 1 : 0;
assign detect_max[267][16] = (mid_1[2151:2144] > mid_2[2159:2152]) ? 1 : 0;
assign detect_max[267][17] = (mid_1[2151:2144] > btm_0[2143:2136]) ? 1 : 0;
assign detect_max[267][18] = (mid_1[2151:2144] > btm_0[2151:2144]) ? 1 : 0;
assign detect_max[267][19] = (mid_1[2151:2144] > btm_0[2159:2152]) ? 1 : 0;
assign detect_max[267][20] = (mid_1[2151:2144] > btm_1[2143:2136]) ? 1 : 0;
assign detect_max[267][21] = (mid_1[2151:2144] > btm_1[2151:2144]) ? 1 : 0;
assign detect_max[267][22] = (mid_1[2151:2144] > btm_1[2159:2152]) ? 1 : 0;
assign detect_max[267][23] = (mid_1[2151:2144] > btm_2[2143:2136]) ? 1 : 0;
assign detect_max[267][24] = (mid_1[2151:2144] > btm_2[2151:2144]) ? 1 : 0;
assign detect_max[267][25] = (mid_1[2151:2144] > btm_2[2159:2152]) ? 1 : 0;

assign detect_max[268][0] = (mid_1[2159:2152] > top_0[2151:2144]) ? 1 : 0;
assign detect_max[268][1] = (mid_1[2159:2152] > top_0[2159:2152]) ? 1 : 0;
assign detect_max[268][2] = (mid_1[2159:2152] > top_0[2167:2160]) ? 1 : 0;
assign detect_max[268][3] = (mid_1[2159:2152] > top_1[2151:2144]) ? 1 : 0;
assign detect_max[268][4] = (mid_1[2159:2152] > top_1[2159:2152]) ? 1 : 0;
assign detect_max[268][5] = (mid_1[2159:2152] > top_1[2167:2160]) ? 1 : 0;
assign detect_max[268][6] = (mid_1[2159:2152] > top_2[2151:2144]) ? 1 : 0;
assign detect_max[268][7] = (mid_1[2159:2152] > top_2[2159:2152]) ? 1 : 0;
assign detect_max[268][8] = (mid_1[2159:2152] > top_2[2167:2160]) ? 1 : 0;
assign detect_max[268][9] = (mid_1[2159:2152] > mid_0[2151:2144]) ? 1 : 0;
assign detect_max[268][10] = (mid_1[2159:2152] > mid_0[2159:2152]) ? 1 : 0;
assign detect_max[268][11] = (mid_1[2159:2152] > mid_0[2167:2160]) ? 1 : 0;
assign detect_max[268][12] = (mid_1[2159:2152] > mid_1[2151:2144]) ? 1 : 0;
assign detect_max[268][13] = (mid_1[2159:2152] > mid_1[2167:2160]) ? 1 : 0;
assign detect_max[268][14] = (mid_1[2159:2152] > mid_2[2151:2144]) ? 1 : 0;
assign detect_max[268][15] = (mid_1[2159:2152] > mid_2[2159:2152]) ? 1 : 0;
assign detect_max[268][16] = (mid_1[2159:2152] > mid_2[2167:2160]) ? 1 : 0;
assign detect_max[268][17] = (mid_1[2159:2152] > btm_0[2151:2144]) ? 1 : 0;
assign detect_max[268][18] = (mid_1[2159:2152] > btm_0[2159:2152]) ? 1 : 0;
assign detect_max[268][19] = (mid_1[2159:2152] > btm_0[2167:2160]) ? 1 : 0;
assign detect_max[268][20] = (mid_1[2159:2152] > btm_1[2151:2144]) ? 1 : 0;
assign detect_max[268][21] = (mid_1[2159:2152] > btm_1[2159:2152]) ? 1 : 0;
assign detect_max[268][22] = (mid_1[2159:2152] > btm_1[2167:2160]) ? 1 : 0;
assign detect_max[268][23] = (mid_1[2159:2152] > btm_2[2151:2144]) ? 1 : 0;
assign detect_max[268][24] = (mid_1[2159:2152] > btm_2[2159:2152]) ? 1 : 0;
assign detect_max[268][25] = (mid_1[2159:2152] > btm_2[2167:2160]) ? 1 : 0;

assign detect_max[269][0] = (mid_1[2167:2160] > top_0[2159:2152]) ? 1 : 0;
assign detect_max[269][1] = (mid_1[2167:2160] > top_0[2167:2160]) ? 1 : 0;
assign detect_max[269][2] = (mid_1[2167:2160] > top_0[2175:2168]) ? 1 : 0;
assign detect_max[269][3] = (mid_1[2167:2160] > top_1[2159:2152]) ? 1 : 0;
assign detect_max[269][4] = (mid_1[2167:2160] > top_1[2167:2160]) ? 1 : 0;
assign detect_max[269][5] = (mid_1[2167:2160] > top_1[2175:2168]) ? 1 : 0;
assign detect_max[269][6] = (mid_1[2167:2160] > top_2[2159:2152]) ? 1 : 0;
assign detect_max[269][7] = (mid_1[2167:2160] > top_2[2167:2160]) ? 1 : 0;
assign detect_max[269][8] = (mid_1[2167:2160] > top_2[2175:2168]) ? 1 : 0;
assign detect_max[269][9] = (mid_1[2167:2160] > mid_0[2159:2152]) ? 1 : 0;
assign detect_max[269][10] = (mid_1[2167:2160] > mid_0[2167:2160]) ? 1 : 0;
assign detect_max[269][11] = (mid_1[2167:2160] > mid_0[2175:2168]) ? 1 : 0;
assign detect_max[269][12] = (mid_1[2167:2160] > mid_1[2159:2152]) ? 1 : 0;
assign detect_max[269][13] = (mid_1[2167:2160] > mid_1[2175:2168]) ? 1 : 0;
assign detect_max[269][14] = (mid_1[2167:2160] > mid_2[2159:2152]) ? 1 : 0;
assign detect_max[269][15] = (mid_1[2167:2160] > mid_2[2167:2160]) ? 1 : 0;
assign detect_max[269][16] = (mid_1[2167:2160] > mid_2[2175:2168]) ? 1 : 0;
assign detect_max[269][17] = (mid_1[2167:2160] > btm_0[2159:2152]) ? 1 : 0;
assign detect_max[269][18] = (mid_1[2167:2160] > btm_0[2167:2160]) ? 1 : 0;
assign detect_max[269][19] = (mid_1[2167:2160] > btm_0[2175:2168]) ? 1 : 0;
assign detect_max[269][20] = (mid_1[2167:2160] > btm_1[2159:2152]) ? 1 : 0;
assign detect_max[269][21] = (mid_1[2167:2160] > btm_1[2167:2160]) ? 1 : 0;
assign detect_max[269][22] = (mid_1[2167:2160] > btm_1[2175:2168]) ? 1 : 0;
assign detect_max[269][23] = (mid_1[2167:2160] > btm_2[2159:2152]) ? 1 : 0;
assign detect_max[269][24] = (mid_1[2167:2160] > btm_2[2167:2160]) ? 1 : 0;
assign detect_max[269][25] = (mid_1[2167:2160] > btm_2[2175:2168]) ? 1 : 0;

assign detect_max[270][0] = (mid_1[2175:2168] > top_0[2167:2160]) ? 1 : 0;
assign detect_max[270][1] = (mid_1[2175:2168] > top_0[2175:2168]) ? 1 : 0;
assign detect_max[270][2] = (mid_1[2175:2168] > top_0[2183:2176]) ? 1 : 0;
assign detect_max[270][3] = (mid_1[2175:2168] > top_1[2167:2160]) ? 1 : 0;
assign detect_max[270][4] = (mid_1[2175:2168] > top_1[2175:2168]) ? 1 : 0;
assign detect_max[270][5] = (mid_1[2175:2168] > top_1[2183:2176]) ? 1 : 0;
assign detect_max[270][6] = (mid_1[2175:2168] > top_2[2167:2160]) ? 1 : 0;
assign detect_max[270][7] = (mid_1[2175:2168] > top_2[2175:2168]) ? 1 : 0;
assign detect_max[270][8] = (mid_1[2175:2168] > top_2[2183:2176]) ? 1 : 0;
assign detect_max[270][9] = (mid_1[2175:2168] > mid_0[2167:2160]) ? 1 : 0;
assign detect_max[270][10] = (mid_1[2175:2168] > mid_0[2175:2168]) ? 1 : 0;
assign detect_max[270][11] = (mid_1[2175:2168] > mid_0[2183:2176]) ? 1 : 0;
assign detect_max[270][12] = (mid_1[2175:2168] > mid_1[2167:2160]) ? 1 : 0;
assign detect_max[270][13] = (mid_1[2175:2168] > mid_1[2183:2176]) ? 1 : 0;
assign detect_max[270][14] = (mid_1[2175:2168] > mid_2[2167:2160]) ? 1 : 0;
assign detect_max[270][15] = (mid_1[2175:2168] > mid_2[2175:2168]) ? 1 : 0;
assign detect_max[270][16] = (mid_1[2175:2168] > mid_2[2183:2176]) ? 1 : 0;
assign detect_max[270][17] = (mid_1[2175:2168] > btm_0[2167:2160]) ? 1 : 0;
assign detect_max[270][18] = (mid_1[2175:2168] > btm_0[2175:2168]) ? 1 : 0;
assign detect_max[270][19] = (mid_1[2175:2168] > btm_0[2183:2176]) ? 1 : 0;
assign detect_max[270][20] = (mid_1[2175:2168] > btm_1[2167:2160]) ? 1 : 0;
assign detect_max[270][21] = (mid_1[2175:2168] > btm_1[2175:2168]) ? 1 : 0;
assign detect_max[270][22] = (mid_1[2175:2168] > btm_1[2183:2176]) ? 1 : 0;
assign detect_max[270][23] = (mid_1[2175:2168] > btm_2[2167:2160]) ? 1 : 0;
assign detect_max[270][24] = (mid_1[2175:2168] > btm_2[2175:2168]) ? 1 : 0;
assign detect_max[270][25] = (mid_1[2175:2168] > btm_2[2183:2176]) ? 1 : 0;

assign detect_max[271][0] = (mid_1[2183:2176] > top_0[2175:2168]) ? 1 : 0;
assign detect_max[271][1] = (mid_1[2183:2176] > top_0[2183:2176]) ? 1 : 0;
assign detect_max[271][2] = (mid_1[2183:2176] > top_0[2191:2184]) ? 1 : 0;
assign detect_max[271][3] = (mid_1[2183:2176] > top_1[2175:2168]) ? 1 : 0;
assign detect_max[271][4] = (mid_1[2183:2176] > top_1[2183:2176]) ? 1 : 0;
assign detect_max[271][5] = (mid_1[2183:2176] > top_1[2191:2184]) ? 1 : 0;
assign detect_max[271][6] = (mid_1[2183:2176] > top_2[2175:2168]) ? 1 : 0;
assign detect_max[271][7] = (mid_1[2183:2176] > top_2[2183:2176]) ? 1 : 0;
assign detect_max[271][8] = (mid_1[2183:2176] > top_2[2191:2184]) ? 1 : 0;
assign detect_max[271][9] = (mid_1[2183:2176] > mid_0[2175:2168]) ? 1 : 0;
assign detect_max[271][10] = (mid_1[2183:2176] > mid_0[2183:2176]) ? 1 : 0;
assign detect_max[271][11] = (mid_1[2183:2176] > mid_0[2191:2184]) ? 1 : 0;
assign detect_max[271][12] = (mid_1[2183:2176] > mid_1[2175:2168]) ? 1 : 0;
assign detect_max[271][13] = (mid_1[2183:2176] > mid_1[2191:2184]) ? 1 : 0;
assign detect_max[271][14] = (mid_1[2183:2176] > mid_2[2175:2168]) ? 1 : 0;
assign detect_max[271][15] = (mid_1[2183:2176] > mid_2[2183:2176]) ? 1 : 0;
assign detect_max[271][16] = (mid_1[2183:2176] > mid_2[2191:2184]) ? 1 : 0;
assign detect_max[271][17] = (mid_1[2183:2176] > btm_0[2175:2168]) ? 1 : 0;
assign detect_max[271][18] = (mid_1[2183:2176] > btm_0[2183:2176]) ? 1 : 0;
assign detect_max[271][19] = (mid_1[2183:2176] > btm_0[2191:2184]) ? 1 : 0;
assign detect_max[271][20] = (mid_1[2183:2176] > btm_1[2175:2168]) ? 1 : 0;
assign detect_max[271][21] = (mid_1[2183:2176] > btm_1[2183:2176]) ? 1 : 0;
assign detect_max[271][22] = (mid_1[2183:2176] > btm_1[2191:2184]) ? 1 : 0;
assign detect_max[271][23] = (mid_1[2183:2176] > btm_2[2175:2168]) ? 1 : 0;
assign detect_max[271][24] = (mid_1[2183:2176] > btm_2[2183:2176]) ? 1 : 0;
assign detect_max[271][25] = (mid_1[2183:2176] > btm_2[2191:2184]) ? 1 : 0;

assign detect_max[272][0] = (mid_1[2191:2184] > top_0[2183:2176]) ? 1 : 0;
assign detect_max[272][1] = (mid_1[2191:2184] > top_0[2191:2184]) ? 1 : 0;
assign detect_max[272][2] = (mid_1[2191:2184] > top_0[2199:2192]) ? 1 : 0;
assign detect_max[272][3] = (mid_1[2191:2184] > top_1[2183:2176]) ? 1 : 0;
assign detect_max[272][4] = (mid_1[2191:2184] > top_1[2191:2184]) ? 1 : 0;
assign detect_max[272][5] = (mid_1[2191:2184] > top_1[2199:2192]) ? 1 : 0;
assign detect_max[272][6] = (mid_1[2191:2184] > top_2[2183:2176]) ? 1 : 0;
assign detect_max[272][7] = (mid_1[2191:2184] > top_2[2191:2184]) ? 1 : 0;
assign detect_max[272][8] = (mid_1[2191:2184] > top_2[2199:2192]) ? 1 : 0;
assign detect_max[272][9] = (mid_1[2191:2184] > mid_0[2183:2176]) ? 1 : 0;
assign detect_max[272][10] = (mid_1[2191:2184] > mid_0[2191:2184]) ? 1 : 0;
assign detect_max[272][11] = (mid_1[2191:2184] > mid_0[2199:2192]) ? 1 : 0;
assign detect_max[272][12] = (mid_1[2191:2184] > mid_1[2183:2176]) ? 1 : 0;
assign detect_max[272][13] = (mid_1[2191:2184] > mid_1[2199:2192]) ? 1 : 0;
assign detect_max[272][14] = (mid_1[2191:2184] > mid_2[2183:2176]) ? 1 : 0;
assign detect_max[272][15] = (mid_1[2191:2184] > mid_2[2191:2184]) ? 1 : 0;
assign detect_max[272][16] = (mid_1[2191:2184] > mid_2[2199:2192]) ? 1 : 0;
assign detect_max[272][17] = (mid_1[2191:2184] > btm_0[2183:2176]) ? 1 : 0;
assign detect_max[272][18] = (mid_1[2191:2184] > btm_0[2191:2184]) ? 1 : 0;
assign detect_max[272][19] = (mid_1[2191:2184] > btm_0[2199:2192]) ? 1 : 0;
assign detect_max[272][20] = (mid_1[2191:2184] > btm_1[2183:2176]) ? 1 : 0;
assign detect_max[272][21] = (mid_1[2191:2184] > btm_1[2191:2184]) ? 1 : 0;
assign detect_max[272][22] = (mid_1[2191:2184] > btm_1[2199:2192]) ? 1 : 0;
assign detect_max[272][23] = (mid_1[2191:2184] > btm_2[2183:2176]) ? 1 : 0;
assign detect_max[272][24] = (mid_1[2191:2184] > btm_2[2191:2184]) ? 1 : 0;
assign detect_max[272][25] = (mid_1[2191:2184] > btm_2[2199:2192]) ? 1 : 0;

assign detect_max[273][0] = (mid_1[2199:2192] > top_0[2191:2184]) ? 1 : 0;
assign detect_max[273][1] = (mid_1[2199:2192] > top_0[2199:2192]) ? 1 : 0;
assign detect_max[273][2] = (mid_1[2199:2192] > top_0[2207:2200]) ? 1 : 0;
assign detect_max[273][3] = (mid_1[2199:2192] > top_1[2191:2184]) ? 1 : 0;
assign detect_max[273][4] = (mid_1[2199:2192] > top_1[2199:2192]) ? 1 : 0;
assign detect_max[273][5] = (mid_1[2199:2192] > top_1[2207:2200]) ? 1 : 0;
assign detect_max[273][6] = (mid_1[2199:2192] > top_2[2191:2184]) ? 1 : 0;
assign detect_max[273][7] = (mid_1[2199:2192] > top_2[2199:2192]) ? 1 : 0;
assign detect_max[273][8] = (mid_1[2199:2192] > top_2[2207:2200]) ? 1 : 0;
assign detect_max[273][9] = (mid_1[2199:2192] > mid_0[2191:2184]) ? 1 : 0;
assign detect_max[273][10] = (mid_1[2199:2192] > mid_0[2199:2192]) ? 1 : 0;
assign detect_max[273][11] = (mid_1[2199:2192] > mid_0[2207:2200]) ? 1 : 0;
assign detect_max[273][12] = (mid_1[2199:2192] > mid_1[2191:2184]) ? 1 : 0;
assign detect_max[273][13] = (mid_1[2199:2192] > mid_1[2207:2200]) ? 1 : 0;
assign detect_max[273][14] = (mid_1[2199:2192] > mid_2[2191:2184]) ? 1 : 0;
assign detect_max[273][15] = (mid_1[2199:2192] > mid_2[2199:2192]) ? 1 : 0;
assign detect_max[273][16] = (mid_1[2199:2192] > mid_2[2207:2200]) ? 1 : 0;
assign detect_max[273][17] = (mid_1[2199:2192] > btm_0[2191:2184]) ? 1 : 0;
assign detect_max[273][18] = (mid_1[2199:2192] > btm_0[2199:2192]) ? 1 : 0;
assign detect_max[273][19] = (mid_1[2199:2192] > btm_0[2207:2200]) ? 1 : 0;
assign detect_max[273][20] = (mid_1[2199:2192] > btm_1[2191:2184]) ? 1 : 0;
assign detect_max[273][21] = (mid_1[2199:2192] > btm_1[2199:2192]) ? 1 : 0;
assign detect_max[273][22] = (mid_1[2199:2192] > btm_1[2207:2200]) ? 1 : 0;
assign detect_max[273][23] = (mid_1[2199:2192] > btm_2[2191:2184]) ? 1 : 0;
assign detect_max[273][24] = (mid_1[2199:2192] > btm_2[2199:2192]) ? 1 : 0;
assign detect_max[273][25] = (mid_1[2199:2192] > btm_2[2207:2200]) ? 1 : 0;

assign detect_max[274][0] = (mid_1[2207:2200] > top_0[2199:2192]) ? 1 : 0;
assign detect_max[274][1] = (mid_1[2207:2200] > top_0[2207:2200]) ? 1 : 0;
assign detect_max[274][2] = (mid_1[2207:2200] > top_0[2215:2208]) ? 1 : 0;
assign detect_max[274][3] = (mid_1[2207:2200] > top_1[2199:2192]) ? 1 : 0;
assign detect_max[274][4] = (mid_1[2207:2200] > top_1[2207:2200]) ? 1 : 0;
assign detect_max[274][5] = (mid_1[2207:2200] > top_1[2215:2208]) ? 1 : 0;
assign detect_max[274][6] = (mid_1[2207:2200] > top_2[2199:2192]) ? 1 : 0;
assign detect_max[274][7] = (mid_1[2207:2200] > top_2[2207:2200]) ? 1 : 0;
assign detect_max[274][8] = (mid_1[2207:2200] > top_2[2215:2208]) ? 1 : 0;
assign detect_max[274][9] = (mid_1[2207:2200] > mid_0[2199:2192]) ? 1 : 0;
assign detect_max[274][10] = (mid_1[2207:2200] > mid_0[2207:2200]) ? 1 : 0;
assign detect_max[274][11] = (mid_1[2207:2200] > mid_0[2215:2208]) ? 1 : 0;
assign detect_max[274][12] = (mid_1[2207:2200] > mid_1[2199:2192]) ? 1 : 0;
assign detect_max[274][13] = (mid_1[2207:2200] > mid_1[2215:2208]) ? 1 : 0;
assign detect_max[274][14] = (mid_1[2207:2200] > mid_2[2199:2192]) ? 1 : 0;
assign detect_max[274][15] = (mid_1[2207:2200] > mid_2[2207:2200]) ? 1 : 0;
assign detect_max[274][16] = (mid_1[2207:2200] > mid_2[2215:2208]) ? 1 : 0;
assign detect_max[274][17] = (mid_1[2207:2200] > btm_0[2199:2192]) ? 1 : 0;
assign detect_max[274][18] = (mid_1[2207:2200] > btm_0[2207:2200]) ? 1 : 0;
assign detect_max[274][19] = (mid_1[2207:2200] > btm_0[2215:2208]) ? 1 : 0;
assign detect_max[274][20] = (mid_1[2207:2200] > btm_1[2199:2192]) ? 1 : 0;
assign detect_max[274][21] = (mid_1[2207:2200] > btm_1[2207:2200]) ? 1 : 0;
assign detect_max[274][22] = (mid_1[2207:2200] > btm_1[2215:2208]) ? 1 : 0;
assign detect_max[274][23] = (mid_1[2207:2200] > btm_2[2199:2192]) ? 1 : 0;
assign detect_max[274][24] = (mid_1[2207:2200] > btm_2[2207:2200]) ? 1 : 0;
assign detect_max[274][25] = (mid_1[2207:2200] > btm_2[2215:2208]) ? 1 : 0;

assign detect_max[275][0] = (mid_1[2215:2208] > top_0[2207:2200]) ? 1 : 0;
assign detect_max[275][1] = (mid_1[2215:2208] > top_0[2215:2208]) ? 1 : 0;
assign detect_max[275][2] = (mid_1[2215:2208] > top_0[2223:2216]) ? 1 : 0;
assign detect_max[275][3] = (mid_1[2215:2208] > top_1[2207:2200]) ? 1 : 0;
assign detect_max[275][4] = (mid_1[2215:2208] > top_1[2215:2208]) ? 1 : 0;
assign detect_max[275][5] = (mid_1[2215:2208] > top_1[2223:2216]) ? 1 : 0;
assign detect_max[275][6] = (mid_1[2215:2208] > top_2[2207:2200]) ? 1 : 0;
assign detect_max[275][7] = (mid_1[2215:2208] > top_2[2215:2208]) ? 1 : 0;
assign detect_max[275][8] = (mid_1[2215:2208] > top_2[2223:2216]) ? 1 : 0;
assign detect_max[275][9] = (mid_1[2215:2208] > mid_0[2207:2200]) ? 1 : 0;
assign detect_max[275][10] = (mid_1[2215:2208] > mid_0[2215:2208]) ? 1 : 0;
assign detect_max[275][11] = (mid_1[2215:2208] > mid_0[2223:2216]) ? 1 : 0;
assign detect_max[275][12] = (mid_1[2215:2208] > mid_1[2207:2200]) ? 1 : 0;
assign detect_max[275][13] = (mid_1[2215:2208] > mid_1[2223:2216]) ? 1 : 0;
assign detect_max[275][14] = (mid_1[2215:2208] > mid_2[2207:2200]) ? 1 : 0;
assign detect_max[275][15] = (mid_1[2215:2208] > mid_2[2215:2208]) ? 1 : 0;
assign detect_max[275][16] = (mid_1[2215:2208] > mid_2[2223:2216]) ? 1 : 0;
assign detect_max[275][17] = (mid_1[2215:2208] > btm_0[2207:2200]) ? 1 : 0;
assign detect_max[275][18] = (mid_1[2215:2208] > btm_0[2215:2208]) ? 1 : 0;
assign detect_max[275][19] = (mid_1[2215:2208] > btm_0[2223:2216]) ? 1 : 0;
assign detect_max[275][20] = (mid_1[2215:2208] > btm_1[2207:2200]) ? 1 : 0;
assign detect_max[275][21] = (mid_1[2215:2208] > btm_1[2215:2208]) ? 1 : 0;
assign detect_max[275][22] = (mid_1[2215:2208] > btm_1[2223:2216]) ? 1 : 0;
assign detect_max[275][23] = (mid_1[2215:2208] > btm_2[2207:2200]) ? 1 : 0;
assign detect_max[275][24] = (mid_1[2215:2208] > btm_2[2215:2208]) ? 1 : 0;
assign detect_max[275][25] = (mid_1[2215:2208] > btm_2[2223:2216]) ? 1 : 0;

assign detect_max[276][0] = (mid_1[2223:2216] > top_0[2215:2208]) ? 1 : 0;
assign detect_max[276][1] = (mid_1[2223:2216] > top_0[2223:2216]) ? 1 : 0;
assign detect_max[276][2] = (mid_1[2223:2216] > top_0[2231:2224]) ? 1 : 0;
assign detect_max[276][3] = (mid_1[2223:2216] > top_1[2215:2208]) ? 1 : 0;
assign detect_max[276][4] = (mid_1[2223:2216] > top_1[2223:2216]) ? 1 : 0;
assign detect_max[276][5] = (mid_1[2223:2216] > top_1[2231:2224]) ? 1 : 0;
assign detect_max[276][6] = (mid_1[2223:2216] > top_2[2215:2208]) ? 1 : 0;
assign detect_max[276][7] = (mid_1[2223:2216] > top_2[2223:2216]) ? 1 : 0;
assign detect_max[276][8] = (mid_1[2223:2216] > top_2[2231:2224]) ? 1 : 0;
assign detect_max[276][9] = (mid_1[2223:2216] > mid_0[2215:2208]) ? 1 : 0;
assign detect_max[276][10] = (mid_1[2223:2216] > mid_0[2223:2216]) ? 1 : 0;
assign detect_max[276][11] = (mid_1[2223:2216] > mid_0[2231:2224]) ? 1 : 0;
assign detect_max[276][12] = (mid_1[2223:2216] > mid_1[2215:2208]) ? 1 : 0;
assign detect_max[276][13] = (mid_1[2223:2216] > mid_1[2231:2224]) ? 1 : 0;
assign detect_max[276][14] = (mid_1[2223:2216] > mid_2[2215:2208]) ? 1 : 0;
assign detect_max[276][15] = (mid_1[2223:2216] > mid_2[2223:2216]) ? 1 : 0;
assign detect_max[276][16] = (mid_1[2223:2216] > mid_2[2231:2224]) ? 1 : 0;
assign detect_max[276][17] = (mid_1[2223:2216] > btm_0[2215:2208]) ? 1 : 0;
assign detect_max[276][18] = (mid_1[2223:2216] > btm_0[2223:2216]) ? 1 : 0;
assign detect_max[276][19] = (mid_1[2223:2216] > btm_0[2231:2224]) ? 1 : 0;
assign detect_max[276][20] = (mid_1[2223:2216] > btm_1[2215:2208]) ? 1 : 0;
assign detect_max[276][21] = (mid_1[2223:2216] > btm_1[2223:2216]) ? 1 : 0;
assign detect_max[276][22] = (mid_1[2223:2216] > btm_1[2231:2224]) ? 1 : 0;
assign detect_max[276][23] = (mid_1[2223:2216] > btm_2[2215:2208]) ? 1 : 0;
assign detect_max[276][24] = (mid_1[2223:2216] > btm_2[2223:2216]) ? 1 : 0;
assign detect_max[276][25] = (mid_1[2223:2216] > btm_2[2231:2224]) ? 1 : 0;

assign detect_max[277][0] = (mid_1[2231:2224] > top_0[2223:2216]) ? 1 : 0;
assign detect_max[277][1] = (mid_1[2231:2224] > top_0[2231:2224]) ? 1 : 0;
assign detect_max[277][2] = (mid_1[2231:2224] > top_0[2239:2232]) ? 1 : 0;
assign detect_max[277][3] = (mid_1[2231:2224] > top_1[2223:2216]) ? 1 : 0;
assign detect_max[277][4] = (mid_1[2231:2224] > top_1[2231:2224]) ? 1 : 0;
assign detect_max[277][5] = (mid_1[2231:2224] > top_1[2239:2232]) ? 1 : 0;
assign detect_max[277][6] = (mid_1[2231:2224] > top_2[2223:2216]) ? 1 : 0;
assign detect_max[277][7] = (mid_1[2231:2224] > top_2[2231:2224]) ? 1 : 0;
assign detect_max[277][8] = (mid_1[2231:2224] > top_2[2239:2232]) ? 1 : 0;
assign detect_max[277][9] = (mid_1[2231:2224] > mid_0[2223:2216]) ? 1 : 0;
assign detect_max[277][10] = (mid_1[2231:2224] > mid_0[2231:2224]) ? 1 : 0;
assign detect_max[277][11] = (mid_1[2231:2224] > mid_0[2239:2232]) ? 1 : 0;
assign detect_max[277][12] = (mid_1[2231:2224] > mid_1[2223:2216]) ? 1 : 0;
assign detect_max[277][13] = (mid_1[2231:2224] > mid_1[2239:2232]) ? 1 : 0;
assign detect_max[277][14] = (mid_1[2231:2224] > mid_2[2223:2216]) ? 1 : 0;
assign detect_max[277][15] = (mid_1[2231:2224] > mid_2[2231:2224]) ? 1 : 0;
assign detect_max[277][16] = (mid_1[2231:2224] > mid_2[2239:2232]) ? 1 : 0;
assign detect_max[277][17] = (mid_1[2231:2224] > btm_0[2223:2216]) ? 1 : 0;
assign detect_max[277][18] = (mid_1[2231:2224] > btm_0[2231:2224]) ? 1 : 0;
assign detect_max[277][19] = (mid_1[2231:2224] > btm_0[2239:2232]) ? 1 : 0;
assign detect_max[277][20] = (mid_1[2231:2224] > btm_1[2223:2216]) ? 1 : 0;
assign detect_max[277][21] = (mid_1[2231:2224] > btm_1[2231:2224]) ? 1 : 0;
assign detect_max[277][22] = (mid_1[2231:2224] > btm_1[2239:2232]) ? 1 : 0;
assign detect_max[277][23] = (mid_1[2231:2224] > btm_2[2223:2216]) ? 1 : 0;
assign detect_max[277][24] = (mid_1[2231:2224] > btm_2[2231:2224]) ? 1 : 0;
assign detect_max[277][25] = (mid_1[2231:2224] > btm_2[2239:2232]) ? 1 : 0;

assign detect_max[278][0] = (mid_1[2239:2232] > top_0[2231:2224]) ? 1 : 0;
assign detect_max[278][1] = (mid_1[2239:2232] > top_0[2239:2232]) ? 1 : 0;
assign detect_max[278][2] = (mid_1[2239:2232] > top_0[2247:2240]) ? 1 : 0;
assign detect_max[278][3] = (mid_1[2239:2232] > top_1[2231:2224]) ? 1 : 0;
assign detect_max[278][4] = (mid_1[2239:2232] > top_1[2239:2232]) ? 1 : 0;
assign detect_max[278][5] = (mid_1[2239:2232] > top_1[2247:2240]) ? 1 : 0;
assign detect_max[278][6] = (mid_1[2239:2232] > top_2[2231:2224]) ? 1 : 0;
assign detect_max[278][7] = (mid_1[2239:2232] > top_2[2239:2232]) ? 1 : 0;
assign detect_max[278][8] = (mid_1[2239:2232] > top_2[2247:2240]) ? 1 : 0;
assign detect_max[278][9] = (mid_1[2239:2232] > mid_0[2231:2224]) ? 1 : 0;
assign detect_max[278][10] = (mid_1[2239:2232] > mid_0[2239:2232]) ? 1 : 0;
assign detect_max[278][11] = (mid_1[2239:2232] > mid_0[2247:2240]) ? 1 : 0;
assign detect_max[278][12] = (mid_1[2239:2232] > mid_1[2231:2224]) ? 1 : 0;
assign detect_max[278][13] = (mid_1[2239:2232] > mid_1[2247:2240]) ? 1 : 0;
assign detect_max[278][14] = (mid_1[2239:2232] > mid_2[2231:2224]) ? 1 : 0;
assign detect_max[278][15] = (mid_1[2239:2232] > mid_2[2239:2232]) ? 1 : 0;
assign detect_max[278][16] = (mid_1[2239:2232] > mid_2[2247:2240]) ? 1 : 0;
assign detect_max[278][17] = (mid_1[2239:2232] > btm_0[2231:2224]) ? 1 : 0;
assign detect_max[278][18] = (mid_1[2239:2232] > btm_0[2239:2232]) ? 1 : 0;
assign detect_max[278][19] = (mid_1[2239:2232] > btm_0[2247:2240]) ? 1 : 0;
assign detect_max[278][20] = (mid_1[2239:2232] > btm_1[2231:2224]) ? 1 : 0;
assign detect_max[278][21] = (mid_1[2239:2232] > btm_1[2239:2232]) ? 1 : 0;
assign detect_max[278][22] = (mid_1[2239:2232] > btm_1[2247:2240]) ? 1 : 0;
assign detect_max[278][23] = (mid_1[2239:2232] > btm_2[2231:2224]) ? 1 : 0;
assign detect_max[278][24] = (mid_1[2239:2232] > btm_2[2239:2232]) ? 1 : 0;
assign detect_max[278][25] = (mid_1[2239:2232] > btm_2[2247:2240]) ? 1 : 0;

assign detect_max[279][0] = (mid_1[2247:2240] > top_0[2239:2232]) ? 1 : 0;
assign detect_max[279][1] = (mid_1[2247:2240] > top_0[2247:2240]) ? 1 : 0;
assign detect_max[279][2] = (mid_1[2247:2240] > top_0[2255:2248]) ? 1 : 0;
assign detect_max[279][3] = (mid_1[2247:2240] > top_1[2239:2232]) ? 1 : 0;
assign detect_max[279][4] = (mid_1[2247:2240] > top_1[2247:2240]) ? 1 : 0;
assign detect_max[279][5] = (mid_1[2247:2240] > top_1[2255:2248]) ? 1 : 0;
assign detect_max[279][6] = (mid_1[2247:2240] > top_2[2239:2232]) ? 1 : 0;
assign detect_max[279][7] = (mid_1[2247:2240] > top_2[2247:2240]) ? 1 : 0;
assign detect_max[279][8] = (mid_1[2247:2240] > top_2[2255:2248]) ? 1 : 0;
assign detect_max[279][9] = (mid_1[2247:2240] > mid_0[2239:2232]) ? 1 : 0;
assign detect_max[279][10] = (mid_1[2247:2240] > mid_0[2247:2240]) ? 1 : 0;
assign detect_max[279][11] = (mid_1[2247:2240] > mid_0[2255:2248]) ? 1 : 0;
assign detect_max[279][12] = (mid_1[2247:2240] > mid_1[2239:2232]) ? 1 : 0;
assign detect_max[279][13] = (mid_1[2247:2240] > mid_1[2255:2248]) ? 1 : 0;
assign detect_max[279][14] = (mid_1[2247:2240] > mid_2[2239:2232]) ? 1 : 0;
assign detect_max[279][15] = (mid_1[2247:2240] > mid_2[2247:2240]) ? 1 : 0;
assign detect_max[279][16] = (mid_1[2247:2240] > mid_2[2255:2248]) ? 1 : 0;
assign detect_max[279][17] = (mid_1[2247:2240] > btm_0[2239:2232]) ? 1 : 0;
assign detect_max[279][18] = (mid_1[2247:2240] > btm_0[2247:2240]) ? 1 : 0;
assign detect_max[279][19] = (mid_1[2247:2240] > btm_0[2255:2248]) ? 1 : 0;
assign detect_max[279][20] = (mid_1[2247:2240] > btm_1[2239:2232]) ? 1 : 0;
assign detect_max[279][21] = (mid_1[2247:2240] > btm_1[2247:2240]) ? 1 : 0;
assign detect_max[279][22] = (mid_1[2247:2240] > btm_1[2255:2248]) ? 1 : 0;
assign detect_max[279][23] = (mid_1[2247:2240] > btm_2[2239:2232]) ? 1 : 0;
assign detect_max[279][24] = (mid_1[2247:2240] > btm_2[2247:2240]) ? 1 : 0;
assign detect_max[279][25] = (mid_1[2247:2240] > btm_2[2255:2248]) ? 1 : 0;

assign detect_max[280][0] = (mid_1[2255:2248] > top_0[2247:2240]) ? 1 : 0;
assign detect_max[280][1] = (mid_1[2255:2248] > top_0[2255:2248]) ? 1 : 0;
assign detect_max[280][2] = (mid_1[2255:2248] > top_0[2263:2256]) ? 1 : 0;
assign detect_max[280][3] = (mid_1[2255:2248] > top_1[2247:2240]) ? 1 : 0;
assign detect_max[280][4] = (mid_1[2255:2248] > top_1[2255:2248]) ? 1 : 0;
assign detect_max[280][5] = (mid_1[2255:2248] > top_1[2263:2256]) ? 1 : 0;
assign detect_max[280][6] = (mid_1[2255:2248] > top_2[2247:2240]) ? 1 : 0;
assign detect_max[280][7] = (mid_1[2255:2248] > top_2[2255:2248]) ? 1 : 0;
assign detect_max[280][8] = (mid_1[2255:2248] > top_2[2263:2256]) ? 1 : 0;
assign detect_max[280][9] = (mid_1[2255:2248] > mid_0[2247:2240]) ? 1 : 0;
assign detect_max[280][10] = (mid_1[2255:2248] > mid_0[2255:2248]) ? 1 : 0;
assign detect_max[280][11] = (mid_1[2255:2248] > mid_0[2263:2256]) ? 1 : 0;
assign detect_max[280][12] = (mid_1[2255:2248] > mid_1[2247:2240]) ? 1 : 0;
assign detect_max[280][13] = (mid_1[2255:2248] > mid_1[2263:2256]) ? 1 : 0;
assign detect_max[280][14] = (mid_1[2255:2248] > mid_2[2247:2240]) ? 1 : 0;
assign detect_max[280][15] = (mid_1[2255:2248] > mid_2[2255:2248]) ? 1 : 0;
assign detect_max[280][16] = (mid_1[2255:2248] > mid_2[2263:2256]) ? 1 : 0;
assign detect_max[280][17] = (mid_1[2255:2248] > btm_0[2247:2240]) ? 1 : 0;
assign detect_max[280][18] = (mid_1[2255:2248] > btm_0[2255:2248]) ? 1 : 0;
assign detect_max[280][19] = (mid_1[2255:2248] > btm_0[2263:2256]) ? 1 : 0;
assign detect_max[280][20] = (mid_1[2255:2248] > btm_1[2247:2240]) ? 1 : 0;
assign detect_max[280][21] = (mid_1[2255:2248] > btm_1[2255:2248]) ? 1 : 0;
assign detect_max[280][22] = (mid_1[2255:2248] > btm_1[2263:2256]) ? 1 : 0;
assign detect_max[280][23] = (mid_1[2255:2248] > btm_2[2247:2240]) ? 1 : 0;
assign detect_max[280][24] = (mid_1[2255:2248] > btm_2[2255:2248]) ? 1 : 0;
assign detect_max[280][25] = (mid_1[2255:2248] > btm_2[2263:2256]) ? 1 : 0;

assign detect_max[281][0] = (mid_1[2263:2256] > top_0[2255:2248]) ? 1 : 0;
assign detect_max[281][1] = (mid_1[2263:2256] > top_0[2263:2256]) ? 1 : 0;
assign detect_max[281][2] = (mid_1[2263:2256] > top_0[2271:2264]) ? 1 : 0;
assign detect_max[281][3] = (mid_1[2263:2256] > top_1[2255:2248]) ? 1 : 0;
assign detect_max[281][4] = (mid_1[2263:2256] > top_1[2263:2256]) ? 1 : 0;
assign detect_max[281][5] = (mid_1[2263:2256] > top_1[2271:2264]) ? 1 : 0;
assign detect_max[281][6] = (mid_1[2263:2256] > top_2[2255:2248]) ? 1 : 0;
assign detect_max[281][7] = (mid_1[2263:2256] > top_2[2263:2256]) ? 1 : 0;
assign detect_max[281][8] = (mid_1[2263:2256] > top_2[2271:2264]) ? 1 : 0;
assign detect_max[281][9] = (mid_1[2263:2256] > mid_0[2255:2248]) ? 1 : 0;
assign detect_max[281][10] = (mid_1[2263:2256] > mid_0[2263:2256]) ? 1 : 0;
assign detect_max[281][11] = (mid_1[2263:2256] > mid_0[2271:2264]) ? 1 : 0;
assign detect_max[281][12] = (mid_1[2263:2256] > mid_1[2255:2248]) ? 1 : 0;
assign detect_max[281][13] = (mid_1[2263:2256] > mid_1[2271:2264]) ? 1 : 0;
assign detect_max[281][14] = (mid_1[2263:2256] > mid_2[2255:2248]) ? 1 : 0;
assign detect_max[281][15] = (mid_1[2263:2256] > mid_2[2263:2256]) ? 1 : 0;
assign detect_max[281][16] = (mid_1[2263:2256] > mid_2[2271:2264]) ? 1 : 0;
assign detect_max[281][17] = (mid_1[2263:2256] > btm_0[2255:2248]) ? 1 : 0;
assign detect_max[281][18] = (mid_1[2263:2256] > btm_0[2263:2256]) ? 1 : 0;
assign detect_max[281][19] = (mid_1[2263:2256] > btm_0[2271:2264]) ? 1 : 0;
assign detect_max[281][20] = (mid_1[2263:2256] > btm_1[2255:2248]) ? 1 : 0;
assign detect_max[281][21] = (mid_1[2263:2256] > btm_1[2263:2256]) ? 1 : 0;
assign detect_max[281][22] = (mid_1[2263:2256] > btm_1[2271:2264]) ? 1 : 0;
assign detect_max[281][23] = (mid_1[2263:2256] > btm_2[2255:2248]) ? 1 : 0;
assign detect_max[281][24] = (mid_1[2263:2256] > btm_2[2263:2256]) ? 1 : 0;
assign detect_max[281][25] = (mid_1[2263:2256] > btm_2[2271:2264]) ? 1 : 0;

assign detect_max[282][0] = (mid_1[2271:2264] > top_0[2263:2256]) ? 1 : 0;
assign detect_max[282][1] = (mid_1[2271:2264] > top_0[2271:2264]) ? 1 : 0;
assign detect_max[282][2] = (mid_1[2271:2264] > top_0[2279:2272]) ? 1 : 0;
assign detect_max[282][3] = (mid_1[2271:2264] > top_1[2263:2256]) ? 1 : 0;
assign detect_max[282][4] = (mid_1[2271:2264] > top_1[2271:2264]) ? 1 : 0;
assign detect_max[282][5] = (mid_1[2271:2264] > top_1[2279:2272]) ? 1 : 0;
assign detect_max[282][6] = (mid_1[2271:2264] > top_2[2263:2256]) ? 1 : 0;
assign detect_max[282][7] = (mid_1[2271:2264] > top_2[2271:2264]) ? 1 : 0;
assign detect_max[282][8] = (mid_1[2271:2264] > top_2[2279:2272]) ? 1 : 0;
assign detect_max[282][9] = (mid_1[2271:2264] > mid_0[2263:2256]) ? 1 : 0;
assign detect_max[282][10] = (mid_1[2271:2264] > mid_0[2271:2264]) ? 1 : 0;
assign detect_max[282][11] = (mid_1[2271:2264] > mid_0[2279:2272]) ? 1 : 0;
assign detect_max[282][12] = (mid_1[2271:2264] > mid_1[2263:2256]) ? 1 : 0;
assign detect_max[282][13] = (mid_1[2271:2264] > mid_1[2279:2272]) ? 1 : 0;
assign detect_max[282][14] = (mid_1[2271:2264] > mid_2[2263:2256]) ? 1 : 0;
assign detect_max[282][15] = (mid_1[2271:2264] > mid_2[2271:2264]) ? 1 : 0;
assign detect_max[282][16] = (mid_1[2271:2264] > mid_2[2279:2272]) ? 1 : 0;
assign detect_max[282][17] = (mid_1[2271:2264] > btm_0[2263:2256]) ? 1 : 0;
assign detect_max[282][18] = (mid_1[2271:2264] > btm_0[2271:2264]) ? 1 : 0;
assign detect_max[282][19] = (mid_1[2271:2264] > btm_0[2279:2272]) ? 1 : 0;
assign detect_max[282][20] = (mid_1[2271:2264] > btm_1[2263:2256]) ? 1 : 0;
assign detect_max[282][21] = (mid_1[2271:2264] > btm_1[2271:2264]) ? 1 : 0;
assign detect_max[282][22] = (mid_1[2271:2264] > btm_1[2279:2272]) ? 1 : 0;
assign detect_max[282][23] = (mid_1[2271:2264] > btm_2[2263:2256]) ? 1 : 0;
assign detect_max[282][24] = (mid_1[2271:2264] > btm_2[2271:2264]) ? 1 : 0;
assign detect_max[282][25] = (mid_1[2271:2264] > btm_2[2279:2272]) ? 1 : 0;

assign detect_max[283][0] = (mid_1[2279:2272] > top_0[2271:2264]) ? 1 : 0;
assign detect_max[283][1] = (mid_1[2279:2272] > top_0[2279:2272]) ? 1 : 0;
assign detect_max[283][2] = (mid_1[2279:2272] > top_0[2287:2280]) ? 1 : 0;
assign detect_max[283][3] = (mid_1[2279:2272] > top_1[2271:2264]) ? 1 : 0;
assign detect_max[283][4] = (mid_1[2279:2272] > top_1[2279:2272]) ? 1 : 0;
assign detect_max[283][5] = (mid_1[2279:2272] > top_1[2287:2280]) ? 1 : 0;
assign detect_max[283][6] = (mid_1[2279:2272] > top_2[2271:2264]) ? 1 : 0;
assign detect_max[283][7] = (mid_1[2279:2272] > top_2[2279:2272]) ? 1 : 0;
assign detect_max[283][8] = (mid_1[2279:2272] > top_2[2287:2280]) ? 1 : 0;
assign detect_max[283][9] = (mid_1[2279:2272] > mid_0[2271:2264]) ? 1 : 0;
assign detect_max[283][10] = (mid_1[2279:2272] > mid_0[2279:2272]) ? 1 : 0;
assign detect_max[283][11] = (mid_1[2279:2272] > mid_0[2287:2280]) ? 1 : 0;
assign detect_max[283][12] = (mid_1[2279:2272] > mid_1[2271:2264]) ? 1 : 0;
assign detect_max[283][13] = (mid_1[2279:2272] > mid_1[2287:2280]) ? 1 : 0;
assign detect_max[283][14] = (mid_1[2279:2272] > mid_2[2271:2264]) ? 1 : 0;
assign detect_max[283][15] = (mid_1[2279:2272] > mid_2[2279:2272]) ? 1 : 0;
assign detect_max[283][16] = (mid_1[2279:2272] > mid_2[2287:2280]) ? 1 : 0;
assign detect_max[283][17] = (mid_1[2279:2272] > btm_0[2271:2264]) ? 1 : 0;
assign detect_max[283][18] = (mid_1[2279:2272] > btm_0[2279:2272]) ? 1 : 0;
assign detect_max[283][19] = (mid_1[2279:2272] > btm_0[2287:2280]) ? 1 : 0;
assign detect_max[283][20] = (mid_1[2279:2272] > btm_1[2271:2264]) ? 1 : 0;
assign detect_max[283][21] = (mid_1[2279:2272] > btm_1[2279:2272]) ? 1 : 0;
assign detect_max[283][22] = (mid_1[2279:2272] > btm_1[2287:2280]) ? 1 : 0;
assign detect_max[283][23] = (mid_1[2279:2272] > btm_2[2271:2264]) ? 1 : 0;
assign detect_max[283][24] = (mid_1[2279:2272] > btm_2[2279:2272]) ? 1 : 0;
assign detect_max[283][25] = (mid_1[2279:2272] > btm_2[2287:2280]) ? 1 : 0;

assign detect_max[284][0] = (mid_1[2287:2280] > top_0[2279:2272]) ? 1 : 0;
assign detect_max[284][1] = (mid_1[2287:2280] > top_0[2287:2280]) ? 1 : 0;
assign detect_max[284][2] = (mid_1[2287:2280] > top_0[2295:2288]) ? 1 : 0;
assign detect_max[284][3] = (mid_1[2287:2280] > top_1[2279:2272]) ? 1 : 0;
assign detect_max[284][4] = (mid_1[2287:2280] > top_1[2287:2280]) ? 1 : 0;
assign detect_max[284][5] = (mid_1[2287:2280] > top_1[2295:2288]) ? 1 : 0;
assign detect_max[284][6] = (mid_1[2287:2280] > top_2[2279:2272]) ? 1 : 0;
assign detect_max[284][7] = (mid_1[2287:2280] > top_2[2287:2280]) ? 1 : 0;
assign detect_max[284][8] = (mid_1[2287:2280] > top_2[2295:2288]) ? 1 : 0;
assign detect_max[284][9] = (mid_1[2287:2280] > mid_0[2279:2272]) ? 1 : 0;
assign detect_max[284][10] = (mid_1[2287:2280] > mid_0[2287:2280]) ? 1 : 0;
assign detect_max[284][11] = (mid_1[2287:2280] > mid_0[2295:2288]) ? 1 : 0;
assign detect_max[284][12] = (mid_1[2287:2280] > mid_1[2279:2272]) ? 1 : 0;
assign detect_max[284][13] = (mid_1[2287:2280] > mid_1[2295:2288]) ? 1 : 0;
assign detect_max[284][14] = (mid_1[2287:2280] > mid_2[2279:2272]) ? 1 : 0;
assign detect_max[284][15] = (mid_1[2287:2280] > mid_2[2287:2280]) ? 1 : 0;
assign detect_max[284][16] = (mid_1[2287:2280] > mid_2[2295:2288]) ? 1 : 0;
assign detect_max[284][17] = (mid_1[2287:2280] > btm_0[2279:2272]) ? 1 : 0;
assign detect_max[284][18] = (mid_1[2287:2280] > btm_0[2287:2280]) ? 1 : 0;
assign detect_max[284][19] = (mid_1[2287:2280] > btm_0[2295:2288]) ? 1 : 0;
assign detect_max[284][20] = (mid_1[2287:2280] > btm_1[2279:2272]) ? 1 : 0;
assign detect_max[284][21] = (mid_1[2287:2280] > btm_1[2287:2280]) ? 1 : 0;
assign detect_max[284][22] = (mid_1[2287:2280] > btm_1[2295:2288]) ? 1 : 0;
assign detect_max[284][23] = (mid_1[2287:2280] > btm_2[2279:2272]) ? 1 : 0;
assign detect_max[284][24] = (mid_1[2287:2280] > btm_2[2287:2280]) ? 1 : 0;
assign detect_max[284][25] = (mid_1[2287:2280] > btm_2[2295:2288]) ? 1 : 0;

assign detect_max[285][0] = (mid_1[2295:2288] > top_0[2287:2280]) ? 1 : 0;
assign detect_max[285][1] = (mid_1[2295:2288] > top_0[2295:2288]) ? 1 : 0;
assign detect_max[285][2] = (mid_1[2295:2288] > top_0[2303:2296]) ? 1 : 0;
assign detect_max[285][3] = (mid_1[2295:2288] > top_1[2287:2280]) ? 1 : 0;
assign detect_max[285][4] = (mid_1[2295:2288] > top_1[2295:2288]) ? 1 : 0;
assign detect_max[285][5] = (mid_1[2295:2288] > top_1[2303:2296]) ? 1 : 0;
assign detect_max[285][6] = (mid_1[2295:2288] > top_2[2287:2280]) ? 1 : 0;
assign detect_max[285][7] = (mid_1[2295:2288] > top_2[2295:2288]) ? 1 : 0;
assign detect_max[285][8] = (mid_1[2295:2288] > top_2[2303:2296]) ? 1 : 0;
assign detect_max[285][9] = (mid_1[2295:2288] > mid_0[2287:2280]) ? 1 : 0;
assign detect_max[285][10] = (mid_1[2295:2288] > mid_0[2295:2288]) ? 1 : 0;
assign detect_max[285][11] = (mid_1[2295:2288] > mid_0[2303:2296]) ? 1 : 0;
assign detect_max[285][12] = (mid_1[2295:2288] > mid_1[2287:2280]) ? 1 : 0;
assign detect_max[285][13] = (mid_1[2295:2288] > mid_1[2303:2296]) ? 1 : 0;
assign detect_max[285][14] = (mid_1[2295:2288] > mid_2[2287:2280]) ? 1 : 0;
assign detect_max[285][15] = (mid_1[2295:2288] > mid_2[2295:2288]) ? 1 : 0;
assign detect_max[285][16] = (mid_1[2295:2288] > mid_2[2303:2296]) ? 1 : 0;
assign detect_max[285][17] = (mid_1[2295:2288] > btm_0[2287:2280]) ? 1 : 0;
assign detect_max[285][18] = (mid_1[2295:2288] > btm_0[2295:2288]) ? 1 : 0;
assign detect_max[285][19] = (mid_1[2295:2288] > btm_0[2303:2296]) ? 1 : 0;
assign detect_max[285][20] = (mid_1[2295:2288] > btm_1[2287:2280]) ? 1 : 0;
assign detect_max[285][21] = (mid_1[2295:2288] > btm_1[2295:2288]) ? 1 : 0;
assign detect_max[285][22] = (mid_1[2295:2288] > btm_1[2303:2296]) ? 1 : 0;
assign detect_max[285][23] = (mid_1[2295:2288] > btm_2[2287:2280]) ? 1 : 0;
assign detect_max[285][24] = (mid_1[2295:2288] > btm_2[2295:2288]) ? 1 : 0;
assign detect_max[285][25] = (mid_1[2295:2288] > btm_2[2303:2296]) ? 1 : 0;

assign detect_max[286][0] = (mid_1[2303:2296] > top_0[2295:2288]) ? 1 : 0;
assign detect_max[286][1] = (mid_1[2303:2296] > top_0[2303:2296]) ? 1 : 0;
assign detect_max[286][2] = (mid_1[2303:2296] > top_0[2311:2304]) ? 1 : 0;
assign detect_max[286][3] = (mid_1[2303:2296] > top_1[2295:2288]) ? 1 : 0;
assign detect_max[286][4] = (mid_1[2303:2296] > top_1[2303:2296]) ? 1 : 0;
assign detect_max[286][5] = (mid_1[2303:2296] > top_1[2311:2304]) ? 1 : 0;
assign detect_max[286][6] = (mid_1[2303:2296] > top_2[2295:2288]) ? 1 : 0;
assign detect_max[286][7] = (mid_1[2303:2296] > top_2[2303:2296]) ? 1 : 0;
assign detect_max[286][8] = (mid_1[2303:2296] > top_2[2311:2304]) ? 1 : 0;
assign detect_max[286][9] = (mid_1[2303:2296] > mid_0[2295:2288]) ? 1 : 0;
assign detect_max[286][10] = (mid_1[2303:2296] > mid_0[2303:2296]) ? 1 : 0;
assign detect_max[286][11] = (mid_1[2303:2296] > mid_0[2311:2304]) ? 1 : 0;
assign detect_max[286][12] = (mid_1[2303:2296] > mid_1[2295:2288]) ? 1 : 0;
assign detect_max[286][13] = (mid_1[2303:2296] > mid_1[2311:2304]) ? 1 : 0;
assign detect_max[286][14] = (mid_1[2303:2296] > mid_2[2295:2288]) ? 1 : 0;
assign detect_max[286][15] = (mid_1[2303:2296] > mid_2[2303:2296]) ? 1 : 0;
assign detect_max[286][16] = (mid_1[2303:2296] > mid_2[2311:2304]) ? 1 : 0;
assign detect_max[286][17] = (mid_1[2303:2296] > btm_0[2295:2288]) ? 1 : 0;
assign detect_max[286][18] = (mid_1[2303:2296] > btm_0[2303:2296]) ? 1 : 0;
assign detect_max[286][19] = (mid_1[2303:2296] > btm_0[2311:2304]) ? 1 : 0;
assign detect_max[286][20] = (mid_1[2303:2296] > btm_1[2295:2288]) ? 1 : 0;
assign detect_max[286][21] = (mid_1[2303:2296] > btm_1[2303:2296]) ? 1 : 0;
assign detect_max[286][22] = (mid_1[2303:2296] > btm_1[2311:2304]) ? 1 : 0;
assign detect_max[286][23] = (mid_1[2303:2296] > btm_2[2295:2288]) ? 1 : 0;
assign detect_max[286][24] = (mid_1[2303:2296] > btm_2[2303:2296]) ? 1 : 0;
assign detect_max[286][25] = (mid_1[2303:2296] > btm_2[2311:2304]) ? 1 : 0;

assign detect_max[287][0] = (mid_1[2311:2304] > top_0[2303:2296]) ? 1 : 0;
assign detect_max[287][1] = (mid_1[2311:2304] > top_0[2311:2304]) ? 1 : 0;
assign detect_max[287][2] = (mid_1[2311:2304] > top_0[2319:2312]) ? 1 : 0;
assign detect_max[287][3] = (mid_1[2311:2304] > top_1[2303:2296]) ? 1 : 0;
assign detect_max[287][4] = (mid_1[2311:2304] > top_1[2311:2304]) ? 1 : 0;
assign detect_max[287][5] = (mid_1[2311:2304] > top_1[2319:2312]) ? 1 : 0;
assign detect_max[287][6] = (mid_1[2311:2304] > top_2[2303:2296]) ? 1 : 0;
assign detect_max[287][7] = (mid_1[2311:2304] > top_2[2311:2304]) ? 1 : 0;
assign detect_max[287][8] = (mid_1[2311:2304] > top_2[2319:2312]) ? 1 : 0;
assign detect_max[287][9] = (mid_1[2311:2304] > mid_0[2303:2296]) ? 1 : 0;
assign detect_max[287][10] = (mid_1[2311:2304] > mid_0[2311:2304]) ? 1 : 0;
assign detect_max[287][11] = (mid_1[2311:2304] > mid_0[2319:2312]) ? 1 : 0;
assign detect_max[287][12] = (mid_1[2311:2304] > mid_1[2303:2296]) ? 1 : 0;
assign detect_max[287][13] = (mid_1[2311:2304] > mid_1[2319:2312]) ? 1 : 0;
assign detect_max[287][14] = (mid_1[2311:2304] > mid_2[2303:2296]) ? 1 : 0;
assign detect_max[287][15] = (mid_1[2311:2304] > mid_2[2311:2304]) ? 1 : 0;
assign detect_max[287][16] = (mid_1[2311:2304] > mid_2[2319:2312]) ? 1 : 0;
assign detect_max[287][17] = (mid_1[2311:2304] > btm_0[2303:2296]) ? 1 : 0;
assign detect_max[287][18] = (mid_1[2311:2304] > btm_0[2311:2304]) ? 1 : 0;
assign detect_max[287][19] = (mid_1[2311:2304] > btm_0[2319:2312]) ? 1 : 0;
assign detect_max[287][20] = (mid_1[2311:2304] > btm_1[2303:2296]) ? 1 : 0;
assign detect_max[287][21] = (mid_1[2311:2304] > btm_1[2311:2304]) ? 1 : 0;
assign detect_max[287][22] = (mid_1[2311:2304] > btm_1[2319:2312]) ? 1 : 0;
assign detect_max[287][23] = (mid_1[2311:2304] > btm_2[2303:2296]) ? 1 : 0;
assign detect_max[287][24] = (mid_1[2311:2304] > btm_2[2311:2304]) ? 1 : 0;
assign detect_max[287][25] = (mid_1[2311:2304] > btm_2[2319:2312]) ? 1 : 0;

assign detect_max[288][0] = (mid_1[2319:2312] > top_0[2311:2304]) ? 1 : 0;
assign detect_max[288][1] = (mid_1[2319:2312] > top_0[2319:2312]) ? 1 : 0;
assign detect_max[288][2] = (mid_1[2319:2312] > top_0[2327:2320]) ? 1 : 0;
assign detect_max[288][3] = (mid_1[2319:2312] > top_1[2311:2304]) ? 1 : 0;
assign detect_max[288][4] = (mid_1[2319:2312] > top_1[2319:2312]) ? 1 : 0;
assign detect_max[288][5] = (mid_1[2319:2312] > top_1[2327:2320]) ? 1 : 0;
assign detect_max[288][6] = (mid_1[2319:2312] > top_2[2311:2304]) ? 1 : 0;
assign detect_max[288][7] = (mid_1[2319:2312] > top_2[2319:2312]) ? 1 : 0;
assign detect_max[288][8] = (mid_1[2319:2312] > top_2[2327:2320]) ? 1 : 0;
assign detect_max[288][9] = (mid_1[2319:2312] > mid_0[2311:2304]) ? 1 : 0;
assign detect_max[288][10] = (mid_1[2319:2312] > mid_0[2319:2312]) ? 1 : 0;
assign detect_max[288][11] = (mid_1[2319:2312] > mid_0[2327:2320]) ? 1 : 0;
assign detect_max[288][12] = (mid_1[2319:2312] > mid_1[2311:2304]) ? 1 : 0;
assign detect_max[288][13] = (mid_1[2319:2312] > mid_1[2327:2320]) ? 1 : 0;
assign detect_max[288][14] = (mid_1[2319:2312] > mid_2[2311:2304]) ? 1 : 0;
assign detect_max[288][15] = (mid_1[2319:2312] > mid_2[2319:2312]) ? 1 : 0;
assign detect_max[288][16] = (mid_1[2319:2312] > mid_2[2327:2320]) ? 1 : 0;
assign detect_max[288][17] = (mid_1[2319:2312] > btm_0[2311:2304]) ? 1 : 0;
assign detect_max[288][18] = (mid_1[2319:2312] > btm_0[2319:2312]) ? 1 : 0;
assign detect_max[288][19] = (mid_1[2319:2312] > btm_0[2327:2320]) ? 1 : 0;
assign detect_max[288][20] = (mid_1[2319:2312] > btm_1[2311:2304]) ? 1 : 0;
assign detect_max[288][21] = (mid_1[2319:2312] > btm_1[2319:2312]) ? 1 : 0;
assign detect_max[288][22] = (mid_1[2319:2312] > btm_1[2327:2320]) ? 1 : 0;
assign detect_max[288][23] = (mid_1[2319:2312] > btm_2[2311:2304]) ? 1 : 0;
assign detect_max[288][24] = (mid_1[2319:2312] > btm_2[2319:2312]) ? 1 : 0;
assign detect_max[288][25] = (mid_1[2319:2312] > btm_2[2327:2320]) ? 1 : 0;

assign detect_max[289][0] = (mid_1[2327:2320] > top_0[2319:2312]) ? 1 : 0;
assign detect_max[289][1] = (mid_1[2327:2320] > top_0[2327:2320]) ? 1 : 0;
assign detect_max[289][2] = (mid_1[2327:2320] > top_0[2335:2328]) ? 1 : 0;
assign detect_max[289][3] = (mid_1[2327:2320] > top_1[2319:2312]) ? 1 : 0;
assign detect_max[289][4] = (mid_1[2327:2320] > top_1[2327:2320]) ? 1 : 0;
assign detect_max[289][5] = (mid_1[2327:2320] > top_1[2335:2328]) ? 1 : 0;
assign detect_max[289][6] = (mid_1[2327:2320] > top_2[2319:2312]) ? 1 : 0;
assign detect_max[289][7] = (mid_1[2327:2320] > top_2[2327:2320]) ? 1 : 0;
assign detect_max[289][8] = (mid_1[2327:2320] > top_2[2335:2328]) ? 1 : 0;
assign detect_max[289][9] = (mid_1[2327:2320] > mid_0[2319:2312]) ? 1 : 0;
assign detect_max[289][10] = (mid_1[2327:2320] > mid_0[2327:2320]) ? 1 : 0;
assign detect_max[289][11] = (mid_1[2327:2320] > mid_0[2335:2328]) ? 1 : 0;
assign detect_max[289][12] = (mid_1[2327:2320] > mid_1[2319:2312]) ? 1 : 0;
assign detect_max[289][13] = (mid_1[2327:2320] > mid_1[2335:2328]) ? 1 : 0;
assign detect_max[289][14] = (mid_1[2327:2320] > mid_2[2319:2312]) ? 1 : 0;
assign detect_max[289][15] = (mid_1[2327:2320] > mid_2[2327:2320]) ? 1 : 0;
assign detect_max[289][16] = (mid_1[2327:2320] > mid_2[2335:2328]) ? 1 : 0;
assign detect_max[289][17] = (mid_1[2327:2320] > btm_0[2319:2312]) ? 1 : 0;
assign detect_max[289][18] = (mid_1[2327:2320] > btm_0[2327:2320]) ? 1 : 0;
assign detect_max[289][19] = (mid_1[2327:2320] > btm_0[2335:2328]) ? 1 : 0;
assign detect_max[289][20] = (mid_1[2327:2320] > btm_1[2319:2312]) ? 1 : 0;
assign detect_max[289][21] = (mid_1[2327:2320] > btm_1[2327:2320]) ? 1 : 0;
assign detect_max[289][22] = (mid_1[2327:2320] > btm_1[2335:2328]) ? 1 : 0;
assign detect_max[289][23] = (mid_1[2327:2320] > btm_2[2319:2312]) ? 1 : 0;
assign detect_max[289][24] = (mid_1[2327:2320] > btm_2[2327:2320]) ? 1 : 0;
assign detect_max[289][25] = (mid_1[2327:2320] > btm_2[2335:2328]) ? 1 : 0;

assign detect_max[290][0] = (mid_1[2335:2328] > top_0[2327:2320]) ? 1 : 0;
assign detect_max[290][1] = (mid_1[2335:2328] > top_0[2335:2328]) ? 1 : 0;
assign detect_max[290][2] = (mid_1[2335:2328] > top_0[2343:2336]) ? 1 : 0;
assign detect_max[290][3] = (mid_1[2335:2328] > top_1[2327:2320]) ? 1 : 0;
assign detect_max[290][4] = (mid_1[2335:2328] > top_1[2335:2328]) ? 1 : 0;
assign detect_max[290][5] = (mid_1[2335:2328] > top_1[2343:2336]) ? 1 : 0;
assign detect_max[290][6] = (mid_1[2335:2328] > top_2[2327:2320]) ? 1 : 0;
assign detect_max[290][7] = (mid_1[2335:2328] > top_2[2335:2328]) ? 1 : 0;
assign detect_max[290][8] = (mid_1[2335:2328] > top_2[2343:2336]) ? 1 : 0;
assign detect_max[290][9] = (mid_1[2335:2328] > mid_0[2327:2320]) ? 1 : 0;
assign detect_max[290][10] = (mid_1[2335:2328] > mid_0[2335:2328]) ? 1 : 0;
assign detect_max[290][11] = (mid_1[2335:2328] > mid_0[2343:2336]) ? 1 : 0;
assign detect_max[290][12] = (mid_1[2335:2328] > mid_1[2327:2320]) ? 1 : 0;
assign detect_max[290][13] = (mid_1[2335:2328] > mid_1[2343:2336]) ? 1 : 0;
assign detect_max[290][14] = (mid_1[2335:2328] > mid_2[2327:2320]) ? 1 : 0;
assign detect_max[290][15] = (mid_1[2335:2328] > mid_2[2335:2328]) ? 1 : 0;
assign detect_max[290][16] = (mid_1[2335:2328] > mid_2[2343:2336]) ? 1 : 0;
assign detect_max[290][17] = (mid_1[2335:2328] > btm_0[2327:2320]) ? 1 : 0;
assign detect_max[290][18] = (mid_1[2335:2328] > btm_0[2335:2328]) ? 1 : 0;
assign detect_max[290][19] = (mid_1[2335:2328] > btm_0[2343:2336]) ? 1 : 0;
assign detect_max[290][20] = (mid_1[2335:2328] > btm_1[2327:2320]) ? 1 : 0;
assign detect_max[290][21] = (mid_1[2335:2328] > btm_1[2335:2328]) ? 1 : 0;
assign detect_max[290][22] = (mid_1[2335:2328] > btm_1[2343:2336]) ? 1 : 0;
assign detect_max[290][23] = (mid_1[2335:2328] > btm_2[2327:2320]) ? 1 : 0;
assign detect_max[290][24] = (mid_1[2335:2328] > btm_2[2335:2328]) ? 1 : 0;
assign detect_max[290][25] = (mid_1[2335:2328] > btm_2[2343:2336]) ? 1 : 0;

assign detect_max[291][0] = (mid_1[2343:2336] > top_0[2335:2328]) ? 1 : 0;
assign detect_max[291][1] = (mid_1[2343:2336] > top_0[2343:2336]) ? 1 : 0;
assign detect_max[291][2] = (mid_1[2343:2336] > top_0[2351:2344]) ? 1 : 0;
assign detect_max[291][3] = (mid_1[2343:2336] > top_1[2335:2328]) ? 1 : 0;
assign detect_max[291][4] = (mid_1[2343:2336] > top_1[2343:2336]) ? 1 : 0;
assign detect_max[291][5] = (mid_1[2343:2336] > top_1[2351:2344]) ? 1 : 0;
assign detect_max[291][6] = (mid_1[2343:2336] > top_2[2335:2328]) ? 1 : 0;
assign detect_max[291][7] = (mid_1[2343:2336] > top_2[2343:2336]) ? 1 : 0;
assign detect_max[291][8] = (mid_1[2343:2336] > top_2[2351:2344]) ? 1 : 0;
assign detect_max[291][9] = (mid_1[2343:2336] > mid_0[2335:2328]) ? 1 : 0;
assign detect_max[291][10] = (mid_1[2343:2336] > mid_0[2343:2336]) ? 1 : 0;
assign detect_max[291][11] = (mid_1[2343:2336] > mid_0[2351:2344]) ? 1 : 0;
assign detect_max[291][12] = (mid_1[2343:2336] > mid_1[2335:2328]) ? 1 : 0;
assign detect_max[291][13] = (mid_1[2343:2336] > mid_1[2351:2344]) ? 1 : 0;
assign detect_max[291][14] = (mid_1[2343:2336] > mid_2[2335:2328]) ? 1 : 0;
assign detect_max[291][15] = (mid_1[2343:2336] > mid_2[2343:2336]) ? 1 : 0;
assign detect_max[291][16] = (mid_1[2343:2336] > mid_2[2351:2344]) ? 1 : 0;
assign detect_max[291][17] = (mid_1[2343:2336] > btm_0[2335:2328]) ? 1 : 0;
assign detect_max[291][18] = (mid_1[2343:2336] > btm_0[2343:2336]) ? 1 : 0;
assign detect_max[291][19] = (mid_1[2343:2336] > btm_0[2351:2344]) ? 1 : 0;
assign detect_max[291][20] = (mid_1[2343:2336] > btm_1[2335:2328]) ? 1 : 0;
assign detect_max[291][21] = (mid_1[2343:2336] > btm_1[2343:2336]) ? 1 : 0;
assign detect_max[291][22] = (mid_1[2343:2336] > btm_1[2351:2344]) ? 1 : 0;
assign detect_max[291][23] = (mid_1[2343:2336] > btm_2[2335:2328]) ? 1 : 0;
assign detect_max[291][24] = (mid_1[2343:2336] > btm_2[2343:2336]) ? 1 : 0;
assign detect_max[291][25] = (mid_1[2343:2336] > btm_2[2351:2344]) ? 1 : 0;

assign detect_max[292][0] = (mid_1[2351:2344] > top_0[2343:2336]) ? 1 : 0;
assign detect_max[292][1] = (mid_1[2351:2344] > top_0[2351:2344]) ? 1 : 0;
assign detect_max[292][2] = (mid_1[2351:2344] > top_0[2359:2352]) ? 1 : 0;
assign detect_max[292][3] = (mid_1[2351:2344] > top_1[2343:2336]) ? 1 : 0;
assign detect_max[292][4] = (mid_1[2351:2344] > top_1[2351:2344]) ? 1 : 0;
assign detect_max[292][5] = (mid_1[2351:2344] > top_1[2359:2352]) ? 1 : 0;
assign detect_max[292][6] = (mid_1[2351:2344] > top_2[2343:2336]) ? 1 : 0;
assign detect_max[292][7] = (mid_1[2351:2344] > top_2[2351:2344]) ? 1 : 0;
assign detect_max[292][8] = (mid_1[2351:2344] > top_2[2359:2352]) ? 1 : 0;
assign detect_max[292][9] = (mid_1[2351:2344] > mid_0[2343:2336]) ? 1 : 0;
assign detect_max[292][10] = (mid_1[2351:2344] > mid_0[2351:2344]) ? 1 : 0;
assign detect_max[292][11] = (mid_1[2351:2344] > mid_0[2359:2352]) ? 1 : 0;
assign detect_max[292][12] = (mid_1[2351:2344] > mid_1[2343:2336]) ? 1 : 0;
assign detect_max[292][13] = (mid_1[2351:2344] > mid_1[2359:2352]) ? 1 : 0;
assign detect_max[292][14] = (mid_1[2351:2344] > mid_2[2343:2336]) ? 1 : 0;
assign detect_max[292][15] = (mid_1[2351:2344] > mid_2[2351:2344]) ? 1 : 0;
assign detect_max[292][16] = (mid_1[2351:2344] > mid_2[2359:2352]) ? 1 : 0;
assign detect_max[292][17] = (mid_1[2351:2344] > btm_0[2343:2336]) ? 1 : 0;
assign detect_max[292][18] = (mid_1[2351:2344] > btm_0[2351:2344]) ? 1 : 0;
assign detect_max[292][19] = (mid_1[2351:2344] > btm_0[2359:2352]) ? 1 : 0;
assign detect_max[292][20] = (mid_1[2351:2344] > btm_1[2343:2336]) ? 1 : 0;
assign detect_max[292][21] = (mid_1[2351:2344] > btm_1[2351:2344]) ? 1 : 0;
assign detect_max[292][22] = (mid_1[2351:2344] > btm_1[2359:2352]) ? 1 : 0;
assign detect_max[292][23] = (mid_1[2351:2344] > btm_2[2343:2336]) ? 1 : 0;
assign detect_max[292][24] = (mid_1[2351:2344] > btm_2[2351:2344]) ? 1 : 0;
assign detect_max[292][25] = (mid_1[2351:2344] > btm_2[2359:2352]) ? 1 : 0;

assign detect_max[293][0] = (mid_1[2359:2352] > top_0[2351:2344]) ? 1 : 0;
assign detect_max[293][1] = (mid_1[2359:2352] > top_0[2359:2352]) ? 1 : 0;
assign detect_max[293][2] = (mid_1[2359:2352] > top_0[2367:2360]) ? 1 : 0;
assign detect_max[293][3] = (mid_1[2359:2352] > top_1[2351:2344]) ? 1 : 0;
assign detect_max[293][4] = (mid_1[2359:2352] > top_1[2359:2352]) ? 1 : 0;
assign detect_max[293][5] = (mid_1[2359:2352] > top_1[2367:2360]) ? 1 : 0;
assign detect_max[293][6] = (mid_1[2359:2352] > top_2[2351:2344]) ? 1 : 0;
assign detect_max[293][7] = (mid_1[2359:2352] > top_2[2359:2352]) ? 1 : 0;
assign detect_max[293][8] = (mid_1[2359:2352] > top_2[2367:2360]) ? 1 : 0;
assign detect_max[293][9] = (mid_1[2359:2352] > mid_0[2351:2344]) ? 1 : 0;
assign detect_max[293][10] = (mid_1[2359:2352] > mid_0[2359:2352]) ? 1 : 0;
assign detect_max[293][11] = (mid_1[2359:2352] > mid_0[2367:2360]) ? 1 : 0;
assign detect_max[293][12] = (mid_1[2359:2352] > mid_1[2351:2344]) ? 1 : 0;
assign detect_max[293][13] = (mid_1[2359:2352] > mid_1[2367:2360]) ? 1 : 0;
assign detect_max[293][14] = (mid_1[2359:2352] > mid_2[2351:2344]) ? 1 : 0;
assign detect_max[293][15] = (mid_1[2359:2352] > mid_2[2359:2352]) ? 1 : 0;
assign detect_max[293][16] = (mid_1[2359:2352] > mid_2[2367:2360]) ? 1 : 0;
assign detect_max[293][17] = (mid_1[2359:2352] > btm_0[2351:2344]) ? 1 : 0;
assign detect_max[293][18] = (mid_1[2359:2352] > btm_0[2359:2352]) ? 1 : 0;
assign detect_max[293][19] = (mid_1[2359:2352] > btm_0[2367:2360]) ? 1 : 0;
assign detect_max[293][20] = (mid_1[2359:2352] > btm_1[2351:2344]) ? 1 : 0;
assign detect_max[293][21] = (mid_1[2359:2352] > btm_1[2359:2352]) ? 1 : 0;
assign detect_max[293][22] = (mid_1[2359:2352] > btm_1[2367:2360]) ? 1 : 0;
assign detect_max[293][23] = (mid_1[2359:2352] > btm_2[2351:2344]) ? 1 : 0;
assign detect_max[293][24] = (mid_1[2359:2352] > btm_2[2359:2352]) ? 1 : 0;
assign detect_max[293][25] = (mid_1[2359:2352] > btm_2[2367:2360]) ? 1 : 0;

assign detect_max[294][0] = (mid_1[2367:2360] > top_0[2359:2352]) ? 1 : 0;
assign detect_max[294][1] = (mid_1[2367:2360] > top_0[2367:2360]) ? 1 : 0;
assign detect_max[294][2] = (mid_1[2367:2360] > top_0[2375:2368]) ? 1 : 0;
assign detect_max[294][3] = (mid_1[2367:2360] > top_1[2359:2352]) ? 1 : 0;
assign detect_max[294][4] = (mid_1[2367:2360] > top_1[2367:2360]) ? 1 : 0;
assign detect_max[294][5] = (mid_1[2367:2360] > top_1[2375:2368]) ? 1 : 0;
assign detect_max[294][6] = (mid_1[2367:2360] > top_2[2359:2352]) ? 1 : 0;
assign detect_max[294][7] = (mid_1[2367:2360] > top_2[2367:2360]) ? 1 : 0;
assign detect_max[294][8] = (mid_1[2367:2360] > top_2[2375:2368]) ? 1 : 0;
assign detect_max[294][9] = (mid_1[2367:2360] > mid_0[2359:2352]) ? 1 : 0;
assign detect_max[294][10] = (mid_1[2367:2360] > mid_0[2367:2360]) ? 1 : 0;
assign detect_max[294][11] = (mid_1[2367:2360] > mid_0[2375:2368]) ? 1 : 0;
assign detect_max[294][12] = (mid_1[2367:2360] > mid_1[2359:2352]) ? 1 : 0;
assign detect_max[294][13] = (mid_1[2367:2360] > mid_1[2375:2368]) ? 1 : 0;
assign detect_max[294][14] = (mid_1[2367:2360] > mid_2[2359:2352]) ? 1 : 0;
assign detect_max[294][15] = (mid_1[2367:2360] > mid_2[2367:2360]) ? 1 : 0;
assign detect_max[294][16] = (mid_1[2367:2360] > mid_2[2375:2368]) ? 1 : 0;
assign detect_max[294][17] = (mid_1[2367:2360] > btm_0[2359:2352]) ? 1 : 0;
assign detect_max[294][18] = (mid_1[2367:2360] > btm_0[2367:2360]) ? 1 : 0;
assign detect_max[294][19] = (mid_1[2367:2360] > btm_0[2375:2368]) ? 1 : 0;
assign detect_max[294][20] = (mid_1[2367:2360] > btm_1[2359:2352]) ? 1 : 0;
assign detect_max[294][21] = (mid_1[2367:2360] > btm_1[2367:2360]) ? 1 : 0;
assign detect_max[294][22] = (mid_1[2367:2360] > btm_1[2375:2368]) ? 1 : 0;
assign detect_max[294][23] = (mid_1[2367:2360] > btm_2[2359:2352]) ? 1 : 0;
assign detect_max[294][24] = (mid_1[2367:2360] > btm_2[2367:2360]) ? 1 : 0;
assign detect_max[294][25] = (mid_1[2367:2360] > btm_2[2375:2368]) ? 1 : 0;

assign detect_max[295][0] = (mid_1[2375:2368] > top_0[2367:2360]) ? 1 : 0;
assign detect_max[295][1] = (mid_1[2375:2368] > top_0[2375:2368]) ? 1 : 0;
assign detect_max[295][2] = (mid_1[2375:2368] > top_0[2383:2376]) ? 1 : 0;
assign detect_max[295][3] = (mid_1[2375:2368] > top_1[2367:2360]) ? 1 : 0;
assign detect_max[295][4] = (mid_1[2375:2368] > top_1[2375:2368]) ? 1 : 0;
assign detect_max[295][5] = (mid_1[2375:2368] > top_1[2383:2376]) ? 1 : 0;
assign detect_max[295][6] = (mid_1[2375:2368] > top_2[2367:2360]) ? 1 : 0;
assign detect_max[295][7] = (mid_1[2375:2368] > top_2[2375:2368]) ? 1 : 0;
assign detect_max[295][8] = (mid_1[2375:2368] > top_2[2383:2376]) ? 1 : 0;
assign detect_max[295][9] = (mid_1[2375:2368] > mid_0[2367:2360]) ? 1 : 0;
assign detect_max[295][10] = (mid_1[2375:2368] > mid_0[2375:2368]) ? 1 : 0;
assign detect_max[295][11] = (mid_1[2375:2368] > mid_0[2383:2376]) ? 1 : 0;
assign detect_max[295][12] = (mid_1[2375:2368] > mid_1[2367:2360]) ? 1 : 0;
assign detect_max[295][13] = (mid_1[2375:2368] > mid_1[2383:2376]) ? 1 : 0;
assign detect_max[295][14] = (mid_1[2375:2368] > mid_2[2367:2360]) ? 1 : 0;
assign detect_max[295][15] = (mid_1[2375:2368] > mid_2[2375:2368]) ? 1 : 0;
assign detect_max[295][16] = (mid_1[2375:2368] > mid_2[2383:2376]) ? 1 : 0;
assign detect_max[295][17] = (mid_1[2375:2368] > btm_0[2367:2360]) ? 1 : 0;
assign detect_max[295][18] = (mid_1[2375:2368] > btm_0[2375:2368]) ? 1 : 0;
assign detect_max[295][19] = (mid_1[2375:2368] > btm_0[2383:2376]) ? 1 : 0;
assign detect_max[295][20] = (mid_1[2375:2368] > btm_1[2367:2360]) ? 1 : 0;
assign detect_max[295][21] = (mid_1[2375:2368] > btm_1[2375:2368]) ? 1 : 0;
assign detect_max[295][22] = (mid_1[2375:2368] > btm_1[2383:2376]) ? 1 : 0;
assign detect_max[295][23] = (mid_1[2375:2368] > btm_2[2367:2360]) ? 1 : 0;
assign detect_max[295][24] = (mid_1[2375:2368] > btm_2[2375:2368]) ? 1 : 0;
assign detect_max[295][25] = (mid_1[2375:2368] > btm_2[2383:2376]) ? 1 : 0;

assign detect_max[296][0] = (mid_1[2383:2376] > top_0[2375:2368]) ? 1 : 0;
assign detect_max[296][1] = (mid_1[2383:2376] > top_0[2383:2376]) ? 1 : 0;
assign detect_max[296][2] = (mid_1[2383:2376] > top_0[2391:2384]) ? 1 : 0;
assign detect_max[296][3] = (mid_1[2383:2376] > top_1[2375:2368]) ? 1 : 0;
assign detect_max[296][4] = (mid_1[2383:2376] > top_1[2383:2376]) ? 1 : 0;
assign detect_max[296][5] = (mid_1[2383:2376] > top_1[2391:2384]) ? 1 : 0;
assign detect_max[296][6] = (mid_1[2383:2376] > top_2[2375:2368]) ? 1 : 0;
assign detect_max[296][7] = (mid_1[2383:2376] > top_2[2383:2376]) ? 1 : 0;
assign detect_max[296][8] = (mid_1[2383:2376] > top_2[2391:2384]) ? 1 : 0;
assign detect_max[296][9] = (mid_1[2383:2376] > mid_0[2375:2368]) ? 1 : 0;
assign detect_max[296][10] = (mid_1[2383:2376] > mid_0[2383:2376]) ? 1 : 0;
assign detect_max[296][11] = (mid_1[2383:2376] > mid_0[2391:2384]) ? 1 : 0;
assign detect_max[296][12] = (mid_1[2383:2376] > mid_1[2375:2368]) ? 1 : 0;
assign detect_max[296][13] = (mid_1[2383:2376] > mid_1[2391:2384]) ? 1 : 0;
assign detect_max[296][14] = (mid_1[2383:2376] > mid_2[2375:2368]) ? 1 : 0;
assign detect_max[296][15] = (mid_1[2383:2376] > mid_2[2383:2376]) ? 1 : 0;
assign detect_max[296][16] = (mid_1[2383:2376] > mid_2[2391:2384]) ? 1 : 0;
assign detect_max[296][17] = (mid_1[2383:2376] > btm_0[2375:2368]) ? 1 : 0;
assign detect_max[296][18] = (mid_1[2383:2376] > btm_0[2383:2376]) ? 1 : 0;
assign detect_max[296][19] = (mid_1[2383:2376] > btm_0[2391:2384]) ? 1 : 0;
assign detect_max[296][20] = (mid_1[2383:2376] > btm_1[2375:2368]) ? 1 : 0;
assign detect_max[296][21] = (mid_1[2383:2376] > btm_1[2383:2376]) ? 1 : 0;
assign detect_max[296][22] = (mid_1[2383:2376] > btm_1[2391:2384]) ? 1 : 0;
assign detect_max[296][23] = (mid_1[2383:2376] > btm_2[2375:2368]) ? 1 : 0;
assign detect_max[296][24] = (mid_1[2383:2376] > btm_2[2383:2376]) ? 1 : 0;
assign detect_max[296][25] = (mid_1[2383:2376] > btm_2[2391:2384]) ? 1 : 0;

assign detect_max[297][0] = (mid_1[2391:2384] > top_0[2383:2376]) ? 1 : 0;
assign detect_max[297][1] = (mid_1[2391:2384] > top_0[2391:2384]) ? 1 : 0;
assign detect_max[297][2] = (mid_1[2391:2384] > top_0[2399:2392]) ? 1 : 0;
assign detect_max[297][3] = (mid_1[2391:2384] > top_1[2383:2376]) ? 1 : 0;
assign detect_max[297][4] = (mid_1[2391:2384] > top_1[2391:2384]) ? 1 : 0;
assign detect_max[297][5] = (mid_1[2391:2384] > top_1[2399:2392]) ? 1 : 0;
assign detect_max[297][6] = (mid_1[2391:2384] > top_2[2383:2376]) ? 1 : 0;
assign detect_max[297][7] = (mid_1[2391:2384] > top_2[2391:2384]) ? 1 : 0;
assign detect_max[297][8] = (mid_1[2391:2384] > top_2[2399:2392]) ? 1 : 0;
assign detect_max[297][9] = (mid_1[2391:2384] > mid_0[2383:2376]) ? 1 : 0;
assign detect_max[297][10] = (mid_1[2391:2384] > mid_0[2391:2384]) ? 1 : 0;
assign detect_max[297][11] = (mid_1[2391:2384] > mid_0[2399:2392]) ? 1 : 0;
assign detect_max[297][12] = (mid_1[2391:2384] > mid_1[2383:2376]) ? 1 : 0;
assign detect_max[297][13] = (mid_1[2391:2384] > mid_1[2399:2392]) ? 1 : 0;
assign detect_max[297][14] = (mid_1[2391:2384] > mid_2[2383:2376]) ? 1 : 0;
assign detect_max[297][15] = (mid_1[2391:2384] > mid_2[2391:2384]) ? 1 : 0;
assign detect_max[297][16] = (mid_1[2391:2384] > mid_2[2399:2392]) ? 1 : 0;
assign detect_max[297][17] = (mid_1[2391:2384] > btm_0[2383:2376]) ? 1 : 0;
assign detect_max[297][18] = (mid_1[2391:2384] > btm_0[2391:2384]) ? 1 : 0;
assign detect_max[297][19] = (mid_1[2391:2384] > btm_0[2399:2392]) ? 1 : 0;
assign detect_max[297][20] = (mid_1[2391:2384] > btm_1[2383:2376]) ? 1 : 0;
assign detect_max[297][21] = (mid_1[2391:2384] > btm_1[2391:2384]) ? 1 : 0;
assign detect_max[297][22] = (mid_1[2391:2384] > btm_1[2399:2392]) ? 1 : 0;
assign detect_max[297][23] = (mid_1[2391:2384] > btm_2[2383:2376]) ? 1 : 0;
assign detect_max[297][24] = (mid_1[2391:2384] > btm_2[2391:2384]) ? 1 : 0;
assign detect_max[297][25] = (mid_1[2391:2384] > btm_2[2399:2392]) ? 1 : 0;

assign detect_max[298][0] = (mid_1[2399:2392] > top_0[2391:2384]) ? 1 : 0;
assign detect_max[298][1] = (mid_1[2399:2392] > top_0[2399:2392]) ? 1 : 0;
assign detect_max[298][2] = (mid_1[2399:2392] > top_0[2407:2400]) ? 1 : 0;
assign detect_max[298][3] = (mid_1[2399:2392] > top_1[2391:2384]) ? 1 : 0;
assign detect_max[298][4] = (mid_1[2399:2392] > top_1[2399:2392]) ? 1 : 0;
assign detect_max[298][5] = (mid_1[2399:2392] > top_1[2407:2400]) ? 1 : 0;
assign detect_max[298][6] = (mid_1[2399:2392] > top_2[2391:2384]) ? 1 : 0;
assign detect_max[298][7] = (mid_1[2399:2392] > top_2[2399:2392]) ? 1 : 0;
assign detect_max[298][8] = (mid_1[2399:2392] > top_2[2407:2400]) ? 1 : 0;
assign detect_max[298][9] = (mid_1[2399:2392] > mid_0[2391:2384]) ? 1 : 0;
assign detect_max[298][10] = (mid_1[2399:2392] > mid_0[2399:2392]) ? 1 : 0;
assign detect_max[298][11] = (mid_1[2399:2392] > mid_0[2407:2400]) ? 1 : 0;
assign detect_max[298][12] = (mid_1[2399:2392] > mid_1[2391:2384]) ? 1 : 0;
assign detect_max[298][13] = (mid_1[2399:2392] > mid_1[2407:2400]) ? 1 : 0;
assign detect_max[298][14] = (mid_1[2399:2392] > mid_2[2391:2384]) ? 1 : 0;
assign detect_max[298][15] = (mid_1[2399:2392] > mid_2[2399:2392]) ? 1 : 0;
assign detect_max[298][16] = (mid_1[2399:2392] > mid_2[2407:2400]) ? 1 : 0;
assign detect_max[298][17] = (mid_1[2399:2392] > btm_0[2391:2384]) ? 1 : 0;
assign detect_max[298][18] = (mid_1[2399:2392] > btm_0[2399:2392]) ? 1 : 0;
assign detect_max[298][19] = (mid_1[2399:2392] > btm_0[2407:2400]) ? 1 : 0;
assign detect_max[298][20] = (mid_1[2399:2392] > btm_1[2391:2384]) ? 1 : 0;
assign detect_max[298][21] = (mid_1[2399:2392] > btm_1[2399:2392]) ? 1 : 0;
assign detect_max[298][22] = (mid_1[2399:2392] > btm_1[2407:2400]) ? 1 : 0;
assign detect_max[298][23] = (mid_1[2399:2392] > btm_2[2391:2384]) ? 1 : 0;
assign detect_max[298][24] = (mid_1[2399:2392] > btm_2[2399:2392]) ? 1 : 0;
assign detect_max[298][25] = (mid_1[2399:2392] > btm_2[2407:2400]) ? 1 : 0;

assign detect_max[299][0] = (mid_1[2407:2400] > top_0[2399:2392]) ? 1 : 0;
assign detect_max[299][1] = (mid_1[2407:2400] > top_0[2407:2400]) ? 1 : 0;
assign detect_max[299][2] = (mid_1[2407:2400] > top_0[2415:2408]) ? 1 : 0;
assign detect_max[299][3] = (mid_1[2407:2400] > top_1[2399:2392]) ? 1 : 0;
assign detect_max[299][4] = (mid_1[2407:2400] > top_1[2407:2400]) ? 1 : 0;
assign detect_max[299][5] = (mid_1[2407:2400] > top_1[2415:2408]) ? 1 : 0;
assign detect_max[299][6] = (mid_1[2407:2400] > top_2[2399:2392]) ? 1 : 0;
assign detect_max[299][7] = (mid_1[2407:2400] > top_2[2407:2400]) ? 1 : 0;
assign detect_max[299][8] = (mid_1[2407:2400] > top_2[2415:2408]) ? 1 : 0;
assign detect_max[299][9] = (mid_1[2407:2400] > mid_0[2399:2392]) ? 1 : 0;
assign detect_max[299][10] = (mid_1[2407:2400] > mid_0[2407:2400]) ? 1 : 0;
assign detect_max[299][11] = (mid_1[2407:2400] > mid_0[2415:2408]) ? 1 : 0;
assign detect_max[299][12] = (mid_1[2407:2400] > mid_1[2399:2392]) ? 1 : 0;
assign detect_max[299][13] = (mid_1[2407:2400] > mid_1[2415:2408]) ? 1 : 0;
assign detect_max[299][14] = (mid_1[2407:2400] > mid_2[2399:2392]) ? 1 : 0;
assign detect_max[299][15] = (mid_1[2407:2400] > mid_2[2407:2400]) ? 1 : 0;
assign detect_max[299][16] = (mid_1[2407:2400] > mid_2[2415:2408]) ? 1 : 0;
assign detect_max[299][17] = (mid_1[2407:2400] > btm_0[2399:2392]) ? 1 : 0;
assign detect_max[299][18] = (mid_1[2407:2400] > btm_0[2407:2400]) ? 1 : 0;
assign detect_max[299][19] = (mid_1[2407:2400] > btm_0[2415:2408]) ? 1 : 0;
assign detect_max[299][20] = (mid_1[2407:2400] > btm_1[2399:2392]) ? 1 : 0;
assign detect_max[299][21] = (mid_1[2407:2400] > btm_1[2407:2400]) ? 1 : 0;
assign detect_max[299][22] = (mid_1[2407:2400] > btm_1[2415:2408]) ? 1 : 0;
assign detect_max[299][23] = (mid_1[2407:2400] > btm_2[2399:2392]) ? 1 : 0;
assign detect_max[299][24] = (mid_1[2407:2400] > btm_2[2407:2400]) ? 1 : 0;
assign detect_max[299][25] = (mid_1[2407:2400] > btm_2[2415:2408]) ? 1 : 0;

assign detect_max[300][0] = (mid_1[2415:2408] > top_0[2407:2400]) ? 1 : 0;
assign detect_max[300][1] = (mid_1[2415:2408] > top_0[2415:2408]) ? 1 : 0;
assign detect_max[300][2] = (mid_1[2415:2408] > top_0[2423:2416]) ? 1 : 0;
assign detect_max[300][3] = (mid_1[2415:2408] > top_1[2407:2400]) ? 1 : 0;
assign detect_max[300][4] = (mid_1[2415:2408] > top_1[2415:2408]) ? 1 : 0;
assign detect_max[300][5] = (mid_1[2415:2408] > top_1[2423:2416]) ? 1 : 0;
assign detect_max[300][6] = (mid_1[2415:2408] > top_2[2407:2400]) ? 1 : 0;
assign detect_max[300][7] = (mid_1[2415:2408] > top_2[2415:2408]) ? 1 : 0;
assign detect_max[300][8] = (mid_1[2415:2408] > top_2[2423:2416]) ? 1 : 0;
assign detect_max[300][9] = (mid_1[2415:2408] > mid_0[2407:2400]) ? 1 : 0;
assign detect_max[300][10] = (mid_1[2415:2408] > mid_0[2415:2408]) ? 1 : 0;
assign detect_max[300][11] = (mid_1[2415:2408] > mid_0[2423:2416]) ? 1 : 0;
assign detect_max[300][12] = (mid_1[2415:2408] > mid_1[2407:2400]) ? 1 : 0;
assign detect_max[300][13] = (mid_1[2415:2408] > mid_1[2423:2416]) ? 1 : 0;
assign detect_max[300][14] = (mid_1[2415:2408] > mid_2[2407:2400]) ? 1 : 0;
assign detect_max[300][15] = (mid_1[2415:2408] > mid_2[2415:2408]) ? 1 : 0;
assign detect_max[300][16] = (mid_1[2415:2408] > mid_2[2423:2416]) ? 1 : 0;
assign detect_max[300][17] = (mid_1[2415:2408] > btm_0[2407:2400]) ? 1 : 0;
assign detect_max[300][18] = (mid_1[2415:2408] > btm_0[2415:2408]) ? 1 : 0;
assign detect_max[300][19] = (mid_1[2415:2408] > btm_0[2423:2416]) ? 1 : 0;
assign detect_max[300][20] = (mid_1[2415:2408] > btm_1[2407:2400]) ? 1 : 0;
assign detect_max[300][21] = (mid_1[2415:2408] > btm_1[2415:2408]) ? 1 : 0;
assign detect_max[300][22] = (mid_1[2415:2408] > btm_1[2423:2416]) ? 1 : 0;
assign detect_max[300][23] = (mid_1[2415:2408] > btm_2[2407:2400]) ? 1 : 0;
assign detect_max[300][24] = (mid_1[2415:2408] > btm_2[2415:2408]) ? 1 : 0;
assign detect_max[300][25] = (mid_1[2415:2408] > btm_2[2423:2416]) ? 1 : 0;

assign detect_max[301][0] = (mid_1[2423:2416] > top_0[2415:2408]) ? 1 : 0;
assign detect_max[301][1] = (mid_1[2423:2416] > top_0[2423:2416]) ? 1 : 0;
assign detect_max[301][2] = (mid_1[2423:2416] > top_0[2431:2424]) ? 1 : 0;
assign detect_max[301][3] = (mid_1[2423:2416] > top_1[2415:2408]) ? 1 : 0;
assign detect_max[301][4] = (mid_1[2423:2416] > top_1[2423:2416]) ? 1 : 0;
assign detect_max[301][5] = (mid_1[2423:2416] > top_1[2431:2424]) ? 1 : 0;
assign detect_max[301][6] = (mid_1[2423:2416] > top_2[2415:2408]) ? 1 : 0;
assign detect_max[301][7] = (mid_1[2423:2416] > top_2[2423:2416]) ? 1 : 0;
assign detect_max[301][8] = (mid_1[2423:2416] > top_2[2431:2424]) ? 1 : 0;
assign detect_max[301][9] = (mid_1[2423:2416] > mid_0[2415:2408]) ? 1 : 0;
assign detect_max[301][10] = (mid_1[2423:2416] > mid_0[2423:2416]) ? 1 : 0;
assign detect_max[301][11] = (mid_1[2423:2416] > mid_0[2431:2424]) ? 1 : 0;
assign detect_max[301][12] = (mid_1[2423:2416] > mid_1[2415:2408]) ? 1 : 0;
assign detect_max[301][13] = (mid_1[2423:2416] > mid_1[2431:2424]) ? 1 : 0;
assign detect_max[301][14] = (mid_1[2423:2416] > mid_2[2415:2408]) ? 1 : 0;
assign detect_max[301][15] = (mid_1[2423:2416] > mid_2[2423:2416]) ? 1 : 0;
assign detect_max[301][16] = (mid_1[2423:2416] > mid_2[2431:2424]) ? 1 : 0;
assign detect_max[301][17] = (mid_1[2423:2416] > btm_0[2415:2408]) ? 1 : 0;
assign detect_max[301][18] = (mid_1[2423:2416] > btm_0[2423:2416]) ? 1 : 0;
assign detect_max[301][19] = (mid_1[2423:2416] > btm_0[2431:2424]) ? 1 : 0;
assign detect_max[301][20] = (mid_1[2423:2416] > btm_1[2415:2408]) ? 1 : 0;
assign detect_max[301][21] = (mid_1[2423:2416] > btm_1[2423:2416]) ? 1 : 0;
assign detect_max[301][22] = (mid_1[2423:2416] > btm_1[2431:2424]) ? 1 : 0;
assign detect_max[301][23] = (mid_1[2423:2416] > btm_2[2415:2408]) ? 1 : 0;
assign detect_max[301][24] = (mid_1[2423:2416] > btm_2[2423:2416]) ? 1 : 0;
assign detect_max[301][25] = (mid_1[2423:2416] > btm_2[2431:2424]) ? 1 : 0;

assign detect_max[302][0] = (mid_1[2431:2424] > top_0[2423:2416]) ? 1 : 0;
assign detect_max[302][1] = (mid_1[2431:2424] > top_0[2431:2424]) ? 1 : 0;
assign detect_max[302][2] = (mid_1[2431:2424] > top_0[2439:2432]) ? 1 : 0;
assign detect_max[302][3] = (mid_1[2431:2424] > top_1[2423:2416]) ? 1 : 0;
assign detect_max[302][4] = (mid_1[2431:2424] > top_1[2431:2424]) ? 1 : 0;
assign detect_max[302][5] = (mid_1[2431:2424] > top_1[2439:2432]) ? 1 : 0;
assign detect_max[302][6] = (mid_1[2431:2424] > top_2[2423:2416]) ? 1 : 0;
assign detect_max[302][7] = (mid_1[2431:2424] > top_2[2431:2424]) ? 1 : 0;
assign detect_max[302][8] = (mid_1[2431:2424] > top_2[2439:2432]) ? 1 : 0;
assign detect_max[302][9] = (mid_1[2431:2424] > mid_0[2423:2416]) ? 1 : 0;
assign detect_max[302][10] = (mid_1[2431:2424] > mid_0[2431:2424]) ? 1 : 0;
assign detect_max[302][11] = (mid_1[2431:2424] > mid_0[2439:2432]) ? 1 : 0;
assign detect_max[302][12] = (mid_1[2431:2424] > mid_1[2423:2416]) ? 1 : 0;
assign detect_max[302][13] = (mid_1[2431:2424] > mid_1[2439:2432]) ? 1 : 0;
assign detect_max[302][14] = (mid_1[2431:2424] > mid_2[2423:2416]) ? 1 : 0;
assign detect_max[302][15] = (mid_1[2431:2424] > mid_2[2431:2424]) ? 1 : 0;
assign detect_max[302][16] = (mid_1[2431:2424] > mid_2[2439:2432]) ? 1 : 0;
assign detect_max[302][17] = (mid_1[2431:2424] > btm_0[2423:2416]) ? 1 : 0;
assign detect_max[302][18] = (mid_1[2431:2424] > btm_0[2431:2424]) ? 1 : 0;
assign detect_max[302][19] = (mid_1[2431:2424] > btm_0[2439:2432]) ? 1 : 0;
assign detect_max[302][20] = (mid_1[2431:2424] > btm_1[2423:2416]) ? 1 : 0;
assign detect_max[302][21] = (mid_1[2431:2424] > btm_1[2431:2424]) ? 1 : 0;
assign detect_max[302][22] = (mid_1[2431:2424] > btm_1[2439:2432]) ? 1 : 0;
assign detect_max[302][23] = (mid_1[2431:2424] > btm_2[2423:2416]) ? 1 : 0;
assign detect_max[302][24] = (mid_1[2431:2424] > btm_2[2431:2424]) ? 1 : 0;
assign detect_max[302][25] = (mid_1[2431:2424] > btm_2[2439:2432]) ? 1 : 0;

assign detect_max[303][0] = (mid_1[2439:2432] > top_0[2431:2424]) ? 1 : 0;
assign detect_max[303][1] = (mid_1[2439:2432] > top_0[2439:2432]) ? 1 : 0;
assign detect_max[303][2] = (mid_1[2439:2432] > top_0[2447:2440]) ? 1 : 0;
assign detect_max[303][3] = (mid_1[2439:2432] > top_1[2431:2424]) ? 1 : 0;
assign detect_max[303][4] = (mid_1[2439:2432] > top_1[2439:2432]) ? 1 : 0;
assign detect_max[303][5] = (mid_1[2439:2432] > top_1[2447:2440]) ? 1 : 0;
assign detect_max[303][6] = (mid_1[2439:2432] > top_2[2431:2424]) ? 1 : 0;
assign detect_max[303][7] = (mid_1[2439:2432] > top_2[2439:2432]) ? 1 : 0;
assign detect_max[303][8] = (mid_1[2439:2432] > top_2[2447:2440]) ? 1 : 0;
assign detect_max[303][9] = (mid_1[2439:2432] > mid_0[2431:2424]) ? 1 : 0;
assign detect_max[303][10] = (mid_1[2439:2432] > mid_0[2439:2432]) ? 1 : 0;
assign detect_max[303][11] = (mid_1[2439:2432] > mid_0[2447:2440]) ? 1 : 0;
assign detect_max[303][12] = (mid_1[2439:2432] > mid_1[2431:2424]) ? 1 : 0;
assign detect_max[303][13] = (mid_1[2439:2432] > mid_1[2447:2440]) ? 1 : 0;
assign detect_max[303][14] = (mid_1[2439:2432] > mid_2[2431:2424]) ? 1 : 0;
assign detect_max[303][15] = (mid_1[2439:2432] > mid_2[2439:2432]) ? 1 : 0;
assign detect_max[303][16] = (mid_1[2439:2432] > mid_2[2447:2440]) ? 1 : 0;
assign detect_max[303][17] = (mid_1[2439:2432] > btm_0[2431:2424]) ? 1 : 0;
assign detect_max[303][18] = (mid_1[2439:2432] > btm_0[2439:2432]) ? 1 : 0;
assign detect_max[303][19] = (mid_1[2439:2432] > btm_0[2447:2440]) ? 1 : 0;
assign detect_max[303][20] = (mid_1[2439:2432] > btm_1[2431:2424]) ? 1 : 0;
assign detect_max[303][21] = (mid_1[2439:2432] > btm_1[2439:2432]) ? 1 : 0;
assign detect_max[303][22] = (mid_1[2439:2432] > btm_1[2447:2440]) ? 1 : 0;
assign detect_max[303][23] = (mid_1[2439:2432] > btm_2[2431:2424]) ? 1 : 0;
assign detect_max[303][24] = (mid_1[2439:2432] > btm_2[2439:2432]) ? 1 : 0;
assign detect_max[303][25] = (mid_1[2439:2432] > btm_2[2447:2440]) ? 1 : 0;

assign detect_max[304][0] = (mid_1[2447:2440] > top_0[2439:2432]) ? 1 : 0;
assign detect_max[304][1] = (mid_1[2447:2440] > top_0[2447:2440]) ? 1 : 0;
assign detect_max[304][2] = (mid_1[2447:2440] > top_0[2455:2448]) ? 1 : 0;
assign detect_max[304][3] = (mid_1[2447:2440] > top_1[2439:2432]) ? 1 : 0;
assign detect_max[304][4] = (mid_1[2447:2440] > top_1[2447:2440]) ? 1 : 0;
assign detect_max[304][5] = (mid_1[2447:2440] > top_1[2455:2448]) ? 1 : 0;
assign detect_max[304][6] = (mid_1[2447:2440] > top_2[2439:2432]) ? 1 : 0;
assign detect_max[304][7] = (mid_1[2447:2440] > top_2[2447:2440]) ? 1 : 0;
assign detect_max[304][8] = (mid_1[2447:2440] > top_2[2455:2448]) ? 1 : 0;
assign detect_max[304][9] = (mid_1[2447:2440] > mid_0[2439:2432]) ? 1 : 0;
assign detect_max[304][10] = (mid_1[2447:2440] > mid_0[2447:2440]) ? 1 : 0;
assign detect_max[304][11] = (mid_1[2447:2440] > mid_0[2455:2448]) ? 1 : 0;
assign detect_max[304][12] = (mid_1[2447:2440] > mid_1[2439:2432]) ? 1 : 0;
assign detect_max[304][13] = (mid_1[2447:2440] > mid_1[2455:2448]) ? 1 : 0;
assign detect_max[304][14] = (mid_1[2447:2440] > mid_2[2439:2432]) ? 1 : 0;
assign detect_max[304][15] = (mid_1[2447:2440] > mid_2[2447:2440]) ? 1 : 0;
assign detect_max[304][16] = (mid_1[2447:2440] > mid_2[2455:2448]) ? 1 : 0;
assign detect_max[304][17] = (mid_1[2447:2440] > btm_0[2439:2432]) ? 1 : 0;
assign detect_max[304][18] = (mid_1[2447:2440] > btm_0[2447:2440]) ? 1 : 0;
assign detect_max[304][19] = (mid_1[2447:2440] > btm_0[2455:2448]) ? 1 : 0;
assign detect_max[304][20] = (mid_1[2447:2440] > btm_1[2439:2432]) ? 1 : 0;
assign detect_max[304][21] = (mid_1[2447:2440] > btm_1[2447:2440]) ? 1 : 0;
assign detect_max[304][22] = (mid_1[2447:2440] > btm_1[2455:2448]) ? 1 : 0;
assign detect_max[304][23] = (mid_1[2447:2440] > btm_2[2439:2432]) ? 1 : 0;
assign detect_max[304][24] = (mid_1[2447:2440] > btm_2[2447:2440]) ? 1 : 0;
assign detect_max[304][25] = (mid_1[2447:2440] > btm_2[2455:2448]) ? 1 : 0;

assign detect_max[305][0] = (mid_1[2455:2448] > top_0[2447:2440]) ? 1 : 0;
assign detect_max[305][1] = (mid_1[2455:2448] > top_0[2455:2448]) ? 1 : 0;
assign detect_max[305][2] = (mid_1[2455:2448] > top_0[2463:2456]) ? 1 : 0;
assign detect_max[305][3] = (mid_1[2455:2448] > top_1[2447:2440]) ? 1 : 0;
assign detect_max[305][4] = (mid_1[2455:2448] > top_1[2455:2448]) ? 1 : 0;
assign detect_max[305][5] = (mid_1[2455:2448] > top_1[2463:2456]) ? 1 : 0;
assign detect_max[305][6] = (mid_1[2455:2448] > top_2[2447:2440]) ? 1 : 0;
assign detect_max[305][7] = (mid_1[2455:2448] > top_2[2455:2448]) ? 1 : 0;
assign detect_max[305][8] = (mid_1[2455:2448] > top_2[2463:2456]) ? 1 : 0;
assign detect_max[305][9] = (mid_1[2455:2448] > mid_0[2447:2440]) ? 1 : 0;
assign detect_max[305][10] = (mid_1[2455:2448] > mid_0[2455:2448]) ? 1 : 0;
assign detect_max[305][11] = (mid_1[2455:2448] > mid_0[2463:2456]) ? 1 : 0;
assign detect_max[305][12] = (mid_1[2455:2448] > mid_1[2447:2440]) ? 1 : 0;
assign detect_max[305][13] = (mid_1[2455:2448] > mid_1[2463:2456]) ? 1 : 0;
assign detect_max[305][14] = (mid_1[2455:2448] > mid_2[2447:2440]) ? 1 : 0;
assign detect_max[305][15] = (mid_1[2455:2448] > mid_2[2455:2448]) ? 1 : 0;
assign detect_max[305][16] = (mid_1[2455:2448] > mid_2[2463:2456]) ? 1 : 0;
assign detect_max[305][17] = (mid_1[2455:2448] > btm_0[2447:2440]) ? 1 : 0;
assign detect_max[305][18] = (mid_1[2455:2448] > btm_0[2455:2448]) ? 1 : 0;
assign detect_max[305][19] = (mid_1[2455:2448] > btm_0[2463:2456]) ? 1 : 0;
assign detect_max[305][20] = (mid_1[2455:2448] > btm_1[2447:2440]) ? 1 : 0;
assign detect_max[305][21] = (mid_1[2455:2448] > btm_1[2455:2448]) ? 1 : 0;
assign detect_max[305][22] = (mid_1[2455:2448] > btm_1[2463:2456]) ? 1 : 0;
assign detect_max[305][23] = (mid_1[2455:2448] > btm_2[2447:2440]) ? 1 : 0;
assign detect_max[305][24] = (mid_1[2455:2448] > btm_2[2455:2448]) ? 1 : 0;
assign detect_max[305][25] = (mid_1[2455:2448] > btm_2[2463:2456]) ? 1 : 0;

assign detect_max[306][0] = (mid_1[2463:2456] > top_0[2455:2448]) ? 1 : 0;
assign detect_max[306][1] = (mid_1[2463:2456] > top_0[2463:2456]) ? 1 : 0;
assign detect_max[306][2] = (mid_1[2463:2456] > top_0[2471:2464]) ? 1 : 0;
assign detect_max[306][3] = (mid_1[2463:2456] > top_1[2455:2448]) ? 1 : 0;
assign detect_max[306][4] = (mid_1[2463:2456] > top_1[2463:2456]) ? 1 : 0;
assign detect_max[306][5] = (mid_1[2463:2456] > top_1[2471:2464]) ? 1 : 0;
assign detect_max[306][6] = (mid_1[2463:2456] > top_2[2455:2448]) ? 1 : 0;
assign detect_max[306][7] = (mid_1[2463:2456] > top_2[2463:2456]) ? 1 : 0;
assign detect_max[306][8] = (mid_1[2463:2456] > top_2[2471:2464]) ? 1 : 0;
assign detect_max[306][9] = (mid_1[2463:2456] > mid_0[2455:2448]) ? 1 : 0;
assign detect_max[306][10] = (mid_1[2463:2456] > mid_0[2463:2456]) ? 1 : 0;
assign detect_max[306][11] = (mid_1[2463:2456] > mid_0[2471:2464]) ? 1 : 0;
assign detect_max[306][12] = (mid_1[2463:2456] > mid_1[2455:2448]) ? 1 : 0;
assign detect_max[306][13] = (mid_1[2463:2456] > mid_1[2471:2464]) ? 1 : 0;
assign detect_max[306][14] = (mid_1[2463:2456] > mid_2[2455:2448]) ? 1 : 0;
assign detect_max[306][15] = (mid_1[2463:2456] > mid_2[2463:2456]) ? 1 : 0;
assign detect_max[306][16] = (mid_1[2463:2456] > mid_2[2471:2464]) ? 1 : 0;
assign detect_max[306][17] = (mid_1[2463:2456] > btm_0[2455:2448]) ? 1 : 0;
assign detect_max[306][18] = (mid_1[2463:2456] > btm_0[2463:2456]) ? 1 : 0;
assign detect_max[306][19] = (mid_1[2463:2456] > btm_0[2471:2464]) ? 1 : 0;
assign detect_max[306][20] = (mid_1[2463:2456] > btm_1[2455:2448]) ? 1 : 0;
assign detect_max[306][21] = (mid_1[2463:2456] > btm_1[2463:2456]) ? 1 : 0;
assign detect_max[306][22] = (mid_1[2463:2456] > btm_1[2471:2464]) ? 1 : 0;
assign detect_max[306][23] = (mid_1[2463:2456] > btm_2[2455:2448]) ? 1 : 0;
assign detect_max[306][24] = (mid_1[2463:2456] > btm_2[2463:2456]) ? 1 : 0;
assign detect_max[306][25] = (mid_1[2463:2456] > btm_2[2471:2464]) ? 1 : 0;

assign detect_max[307][0] = (mid_1[2471:2464] > top_0[2463:2456]) ? 1 : 0;
assign detect_max[307][1] = (mid_1[2471:2464] > top_0[2471:2464]) ? 1 : 0;
assign detect_max[307][2] = (mid_1[2471:2464] > top_0[2479:2472]) ? 1 : 0;
assign detect_max[307][3] = (mid_1[2471:2464] > top_1[2463:2456]) ? 1 : 0;
assign detect_max[307][4] = (mid_1[2471:2464] > top_1[2471:2464]) ? 1 : 0;
assign detect_max[307][5] = (mid_1[2471:2464] > top_1[2479:2472]) ? 1 : 0;
assign detect_max[307][6] = (mid_1[2471:2464] > top_2[2463:2456]) ? 1 : 0;
assign detect_max[307][7] = (mid_1[2471:2464] > top_2[2471:2464]) ? 1 : 0;
assign detect_max[307][8] = (mid_1[2471:2464] > top_2[2479:2472]) ? 1 : 0;
assign detect_max[307][9] = (mid_1[2471:2464] > mid_0[2463:2456]) ? 1 : 0;
assign detect_max[307][10] = (mid_1[2471:2464] > mid_0[2471:2464]) ? 1 : 0;
assign detect_max[307][11] = (mid_1[2471:2464] > mid_0[2479:2472]) ? 1 : 0;
assign detect_max[307][12] = (mid_1[2471:2464] > mid_1[2463:2456]) ? 1 : 0;
assign detect_max[307][13] = (mid_1[2471:2464] > mid_1[2479:2472]) ? 1 : 0;
assign detect_max[307][14] = (mid_1[2471:2464] > mid_2[2463:2456]) ? 1 : 0;
assign detect_max[307][15] = (mid_1[2471:2464] > mid_2[2471:2464]) ? 1 : 0;
assign detect_max[307][16] = (mid_1[2471:2464] > mid_2[2479:2472]) ? 1 : 0;
assign detect_max[307][17] = (mid_1[2471:2464] > btm_0[2463:2456]) ? 1 : 0;
assign detect_max[307][18] = (mid_1[2471:2464] > btm_0[2471:2464]) ? 1 : 0;
assign detect_max[307][19] = (mid_1[2471:2464] > btm_0[2479:2472]) ? 1 : 0;
assign detect_max[307][20] = (mid_1[2471:2464] > btm_1[2463:2456]) ? 1 : 0;
assign detect_max[307][21] = (mid_1[2471:2464] > btm_1[2471:2464]) ? 1 : 0;
assign detect_max[307][22] = (mid_1[2471:2464] > btm_1[2479:2472]) ? 1 : 0;
assign detect_max[307][23] = (mid_1[2471:2464] > btm_2[2463:2456]) ? 1 : 0;
assign detect_max[307][24] = (mid_1[2471:2464] > btm_2[2471:2464]) ? 1 : 0;
assign detect_max[307][25] = (mid_1[2471:2464] > btm_2[2479:2472]) ? 1 : 0;

assign detect_max[308][0] = (mid_1[2479:2472] > top_0[2471:2464]) ? 1 : 0;
assign detect_max[308][1] = (mid_1[2479:2472] > top_0[2479:2472]) ? 1 : 0;
assign detect_max[308][2] = (mid_1[2479:2472] > top_0[2487:2480]) ? 1 : 0;
assign detect_max[308][3] = (mid_1[2479:2472] > top_1[2471:2464]) ? 1 : 0;
assign detect_max[308][4] = (mid_1[2479:2472] > top_1[2479:2472]) ? 1 : 0;
assign detect_max[308][5] = (mid_1[2479:2472] > top_1[2487:2480]) ? 1 : 0;
assign detect_max[308][6] = (mid_1[2479:2472] > top_2[2471:2464]) ? 1 : 0;
assign detect_max[308][7] = (mid_1[2479:2472] > top_2[2479:2472]) ? 1 : 0;
assign detect_max[308][8] = (mid_1[2479:2472] > top_2[2487:2480]) ? 1 : 0;
assign detect_max[308][9] = (mid_1[2479:2472] > mid_0[2471:2464]) ? 1 : 0;
assign detect_max[308][10] = (mid_1[2479:2472] > mid_0[2479:2472]) ? 1 : 0;
assign detect_max[308][11] = (mid_1[2479:2472] > mid_0[2487:2480]) ? 1 : 0;
assign detect_max[308][12] = (mid_1[2479:2472] > mid_1[2471:2464]) ? 1 : 0;
assign detect_max[308][13] = (mid_1[2479:2472] > mid_1[2487:2480]) ? 1 : 0;
assign detect_max[308][14] = (mid_1[2479:2472] > mid_2[2471:2464]) ? 1 : 0;
assign detect_max[308][15] = (mid_1[2479:2472] > mid_2[2479:2472]) ? 1 : 0;
assign detect_max[308][16] = (mid_1[2479:2472] > mid_2[2487:2480]) ? 1 : 0;
assign detect_max[308][17] = (mid_1[2479:2472] > btm_0[2471:2464]) ? 1 : 0;
assign detect_max[308][18] = (mid_1[2479:2472] > btm_0[2479:2472]) ? 1 : 0;
assign detect_max[308][19] = (mid_1[2479:2472] > btm_0[2487:2480]) ? 1 : 0;
assign detect_max[308][20] = (mid_1[2479:2472] > btm_1[2471:2464]) ? 1 : 0;
assign detect_max[308][21] = (mid_1[2479:2472] > btm_1[2479:2472]) ? 1 : 0;
assign detect_max[308][22] = (mid_1[2479:2472] > btm_1[2487:2480]) ? 1 : 0;
assign detect_max[308][23] = (mid_1[2479:2472] > btm_2[2471:2464]) ? 1 : 0;
assign detect_max[308][24] = (mid_1[2479:2472] > btm_2[2479:2472]) ? 1 : 0;
assign detect_max[308][25] = (mid_1[2479:2472] > btm_2[2487:2480]) ? 1 : 0;

assign detect_max[309][0] = (mid_1[2487:2480] > top_0[2479:2472]) ? 1 : 0;
assign detect_max[309][1] = (mid_1[2487:2480] > top_0[2487:2480]) ? 1 : 0;
assign detect_max[309][2] = (mid_1[2487:2480] > top_0[2495:2488]) ? 1 : 0;
assign detect_max[309][3] = (mid_1[2487:2480] > top_1[2479:2472]) ? 1 : 0;
assign detect_max[309][4] = (mid_1[2487:2480] > top_1[2487:2480]) ? 1 : 0;
assign detect_max[309][5] = (mid_1[2487:2480] > top_1[2495:2488]) ? 1 : 0;
assign detect_max[309][6] = (mid_1[2487:2480] > top_2[2479:2472]) ? 1 : 0;
assign detect_max[309][7] = (mid_1[2487:2480] > top_2[2487:2480]) ? 1 : 0;
assign detect_max[309][8] = (mid_1[2487:2480] > top_2[2495:2488]) ? 1 : 0;
assign detect_max[309][9] = (mid_1[2487:2480] > mid_0[2479:2472]) ? 1 : 0;
assign detect_max[309][10] = (mid_1[2487:2480] > mid_0[2487:2480]) ? 1 : 0;
assign detect_max[309][11] = (mid_1[2487:2480] > mid_0[2495:2488]) ? 1 : 0;
assign detect_max[309][12] = (mid_1[2487:2480] > mid_1[2479:2472]) ? 1 : 0;
assign detect_max[309][13] = (mid_1[2487:2480] > mid_1[2495:2488]) ? 1 : 0;
assign detect_max[309][14] = (mid_1[2487:2480] > mid_2[2479:2472]) ? 1 : 0;
assign detect_max[309][15] = (mid_1[2487:2480] > mid_2[2487:2480]) ? 1 : 0;
assign detect_max[309][16] = (mid_1[2487:2480] > mid_2[2495:2488]) ? 1 : 0;
assign detect_max[309][17] = (mid_1[2487:2480] > btm_0[2479:2472]) ? 1 : 0;
assign detect_max[309][18] = (mid_1[2487:2480] > btm_0[2487:2480]) ? 1 : 0;
assign detect_max[309][19] = (mid_1[2487:2480] > btm_0[2495:2488]) ? 1 : 0;
assign detect_max[309][20] = (mid_1[2487:2480] > btm_1[2479:2472]) ? 1 : 0;
assign detect_max[309][21] = (mid_1[2487:2480] > btm_1[2487:2480]) ? 1 : 0;
assign detect_max[309][22] = (mid_1[2487:2480] > btm_1[2495:2488]) ? 1 : 0;
assign detect_max[309][23] = (mid_1[2487:2480] > btm_2[2479:2472]) ? 1 : 0;
assign detect_max[309][24] = (mid_1[2487:2480] > btm_2[2487:2480]) ? 1 : 0;
assign detect_max[309][25] = (mid_1[2487:2480] > btm_2[2495:2488]) ? 1 : 0;

assign detect_max[310][0] = (mid_1[2495:2488] > top_0[2487:2480]) ? 1 : 0;
assign detect_max[310][1] = (mid_1[2495:2488] > top_0[2495:2488]) ? 1 : 0;
assign detect_max[310][2] = (mid_1[2495:2488] > top_0[2503:2496]) ? 1 : 0;
assign detect_max[310][3] = (mid_1[2495:2488] > top_1[2487:2480]) ? 1 : 0;
assign detect_max[310][4] = (mid_1[2495:2488] > top_1[2495:2488]) ? 1 : 0;
assign detect_max[310][5] = (mid_1[2495:2488] > top_1[2503:2496]) ? 1 : 0;
assign detect_max[310][6] = (mid_1[2495:2488] > top_2[2487:2480]) ? 1 : 0;
assign detect_max[310][7] = (mid_1[2495:2488] > top_2[2495:2488]) ? 1 : 0;
assign detect_max[310][8] = (mid_1[2495:2488] > top_2[2503:2496]) ? 1 : 0;
assign detect_max[310][9] = (mid_1[2495:2488] > mid_0[2487:2480]) ? 1 : 0;
assign detect_max[310][10] = (mid_1[2495:2488] > mid_0[2495:2488]) ? 1 : 0;
assign detect_max[310][11] = (mid_1[2495:2488] > mid_0[2503:2496]) ? 1 : 0;
assign detect_max[310][12] = (mid_1[2495:2488] > mid_1[2487:2480]) ? 1 : 0;
assign detect_max[310][13] = (mid_1[2495:2488] > mid_1[2503:2496]) ? 1 : 0;
assign detect_max[310][14] = (mid_1[2495:2488] > mid_2[2487:2480]) ? 1 : 0;
assign detect_max[310][15] = (mid_1[2495:2488] > mid_2[2495:2488]) ? 1 : 0;
assign detect_max[310][16] = (mid_1[2495:2488] > mid_2[2503:2496]) ? 1 : 0;
assign detect_max[310][17] = (mid_1[2495:2488] > btm_0[2487:2480]) ? 1 : 0;
assign detect_max[310][18] = (mid_1[2495:2488] > btm_0[2495:2488]) ? 1 : 0;
assign detect_max[310][19] = (mid_1[2495:2488] > btm_0[2503:2496]) ? 1 : 0;
assign detect_max[310][20] = (mid_1[2495:2488] > btm_1[2487:2480]) ? 1 : 0;
assign detect_max[310][21] = (mid_1[2495:2488] > btm_1[2495:2488]) ? 1 : 0;
assign detect_max[310][22] = (mid_1[2495:2488] > btm_1[2503:2496]) ? 1 : 0;
assign detect_max[310][23] = (mid_1[2495:2488] > btm_2[2487:2480]) ? 1 : 0;
assign detect_max[310][24] = (mid_1[2495:2488] > btm_2[2495:2488]) ? 1 : 0;
assign detect_max[310][25] = (mid_1[2495:2488] > btm_2[2503:2496]) ? 1 : 0;

assign detect_max[311][0] = (mid_1[2503:2496] > top_0[2495:2488]) ? 1 : 0;
assign detect_max[311][1] = (mid_1[2503:2496] > top_0[2503:2496]) ? 1 : 0;
assign detect_max[311][2] = (mid_1[2503:2496] > top_0[2511:2504]) ? 1 : 0;
assign detect_max[311][3] = (mid_1[2503:2496] > top_1[2495:2488]) ? 1 : 0;
assign detect_max[311][4] = (mid_1[2503:2496] > top_1[2503:2496]) ? 1 : 0;
assign detect_max[311][5] = (mid_1[2503:2496] > top_1[2511:2504]) ? 1 : 0;
assign detect_max[311][6] = (mid_1[2503:2496] > top_2[2495:2488]) ? 1 : 0;
assign detect_max[311][7] = (mid_1[2503:2496] > top_2[2503:2496]) ? 1 : 0;
assign detect_max[311][8] = (mid_1[2503:2496] > top_2[2511:2504]) ? 1 : 0;
assign detect_max[311][9] = (mid_1[2503:2496] > mid_0[2495:2488]) ? 1 : 0;
assign detect_max[311][10] = (mid_1[2503:2496] > mid_0[2503:2496]) ? 1 : 0;
assign detect_max[311][11] = (mid_1[2503:2496] > mid_0[2511:2504]) ? 1 : 0;
assign detect_max[311][12] = (mid_1[2503:2496] > mid_1[2495:2488]) ? 1 : 0;
assign detect_max[311][13] = (mid_1[2503:2496] > mid_1[2511:2504]) ? 1 : 0;
assign detect_max[311][14] = (mid_1[2503:2496] > mid_2[2495:2488]) ? 1 : 0;
assign detect_max[311][15] = (mid_1[2503:2496] > mid_2[2503:2496]) ? 1 : 0;
assign detect_max[311][16] = (mid_1[2503:2496] > mid_2[2511:2504]) ? 1 : 0;
assign detect_max[311][17] = (mid_1[2503:2496] > btm_0[2495:2488]) ? 1 : 0;
assign detect_max[311][18] = (mid_1[2503:2496] > btm_0[2503:2496]) ? 1 : 0;
assign detect_max[311][19] = (mid_1[2503:2496] > btm_0[2511:2504]) ? 1 : 0;
assign detect_max[311][20] = (mid_1[2503:2496] > btm_1[2495:2488]) ? 1 : 0;
assign detect_max[311][21] = (mid_1[2503:2496] > btm_1[2503:2496]) ? 1 : 0;
assign detect_max[311][22] = (mid_1[2503:2496] > btm_1[2511:2504]) ? 1 : 0;
assign detect_max[311][23] = (mid_1[2503:2496] > btm_2[2495:2488]) ? 1 : 0;
assign detect_max[311][24] = (mid_1[2503:2496] > btm_2[2503:2496]) ? 1 : 0;
assign detect_max[311][25] = (mid_1[2503:2496] > btm_2[2511:2504]) ? 1 : 0;

assign detect_max[312][0] = (mid_1[2511:2504] > top_0[2503:2496]) ? 1 : 0;
assign detect_max[312][1] = (mid_1[2511:2504] > top_0[2511:2504]) ? 1 : 0;
assign detect_max[312][2] = (mid_1[2511:2504] > top_0[2519:2512]) ? 1 : 0;
assign detect_max[312][3] = (mid_1[2511:2504] > top_1[2503:2496]) ? 1 : 0;
assign detect_max[312][4] = (mid_1[2511:2504] > top_1[2511:2504]) ? 1 : 0;
assign detect_max[312][5] = (mid_1[2511:2504] > top_1[2519:2512]) ? 1 : 0;
assign detect_max[312][6] = (mid_1[2511:2504] > top_2[2503:2496]) ? 1 : 0;
assign detect_max[312][7] = (mid_1[2511:2504] > top_2[2511:2504]) ? 1 : 0;
assign detect_max[312][8] = (mid_1[2511:2504] > top_2[2519:2512]) ? 1 : 0;
assign detect_max[312][9] = (mid_1[2511:2504] > mid_0[2503:2496]) ? 1 : 0;
assign detect_max[312][10] = (mid_1[2511:2504] > mid_0[2511:2504]) ? 1 : 0;
assign detect_max[312][11] = (mid_1[2511:2504] > mid_0[2519:2512]) ? 1 : 0;
assign detect_max[312][12] = (mid_1[2511:2504] > mid_1[2503:2496]) ? 1 : 0;
assign detect_max[312][13] = (mid_1[2511:2504] > mid_1[2519:2512]) ? 1 : 0;
assign detect_max[312][14] = (mid_1[2511:2504] > mid_2[2503:2496]) ? 1 : 0;
assign detect_max[312][15] = (mid_1[2511:2504] > mid_2[2511:2504]) ? 1 : 0;
assign detect_max[312][16] = (mid_1[2511:2504] > mid_2[2519:2512]) ? 1 : 0;
assign detect_max[312][17] = (mid_1[2511:2504] > btm_0[2503:2496]) ? 1 : 0;
assign detect_max[312][18] = (mid_1[2511:2504] > btm_0[2511:2504]) ? 1 : 0;
assign detect_max[312][19] = (mid_1[2511:2504] > btm_0[2519:2512]) ? 1 : 0;
assign detect_max[312][20] = (mid_1[2511:2504] > btm_1[2503:2496]) ? 1 : 0;
assign detect_max[312][21] = (mid_1[2511:2504] > btm_1[2511:2504]) ? 1 : 0;
assign detect_max[312][22] = (mid_1[2511:2504] > btm_1[2519:2512]) ? 1 : 0;
assign detect_max[312][23] = (mid_1[2511:2504] > btm_2[2503:2496]) ? 1 : 0;
assign detect_max[312][24] = (mid_1[2511:2504] > btm_2[2511:2504]) ? 1 : 0;
assign detect_max[312][25] = (mid_1[2511:2504] > btm_2[2519:2512]) ? 1 : 0;

assign detect_max[313][0] = (mid_1[2519:2512] > top_0[2511:2504]) ? 1 : 0;
assign detect_max[313][1] = (mid_1[2519:2512] > top_0[2519:2512]) ? 1 : 0;
assign detect_max[313][2] = (mid_1[2519:2512] > top_0[2527:2520]) ? 1 : 0;
assign detect_max[313][3] = (mid_1[2519:2512] > top_1[2511:2504]) ? 1 : 0;
assign detect_max[313][4] = (mid_1[2519:2512] > top_1[2519:2512]) ? 1 : 0;
assign detect_max[313][5] = (mid_1[2519:2512] > top_1[2527:2520]) ? 1 : 0;
assign detect_max[313][6] = (mid_1[2519:2512] > top_2[2511:2504]) ? 1 : 0;
assign detect_max[313][7] = (mid_1[2519:2512] > top_2[2519:2512]) ? 1 : 0;
assign detect_max[313][8] = (mid_1[2519:2512] > top_2[2527:2520]) ? 1 : 0;
assign detect_max[313][9] = (mid_1[2519:2512] > mid_0[2511:2504]) ? 1 : 0;
assign detect_max[313][10] = (mid_1[2519:2512] > mid_0[2519:2512]) ? 1 : 0;
assign detect_max[313][11] = (mid_1[2519:2512] > mid_0[2527:2520]) ? 1 : 0;
assign detect_max[313][12] = (mid_1[2519:2512] > mid_1[2511:2504]) ? 1 : 0;
assign detect_max[313][13] = (mid_1[2519:2512] > mid_1[2527:2520]) ? 1 : 0;
assign detect_max[313][14] = (mid_1[2519:2512] > mid_2[2511:2504]) ? 1 : 0;
assign detect_max[313][15] = (mid_1[2519:2512] > mid_2[2519:2512]) ? 1 : 0;
assign detect_max[313][16] = (mid_1[2519:2512] > mid_2[2527:2520]) ? 1 : 0;
assign detect_max[313][17] = (mid_1[2519:2512] > btm_0[2511:2504]) ? 1 : 0;
assign detect_max[313][18] = (mid_1[2519:2512] > btm_0[2519:2512]) ? 1 : 0;
assign detect_max[313][19] = (mid_1[2519:2512] > btm_0[2527:2520]) ? 1 : 0;
assign detect_max[313][20] = (mid_1[2519:2512] > btm_1[2511:2504]) ? 1 : 0;
assign detect_max[313][21] = (mid_1[2519:2512] > btm_1[2519:2512]) ? 1 : 0;
assign detect_max[313][22] = (mid_1[2519:2512] > btm_1[2527:2520]) ? 1 : 0;
assign detect_max[313][23] = (mid_1[2519:2512] > btm_2[2511:2504]) ? 1 : 0;
assign detect_max[313][24] = (mid_1[2519:2512] > btm_2[2519:2512]) ? 1 : 0;
assign detect_max[313][25] = (mid_1[2519:2512] > btm_2[2527:2520]) ? 1 : 0;

assign detect_max[314][0] = (mid_1[2527:2520] > top_0[2519:2512]) ? 1 : 0;
assign detect_max[314][1] = (mid_1[2527:2520] > top_0[2527:2520]) ? 1 : 0;
assign detect_max[314][2] = (mid_1[2527:2520] > top_0[2535:2528]) ? 1 : 0;
assign detect_max[314][3] = (mid_1[2527:2520] > top_1[2519:2512]) ? 1 : 0;
assign detect_max[314][4] = (mid_1[2527:2520] > top_1[2527:2520]) ? 1 : 0;
assign detect_max[314][5] = (mid_1[2527:2520] > top_1[2535:2528]) ? 1 : 0;
assign detect_max[314][6] = (mid_1[2527:2520] > top_2[2519:2512]) ? 1 : 0;
assign detect_max[314][7] = (mid_1[2527:2520] > top_2[2527:2520]) ? 1 : 0;
assign detect_max[314][8] = (mid_1[2527:2520] > top_2[2535:2528]) ? 1 : 0;
assign detect_max[314][9] = (mid_1[2527:2520] > mid_0[2519:2512]) ? 1 : 0;
assign detect_max[314][10] = (mid_1[2527:2520] > mid_0[2527:2520]) ? 1 : 0;
assign detect_max[314][11] = (mid_1[2527:2520] > mid_0[2535:2528]) ? 1 : 0;
assign detect_max[314][12] = (mid_1[2527:2520] > mid_1[2519:2512]) ? 1 : 0;
assign detect_max[314][13] = (mid_1[2527:2520] > mid_1[2535:2528]) ? 1 : 0;
assign detect_max[314][14] = (mid_1[2527:2520] > mid_2[2519:2512]) ? 1 : 0;
assign detect_max[314][15] = (mid_1[2527:2520] > mid_2[2527:2520]) ? 1 : 0;
assign detect_max[314][16] = (mid_1[2527:2520] > mid_2[2535:2528]) ? 1 : 0;
assign detect_max[314][17] = (mid_1[2527:2520] > btm_0[2519:2512]) ? 1 : 0;
assign detect_max[314][18] = (mid_1[2527:2520] > btm_0[2527:2520]) ? 1 : 0;
assign detect_max[314][19] = (mid_1[2527:2520] > btm_0[2535:2528]) ? 1 : 0;
assign detect_max[314][20] = (mid_1[2527:2520] > btm_1[2519:2512]) ? 1 : 0;
assign detect_max[314][21] = (mid_1[2527:2520] > btm_1[2527:2520]) ? 1 : 0;
assign detect_max[314][22] = (mid_1[2527:2520] > btm_1[2535:2528]) ? 1 : 0;
assign detect_max[314][23] = (mid_1[2527:2520] > btm_2[2519:2512]) ? 1 : 0;
assign detect_max[314][24] = (mid_1[2527:2520] > btm_2[2527:2520]) ? 1 : 0;
assign detect_max[314][25] = (mid_1[2527:2520] > btm_2[2535:2528]) ? 1 : 0;

assign detect_max[315][0] = (mid_1[2535:2528] > top_0[2527:2520]) ? 1 : 0;
assign detect_max[315][1] = (mid_1[2535:2528] > top_0[2535:2528]) ? 1 : 0;
assign detect_max[315][2] = (mid_1[2535:2528] > top_0[2543:2536]) ? 1 : 0;
assign detect_max[315][3] = (mid_1[2535:2528] > top_1[2527:2520]) ? 1 : 0;
assign detect_max[315][4] = (mid_1[2535:2528] > top_1[2535:2528]) ? 1 : 0;
assign detect_max[315][5] = (mid_1[2535:2528] > top_1[2543:2536]) ? 1 : 0;
assign detect_max[315][6] = (mid_1[2535:2528] > top_2[2527:2520]) ? 1 : 0;
assign detect_max[315][7] = (mid_1[2535:2528] > top_2[2535:2528]) ? 1 : 0;
assign detect_max[315][8] = (mid_1[2535:2528] > top_2[2543:2536]) ? 1 : 0;
assign detect_max[315][9] = (mid_1[2535:2528] > mid_0[2527:2520]) ? 1 : 0;
assign detect_max[315][10] = (mid_1[2535:2528] > mid_0[2535:2528]) ? 1 : 0;
assign detect_max[315][11] = (mid_1[2535:2528] > mid_0[2543:2536]) ? 1 : 0;
assign detect_max[315][12] = (mid_1[2535:2528] > mid_1[2527:2520]) ? 1 : 0;
assign detect_max[315][13] = (mid_1[2535:2528] > mid_1[2543:2536]) ? 1 : 0;
assign detect_max[315][14] = (mid_1[2535:2528] > mid_2[2527:2520]) ? 1 : 0;
assign detect_max[315][15] = (mid_1[2535:2528] > mid_2[2535:2528]) ? 1 : 0;
assign detect_max[315][16] = (mid_1[2535:2528] > mid_2[2543:2536]) ? 1 : 0;
assign detect_max[315][17] = (mid_1[2535:2528] > btm_0[2527:2520]) ? 1 : 0;
assign detect_max[315][18] = (mid_1[2535:2528] > btm_0[2535:2528]) ? 1 : 0;
assign detect_max[315][19] = (mid_1[2535:2528] > btm_0[2543:2536]) ? 1 : 0;
assign detect_max[315][20] = (mid_1[2535:2528] > btm_1[2527:2520]) ? 1 : 0;
assign detect_max[315][21] = (mid_1[2535:2528] > btm_1[2535:2528]) ? 1 : 0;
assign detect_max[315][22] = (mid_1[2535:2528] > btm_1[2543:2536]) ? 1 : 0;
assign detect_max[315][23] = (mid_1[2535:2528] > btm_2[2527:2520]) ? 1 : 0;
assign detect_max[315][24] = (mid_1[2535:2528] > btm_2[2535:2528]) ? 1 : 0;
assign detect_max[315][25] = (mid_1[2535:2528] > btm_2[2543:2536]) ? 1 : 0;

assign detect_max[316][0] = (mid_1[2543:2536] > top_0[2535:2528]) ? 1 : 0;
assign detect_max[316][1] = (mid_1[2543:2536] > top_0[2543:2536]) ? 1 : 0;
assign detect_max[316][2] = (mid_1[2543:2536] > top_0[2551:2544]) ? 1 : 0;
assign detect_max[316][3] = (mid_1[2543:2536] > top_1[2535:2528]) ? 1 : 0;
assign detect_max[316][4] = (mid_1[2543:2536] > top_1[2543:2536]) ? 1 : 0;
assign detect_max[316][5] = (mid_1[2543:2536] > top_1[2551:2544]) ? 1 : 0;
assign detect_max[316][6] = (mid_1[2543:2536] > top_2[2535:2528]) ? 1 : 0;
assign detect_max[316][7] = (mid_1[2543:2536] > top_2[2543:2536]) ? 1 : 0;
assign detect_max[316][8] = (mid_1[2543:2536] > top_2[2551:2544]) ? 1 : 0;
assign detect_max[316][9] = (mid_1[2543:2536] > mid_0[2535:2528]) ? 1 : 0;
assign detect_max[316][10] = (mid_1[2543:2536] > mid_0[2543:2536]) ? 1 : 0;
assign detect_max[316][11] = (mid_1[2543:2536] > mid_0[2551:2544]) ? 1 : 0;
assign detect_max[316][12] = (mid_1[2543:2536] > mid_1[2535:2528]) ? 1 : 0;
assign detect_max[316][13] = (mid_1[2543:2536] > mid_1[2551:2544]) ? 1 : 0;
assign detect_max[316][14] = (mid_1[2543:2536] > mid_2[2535:2528]) ? 1 : 0;
assign detect_max[316][15] = (mid_1[2543:2536] > mid_2[2543:2536]) ? 1 : 0;
assign detect_max[316][16] = (mid_1[2543:2536] > mid_2[2551:2544]) ? 1 : 0;
assign detect_max[316][17] = (mid_1[2543:2536] > btm_0[2535:2528]) ? 1 : 0;
assign detect_max[316][18] = (mid_1[2543:2536] > btm_0[2543:2536]) ? 1 : 0;
assign detect_max[316][19] = (mid_1[2543:2536] > btm_0[2551:2544]) ? 1 : 0;
assign detect_max[316][20] = (mid_1[2543:2536] > btm_1[2535:2528]) ? 1 : 0;
assign detect_max[316][21] = (mid_1[2543:2536] > btm_1[2543:2536]) ? 1 : 0;
assign detect_max[316][22] = (mid_1[2543:2536] > btm_1[2551:2544]) ? 1 : 0;
assign detect_max[316][23] = (mid_1[2543:2536] > btm_2[2535:2528]) ? 1 : 0;
assign detect_max[316][24] = (mid_1[2543:2536] > btm_2[2543:2536]) ? 1 : 0;
assign detect_max[316][25] = (mid_1[2543:2536] > btm_2[2551:2544]) ? 1 : 0;

assign detect_max[317][0] = (mid_1[2551:2544] > top_0[2543:2536]) ? 1 : 0;
assign detect_max[317][1] = (mid_1[2551:2544] > top_0[2551:2544]) ? 1 : 0;
assign detect_max[317][2] = (mid_1[2551:2544] > top_0[2559:2552]) ? 1 : 0;
assign detect_max[317][3] = (mid_1[2551:2544] > top_1[2543:2536]) ? 1 : 0;
assign detect_max[317][4] = (mid_1[2551:2544] > top_1[2551:2544]) ? 1 : 0;
assign detect_max[317][5] = (mid_1[2551:2544] > top_1[2559:2552]) ? 1 : 0;
assign detect_max[317][6] = (mid_1[2551:2544] > top_2[2543:2536]) ? 1 : 0;
assign detect_max[317][7] = (mid_1[2551:2544] > top_2[2551:2544]) ? 1 : 0;
assign detect_max[317][8] = (mid_1[2551:2544] > top_2[2559:2552]) ? 1 : 0;
assign detect_max[317][9] = (mid_1[2551:2544] > mid_0[2543:2536]) ? 1 : 0;
assign detect_max[317][10] = (mid_1[2551:2544] > mid_0[2551:2544]) ? 1 : 0;
assign detect_max[317][11] = (mid_1[2551:2544] > mid_0[2559:2552]) ? 1 : 0;
assign detect_max[317][12] = (mid_1[2551:2544] > mid_1[2543:2536]) ? 1 : 0;
assign detect_max[317][13] = (mid_1[2551:2544] > mid_1[2559:2552]) ? 1 : 0;
assign detect_max[317][14] = (mid_1[2551:2544] > mid_2[2543:2536]) ? 1 : 0;
assign detect_max[317][15] = (mid_1[2551:2544] > mid_2[2551:2544]) ? 1 : 0;
assign detect_max[317][16] = (mid_1[2551:2544] > mid_2[2559:2552]) ? 1 : 0;
assign detect_max[317][17] = (mid_1[2551:2544] > btm_0[2543:2536]) ? 1 : 0;
assign detect_max[317][18] = (mid_1[2551:2544] > btm_0[2551:2544]) ? 1 : 0;
assign detect_max[317][19] = (mid_1[2551:2544] > btm_0[2559:2552]) ? 1 : 0;
assign detect_max[317][20] = (mid_1[2551:2544] > btm_1[2543:2536]) ? 1 : 0;
assign detect_max[317][21] = (mid_1[2551:2544] > btm_1[2551:2544]) ? 1 : 0;
assign detect_max[317][22] = (mid_1[2551:2544] > btm_1[2559:2552]) ? 1 : 0;
assign detect_max[317][23] = (mid_1[2551:2544] > btm_2[2543:2536]) ? 1 : 0;
assign detect_max[317][24] = (mid_1[2551:2544] > btm_2[2551:2544]) ? 1 : 0;
assign detect_max[317][25] = (mid_1[2551:2544] > btm_2[2559:2552]) ? 1 : 0;

assign detect_max[318][0] = (mid_1[2559:2552] > top_0[2551:2544]) ? 1 : 0;
assign detect_max[318][1] = (mid_1[2559:2552] > top_0[2559:2552]) ? 1 : 0;
assign detect_max[318][2] = (mid_1[2559:2552] > top_0[2567:2560]) ? 1 : 0;
assign detect_max[318][3] = (mid_1[2559:2552] > top_1[2551:2544]) ? 1 : 0;
assign detect_max[318][4] = (mid_1[2559:2552] > top_1[2559:2552]) ? 1 : 0;
assign detect_max[318][5] = (mid_1[2559:2552] > top_1[2567:2560]) ? 1 : 0;
assign detect_max[318][6] = (mid_1[2559:2552] > top_2[2551:2544]) ? 1 : 0;
assign detect_max[318][7] = (mid_1[2559:2552] > top_2[2559:2552]) ? 1 : 0;
assign detect_max[318][8] = (mid_1[2559:2552] > top_2[2567:2560]) ? 1 : 0;
assign detect_max[318][9] = (mid_1[2559:2552] > mid_0[2551:2544]) ? 1 : 0;
assign detect_max[318][10] = (mid_1[2559:2552] > mid_0[2559:2552]) ? 1 : 0;
assign detect_max[318][11] = (mid_1[2559:2552] > mid_0[2567:2560]) ? 1 : 0;
assign detect_max[318][12] = (mid_1[2559:2552] > mid_1[2551:2544]) ? 1 : 0;
assign detect_max[318][13] = (mid_1[2559:2552] > mid_1[2567:2560]) ? 1 : 0;
assign detect_max[318][14] = (mid_1[2559:2552] > mid_2[2551:2544]) ? 1 : 0;
assign detect_max[318][15] = (mid_1[2559:2552] > mid_2[2559:2552]) ? 1 : 0;
assign detect_max[318][16] = (mid_1[2559:2552] > mid_2[2567:2560]) ? 1 : 0;
assign detect_max[318][17] = (mid_1[2559:2552] > btm_0[2551:2544]) ? 1 : 0;
assign detect_max[318][18] = (mid_1[2559:2552] > btm_0[2559:2552]) ? 1 : 0;
assign detect_max[318][19] = (mid_1[2559:2552] > btm_0[2567:2560]) ? 1 : 0;
assign detect_max[318][20] = (mid_1[2559:2552] > btm_1[2551:2544]) ? 1 : 0;
assign detect_max[318][21] = (mid_1[2559:2552] > btm_1[2559:2552]) ? 1 : 0;
assign detect_max[318][22] = (mid_1[2559:2552] > btm_1[2567:2560]) ? 1 : 0;
assign detect_max[318][23] = (mid_1[2559:2552] > btm_2[2551:2544]) ? 1 : 0;
assign detect_max[318][24] = (mid_1[2559:2552] > btm_2[2559:2552]) ? 1 : 0;
assign detect_max[318][25] = (mid_1[2559:2552] > btm_2[2567:2560]) ? 1 : 0;

assign detect_max[319][0] = (mid_1[2567:2560] > top_0[2559:2552]) ? 1 : 0;
assign detect_max[319][1] = (mid_1[2567:2560] > top_0[2567:2560]) ? 1 : 0;
assign detect_max[319][2] = (mid_1[2567:2560] > top_0[2575:2568]) ? 1 : 0;
assign detect_max[319][3] = (mid_1[2567:2560] > top_1[2559:2552]) ? 1 : 0;
assign detect_max[319][4] = (mid_1[2567:2560] > top_1[2567:2560]) ? 1 : 0;
assign detect_max[319][5] = (mid_1[2567:2560] > top_1[2575:2568]) ? 1 : 0;
assign detect_max[319][6] = (mid_1[2567:2560] > top_2[2559:2552]) ? 1 : 0;
assign detect_max[319][7] = (mid_1[2567:2560] > top_2[2567:2560]) ? 1 : 0;
assign detect_max[319][8] = (mid_1[2567:2560] > top_2[2575:2568]) ? 1 : 0;
assign detect_max[319][9] = (mid_1[2567:2560] > mid_0[2559:2552]) ? 1 : 0;
assign detect_max[319][10] = (mid_1[2567:2560] > mid_0[2567:2560]) ? 1 : 0;
assign detect_max[319][11] = (mid_1[2567:2560] > mid_0[2575:2568]) ? 1 : 0;
assign detect_max[319][12] = (mid_1[2567:2560] > mid_1[2559:2552]) ? 1 : 0;
assign detect_max[319][13] = (mid_1[2567:2560] > mid_1[2575:2568]) ? 1 : 0;
assign detect_max[319][14] = (mid_1[2567:2560] > mid_2[2559:2552]) ? 1 : 0;
assign detect_max[319][15] = (mid_1[2567:2560] > mid_2[2567:2560]) ? 1 : 0;
assign detect_max[319][16] = (mid_1[2567:2560] > mid_2[2575:2568]) ? 1 : 0;
assign detect_max[319][17] = (mid_1[2567:2560] > btm_0[2559:2552]) ? 1 : 0;
assign detect_max[319][18] = (mid_1[2567:2560] > btm_0[2567:2560]) ? 1 : 0;
assign detect_max[319][19] = (mid_1[2567:2560] > btm_0[2575:2568]) ? 1 : 0;
assign detect_max[319][20] = (mid_1[2567:2560] > btm_1[2559:2552]) ? 1 : 0;
assign detect_max[319][21] = (mid_1[2567:2560] > btm_1[2567:2560]) ? 1 : 0;
assign detect_max[319][22] = (mid_1[2567:2560] > btm_1[2575:2568]) ? 1 : 0;
assign detect_max[319][23] = (mid_1[2567:2560] > btm_2[2559:2552]) ? 1 : 0;
assign detect_max[319][24] = (mid_1[2567:2560] > btm_2[2567:2560]) ? 1 : 0;
assign detect_max[319][25] = (mid_1[2567:2560] > btm_2[2575:2568]) ? 1 : 0;

assign detect_max[320][0] = (mid_1[2575:2568] > top_0[2567:2560]) ? 1 : 0;
assign detect_max[320][1] = (mid_1[2575:2568] > top_0[2575:2568]) ? 1 : 0;
assign detect_max[320][2] = (mid_1[2575:2568] > top_0[2583:2576]) ? 1 : 0;
assign detect_max[320][3] = (mid_1[2575:2568] > top_1[2567:2560]) ? 1 : 0;
assign detect_max[320][4] = (mid_1[2575:2568] > top_1[2575:2568]) ? 1 : 0;
assign detect_max[320][5] = (mid_1[2575:2568] > top_1[2583:2576]) ? 1 : 0;
assign detect_max[320][6] = (mid_1[2575:2568] > top_2[2567:2560]) ? 1 : 0;
assign detect_max[320][7] = (mid_1[2575:2568] > top_2[2575:2568]) ? 1 : 0;
assign detect_max[320][8] = (mid_1[2575:2568] > top_2[2583:2576]) ? 1 : 0;
assign detect_max[320][9] = (mid_1[2575:2568] > mid_0[2567:2560]) ? 1 : 0;
assign detect_max[320][10] = (mid_1[2575:2568] > mid_0[2575:2568]) ? 1 : 0;
assign detect_max[320][11] = (mid_1[2575:2568] > mid_0[2583:2576]) ? 1 : 0;
assign detect_max[320][12] = (mid_1[2575:2568] > mid_1[2567:2560]) ? 1 : 0;
assign detect_max[320][13] = (mid_1[2575:2568] > mid_1[2583:2576]) ? 1 : 0;
assign detect_max[320][14] = (mid_1[2575:2568] > mid_2[2567:2560]) ? 1 : 0;
assign detect_max[320][15] = (mid_1[2575:2568] > mid_2[2575:2568]) ? 1 : 0;
assign detect_max[320][16] = (mid_1[2575:2568] > mid_2[2583:2576]) ? 1 : 0;
assign detect_max[320][17] = (mid_1[2575:2568] > btm_0[2567:2560]) ? 1 : 0;
assign detect_max[320][18] = (mid_1[2575:2568] > btm_0[2575:2568]) ? 1 : 0;
assign detect_max[320][19] = (mid_1[2575:2568] > btm_0[2583:2576]) ? 1 : 0;
assign detect_max[320][20] = (mid_1[2575:2568] > btm_1[2567:2560]) ? 1 : 0;
assign detect_max[320][21] = (mid_1[2575:2568] > btm_1[2575:2568]) ? 1 : 0;
assign detect_max[320][22] = (mid_1[2575:2568] > btm_1[2583:2576]) ? 1 : 0;
assign detect_max[320][23] = (mid_1[2575:2568] > btm_2[2567:2560]) ? 1 : 0;
assign detect_max[320][24] = (mid_1[2575:2568] > btm_2[2575:2568]) ? 1 : 0;
assign detect_max[320][25] = (mid_1[2575:2568] > btm_2[2583:2576]) ? 1 : 0;

assign detect_max[321][0] = (mid_1[2583:2576] > top_0[2575:2568]) ? 1 : 0;
assign detect_max[321][1] = (mid_1[2583:2576] > top_0[2583:2576]) ? 1 : 0;
assign detect_max[321][2] = (mid_1[2583:2576] > top_0[2591:2584]) ? 1 : 0;
assign detect_max[321][3] = (mid_1[2583:2576] > top_1[2575:2568]) ? 1 : 0;
assign detect_max[321][4] = (mid_1[2583:2576] > top_1[2583:2576]) ? 1 : 0;
assign detect_max[321][5] = (mid_1[2583:2576] > top_1[2591:2584]) ? 1 : 0;
assign detect_max[321][6] = (mid_1[2583:2576] > top_2[2575:2568]) ? 1 : 0;
assign detect_max[321][7] = (mid_1[2583:2576] > top_2[2583:2576]) ? 1 : 0;
assign detect_max[321][8] = (mid_1[2583:2576] > top_2[2591:2584]) ? 1 : 0;
assign detect_max[321][9] = (mid_1[2583:2576] > mid_0[2575:2568]) ? 1 : 0;
assign detect_max[321][10] = (mid_1[2583:2576] > mid_0[2583:2576]) ? 1 : 0;
assign detect_max[321][11] = (mid_1[2583:2576] > mid_0[2591:2584]) ? 1 : 0;
assign detect_max[321][12] = (mid_1[2583:2576] > mid_1[2575:2568]) ? 1 : 0;
assign detect_max[321][13] = (mid_1[2583:2576] > mid_1[2591:2584]) ? 1 : 0;
assign detect_max[321][14] = (mid_1[2583:2576] > mid_2[2575:2568]) ? 1 : 0;
assign detect_max[321][15] = (mid_1[2583:2576] > mid_2[2583:2576]) ? 1 : 0;
assign detect_max[321][16] = (mid_1[2583:2576] > mid_2[2591:2584]) ? 1 : 0;
assign detect_max[321][17] = (mid_1[2583:2576] > btm_0[2575:2568]) ? 1 : 0;
assign detect_max[321][18] = (mid_1[2583:2576] > btm_0[2583:2576]) ? 1 : 0;
assign detect_max[321][19] = (mid_1[2583:2576] > btm_0[2591:2584]) ? 1 : 0;
assign detect_max[321][20] = (mid_1[2583:2576] > btm_1[2575:2568]) ? 1 : 0;
assign detect_max[321][21] = (mid_1[2583:2576] > btm_1[2583:2576]) ? 1 : 0;
assign detect_max[321][22] = (mid_1[2583:2576] > btm_1[2591:2584]) ? 1 : 0;
assign detect_max[321][23] = (mid_1[2583:2576] > btm_2[2575:2568]) ? 1 : 0;
assign detect_max[321][24] = (mid_1[2583:2576] > btm_2[2583:2576]) ? 1 : 0;
assign detect_max[321][25] = (mid_1[2583:2576] > btm_2[2591:2584]) ? 1 : 0;

assign detect_max[322][0] = (mid_1[2591:2584] > top_0[2583:2576]) ? 1 : 0;
assign detect_max[322][1] = (mid_1[2591:2584] > top_0[2591:2584]) ? 1 : 0;
assign detect_max[322][2] = (mid_1[2591:2584] > top_0[2599:2592]) ? 1 : 0;
assign detect_max[322][3] = (mid_1[2591:2584] > top_1[2583:2576]) ? 1 : 0;
assign detect_max[322][4] = (mid_1[2591:2584] > top_1[2591:2584]) ? 1 : 0;
assign detect_max[322][5] = (mid_1[2591:2584] > top_1[2599:2592]) ? 1 : 0;
assign detect_max[322][6] = (mid_1[2591:2584] > top_2[2583:2576]) ? 1 : 0;
assign detect_max[322][7] = (mid_1[2591:2584] > top_2[2591:2584]) ? 1 : 0;
assign detect_max[322][8] = (mid_1[2591:2584] > top_2[2599:2592]) ? 1 : 0;
assign detect_max[322][9] = (mid_1[2591:2584] > mid_0[2583:2576]) ? 1 : 0;
assign detect_max[322][10] = (mid_1[2591:2584] > mid_0[2591:2584]) ? 1 : 0;
assign detect_max[322][11] = (mid_1[2591:2584] > mid_0[2599:2592]) ? 1 : 0;
assign detect_max[322][12] = (mid_1[2591:2584] > mid_1[2583:2576]) ? 1 : 0;
assign detect_max[322][13] = (mid_1[2591:2584] > mid_1[2599:2592]) ? 1 : 0;
assign detect_max[322][14] = (mid_1[2591:2584] > mid_2[2583:2576]) ? 1 : 0;
assign detect_max[322][15] = (mid_1[2591:2584] > mid_2[2591:2584]) ? 1 : 0;
assign detect_max[322][16] = (mid_1[2591:2584] > mid_2[2599:2592]) ? 1 : 0;
assign detect_max[322][17] = (mid_1[2591:2584] > btm_0[2583:2576]) ? 1 : 0;
assign detect_max[322][18] = (mid_1[2591:2584] > btm_0[2591:2584]) ? 1 : 0;
assign detect_max[322][19] = (mid_1[2591:2584] > btm_0[2599:2592]) ? 1 : 0;
assign detect_max[322][20] = (mid_1[2591:2584] > btm_1[2583:2576]) ? 1 : 0;
assign detect_max[322][21] = (mid_1[2591:2584] > btm_1[2591:2584]) ? 1 : 0;
assign detect_max[322][22] = (mid_1[2591:2584] > btm_1[2599:2592]) ? 1 : 0;
assign detect_max[322][23] = (mid_1[2591:2584] > btm_2[2583:2576]) ? 1 : 0;
assign detect_max[322][24] = (mid_1[2591:2584] > btm_2[2591:2584]) ? 1 : 0;
assign detect_max[322][25] = (mid_1[2591:2584] > btm_2[2599:2592]) ? 1 : 0;

assign detect_max[323][0] = (mid_1[2599:2592] > top_0[2591:2584]) ? 1 : 0;
assign detect_max[323][1] = (mid_1[2599:2592] > top_0[2599:2592]) ? 1 : 0;
assign detect_max[323][2] = (mid_1[2599:2592] > top_0[2607:2600]) ? 1 : 0;
assign detect_max[323][3] = (mid_1[2599:2592] > top_1[2591:2584]) ? 1 : 0;
assign detect_max[323][4] = (mid_1[2599:2592] > top_1[2599:2592]) ? 1 : 0;
assign detect_max[323][5] = (mid_1[2599:2592] > top_1[2607:2600]) ? 1 : 0;
assign detect_max[323][6] = (mid_1[2599:2592] > top_2[2591:2584]) ? 1 : 0;
assign detect_max[323][7] = (mid_1[2599:2592] > top_2[2599:2592]) ? 1 : 0;
assign detect_max[323][8] = (mid_1[2599:2592] > top_2[2607:2600]) ? 1 : 0;
assign detect_max[323][9] = (mid_1[2599:2592] > mid_0[2591:2584]) ? 1 : 0;
assign detect_max[323][10] = (mid_1[2599:2592] > mid_0[2599:2592]) ? 1 : 0;
assign detect_max[323][11] = (mid_1[2599:2592] > mid_0[2607:2600]) ? 1 : 0;
assign detect_max[323][12] = (mid_1[2599:2592] > mid_1[2591:2584]) ? 1 : 0;
assign detect_max[323][13] = (mid_1[2599:2592] > mid_1[2607:2600]) ? 1 : 0;
assign detect_max[323][14] = (mid_1[2599:2592] > mid_2[2591:2584]) ? 1 : 0;
assign detect_max[323][15] = (mid_1[2599:2592] > mid_2[2599:2592]) ? 1 : 0;
assign detect_max[323][16] = (mid_1[2599:2592] > mid_2[2607:2600]) ? 1 : 0;
assign detect_max[323][17] = (mid_1[2599:2592] > btm_0[2591:2584]) ? 1 : 0;
assign detect_max[323][18] = (mid_1[2599:2592] > btm_0[2599:2592]) ? 1 : 0;
assign detect_max[323][19] = (mid_1[2599:2592] > btm_0[2607:2600]) ? 1 : 0;
assign detect_max[323][20] = (mid_1[2599:2592] > btm_1[2591:2584]) ? 1 : 0;
assign detect_max[323][21] = (mid_1[2599:2592] > btm_1[2599:2592]) ? 1 : 0;
assign detect_max[323][22] = (mid_1[2599:2592] > btm_1[2607:2600]) ? 1 : 0;
assign detect_max[323][23] = (mid_1[2599:2592] > btm_2[2591:2584]) ? 1 : 0;
assign detect_max[323][24] = (mid_1[2599:2592] > btm_2[2599:2592]) ? 1 : 0;
assign detect_max[323][25] = (mid_1[2599:2592] > btm_2[2607:2600]) ? 1 : 0;

assign detect_max[324][0] = (mid_1[2607:2600] > top_0[2599:2592]) ? 1 : 0;
assign detect_max[324][1] = (mid_1[2607:2600] > top_0[2607:2600]) ? 1 : 0;
assign detect_max[324][2] = (mid_1[2607:2600] > top_0[2615:2608]) ? 1 : 0;
assign detect_max[324][3] = (mid_1[2607:2600] > top_1[2599:2592]) ? 1 : 0;
assign detect_max[324][4] = (mid_1[2607:2600] > top_1[2607:2600]) ? 1 : 0;
assign detect_max[324][5] = (mid_1[2607:2600] > top_1[2615:2608]) ? 1 : 0;
assign detect_max[324][6] = (mid_1[2607:2600] > top_2[2599:2592]) ? 1 : 0;
assign detect_max[324][7] = (mid_1[2607:2600] > top_2[2607:2600]) ? 1 : 0;
assign detect_max[324][8] = (mid_1[2607:2600] > top_2[2615:2608]) ? 1 : 0;
assign detect_max[324][9] = (mid_1[2607:2600] > mid_0[2599:2592]) ? 1 : 0;
assign detect_max[324][10] = (mid_1[2607:2600] > mid_0[2607:2600]) ? 1 : 0;
assign detect_max[324][11] = (mid_1[2607:2600] > mid_0[2615:2608]) ? 1 : 0;
assign detect_max[324][12] = (mid_1[2607:2600] > mid_1[2599:2592]) ? 1 : 0;
assign detect_max[324][13] = (mid_1[2607:2600] > mid_1[2615:2608]) ? 1 : 0;
assign detect_max[324][14] = (mid_1[2607:2600] > mid_2[2599:2592]) ? 1 : 0;
assign detect_max[324][15] = (mid_1[2607:2600] > mid_2[2607:2600]) ? 1 : 0;
assign detect_max[324][16] = (mid_1[2607:2600] > mid_2[2615:2608]) ? 1 : 0;
assign detect_max[324][17] = (mid_1[2607:2600] > btm_0[2599:2592]) ? 1 : 0;
assign detect_max[324][18] = (mid_1[2607:2600] > btm_0[2607:2600]) ? 1 : 0;
assign detect_max[324][19] = (mid_1[2607:2600] > btm_0[2615:2608]) ? 1 : 0;
assign detect_max[324][20] = (mid_1[2607:2600] > btm_1[2599:2592]) ? 1 : 0;
assign detect_max[324][21] = (mid_1[2607:2600] > btm_1[2607:2600]) ? 1 : 0;
assign detect_max[324][22] = (mid_1[2607:2600] > btm_1[2615:2608]) ? 1 : 0;
assign detect_max[324][23] = (mid_1[2607:2600] > btm_2[2599:2592]) ? 1 : 0;
assign detect_max[324][24] = (mid_1[2607:2600] > btm_2[2607:2600]) ? 1 : 0;
assign detect_max[324][25] = (mid_1[2607:2600] > btm_2[2615:2608]) ? 1 : 0;

assign detect_max[325][0] = (mid_1[2615:2608] > top_0[2607:2600]) ? 1 : 0;
assign detect_max[325][1] = (mid_1[2615:2608] > top_0[2615:2608]) ? 1 : 0;
assign detect_max[325][2] = (mid_1[2615:2608] > top_0[2623:2616]) ? 1 : 0;
assign detect_max[325][3] = (mid_1[2615:2608] > top_1[2607:2600]) ? 1 : 0;
assign detect_max[325][4] = (mid_1[2615:2608] > top_1[2615:2608]) ? 1 : 0;
assign detect_max[325][5] = (mid_1[2615:2608] > top_1[2623:2616]) ? 1 : 0;
assign detect_max[325][6] = (mid_1[2615:2608] > top_2[2607:2600]) ? 1 : 0;
assign detect_max[325][7] = (mid_1[2615:2608] > top_2[2615:2608]) ? 1 : 0;
assign detect_max[325][8] = (mid_1[2615:2608] > top_2[2623:2616]) ? 1 : 0;
assign detect_max[325][9] = (mid_1[2615:2608] > mid_0[2607:2600]) ? 1 : 0;
assign detect_max[325][10] = (mid_1[2615:2608] > mid_0[2615:2608]) ? 1 : 0;
assign detect_max[325][11] = (mid_1[2615:2608] > mid_0[2623:2616]) ? 1 : 0;
assign detect_max[325][12] = (mid_1[2615:2608] > mid_1[2607:2600]) ? 1 : 0;
assign detect_max[325][13] = (mid_1[2615:2608] > mid_1[2623:2616]) ? 1 : 0;
assign detect_max[325][14] = (mid_1[2615:2608] > mid_2[2607:2600]) ? 1 : 0;
assign detect_max[325][15] = (mid_1[2615:2608] > mid_2[2615:2608]) ? 1 : 0;
assign detect_max[325][16] = (mid_1[2615:2608] > mid_2[2623:2616]) ? 1 : 0;
assign detect_max[325][17] = (mid_1[2615:2608] > btm_0[2607:2600]) ? 1 : 0;
assign detect_max[325][18] = (mid_1[2615:2608] > btm_0[2615:2608]) ? 1 : 0;
assign detect_max[325][19] = (mid_1[2615:2608] > btm_0[2623:2616]) ? 1 : 0;
assign detect_max[325][20] = (mid_1[2615:2608] > btm_1[2607:2600]) ? 1 : 0;
assign detect_max[325][21] = (mid_1[2615:2608] > btm_1[2615:2608]) ? 1 : 0;
assign detect_max[325][22] = (mid_1[2615:2608] > btm_1[2623:2616]) ? 1 : 0;
assign detect_max[325][23] = (mid_1[2615:2608] > btm_2[2607:2600]) ? 1 : 0;
assign detect_max[325][24] = (mid_1[2615:2608] > btm_2[2615:2608]) ? 1 : 0;
assign detect_max[325][25] = (mid_1[2615:2608] > btm_2[2623:2616]) ? 1 : 0;

assign detect_max[326][0] = (mid_1[2623:2616] > top_0[2615:2608]) ? 1 : 0;
assign detect_max[326][1] = (mid_1[2623:2616] > top_0[2623:2616]) ? 1 : 0;
assign detect_max[326][2] = (mid_1[2623:2616] > top_0[2631:2624]) ? 1 : 0;
assign detect_max[326][3] = (mid_1[2623:2616] > top_1[2615:2608]) ? 1 : 0;
assign detect_max[326][4] = (mid_1[2623:2616] > top_1[2623:2616]) ? 1 : 0;
assign detect_max[326][5] = (mid_1[2623:2616] > top_1[2631:2624]) ? 1 : 0;
assign detect_max[326][6] = (mid_1[2623:2616] > top_2[2615:2608]) ? 1 : 0;
assign detect_max[326][7] = (mid_1[2623:2616] > top_2[2623:2616]) ? 1 : 0;
assign detect_max[326][8] = (mid_1[2623:2616] > top_2[2631:2624]) ? 1 : 0;
assign detect_max[326][9] = (mid_1[2623:2616] > mid_0[2615:2608]) ? 1 : 0;
assign detect_max[326][10] = (mid_1[2623:2616] > mid_0[2623:2616]) ? 1 : 0;
assign detect_max[326][11] = (mid_1[2623:2616] > mid_0[2631:2624]) ? 1 : 0;
assign detect_max[326][12] = (mid_1[2623:2616] > mid_1[2615:2608]) ? 1 : 0;
assign detect_max[326][13] = (mid_1[2623:2616] > mid_1[2631:2624]) ? 1 : 0;
assign detect_max[326][14] = (mid_1[2623:2616] > mid_2[2615:2608]) ? 1 : 0;
assign detect_max[326][15] = (mid_1[2623:2616] > mid_2[2623:2616]) ? 1 : 0;
assign detect_max[326][16] = (mid_1[2623:2616] > mid_2[2631:2624]) ? 1 : 0;
assign detect_max[326][17] = (mid_1[2623:2616] > btm_0[2615:2608]) ? 1 : 0;
assign detect_max[326][18] = (mid_1[2623:2616] > btm_0[2623:2616]) ? 1 : 0;
assign detect_max[326][19] = (mid_1[2623:2616] > btm_0[2631:2624]) ? 1 : 0;
assign detect_max[326][20] = (mid_1[2623:2616] > btm_1[2615:2608]) ? 1 : 0;
assign detect_max[326][21] = (mid_1[2623:2616] > btm_1[2623:2616]) ? 1 : 0;
assign detect_max[326][22] = (mid_1[2623:2616] > btm_1[2631:2624]) ? 1 : 0;
assign detect_max[326][23] = (mid_1[2623:2616] > btm_2[2615:2608]) ? 1 : 0;
assign detect_max[326][24] = (mid_1[2623:2616] > btm_2[2623:2616]) ? 1 : 0;
assign detect_max[326][25] = (mid_1[2623:2616] > btm_2[2631:2624]) ? 1 : 0;

assign detect_max[327][0] = (mid_1[2631:2624] > top_0[2623:2616]) ? 1 : 0;
assign detect_max[327][1] = (mid_1[2631:2624] > top_0[2631:2624]) ? 1 : 0;
assign detect_max[327][2] = (mid_1[2631:2624] > top_0[2639:2632]) ? 1 : 0;
assign detect_max[327][3] = (mid_1[2631:2624] > top_1[2623:2616]) ? 1 : 0;
assign detect_max[327][4] = (mid_1[2631:2624] > top_1[2631:2624]) ? 1 : 0;
assign detect_max[327][5] = (mid_1[2631:2624] > top_1[2639:2632]) ? 1 : 0;
assign detect_max[327][6] = (mid_1[2631:2624] > top_2[2623:2616]) ? 1 : 0;
assign detect_max[327][7] = (mid_1[2631:2624] > top_2[2631:2624]) ? 1 : 0;
assign detect_max[327][8] = (mid_1[2631:2624] > top_2[2639:2632]) ? 1 : 0;
assign detect_max[327][9] = (mid_1[2631:2624] > mid_0[2623:2616]) ? 1 : 0;
assign detect_max[327][10] = (mid_1[2631:2624] > mid_0[2631:2624]) ? 1 : 0;
assign detect_max[327][11] = (mid_1[2631:2624] > mid_0[2639:2632]) ? 1 : 0;
assign detect_max[327][12] = (mid_1[2631:2624] > mid_1[2623:2616]) ? 1 : 0;
assign detect_max[327][13] = (mid_1[2631:2624] > mid_1[2639:2632]) ? 1 : 0;
assign detect_max[327][14] = (mid_1[2631:2624] > mid_2[2623:2616]) ? 1 : 0;
assign detect_max[327][15] = (mid_1[2631:2624] > mid_2[2631:2624]) ? 1 : 0;
assign detect_max[327][16] = (mid_1[2631:2624] > mid_2[2639:2632]) ? 1 : 0;
assign detect_max[327][17] = (mid_1[2631:2624] > btm_0[2623:2616]) ? 1 : 0;
assign detect_max[327][18] = (mid_1[2631:2624] > btm_0[2631:2624]) ? 1 : 0;
assign detect_max[327][19] = (mid_1[2631:2624] > btm_0[2639:2632]) ? 1 : 0;
assign detect_max[327][20] = (mid_1[2631:2624] > btm_1[2623:2616]) ? 1 : 0;
assign detect_max[327][21] = (mid_1[2631:2624] > btm_1[2631:2624]) ? 1 : 0;
assign detect_max[327][22] = (mid_1[2631:2624] > btm_1[2639:2632]) ? 1 : 0;
assign detect_max[327][23] = (mid_1[2631:2624] > btm_2[2623:2616]) ? 1 : 0;
assign detect_max[327][24] = (mid_1[2631:2624] > btm_2[2631:2624]) ? 1 : 0;
assign detect_max[327][25] = (mid_1[2631:2624] > btm_2[2639:2632]) ? 1 : 0;

assign detect_max[328][0] = (mid_1[2639:2632] > top_0[2631:2624]) ? 1 : 0;
assign detect_max[328][1] = (mid_1[2639:2632] > top_0[2639:2632]) ? 1 : 0;
assign detect_max[328][2] = (mid_1[2639:2632] > top_0[2647:2640]) ? 1 : 0;
assign detect_max[328][3] = (mid_1[2639:2632] > top_1[2631:2624]) ? 1 : 0;
assign detect_max[328][4] = (mid_1[2639:2632] > top_1[2639:2632]) ? 1 : 0;
assign detect_max[328][5] = (mid_1[2639:2632] > top_1[2647:2640]) ? 1 : 0;
assign detect_max[328][6] = (mid_1[2639:2632] > top_2[2631:2624]) ? 1 : 0;
assign detect_max[328][7] = (mid_1[2639:2632] > top_2[2639:2632]) ? 1 : 0;
assign detect_max[328][8] = (mid_1[2639:2632] > top_2[2647:2640]) ? 1 : 0;
assign detect_max[328][9] = (mid_1[2639:2632] > mid_0[2631:2624]) ? 1 : 0;
assign detect_max[328][10] = (mid_1[2639:2632] > mid_0[2639:2632]) ? 1 : 0;
assign detect_max[328][11] = (mid_1[2639:2632] > mid_0[2647:2640]) ? 1 : 0;
assign detect_max[328][12] = (mid_1[2639:2632] > mid_1[2631:2624]) ? 1 : 0;
assign detect_max[328][13] = (mid_1[2639:2632] > mid_1[2647:2640]) ? 1 : 0;
assign detect_max[328][14] = (mid_1[2639:2632] > mid_2[2631:2624]) ? 1 : 0;
assign detect_max[328][15] = (mid_1[2639:2632] > mid_2[2639:2632]) ? 1 : 0;
assign detect_max[328][16] = (mid_1[2639:2632] > mid_2[2647:2640]) ? 1 : 0;
assign detect_max[328][17] = (mid_1[2639:2632] > btm_0[2631:2624]) ? 1 : 0;
assign detect_max[328][18] = (mid_1[2639:2632] > btm_0[2639:2632]) ? 1 : 0;
assign detect_max[328][19] = (mid_1[2639:2632] > btm_0[2647:2640]) ? 1 : 0;
assign detect_max[328][20] = (mid_1[2639:2632] > btm_1[2631:2624]) ? 1 : 0;
assign detect_max[328][21] = (mid_1[2639:2632] > btm_1[2639:2632]) ? 1 : 0;
assign detect_max[328][22] = (mid_1[2639:2632] > btm_1[2647:2640]) ? 1 : 0;
assign detect_max[328][23] = (mid_1[2639:2632] > btm_2[2631:2624]) ? 1 : 0;
assign detect_max[328][24] = (mid_1[2639:2632] > btm_2[2639:2632]) ? 1 : 0;
assign detect_max[328][25] = (mid_1[2639:2632] > btm_2[2647:2640]) ? 1 : 0;

assign detect_max[329][0] = (mid_1[2647:2640] > top_0[2639:2632]) ? 1 : 0;
assign detect_max[329][1] = (mid_1[2647:2640] > top_0[2647:2640]) ? 1 : 0;
assign detect_max[329][2] = (mid_1[2647:2640] > top_0[2655:2648]) ? 1 : 0;
assign detect_max[329][3] = (mid_1[2647:2640] > top_1[2639:2632]) ? 1 : 0;
assign detect_max[329][4] = (mid_1[2647:2640] > top_1[2647:2640]) ? 1 : 0;
assign detect_max[329][5] = (mid_1[2647:2640] > top_1[2655:2648]) ? 1 : 0;
assign detect_max[329][6] = (mid_1[2647:2640] > top_2[2639:2632]) ? 1 : 0;
assign detect_max[329][7] = (mid_1[2647:2640] > top_2[2647:2640]) ? 1 : 0;
assign detect_max[329][8] = (mid_1[2647:2640] > top_2[2655:2648]) ? 1 : 0;
assign detect_max[329][9] = (mid_1[2647:2640] > mid_0[2639:2632]) ? 1 : 0;
assign detect_max[329][10] = (mid_1[2647:2640] > mid_0[2647:2640]) ? 1 : 0;
assign detect_max[329][11] = (mid_1[2647:2640] > mid_0[2655:2648]) ? 1 : 0;
assign detect_max[329][12] = (mid_1[2647:2640] > mid_1[2639:2632]) ? 1 : 0;
assign detect_max[329][13] = (mid_1[2647:2640] > mid_1[2655:2648]) ? 1 : 0;
assign detect_max[329][14] = (mid_1[2647:2640] > mid_2[2639:2632]) ? 1 : 0;
assign detect_max[329][15] = (mid_1[2647:2640] > mid_2[2647:2640]) ? 1 : 0;
assign detect_max[329][16] = (mid_1[2647:2640] > mid_2[2655:2648]) ? 1 : 0;
assign detect_max[329][17] = (mid_1[2647:2640] > btm_0[2639:2632]) ? 1 : 0;
assign detect_max[329][18] = (mid_1[2647:2640] > btm_0[2647:2640]) ? 1 : 0;
assign detect_max[329][19] = (mid_1[2647:2640] > btm_0[2655:2648]) ? 1 : 0;
assign detect_max[329][20] = (mid_1[2647:2640] > btm_1[2639:2632]) ? 1 : 0;
assign detect_max[329][21] = (mid_1[2647:2640] > btm_1[2647:2640]) ? 1 : 0;
assign detect_max[329][22] = (mid_1[2647:2640] > btm_1[2655:2648]) ? 1 : 0;
assign detect_max[329][23] = (mid_1[2647:2640] > btm_2[2639:2632]) ? 1 : 0;
assign detect_max[329][24] = (mid_1[2647:2640] > btm_2[2647:2640]) ? 1 : 0;
assign detect_max[329][25] = (mid_1[2647:2640] > btm_2[2655:2648]) ? 1 : 0;

assign detect_max[330][0] = (mid_1[2655:2648] > top_0[2647:2640]) ? 1 : 0;
assign detect_max[330][1] = (mid_1[2655:2648] > top_0[2655:2648]) ? 1 : 0;
assign detect_max[330][2] = (mid_1[2655:2648] > top_0[2663:2656]) ? 1 : 0;
assign detect_max[330][3] = (mid_1[2655:2648] > top_1[2647:2640]) ? 1 : 0;
assign detect_max[330][4] = (mid_1[2655:2648] > top_1[2655:2648]) ? 1 : 0;
assign detect_max[330][5] = (mid_1[2655:2648] > top_1[2663:2656]) ? 1 : 0;
assign detect_max[330][6] = (mid_1[2655:2648] > top_2[2647:2640]) ? 1 : 0;
assign detect_max[330][7] = (mid_1[2655:2648] > top_2[2655:2648]) ? 1 : 0;
assign detect_max[330][8] = (mid_1[2655:2648] > top_2[2663:2656]) ? 1 : 0;
assign detect_max[330][9] = (mid_1[2655:2648] > mid_0[2647:2640]) ? 1 : 0;
assign detect_max[330][10] = (mid_1[2655:2648] > mid_0[2655:2648]) ? 1 : 0;
assign detect_max[330][11] = (mid_1[2655:2648] > mid_0[2663:2656]) ? 1 : 0;
assign detect_max[330][12] = (mid_1[2655:2648] > mid_1[2647:2640]) ? 1 : 0;
assign detect_max[330][13] = (mid_1[2655:2648] > mid_1[2663:2656]) ? 1 : 0;
assign detect_max[330][14] = (mid_1[2655:2648] > mid_2[2647:2640]) ? 1 : 0;
assign detect_max[330][15] = (mid_1[2655:2648] > mid_2[2655:2648]) ? 1 : 0;
assign detect_max[330][16] = (mid_1[2655:2648] > mid_2[2663:2656]) ? 1 : 0;
assign detect_max[330][17] = (mid_1[2655:2648] > btm_0[2647:2640]) ? 1 : 0;
assign detect_max[330][18] = (mid_1[2655:2648] > btm_0[2655:2648]) ? 1 : 0;
assign detect_max[330][19] = (mid_1[2655:2648] > btm_0[2663:2656]) ? 1 : 0;
assign detect_max[330][20] = (mid_1[2655:2648] > btm_1[2647:2640]) ? 1 : 0;
assign detect_max[330][21] = (mid_1[2655:2648] > btm_1[2655:2648]) ? 1 : 0;
assign detect_max[330][22] = (mid_1[2655:2648] > btm_1[2663:2656]) ? 1 : 0;
assign detect_max[330][23] = (mid_1[2655:2648] > btm_2[2647:2640]) ? 1 : 0;
assign detect_max[330][24] = (mid_1[2655:2648] > btm_2[2655:2648]) ? 1 : 0;
assign detect_max[330][25] = (mid_1[2655:2648] > btm_2[2663:2656]) ? 1 : 0;

assign detect_max[331][0] = (mid_1[2663:2656] > top_0[2655:2648]) ? 1 : 0;
assign detect_max[331][1] = (mid_1[2663:2656] > top_0[2663:2656]) ? 1 : 0;
assign detect_max[331][2] = (mid_1[2663:2656] > top_0[2671:2664]) ? 1 : 0;
assign detect_max[331][3] = (mid_1[2663:2656] > top_1[2655:2648]) ? 1 : 0;
assign detect_max[331][4] = (mid_1[2663:2656] > top_1[2663:2656]) ? 1 : 0;
assign detect_max[331][5] = (mid_1[2663:2656] > top_1[2671:2664]) ? 1 : 0;
assign detect_max[331][6] = (mid_1[2663:2656] > top_2[2655:2648]) ? 1 : 0;
assign detect_max[331][7] = (mid_1[2663:2656] > top_2[2663:2656]) ? 1 : 0;
assign detect_max[331][8] = (mid_1[2663:2656] > top_2[2671:2664]) ? 1 : 0;
assign detect_max[331][9] = (mid_1[2663:2656] > mid_0[2655:2648]) ? 1 : 0;
assign detect_max[331][10] = (mid_1[2663:2656] > mid_0[2663:2656]) ? 1 : 0;
assign detect_max[331][11] = (mid_1[2663:2656] > mid_0[2671:2664]) ? 1 : 0;
assign detect_max[331][12] = (mid_1[2663:2656] > mid_1[2655:2648]) ? 1 : 0;
assign detect_max[331][13] = (mid_1[2663:2656] > mid_1[2671:2664]) ? 1 : 0;
assign detect_max[331][14] = (mid_1[2663:2656] > mid_2[2655:2648]) ? 1 : 0;
assign detect_max[331][15] = (mid_1[2663:2656] > mid_2[2663:2656]) ? 1 : 0;
assign detect_max[331][16] = (mid_1[2663:2656] > mid_2[2671:2664]) ? 1 : 0;
assign detect_max[331][17] = (mid_1[2663:2656] > btm_0[2655:2648]) ? 1 : 0;
assign detect_max[331][18] = (mid_1[2663:2656] > btm_0[2663:2656]) ? 1 : 0;
assign detect_max[331][19] = (mid_1[2663:2656] > btm_0[2671:2664]) ? 1 : 0;
assign detect_max[331][20] = (mid_1[2663:2656] > btm_1[2655:2648]) ? 1 : 0;
assign detect_max[331][21] = (mid_1[2663:2656] > btm_1[2663:2656]) ? 1 : 0;
assign detect_max[331][22] = (mid_1[2663:2656] > btm_1[2671:2664]) ? 1 : 0;
assign detect_max[331][23] = (mid_1[2663:2656] > btm_2[2655:2648]) ? 1 : 0;
assign detect_max[331][24] = (mid_1[2663:2656] > btm_2[2663:2656]) ? 1 : 0;
assign detect_max[331][25] = (mid_1[2663:2656] > btm_2[2671:2664]) ? 1 : 0;

assign detect_max[332][0] = (mid_1[2671:2664] > top_0[2663:2656]) ? 1 : 0;
assign detect_max[332][1] = (mid_1[2671:2664] > top_0[2671:2664]) ? 1 : 0;
assign detect_max[332][2] = (mid_1[2671:2664] > top_0[2679:2672]) ? 1 : 0;
assign detect_max[332][3] = (mid_1[2671:2664] > top_1[2663:2656]) ? 1 : 0;
assign detect_max[332][4] = (mid_1[2671:2664] > top_1[2671:2664]) ? 1 : 0;
assign detect_max[332][5] = (mid_1[2671:2664] > top_1[2679:2672]) ? 1 : 0;
assign detect_max[332][6] = (mid_1[2671:2664] > top_2[2663:2656]) ? 1 : 0;
assign detect_max[332][7] = (mid_1[2671:2664] > top_2[2671:2664]) ? 1 : 0;
assign detect_max[332][8] = (mid_1[2671:2664] > top_2[2679:2672]) ? 1 : 0;
assign detect_max[332][9] = (mid_1[2671:2664] > mid_0[2663:2656]) ? 1 : 0;
assign detect_max[332][10] = (mid_1[2671:2664] > mid_0[2671:2664]) ? 1 : 0;
assign detect_max[332][11] = (mid_1[2671:2664] > mid_0[2679:2672]) ? 1 : 0;
assign detect_max[332][12] = (mid_1[2671:2664] > mid_1[2663:2656]) ? 1 : 0;
assign detect_max[332][13] = (mid_1[2671:2664] > mid_1[2679:2672]) ? 1 : 0;
assign detect_max[332][14] = (mid_1[2671:2664] > mid_2[2663:2656]) ? 1 : 0;
assign detect_max[332][15] = (mid_1[2671:2664] > mid_2[2671:2664]) ? 1 : 0;
assign detect_max[332][16] = (mid_1[2671:2664] > mid_2[2679:2672]) ? 1 : 0;
assign detect_max[332][17] = (mid_1[2671:2664] > btm_0[2663:2656]) ? 1 : 0;
assign detect_max[332][18] = (mid_1[2671:2664] > btm_0[2671:2664]) ? 1 : 0;
assign detect_max[332][19] = (mid_1[2671:2664] > btm_0[2679:2672]) ? 1 : 0;
assign detect_max[332][20] = (mid_1[2671:2664] > btm_1[2663:2656]) ? 1 : 0;
assign detect_max[332][21] = (mid_1[2671:2664] > btm_1[2671:2664]) ? 1 : 0;
assign detect_max[332][22] = (mid_1[2671:2664] > btm_1[2679:2672]) ? 1 : 0;
assign detect_max[332][23] = (mid_1[2671:2664] > btm_2[2663:2656]) ? 1 : 0;
assign detect_max[332][24] = (mid_1[2671:2664] > btm_2[2671:2664]) ? 1 : 0;
assign detect_max[332][25] = (mid_1[2671:2664] > btm_2[2679:2672]) ? 1 : 0;

assign detect_max[333][0] = (mid_1[2679:2672] > top_0[2671:2664]) ? 1 : 0;
assign detect_max[333][1] = (mid_1[2679:2672] > top_0[2679:2672]) ? 1 : 0;
assign detect_max[333][2] = (mid_1[2679:2672] > top_0[2687:2680]) ? 1 : 0;
assign detect_max[333][3] = (mid_1[2679:2672] > top_1[2671:2664]) ? 1 : 0;
assign detect_max[333][4] = (mid_1[2679:2672] > top_1[2679:2672]) ? 1 : 0;
assign detect_max[333][5] = (mid_1[2679:2672] > top_1[2687:2680]) ? 1 : 0;
assign detect_max[333][6] = (mid_1[2679:2672] > top_2[2671:2664]) ? 1 : 0;
assign detect_max[333][7] = (mid_1[2679:2672] > top_2[2679:2672]) ? 1 : 0;
assign detect_max[333][8] = (mid_1[2679:2672] > top_2[2687:2680]) ? 1 : 0;
assign detect_max[333][9] = (mid_1[2679:2672] > mid_0[2671:2664]) ? 1 : 0;
assign detect_max[333][10] = (mid_1[2679:2672] > mid_0[2679:2672]) ? 1 : 0;
assign detect_max[333][11] = (mid_1[2679:2672] > mid_0[2687:2680]) ? 1 : 0;
assign detect_max[333][12] = (mid_1[2679:2672] > mid_1[2671:2664]) ? 1 : 0;
assign detect_max[333][13] = (mid_1[2679:2672] > mid_1[2687:2680]) ? 1 : 0;
assign detect_max[333][14] = (mid_1[2679:2672] > mid_2[2671:2664]) ? 1 : 0;
assign detect_max[333][15] = (mid_1[2679:2672] > mid_2[2679:2672]) ? 1 : 0;
assign detect_max[333][16] = (mid_1[2679:2672] > mid_2[2687:2680]) ? 1 : 0;
assign detect_max[333][17] = (mid_1[2679:2672] > btm_0[2671:2664]) ? 1 : 0;
assign detect_max[333][18] = (mid_1[2679:2672] > btm_0[2679:2672]) ? 1 : 0;
assign detect_max[333][19] = (mid_1[2679:2672] > btm_0[2687:2680]) ? 1 : 0;
assign detect_max[333][20] = (mid_1[2679:2672] > btm_1[2671:2664]) ? 1 : 0;
assign detect_max[333][21] = (mid_1[2679:2672] > btm_1[2679:2672]) ? 1 : 0;
assign detect_max[333][22] = (mid_1[2679:2672] > btm_1[2687:2680]) ? 1 : 0;
assign detect_max[333][23] = (mid_1[2679:2672] > btm_2[2671:2664]) ? 1 : 0;
assign detect_max[333][24] = (mid_1[2679:2672] > btm_2[2679:2672]) ? 1 : 0;
assign detect_max[333][25] = (mid_1[2679:2672] > btm_2[2687:2680]) ? 1 : 0;

assign detect_max[334][0] = (mid_1[2687:2680] > top_0[2679:2672]) ? 1 : 0;
assign detect_max[334][1] = (mid_1[2687:2680] > top_0[2687:2680]) ? 1 : 0;
assign detect_max[334][2] = (mid_1[2687:2680] > top_0[2695:2688]) ? 1 : 0;
assign detect_max[334][3] = (mid_1[2687:2680] > top_1[2679:2672]) ? 1 : 0;
assign detect_max[334][4] = (mid_1[2687:2680] > top_1[2687:2680]) ? 1 : 0;
assign detect_max[334][5] = (mid_1[2687:2680] > top_1[2695:2688]) ? 1 : 0;
assign detect_max[334][6] = (mid_1[2687:2680] > top_2[2679:2672]) ? 1 : 0;
assign detect_max[334][7] = (mid_1[2687:2680] > top_2[2687:2680]) ? 1 : 0;
assign detect_max[334][8] = (mid_1[2687:2680] > top_2[2695:2688]) ? 1 : 0;
assign detect_max[334][9] = (mid_1[2687:2680] > mid_0[2679:2672]) ? 1 : 0;
assign detect_max[334][10] = (mid_1[2687:2680] > mid_0[2687:2680]) ? 1 : 0;
assign detect_max[334][11] = (mid_1[2687:2680] > mid_0[2695:2688]) ? 1 : 0;
assign detect_max[334][12] = (mid_1[2687:2680] > mid_1[2679:2672]) ? 1 : 0;
assign detect_max[334][13] = (mid_1[2687:2680] > mid_1[2695:2688]) ? 1 : 0;
assign detect_max[334][14] = (mid_1[2687:2680] > mid_2[2679:2672]) ? 1 : 0;
assign detect_max[334][15] = (mid_1[2687:2680] > mid_2[2687:2680]) ? 1 : 0;
assign detect_max[334][16] = (mid_1[2687:2680] > mid_2[2695:2688]) ? 1 : 0;
assign detect_max[334][17] = (mid_1[2687:2680] > btm_0[2679:2672]) ? 1 : 0;
assign detect_max[334][18] = (mid_1[2687:2680] > btm_0[2687:2680]) ? 1 : 0;
assign detect_max[334][19] = (mid_1[2687:2680] > btm_0[2695:2688]) ? 1 : 0;
assign detect_max[334][20] = (mid_1[2687:2680] > btm_1[2679:2672]) ? 1 : 0;
assign detect_max[334][21] = (mid_1[2687:2680] > btm_1[2687:2680]) ? 1 : 0;
assign detect_max[334][22] = (mid_1[2687:2680] > btm_1[2695:2688]) ? 1 : 0;
assign detect_max[334][23] = (mid_1[2687:2680] > btm_2[2679:2672]) ? 1 : 0;
assign detect_max[334][24] = (mid_1[2687:2680] > btm_2[2687:2680]) ? 1 : 0;
assign detect_max[334][25] = (mid_1[2687:2680] > btm_2[2695:2688]) ? 1 : 0;

assign detect_max[335][0] = (mid_1[2695:2688] > top_0[2687:2680]) ? 1 : 0;
assign detect_max[335][1] = (mid_1[2695:2688] > top_0[2695:2688]) ? 1 : 0;
assign detect_max[335][2] = (mid_1[2695:2688] > top_0[2703:2696]) ? 1 : 0;
assign detect_max[335][3] = (mid_1[2695:2688] > top_1[2687:2680]) ? 1 : 0;
assign detect_max[335][4] = (mid_1[2695:2688] > top_1[2695:2688]) ? 1 : 0;
assign detect_max[335][5] = (mid_1[2695:2688] > top_1[2703:2696]) ? 1 : 0;
assign detect_max[335][6] = (mid_1[2695:2688] > top_2[2687:2680]) ? 1 : 0;
assign detect_max[335][7] = (mid_1[2695:2688] > top_2[2695:2688]) ? 1 : 0;
assign detect_max[335][8] = (mid_1[2695:2688] > top_2[2703:2696]) ? 1 : 0;
assign detect_max[335][9] = (mid_1[2695:2688] > mid_0[2687:2680]) ? 1 : 0;
assign detect_max[335][10] = (mid_1[2695:2688] > mid_0[2695:2688]) ? 1 : 0;
assign detect_max[335][11] = (mid_1[2695:2688] > mid_0[2703:2696]) ? 1 : 0;
assign detect_max[335][12] = (mid_1[2695:2688] > mid_1[2687:2680]) ? 1 : 0;
assign detect_max[335][13] = (mid_1[2695:2688] > mid_1[2703:2696]) ? 1 : 0;
assign detect_max[335][14] = (mid_1[2695:2688] > mid_2[2687:2680]) ? 1 : 0;
assign detect_max[335][15] = (mid_1[2695:2688] > mid_2[2695:2688]) ? 1 : 0;
assign detect_max[335][16] = (mid_1[2695:2688] > mid_2[2703:2696]) ? 1 : 0;
assign detect_max[335][17] = (mid_1[2695:2688] > btm_0[2687:2680]) ? 1 : 0;
assign detect_max[335][18] = (mid_1[2695:2688] > btm_0[2695:2688]) ? 1 : 0;
assign detect_max[335][19] = (mid_1[2695:2688] > btm_0[2703:2696]) ? 1 : 0;
assign detect_max[335][20] = (mid_1[2695:2688] > btm_1[2687:2680]) ? 1 : 0;
assign detect_max[335][21] = (mid_1[2695:2688] > btm_1[2695:2688]) ? 1 : 0;
assign detect_max[335][22] = (mid_1[2695:2688] > btm_1[2703:2696]) ? 1 : 0;
assign detect_max[335][23] = (mid_1[2695:2688] > btm_2[2687:2680]) ? 1 : 0;
assign detect_max[335][24] = (mid_1[2695:2688] > btm_2[2695:2688]) ? 1 : 0;
assign detect_max[335][25] = (mid_1[2695:2688] > btm_2[2703:2696]) ? 1 : 0;

assign detect_max[336][0] = (mid_1[2703:2696] > top_0[2695:2688]) ? 1 : 0;
assign detect_max[336][1] = (mid_1[2703:2696] > top_0[2703:2696]) ? 1 : 0;
assign detect_max[336][2] = (mid_1[2703:2696] > top_0[2711:2704]) ? 1 : 0;
assign detect_max[336][3] = (mid_1[2703:2696] > top_1[2695:2688]) ? 1 : 0;
assign detect_max[336][4] = (mid_1[2703:2696] > top_1[2703:2696]) ? 1 : 0;
assign detect_max[336][5] = (mid_1[2703:2696] > top_1[2711:2704]) ? 1 : 0;
assign detect_max[336][6] = (mid_1[2703:2696] > top_2[2695:2688]) ? 1 : 0;
assign detect_max[336][7] = (mid_1[2703:2696] > top_2[2703:2696]) ? 1 : 0;
assign detect_max[336][8] = (mid_1[2703:2696] > top_2[2711:2704]) ? 1 : 0;
assign detect_max[336][9] = (mid_1[2703:2696] > mid_0[2695:2688]) ? 1 : 0;
assign detect_max[336][10] = (mid_1[2703:2696] > mid_0[2703:2696]) ? 1 : 0;
assign detect_max[336][11] = (mid_1[2703:2696] > mid_0[2711:2704]) ? 1 : 0;
assign detect_max[336][12] = (mid_1[2703:2696] > mid_1[2695:2688]) ? 1 : 0;
assign detect_max[336][13] = (mid_1[2703:2696] > mid_1[2711:2704]) ? 1 : 0;
assign detect_max[336][14] = (mid_1[2703:2696] > mid_2[2695:2688]) ? 1 : 0;
assign detect_max[336][15] = (mid_1[2703:2696] > mid_2[2703:2696]) ? 1 : 0;
assign detect_max[336][16] = (mid_1[2703:2696] > mid_2[2711:2704]) ? 1 : 0;
assign detect_max[336][17] = (mid_1[2703:2696] > btm_0[2695:2688]) ? 1 : 0;
assign detect_max[336][18] = (mid_1[2703:2696] > btm_0[2703:2696]) ? 1 : 0;
assign detect_max[336][19] = (mid_1[2703:2696] > btm_0[2711:2704]) ? 1 : 0;
assign detect_max[336][20] = (mid_1[2703:2696] > btm_1[2695:2688]) ? 1 : 0;
assign detect_max[336][21] = (mid_1[2703:2696] > btm_1[2703:2696]) ? 1 : 0;
assign detect_max[336][22] = (mid_1[2703:2696] > btm_1[2711:2704]) ? 1 : 0;
assign detect_max[336][23] = (mid_1[2703:2696] > btm_2[2695:2688]) ? 1 : 0;
assign detect_max[336][24] = (mid_1[2703:2696] > btm_2[2703:2696]) ? 1 : 0;
assign detect_max[336][25] = (mid_1[2703:2696] > btm_2[2711:2704]) ? 1 : 0;

assign detect_max[337][0] = (mid_1[2711:2704] > top_0[2703:2696]) ? 1 : 0;
assign detect_max[337][1] = (mid_1[2711:2704] > top_0[2711:2704]) ? 1 : 0;
assign detect_max[337][2] = (mid_1[2711:2704] > top_0[2719:2712]) ? 1 : 0;
assign detect_max[337][3] = (mid_1[2711:2704] > top_1[2703:2696]) ? 1 : 0;
assign detect_max[337][4] = (mid_1[2711:2704] > top_1[2711:2704]) ? 1 : 0;
assign detect_max[337][5] = (mid_1[2711:2704] > top_1[2719:2712]) ? 1 : 0;
assign detect_max[337][6] = (mid_1[2711:2704] > top_2[2703:2696]) ? 1 : 0;
assign detect_max[337][7] = (mid_1[2711:2704] > top_2[2711:2704]) ? 1 : 0;
assign detect_max[337][8] = (mid_1[2711:2704] > top_2[2719:2712]) ? 1 : 0;
assign detect_max[337][9] = (mid_1[2711:2704] > mid_0[2703:2696]) ? 1 : 0;
assign detect_max[337][10] = (mid_1[2711:2704] > mid_0[2711:2704]) ? 1 : 0;
assign detect_max[337][11] = (mid_1[2711:2704] > mid_0[2719:2712]) ? 1 : 0;
assign detect_max[337][12] = (mid_1[2711:2704] > mid_1[2703:2696]) ? 1 : 0;
assign detect_max[337][13] = (mid_1[2711:2704] > mid_1[2719:2712]) ? 1 : 0;
assign detect_max[337][14] = (mid_1[2711:2704] > mid_2[2703:2696]) ? 1 : 0;
assign detect_max[337][15] = (mid_1[2711:2704] > mid_2[2711:2704]) ? 1 : 0;
assign detect_max[337][16] = (mid_1[2711:2704] > mid_2[2719:2712]) ? 1 : 0;
assign detect_max[337][17] = (mid_1[2711:2704] > btm_0[2703:2696]) ? 1 : 0;
assign detect_max[337][18] = (mid_1[2711:2704] > btm_0[2711:2704]) ? 1 : 0;
assign detect_max[337][19] = (mid_1[2711:2704] > btm_0[2719:2712]) ? 1 : 0;
assign detect_max[337][20] = (mid_1[2711:2704] > btm_1[2703:2696]) ? 1 : 0;
assign detect_max[337][21] = (mid_1[2711:2704] > btm_1[2711:2704]) ? 1 : 0;
assign detect_max[337][22] = (mid_1[2711:2704] > btm_1[2719:2712]) ? 1 : 0;
assign detect_max[337][23] = (mid_1[2711:2704] > btm_2[2703:2696]) ? 1 : 0;
assign detect_max[337][24] = (mid_1[2711:2704] > btm_2[2711:2704]) ? 1 : 0;
assign detect_max[337][25] = (mid_1[2711:2704] > btm_2[2719:2712]) ? 1 : 0;

assign detect_max[338][0] = (mid_1[2719:2712] > top_0[2711:2704]) ? 1 : 0;
assign detect_max[338][1] = (mid_1[2719:2712] > top_0[2719:2712]) ? 1 : 0;
assign detect_max[338][2] = (mid_1[2719:2712] > top_0[2727:2720]) ? 1 : 0;
assign detect_max[338][3] = (mid_1[2719:2712] > top_1[2711:2704]) ? 1 : 0;
assign detect_max[338][4] = (mid_1[2719:2712] > top_1[2719:2712]) ? 1 : 0;
assign detect_max[338][5] = (mid_1[2719:2712] > top_1[2727:2720]) ? 1 : 0;
assign detect_max[338][6] = (mid_1[2719:2712] > top_2[2711:2704]) ? 1 : 0;
assign detect_max[338][7] = (mid_1[2719:2712] > top_2[2719:2712]) ? 1 : 0;
assign detect_max[338][8] = (mid_1[2719:2712] > top_2[2727:2720]) ? 1 : 0;
assign detect_max[338][9] = (mid_1[2719:2712] > mid_0[2711:2704]) ? 1 : 0;
assign detect_max[338][10] = (mid_1[2719:2712] > mid_0[2719:2712]) ? 1 : 0;
assign detect_max[338][11] = (mid_1[2719:2712] > mid_0[2727:2720]) ? 1 : 0;
assign detect_max[338][12] = (mid_1[2719:2712] > mid_1[2711:2704]) ? 1 : 0;
assign detect_max[338][13] = (mid_1[2719:2712] > mid_1[2727:2720]) ? 1 : 0;
assign detect_max[338][14] = (mid_1[2719:2712] > mid_2[2711:2704]) ? 1 : 0;
assign detect_max[338][15] = (mid_1[2719:2712] > mid_2[2719:2712]) ? 1 : 0;
assign detect_max[338][16] = (mid_1[2719:2712] > mid_2[2727:2720]) ? 1 : 0;
assign detect_max[338][17] = (mid_1[2719:2712] > btm_0[2711:2704]) ? 1 : 0;
assign detect_max[338][18] = (mid_1[2719:2712] > btm_0[2719:2712]) ? 1 : 0;
assign detect_max[338][19] = (mid_1[2719:2712] > btm_0[2727:2720]) ? 1 : 0;
assign detect_max[338][20] = (mid_1[2719:2712] > btm_1[2711:2704]) ? 1 : 0;
assign detect_max[338][21] = (mid_1[2719:2712] > btm_1[2719:2712]) ? 1 : 0;
assign detect_max[338][22] = (mid_1[2719:2712] > btm_1[2727:2720]) ? 1 : 0;
assign detect_max[338][23] = (mid_1[2719:2712] > btm_2[2711:2704]) ? 1 : 0;
assign detect_max[338][24] = (mid_1[2719:2712] > btm_2[2719:2712]) ? 1 : 0;
assign detect_max[338][25] = (mid_1[2719:2712] > btm_2[2727:2720]) ? 1 : 0;

assign detect_max[339][0] = (mid_1[2727:2720] > top_0[2719:2712]) ? 1 : 0;
assign detect_max[339][1] = (mid_1[2727:2720] > top_0[2727:2720]) ? 1 : 0;
assign detect_max[339][2] = (mid_1[2727:2720] > top_0[2735:2728]) ? 1 : 0;
assign detect_max[339][3] = (mid_1[2727:2720] > top_1[2719:2712]) ? 1 : 0;
assign detect_max[339][4] = (mid_1[2727:2720] > top_1[2727:2720]) ? 1 : 0;
assign detect_max[339][5] = (mid_1[2727:2720] > top_1[2735:2728]) ? 1 : 0;
assign detect_max[339][6] = (mid_1[2727:2720] > top_2[2719:2712]) ? 1 : 0;
assign detect_max[339][7] = (mid_1[2727:2720] > top_2[2727:2720]) ? 1 : 0;
assign detect_max[339][8] = (mid_1[2727:2720] > top_2[2735:2728]) ? 1 : 0;
assign detect_max[339][9] = (mid_1[2727:2720] > mid_0[2719:2712]) ? 1 : 0;
assign detect_max[339][10] = (mid_1[2727:2720] > mid_0[2727:2720]) ? 1 : 0;
assign detect_max[339][11] = (mid_1[2727:2720] > mid_0[2735:2728]) ? 1 : 0;
assign detect_max[339][12] = (mid_1[2727:2720] > mid_1[2719:2712]) ? 1 : 0;
assign detect_max[339][13] = (mid_1[2727:2720] > mid_1[2735:2728]) ? 1 : 0;
assign detect_max[339][14] = (mid_1[2727:2720] > mid_2[2719:2712]) ? 1 : 0;
assign detect_max[339][15] = (mid_1[2727:2720] > mid_2[2727:2720]) ? 1 : 0;
assign detect_max[339][16] = (mid_1[2727:2720] > mid_2[2735:2728]) ? 1 : 0;
assign detect_max[339][17] = (mid_1[2727:2720] > btm_0[2719:2712]) ? 1 : 0;
assign detect_max[339][18] = (mid_1[2727:2720] > btm_0[2727:2720]) ? 1 : 0;
assign detect_max[339][19] = (mid_1[2727:2720] > btm_0[2735:2728]) ? 1 : 0;
assign detect_max[339][20] = (mid_1[2727:2720] > btm_1[2719:2712]) ? 1 : 0;
assign detect_max[339][21] = (mid_1[2727:2720] > btm_1[2727:2720]) ? 1 : 0;
assign detect_max[339][22] = (mid_1[2727:2720] > btm_1[2735:2728]) ? 1 : 0;
assign detect_max[339][23] = (mid_1[2727:2720] > btm_2[2719:2712]) ? 1 : 0;
assign detect_max[339][24] = (mid_1[2727:2720] > btm_2[2727:2720]) ? 1 : 0;
assign detect_max[339][25] = (mid_1[2727:2720] > btm_2[2735:2728]) ? 1 : 0;

assign detect_max[340][0] = (mid_1[2735:2728] > top_0[2727:2720]) ? 1 : 0;
assign detect_max[340][1] = (mid_1[2735:2728] > top_0[2735:2728]) ? 1 : 0;
assign detect_max[340][2] = (mid_1[2735:2728] > top_0[2743:2736]) ? 1 : 0;
assign detect_max[340][3] = (mid_1[2735:2728] > top_1[2727:2720]) ? 1 : 0;
assign detect_max[340][4] = (mid_1[2735:2728] > top_1[2735:2728]) ? 1 : 0;
assign detect_max[340][5] = (mid_1[2735:2728] > top_1[2743:2736]) ? 1 : 0;
assign detect_max[340][6] = (mid_1[2735:2728] > top_2[2727:2720]) ? 1 : 0;
assign detect_max[340][7] = (mid_1[2735:2728] > top_2[2735:2728]) ? 1 : 0;
assign detect_max[340][8] = (mid_1[2735:2728] > top_2[2743:2736]) ? 1 : 0;
assign detect_max[340][9] = (mid_1[2735:2728] > mid_0[2727:2720]) ? 1 : 0;
assign detect_max[340][10] = (mid_1[2735:2728] > mid_0[2735:2728]) ? 1 : 0;
assign detect_max[340][11] = (mid_1[2735:2728] > mid_0[2743:2736]) ? 1 : 0;
assign detect_max[340][12] = (mid_1[2735:2728] > mid_1[2727:2720]) ? 1 : 0;
assign detect_max[340][13] = (mid_1[2735:2728] > mid_1[2743:2736]) ? 1 : 0;
assign detect_max[340][14] = (mid_1[2735:2728] > mid_2[2727:2720]) ? 1 : 0;
assign detect_max[340][15] = (mid_1[2735:2728] > mid_2[2735:2728]) ? 1 : 0;
assign detect_max[340][16] = (mid_1[2735:2728] > mid_2[2743:2736]) ? 1 : 0;
assign detect_max[340][17] = (mid_1[2735:2728] > btm_0[2727:2720]) ? 1 : 0;
assign detect_max[340][18] = (mid_1[2735:2728] > btm_0[2735:2728]) ? 1 : 0;
assign detect_max[340][19] = (mid_1[2735:2728] > btm_0[2743:2736]) ? 1 : 0;
assign detect_max[340][20] = (mid_1[2735:2728] > btm_1[2727:2720]) ? 1 : 0;
assign detect_max[340][21] = (mid_1[2735:2728] > btm_1[2735:2728]) ? 1 : 0;
assign detect_max[340][22] = (mid_1[2735:2728] > btm_1[2743:2736]) ? 1 : 0;
assign detect_max[340][23] = (mid_1[2735:2728] > btm_2[2727:2720]) ? 1 : 0;
assign detect_max[340][24] = (mid_1[2735:2728] > btm_2[2735:2728]) ? 1 : 0;
assign detect_max[340][25] = (mid_1[2735:2728] > btm_2[2743:2736]) ? 1 : 0;

assign detect_max[341][0] = (mid_1[2743:2736] > top_0[2735:2728]) ? 1 : 0;
assign detect_max[341][1] = (mid_1[2743:2736] > top_0[2743:2736]) ? 1 : 0;
assign detect_max[341][2] = (mid_1[2743:2736] > top_0[2751:2744]) ? 1 : 0;
assign detect_max[341][3] = (mid_1[2743:2736] > top_1[2735:2728]) ? 1 : 0;
assign detect_max[341][4] = (mid_1[2743:2736] > top_1[2743:2736]) ? 1 : 0;
assign detect_max[341][5] = (mid_1[2743:2736] > top_1[2751:2744]) ? 1 : 0;
assign detect_max[341][6] = (mid_1[2743:2736] > top_2[2735:2728]) ? 1 : 0;
assign detect_max[341][7] = (mid_1[2743:2736] > top_2[2743:2736]) ? 1 : 0;
assign detect_max[341][8] = (mid_1[2743:2736] > top_2[2751:2744]) ? 1 : 0;
assign detect_max[341][9] = (mid_1[2743:2736] > mid_0[2735:2728]) ? 1 : 0;
assign detect_max[341][10] = (mid_1[2743:2736] > mid_0[2743:2736]) ? 1 : 0;
assign detect_max[341][11] = (mid_1[2743:2736] > mid_0[2751:2744]) ? 1 : 0;
assign detect_max[341][12] = (mid_1[2743:2736] > mid_1[2735:2728]) ? 1 : 0;
assign detect_max[341][13] = (mid_1[2743:2736] > mid_1[2751:2744]) ? 1 : 0;
assign detect_max[341][14] = (mid_1[2743:2736] > mid_2[2735:2728]) ? 1 : 0;
assign detect_max[341][15] = (mid_1[2743:2736] > mid_2[2743:2736]) ? 1 : 0;
assign detect_max[341][16] = (mid_1[2743:2736] > mid_2[2751:2744]) ? 1 : 0;
assign detect_max[341][17] = (mid_1[2743:2736] > btm_0[2735:2728]) ? 1 : 0;
assign detect_max[341][18] = (mid_1[2743:2736] > btm_0[2743:2736]) ? 1 : 0;
assign detect_max[341][19] = (mid_1[2743:2736] > btm_0[2751:2744]) ? 1 : 0;
assign detect_max[341][20] = (mid_1[2743:2736] > btm_1[2735:2728]) ? 1 : 0;
assign detect_max[341][21] = (mid_1[2743:2736] > btm_1[2743:2736]) ? 1 : 0;
assign detect_max[341][22] = (mid_1[2743:2736] > btm_1[2751:2744]) ? 1 : 0;
assign detect_max[341][23] = (mid_1[2743:2736] > btm_2[2735:2728]) ? 1 : 0;
assign detect_max[341][24] = (mid_1[2743:2736] > btm_2[2743:2736]) ? 1 : 0;
assign detect_max[341][25] = (mid_1[2743:2736] > btm_2[2751:2744]) ? 1 : 0;

assign detect_max[342][0] = (mid_1[2751:2744] > top_0[2743:2736]) ? 1 : 0;
assign detect_max[342][1] = (mid_1[2751:2744] > top_0[2751:2744]) ? 1 : 0;
assign detect_max[342][2] = (mid_1[2751:2744] > top_0[2759:2752]) ? 1 : 0;
assign detect_max[342][3] = (mid_1[2751:2744] > top_1[2743:2736]) ? 1 : 0;
assign detect_max[342][4] = (mid_1[2751:2744] > top_1[2751:2744]) ? 1 : 0;
assign detect_max[342][5] = (mid_1[2751:2744] > top_1[2759:2752]) ? 1 : 0;
assign detect_max[342][6] = (mid_1[2751:2744] > top_2[2743:2736]) ? 1 : 0;
assign detect_max[342][7] = (mid_1[2751:2744] > top_2[2751:2744]) ? 1 : 0;
assign detect_max[342][8] = (mid_1[2751:2744] > top_2[2759:2752]) ? 1 : 0;
assign detect_max[342][9] = (mid_1[2751:2744] > mid_0[2743:2736]) ? 1 : 0;
assign detect_max[342][10] = (mid_1[2751:2744] > mid_0[2751:2744]) ? 1 : 0;
assign detect_max[342][11] = (mid_1[2751:2744] > mid_0[2759:2752]) ? 1 : 0;
assign detect_max[342][12] = (mid_1[2751:2744] > mid_1[2743:2736]) ? 1 : 0;
assign detect_max[342][13] = (mid_1[2751:2744] > mid_1[2759:2752]) ? 1 : 0;
assign detect_max[342][14] = (mid_1[2751:2744] > mid_2[2743:2736]) ? 1 : 0;
assign detect_max[342][15] = (mid_1[2751:2744] > mid_2[2751:2744]) ? 1 : 0;
assign detect_max[342][16] = (mid_1[2751:2744] > mid_2[2759:2752]) ? 1 : 0;
assign detect_max[342][17] = (mid_1[2751:2744] > btm_0[2743:2736]) ? 1 : 0;
assign detect_max[342][18] = (mid_1[2751:2744] > btm_0[2751:2744]) ? 1 : 0;
assign detect_max[342][19] = (mid_1[2751:2744] > btm_0[2759:2752]) ? 1 : 0;
assign detect_max[342][20] = (mid_1[2751:2744] > btm_1[2743:2736]) ? 1 : 0;
assign detect_max[342][21] = (mid_1[2751:2744] > btm_1[2751:2744]) ? 1 : 0;
assign detect_max[342][22] = (mid_1[2751:2744] > btm_1[2759:2752]) ? 1 : 0;
assign detect_max[342][23] = (mid_1[2751:2744] > btm_2[2743:2736]) ? 1 : 0;
assign detect_max[342][24] = (mid_1[2751:2744] > btm_2[2751:2744]) ? 1 : 0;
assign detect_max[342][25] = (mid_1[2751:2744] > btm_2[2759:2752]) ? 1 : 0;

assign detect_max[343][0] = (mid_1[2759:2752] > top_0[2751:2744]) ? 1 : 0;
assign detect_max[343][1] = (mid_1[2759:2752] > top_0[2759:2752]) ? 1 : 0;
assign detect_max[343][2] = (mid_1[2759:2752] > top_0[2767:2760]) ? 1 : 0;
assign detect_max[343][3] = (mid_1[2759:2752] > top_1[2751:2744]) ? 1 : 0;
assign detect_max[343][4] = (mid_1[2759:2752] > top_1[2759:2752]) ? 1 : 0;
assign detect_max[343][5] = (mid_1[2759:2752] > top_1[2767:2760]) ? 1 : 0;
assign detect_max[343][6] = (mid_1[2759:2752] > top_2[2751:2744]) ? 1 : 0;
assign detect_max[343][7] = (mid_1[2759:2752] > top_2[2759:2752]) ? 1 : 0;
assign detect_max[343][8] = (mid_1[2759:2752] > top_2[2767:2760]) ? 1 : 0;
assign detect_max[343][9] = (mid_1[2759:2752] > mid_0[2751:2744]) ? 1 : 0;
assign detect_max[343][10] = (mid_1[2759:2752] > mid_0[2759:2752]) ? 1 : 0;
assign detect_max[343][11] = (mid_1[2759:2752] > mid_0[2767:2760]) ? 1 : 0;
assign detect_max[343][12] = (mid_1[2759:2752] > mid_1[2751:2744]) ? 1 : 0;
assign detect_max[343][13] = (mid_1[2759:2752] > mid_1[2767:2760]) ? 1 : 0;
assign detect_max[343][14] = (mid_1[2759:2752] > mid_2[2751:2744]) ? 1 : 0;
assign detect_max[343][15] = (mid_1[2759:2752] > mid_2[2759:2752]) ? 1 : 0;
assign detect_max[343][16] = (mid_1[2759:2752] > mid_2[2767:2760]) ? 1 : 0;
assign detect_max[343][17] = (mid_1[2759:2752] > btm_0[2751:2744]) ? 1 : 0;
assign detect_max[343][18] = (mid_1[2759:2752] > btm_0[2759:2752]) ? 1 : 0;
assign detect_max[343][19] = (mid_1[2759:2752] > btm_0[2767:2760]) ? 1 : 0;
assign detect_max[343][20] = (mid_1[2759:2752] > btm_1[2751:2744]) ? 1 : 0;
assign detect_max[343][21] = (mid_1[2759:2752] > btm_1[2759:2752]) ? 1 : 0;
assign detect_max[343][22] = (mid_1[2759:2752] > btm_1[2767:2760]) ? 1 : 0;
assign detect_max[343][23] = (mid_1[2759:2752] > btm_2[2751:2744]) ? 1 : 0;
assign detect_max[343][24] = (mid_1[2759:2752] > btm_2[2759:2752]) ? 1 : 0;
assign detect_max[343][25] = (mid_1[2759:2752] > btm_2[2767:2760]) ? 1 : 0;

assign detect_max[344][0] = (mid_1[2767:2760] > top_0[2759:2752]) ? 1 : 0;
assign detect_max[344][1] = (mid_1[2767:2760] > top_0[2767:2760]) ? 1 : 0;
assign detect_max[344][2] = (mid_1[2767:2760] > top_0[2775:2768]) ? 1 : 0;
assign detect_max[344][3] = (mid_1[2767:2760] > top_1[2759:2752]) ? 1 : 0;
assign detect_max[344][4] = (mid_1[2767:2760] > top_1[2767:2760]) ? 1 : 0;
assign detect_max[344][5] = (mid_1[2767:2760] > top_1[2775:2768]) ? 1 : 0;
assign detect_max[344][6] = (mid_1[2767:2760] > top_2[2759:2752]) ? 1 : 0;
assign detect_max[344][7] = (mid_1[2767:2760] > top_2[2767:2760]) ? 1 : 0;
assign detect_max[344][8] = (mid_1[2767:2760] > top_2[2775:2768]) ? 1 : 0;
assign detect_max[344][9] = (mid_1[2767:2760] > mid_0[2759:2752]) ? 1 : 0;
assign detect_max[344][10] = (mid_1[2767:2760] > mid_0[2767:2760]) ? 1 : 0;
assign detect_max[344][11] = (mid_1[2767:2760] > mid_0[2775:2768]) ? 1 : 0;
assign detect_max[344][12] = (mid_1[2767:2760] > mid_1[2759:2752]) ? 1 : 0;
assign detect_max[344][13] = (mid_1[2767:2760] > mid_1[2775:2768]) ? 1 : 0;
assign detect_max[344][14] = (mid_1[2767:2760] > mid_2[2759:2752]) ? 1 : 0;
assign detect_max[344][15] = (mid_1[2767:2760] > mid_2[2767:2760]) ? 1 : 0;
assign detect_max[344][16] = (mid_1[2767:2760] > mid_2[2775:2768]) ? 1 : 0;
assign detect_max[344][17] = (mid_1[2767:2760] > btm_0[2759:2752]) ? 1 : 0;
assign detect_max[344][18] = (mid_1[2767:2760] > btm_0[2767:2760]) ? 1 : 0;
assign detect_max[344][19] = (mid_1[2767:2760] > btm_0[2775:2768]) ? 1 : 0;
assign detect_max[344][20] = (mid_1[2767:2760] > btm_1[2759:2752]) ? 1 : 0;
assign detect_max[344][21] = (mid_1[2767:2760] > btm_1[2767:2760]) ? 1 : 0;
assign detect_max[344][22] = (mid_1[2767:2760] > btm_1[2775:2768]) ? 1 : 0;
assign detect_max[344][23] = (mid_1[2767:2760] > btm_2[2759:2752]) ? 1 : 0;
assign detect_max[344][24] = (mid_1[2767:2760] > btm_2[2767:2760]) ? 1 : 0;
assign detect_max[344][25] = (mid_1[2767:2760] > btm_2[2775:2768]) ? 1 : 0;

assign detect_max[345][0] = (mid_1[2775:2768] > top_0[2767:2760]) ? 1 : 0;
assign detect_max[345][1] = (mid_1[2775:2768] > top_0[2775:2768]) ? 1 : 0;
assign detect_max[345][2] = (mid_1[2775:2768] > top_0[2783:2776]) ? 1 : 0;
assign detect_max[345][3] = (mid_1[2775:2768] > top_1[2767:2760]) ? 1 : 0;
assign detect_max[345][4] = (mid_1[2775:2768] > top_1[2775:2768]) ? 1 : 0;
assign detect_max[345][5] = (mid_1[2775:2768] > top_1[2783:2776]) ? 1 : 0;
assign detect_max[345][6] = (mid_1[2775:2768] > top_2[2767:2760]) ? 1 : 0;
assign detect_max[345][7] = (mid_1[2775:2768] > top_2[2775:2768]) ? 1 : 0;
assign detect_max[345][8] = (mid_1[2775:2768] > top_2[2783:2776]) ? 1 : 0;
assign detect_max[345][9] = (mid_1[2775:2768] > mid_0[2767:2760]) ? 1 : 0;
assign detect_max[345][10] = (mid_1[2775:2768] > mid_0[2775:2768]) ? 1 : 0;
assign detect_max[345][11] = (mid_1[2775:2768] > mid_0[2783:2776]) ? 1 : 0;
assign detect_max[345][12] = (mid_1[2775:2768] > mid_1[2767:2760]) ? 1 : 0;
assign detect_max[345][13] = (mid_1[2775:2768] > mid_1[2783:2776]) ? 1 : 0;
assign detect_max[345][14] = (mid_1[2775:2768] > mid_2[2767:2760]) ? 1 : 0;
assign detect_max[345][15] = (mid_1[2775:2768] > mid_2[2775:2768]) ? 1 : 0;
assign detect_max[345][16] = (mid_1[2775:2768] > mid_2[2783:2776]) ? 1 : 0;
assign detect_max[345][17] = (mid_1[2775:2768] > btm_0[2767:2760]) ? 1 : 0;
assign detect_max[345][18] = (mid_1[2775:2768] > btm_0[2775:2768]) ? 1 : 0;
assign detect_max[345][19] = (mid_1[2775:2768] > btm_0[2783:2776]) ? 1 : 0;
assign detect_max[345][20] = (mid_1[2775:2768] > btm_1[2767:2760]) ? 1 : 0;
assign detect_max[345][21] = (mid_1[2775:2768] > btm_1[2775:2768]) ? 1 : 0;
assign detect_max[345][22] = (mid_1[2775:2768] > btm_1[2783:2776]) ? 1 : 0;
assign detect_max[345][23] = (mid_1[2775:2768] > btm_2[2767:2760]) ? 1 : 0;
assign detect_max[345][24] = (mid_1[2775:2768] > btm_2[2775:2768]) ? 1 : 0;
assign detect_max[345][25] = (mid_1[2775:2768] > btm_2[2783:2776]) ? 1 : 0;

assign detect_max[346][0] = (mid_1[2783:2776] > top_0[2775:2768]) ? 1 : 0;
assign detect_max[346][1] = (mid_1[2783:2776] > top_0[2783:2776]) ? 1 : 0;
assign detect_max[346][2] = (mid_1[2783:2776] > top_0[2791:2784]) ? 1 : 0;
assign detect_max[346][3] = (mid_1[2783:2776] > top_1[2775:2768]) ? 1 : 0;
assign detect_max[346][4] = (mid_1[2783:2776] > top_1[2783:2776]) ? 1 : 0;
assign detect_max[346][5] = (mid_1[2783:2776] > top_1[2791:2784]) ? 1 : 0;
assign detect_max[346][6] = (mid_1[2783:2776] > top_2[2775:2768]) ? 1 : 0;
assign detect_max[346][7] = (mid_1[2783:2776] > top_2[2783:2776]) ? 1 : 0;
assign detect_max[346][8] = (mid_1[2783:2776] > top_2[2791:2784]) ? 1 : 0;
assign detect_max[346][9] = (mid_1[2783:2776] > mid_0[2775:2768]) ? 1 : 0;
assign detect_max[346][10] = (mid_1[2783:2776] > mid_0[2783:2776]) ? 1 : 0;
assign detect_max[346][11] = (mid_1[2783:2776] > mid_0[2791:2784]) ? 1 : 0;
assign detect_max[346][12] = (mid_1[2783:2776] > mid_1[2775:2768]) ? 1 : 0;
assign detect_max[346][13] = (mid_1[2783:2776] > mid_1[2791:2784]) ? 1 : 0;
assign detect_max[346][14] = (mid_1[2783:2776] > mid_2[2775:2768]) ? 1 : 0;
assign detect_max[346][15] = (mid_1[2783:2776] > mid_2[2783:2776]) ? 1 : 0;
assign detect_max[346][16] = (mid_1[2783:2776] > mid_2[2791:2784]) ? 1 : 0;
assign detect_max[346][17] = (mid_1[2783:2776] > btm_0[2775:2768]) ? 1 : 0;
assign detect_max[346][18] = (mid_1[2783:2776] > btm_0[2783:2776]) ? 1 : 0;
assign detect_max[346][19] = (mid_1[2783:2776] > btm_0[2791:2784]) ? 1 : 0;
assign detect_max[346][20] = (mid_1[2783:2776] > btm_1[2775:2768]) ? 1 : 0;
assign detect_max[346][21] = (mid_1[2783:2776] > btm_1[2783:2776]) ? 1 : 0;
assign detect_max[346][22] = (mid_1[2783:2776] > btm_1[2791:2784]) ? 1 : 0;
assign detect_max[346][23] = (mid_1[2783:2776] > btm_2[2775:2768]) ? 1 : 0;
assign detect_max[346][24] = (mid_1[2783:2776] > btm_2[2783:2776]) ? 1 : 0;
assign detect_max[346][25] = (mid_1[2783:2776] > btm_2[2791:2784]) ? 1 : 0;

assign detect_max[347][0] = (mid_1[2791:2784] > top_0[2783:2776]) ? 1 : 0;
assign detect_max[347][1] = (mid_1[2791:2784] > top_0[2791:2784]) ? 1 : 0;
assign detect_max[347][2] = (mid_1[2791:2784] > top_0[2799:2792]) ? 1 : 0;
assign detect_max[347][3] = (mid_1[2791:2784] > top_1[2783:2776]) ? 1 : 0;
assign detect_max[347][4] = (mid_1[2791:2784] > top_1[2791:2784]) ? 1 : 0;
assign detect_max[347][5] = (mid_1[2791:2784] > top_1[2799:2792]) ? 1 : 0;
assign detect_max[347][6] = (mid_1[2791:2784] > top_2[2783:2776]) ? 1 : 0;
assign detect_max[347][7] = (mid_1[2791:2784] > top_2[2791:2784]) ? 1 : 0;
assign detect_max[347][8] = (mid_1[2791:2784] > top_2[2799:2792]) ? 1 : 0;
assign detect_max[347][9] = (mid_1[2791:2784] > mid_0[2783:2776]) ? 1 : 0;
assign detect_max[347][10] = (mid_1[2791:2784] > mid_0[2791:2784]) ? 1 : 0;
assign detect_max[347][11] = (mid_1[2791:2784] > mid_0[2799:2792]) ? 1 : 0;
assign detect_max[347][12] = (mid_1[2791:2784] > mid_1[2783:2776]) ? 1 : 0;
assign detect_max[347][13] = (mid_1[2791:2784] > mid_1[2799:2792]) ? 1 : 0;
assign detect_max[347][14] = (mid_1[2791:2784] > mid_2[2783:2776]) ? 1 : 0;
assign detect_max[347][15] = (mid_1[2791:2784] > mid_2[2791:2784]) ? 1 : 0;
assign detect_max[347][16] = (mid_1[2791:2784] > mid_2[2799:2792]) ? 1 : 0;
assign detect_max[347][17] = (mid_1[2791:2784] > btm_0[2783:2776]) ? 1 : 0;
assign detect_max[347][18] = (mid_1[2791:2784] > btm_0[2791:2784]) ? 1 : 0;
assign detect_max[347][19] = (mid_1[2791:2784] > btm_0[2799:2792]) ? 1 : 0;
assign detect_max[347][20] = (mid_1[2791:2784] > btm_1[2783:2776]) ? 1 : 0;
assign detect_max[347][21] = (mid_1[2791:2784] > btm_1[2791:2784]) ? 1 : 0;
assign detect_max[347][22] = (mid_1[2791:2784] > btm_1[2799:2792]) ? 1 : 0;
assign detect_max[347][23] = (mid_1[2791:2784] > btm_2[2783:2776]) ? 1 : 0;
assign detect_max[347][24] = (mid_1[2791:2784] > btm_2[2791:2784]) ? 1 : 0;
assign detect_max[347][25] = (mid_1[2791:2784] > btm_2[2799:2792]) ? 1 : 0;

assign detect_max[348][0] = (mid_1[2799:2792] > top_0[2791:2784]) ? 1 : 0;
assign detect_max[348][1] = (mid_1[2799:2792] > top_0[2799:2792]) ? 1 : 0;
assign detect_max[348][2] = (mid_1[2799:2792] > top_0[2807:2800]) ? 1 : 0;
assign detect_max[348][3] = (mid_1[2799:2792] > top_1[2791:2784]) ? 1 : 0;
assign detect_max[348][4] = (mid_1[2799:2792] > top_1[2799:2792]) ? 1 : 0;
assign detect_max[348][5] = (mid_1[2799:2792] > top_1[2807:2800]) ? 1 : 0;
assign detect_max[348][6] = (mid_1[2799:2792] > top_2[2791:2784]) ? 1 : 0;
assign detect_max[348][7] = (mid_1[2799:2792] > top_2[2799:2792]) ? 1 : 0;
assign detect_max[348][8] = (mid_1[2799:2792] > top_2[2807:2800]) ? 1 : 0;
assign detect_max[348][9] = (mid_1[2799:2792] > mid_0[2791:2784]) ? 1 : 0;
assign detect_max[348][10] = (mid_1[2799:2792] > mid_0[2799:2792]) ? 1 : 0;
assign detect_max[348][11] = (mid_1[2799:2792] > mid_0[2807:2800]) ? 1 : 0;
assign detect_max[348][12] = (mid_1[2799:2792] > mid_1[2791:2784]) ? 1 : 0;
assign detect_max[348][13] = (mid_1[2799:2792] > mid_1[2807:2800]) ? 1 : 0;
assign detect_max[348][14] = (mid_1[2799:2792] > mid_2[2791:2784]) ? 1 : 0;
assign detect_max[348][15] = (mid_1[2799:2792] > mid_2[2799:2792]) ? 1 : 0;
assign detect_max[348][16] = (mid_1[2799:2792] > mid_2[2807:2800]) ? 1 : 0;
assign detect_max[348][17] = (mid_1[2799:2792] > btm_0[2791:2784]) ? 1 : 0;
assign detect_max[348][18] = (mid_1[2799:2792] > btm_0[2799:2792]) ? 1 : 0;
assign detect_max[348][19] = (mid_1[2799:2792] > btm_0[2807:2800]) ? 1 : 0;
assign detect_max[348][20] = (mid_1[2799:2792] > btm_1[2791:2784]) ? 1 : 0;
assign detect_max[348][21] = (mid_1[2799:2792] > btm_1[2799:2792]) ? 1 : 0;
assign detect_max[348][22] = (mid_1[2799:2792] > btm_1[2807:2800]) ? 1 : 0;
assign detect_max[348][23] = (mid_1[2799:2792] > btm_2[2791:2784]) ? 1 : 0;
assign detect_max[348][24] = (mid_1[2799:2792] > btm_2[2799:2792]) ? 1 : 0;
assign detect_max[348][25] = (mid_1[2799:2792] > btm_2[2807:2800]) ? 1 : 0;

assign detect_max[349][0] = (mid_1[2807:2800] > top_0[2799:2792]) ? 1 : 0;
assign detect_max[349][1] = (mid_1[2807:2800] > top_0[2807:2800]) ? 1 : 0;
assign detect_max[349][2] = (mid_1[2807:2800] > top_0[2815:2808]) ? 1 : 0;
assign detect_max[349][3] = (mid_1[2807:2800] > top_1[2799:2792]) ? 1 : 0;
assign detect_max[349][4] = (mid_1[2807:2800] > top_1[2807:2800]) ? 1 : 0;
assign detect_max[349][5] = (mid_1[2807:2800] > top_1[2815:2808]) ? 1 : 0;
assign detect_max[349][6] = (mid_1[2807:2800] > top_2[2799:2792]) ? 1 : 0;
assign detect_max[349][7] = (mid_1[2807:2800] > top_2[2807:2800]) ? 1 : 0;
assign detect_max[349][8] = (mid_1[2807:2800] > top_2[2815:2808]) ? 1 : 0;
assign detect_max[349][9] = (mid_1[2807:2800] > mid_0[2799:2792]) ? 1 : 0;
assign detect_max[349][10] = (mid_1[2807:2800] > mid_0[2807:2800]) ? 1 : 0;
assign detect_max[349][11] = (mid_1[2807:2800] > mid_0[2815:2808]) ? 1 : 0;
assign detect_max[349][12] = (mid_1[2807:2800] > mid_1[2799:2792]) ? 1 : 0;
assign detect_max[349][13] = (mid_1[2807:2800] > mid_1[2815:2808]) ? 1 : 0;
assign detect_max[349][14] = (mid_1[2807:2800] > mid_2[2799:2792]) ? 1 : 0;
assign detect_max[349][15] = (mid_1[2807:2800] > mid_2[2807:2800]) ? 1 : 0;
assign detect_max[349][16] = (mid_1[2807:2800] > mid_2[2815:2808]) ? 1 : 0;
assign detect_max[349][17] = (mid_1[2807:2800] > btm_0[2799:2792]) ? 1 : 0;
assign detect_max[349][18] = (mid_1[2807:2800] > btm_0[2807:2800]) ? 1 : 0;
assign detect_max[349][19] = (mid_1[2807:2800] > btm_0[2815:2808]) ? 1 : 0;
assign detect_max[349][20] = (mid_1[2807:2800] > btm_1[2799:2792]) ? 1 : 0;
assign detect_max[349][21] = (mid_1[2807:2800] > btm_1[2807:2800]) ? 1 : 0;
assign detect_max[349][22] = (mid_1[2807:2800] > btm_1[2815:2808]) ? 1 : 0;
assign detect_max[349][23] = (mid_1[2807:2800] > btm_2[2799:2792]) ? 1 : 0;
assign detect_max[349][24] = (mid_1[2807:2800] > btm_2[2807:2800]) ? 1 : 0;
assign detect_max[349][25] = (mid_1[2807:2800] > btm_2[2815:2808]) ? 1 : 0;

assign detect_max[350][0] = (mid_1[2815:2808] > top_0[2807:2800]) ? 1 : 0;
assign detect_max[350][1] = (mid_1[2815:2808] > top_0[2815:2808]) ? 1 : 0;
assign detect_max[350][2] = (mid_1[2815:2808] > top_0[2823:2816]) ? 1 : 0;
assign detect_max[350][3] = (mid_1[2815:2808] > top_1[2807:2800]) ? 1 : 0;
assign detect_max[350][4] = (mid_1[2815:2808] > top_1[2815:2808]) ? 1 : 0;
assign detect_max[350][5] = (mid_1[2815:2808] > top_1[2823:2816]) ? 1 : 0;
assign detect_max[350][6] = (mid_1[2815:2808] > top_2[2807:2800]) ? 1 : 0;
assign detect_max[350][7] = (mid_1[2815:2808] > top_2[2815:2808]) ? 1 : 0;
assign detect_max[350][8] = (mid_1[2815:2808] > top_2[2823:2816]) ? 1 : 0;
assign detect_max[350][9] = (mid_1[2815:2808] > mid_0[2807:2800]) ? 1 : 0;
assign detect_max[350][10] = (mid_1[2815:2808] > mid_0[2815:2808]) ? 1 : 0;
assign detect_max[350][11] = (mid_1[2815:2808] > mid_0[2823:2816]) ? 1 : 0;
assign detect_max[350][12] = (mid_1[2815:2808] > mid_1[2807:2800]) ? 1 : 0;
assign detect_max[350][13] = (mid_1[2815:2808] > mid_1[2823:2816]) ? 1 : 0;
assign detect_max[350][14] = (mid_1[2815:2808] > mid_2[2807:2800]) ? 1 : 0;
assign detect_max[350][15] = (mid_1[2815:2808] > mid_2[2815:2808]) ? 1 : 0;
assign detect_max[350][16] = (mid_1[2815:2808] > mid_2[2823:2816]) ? 1 : 0;
assign detect_max[350][17] = (mid_1[2815:2808] > btm_0[2807:2800]) ? 1 : 0;
assign detect_max[350][18] = (mid_1[2815:2808] > btm_0[2815:2808]) ? 1 : 0;
assign detect_max[350][19] = (mid_1[2815:2808] > btm_0[2823:2816]) ? 1 : 0;
assign detect_max[350][20] = (mid_1[2815:2808] > btm_1[2807:2800]) ? 1 : 0;
assign detect_max[350][21] = (mid_1[2815:2808] > btm_1[2815:2808]) ? 1 : 0;
assign detect_max[350][22] = (mid_1[2815:2808] > btm_1[2823:2816]) ? 1 : 0;
assign detect_max[350][23] = (mid_1[2815:2808] > btm_2[2807:2800]) ? 1 : 0;
assign detect_max[350][24] = (mid_1[2815:2808] > btm_2[2815:2808]) ? 1 : 0;
assign detect_max[350][25] = (mid_1[2815:2808] > btm_2[2823:2816]) ? 1 : 0;

assign detect_max[351][0] = (mid_1[2823:2816] > top_0[2815:2808]) ? 1 : 0;
assign detect_max[351][1] = (mid_1[2823:2816] > top_0[2823:2816]) ? 1 : 0;
assign detect_max[351][2] = (mid_1[2823:2816] > top_0[2831:2824]) ? 1 : 0;
assign detect_max[351][3] = (mid_1[2823:2816] > top_1[2815:2808]) ? 1 : 0;
assign detect_max[351][4] = (mid_1[2823:2816] > top_1[2823:2816]) ? 1 : 0;
assign detect_max[351][5] = (mid_1[2823:2816] > top_1[2831:2824]) ? 1 : 0;
assign detect_max[351][6] = (mid_1[2823:2816] > top_2[2815:2808]) ? 1 : 0;
assign detect_max[351][7] = (mid_1[2823:2816] > top_2[2823:2816]) ? 1 : 0;
assign detect_max[351][8] = (mid_1[2823:2816] > top_2[2831:2824]) ? 1 : 0;
assign detect_max[351][9] = (mid_1[2823:2816] > mid_0[2815:2808]) ? 1 : 0;
assign detect_max[351][10] = (mid_1[2823:2816] > mid_0[2823:2816]) ? 1 : 0;
assign detect_max[351][11] = (mid_1[2823:2816] > mid_0[2831:2824]) ? 1 : 0;
assign detect_max[351][12] = (mid_1[2823:2816] > mid_1[2815:2808]) ? 1 : 0;
assign detect_max[351][13] = (mid_1[2823:2816] > mid_1[2831:2824]) ? 1 : 0;
assign detect_max[351][14] = (mid_1[2823:2816] > mid_2[2815:2808]) ? 1 : 0;
assign detect_max[351][15] = (mid_1[2823:2816] > mid_2[2823:2816]) ? 1 : 0;
assign detect_max[351][16] = (mid_1[2823:2816] > mid_2[2831:2824]) ? 1 : 0;
assign detect_max[351][17] = (mid_1[2823:2816] > btm_0[2815:2808]) ? 1 : 0;
assign detect_max[351][18] = (mid_1[2823:2816] > btm_0[2823:2816]) ? 1 : 0;
assign detect_max[351][19] = (mid_1[2823:2816] > btm_0[2831:2824]) ? 1 : 0;
assign detect_max[351][20] = (mid_1[2823:2816] > btm_1[2815:2808]) ? 1 : 0;
assign detect_max[351][21] = (mid_1[2823:2816] > btm_1[2823:2816]) ? 1 : 0;
assign detect_max[351][22] = (mid_1[2823:2816] > btm_1[2831:2824]) ? 1 : 0;
assign detect_max[351][23] = (mid_1[2823:2816] > btm_2[2815:2808]) ? 1 : 0;
assign detect_max[351][24] = (mid_1[2823:2816] > btm_2[2823:2816]) ? 1 : 0;
assign detect_max[351][25] = (mid_1[2823:2816] > btm_2[2831:2824]) ? 1 : 0;

assign detect_max[352][0] = (mid_1[2831:2824] > top_0[2823:2816]) ? 1 : 0;
assign detect_max[352][1] = (mid_1[2831:2824] > top_0[2831:2824]) ? 1 : 0;
assign detect_max[352][2] = (mid_1[2831:2824] > top_0[2839:2832]) ? 1 : 0;
assign detect_max[352][3] = (mid_1[2831:2824] > top_1[2823:2816]) ? 1 : 0;
assign detect_max[352][4] = (mid_1[2831:2824] > top_1[2831:2824]) ? 1 : 0;
assign detect_max[352][5] = (mid_1[2831:2824] > top_1[2839:2832]) ? 1 : 0;
assign detect_max[352][6] = (mid_1[2831:2824] > top_2[2823:2816]) ? 1 : 0;
assign detect_max[352][7] = (mid_1[2831:2824] > top_2[2831:2824]) ? 1 : 0;
assign detect_max[352][8] = (mid_1[2831:2824] > top_2[2839:2832]) ? 1 : 0;
assign detect_max[352][9] = (mid_1[2831:2824] > mid_0[2823:2816]) ? 1 : 0;
assign detect_max[352][10] = (mid_1[2831:2824] > mid_0[2831:2824]) ? 1 : 0;
assign detect_max[352][11] = (mid_1[2831:2824] > mid_0[2839:2832]) ? 1 : 0;
assign detect_max[352][12] = (mid_1[2831:2824] > mid_1[2823:2816]) ? 1 : 0;
assign detect_max[352][13] = (mid_1[2831:2824] > mid_1[2839:2832]) ? 1 : 0;
assign detect_max[352][14] = (mid_1[2831:2824] > mid_2[2823:2816]) ? 1 : 0;
assign detect_max[352][15] = (mid_1[2831:2824] > mid_2[2831:2824]) ? 1 : 0;
assign detect_max[352][16] = (mid_1[2831:2824] > mid_2[2839:2832]) ? 1 : 0;
assign detect_max[352][17] = (mid_1[2831:2824] > btm_0[2823:2816]) ? 1 : 0;
assign detect_max[352][18] = (mid_1[2831:2824] > btm_0[2831:2824]) ? 1 : 0;
assign detect_max[352][19] = (mid_1[2831:2824] > btm_0[2839:2832]) ? 1 : 0;
assign detect_max[352][20] = (mid_1[2831:2824] > btm_1[2823:2816]) ? 1 : 0;
assign detect_max[352][21] = (mid_1[2831:2824] > btm_1[2831:2824]) ? 1 : 0;
assign detect_max[352][22] = (mid_1[2831:2824] > btm_1[2839:2832]) ? 1 : 0;
assign detect_max[352][23] = (mid_1[2831:2824] > btm_2[2823:2816]) ? 1 : 0;
assign detect_max[352][24] = (mid_1[2831:2824] > btm_2[2831:2824]) ? 1 : 0;
assign detect_max[352][25] = (mid_1[2831:2824] > btm_2[2839:2832]) ? 1 : 0;

assign detect_max[353][0] = (mid_1[2839:2832] > top_0[2831:2824]) ? 1 : 0;
assign detect_max[353][1] = (mid_1[2839:2832] > top_0[2839:2832]) ? 1 : 0;
assign detect_max[353][2] = (mid_1[2839:2832] > top_0[2847:2840]) ? 1 : 0;
assign detect_max[353][3] = (mid_1[2839:2832] > top_1[2831:2824]) ? 1 : 0;
assign detect_max[353][4] = (mid_1[2839:2832] > top_1[2839:2832]) ? 1 : 0;
assign detect_max[353][5] = (mid_1[2839:2832] > top_1[2847:2840]) ? 1 : 0;
assign detect_max[353][6] = (mid_1[2839:2832] > top_2[2831:2824]) ? 1 : 0;
assign detect_max[353][7] = (mid_1[2839:2832] > top_2[2839:2832]) ? 1 : 0;
assign detect_max[353][8] = (mid_1[2839:2832] > top_2[2847:2840]) ? 1 : 0;
assign detect_max[353][9] = (mid_1[2839:2832] > mid_0[2831:2824]) ? 1 : 0;
assign detect_max[353][10] = (mid_1[2839:2832] > mid_0[2839:2832]) ? 1 : 0;
assign detect_max[353][11] = (mid_1[2839:2832] > mid_0[2847:2840]) ? 1 : 0;
assign detect_max[353][12] = (mid_1[2839:2832] > mid_1[2831:2824]) ? 1 : 0;
assign detect_max[353][13] = (mid_1[2839:2832] > mid_1[2847:2840]) ? 1 : 0;
assign detect_max[353][14] = (mid_1[2839:2832] > mid_2[2831:2824]) ? 1 : 0;
assign detect_max[353][15] = (mid_1[2839:2832] > mid_2[2839:2832]) ? 1 : 0;
assign detect_max[353][16] = (mid_1[2839:2832] > mid_2[2847:2840]) ? 1 : 0;
assign detect_max[353][17] = (mid_1[2839:2832] > btm_0[2831:2824]) ? 1 : 0;
assign detect_max[353][18] = (mid_1[2839:2832] > btm_0[2839:2832]) ? 1 : 0;
assign detect_max[353][19] = (mid_1[2839:2832] > btm_0[2847:2840]) ? 1 : 0;
assign detect_max[353][20] = (mid_1[2839:2832] > btm_1[2831:2824]) ? 1 : 0;
assign detect_max[353][21] = (mid_1[2839:2832] > btm_1[2839:2832]) ? 1 : 0;
assign detect_max[353][22] = (mid_1[2839:2832] > btm_1[2847:2840]) ? 1 : 0;
assign detect_max[353][23] = (mid_1[2839:2832] > btm_2[2831:2824]) ? 1 : 0;
assign detect_max[353][24] = (mid_1[2839:2832] > btm_2[2839:2832]) ? 1 : 0;
assign detect_max[353][25] = (mid_1[2839:2832] > btm_2[2847:2840]) ? 1 : 0;

assign detect_max[354][0] = (mid_1[2847:2840] > top_0[2839:2832]) ? 1 : 0;
assign detect_max[354][1] = (mid_1[2847:2840] > top_0[2847:2840]) ? 1 : 0;
assign detect_max[354][2] = (mid_1[2847:2840] > top_0[2855:2848]) ? 1 : 0;
assign detect_max[354][3] = (mid_1[2847:2840] > top_1[2839:2832]) ? 1 : 0;
assign detect_max[354][4] = (mid_1[2847:2840] > top_1[2847:2840]) ? 1 : 0;
assign detect_max[354][5] = (mid_1[2847:2840] > top_1[2855:2848]) ? 1 : 0;
assign detect_max[354][6] = (mid_1[2847:2840] > top_2[2839:2832]) ? 1 : 0;
assign detect_max[354][7] = (mid_1[2847:2840] > top_2[2847:2840]) ? 1 : 0;
assign detect_max[354][8] = (mid_1[2847:2840] > top_2[2855:2848]) ? 1 : 0;
assign detect_max[354][9] = (mid_1[2847:2840] > mid_0[2839:2832]) ? 1 : 0;
assign detect_max[354][10] = (mid_1[2847:2840] > mid_0[2847:2840]) ? 1 : 0;
assign detect_max[354][11] = (mid_1[2847:2840] > mid_0[2855:2848]) ? 1 : 0;
assign detect_max[354][12] = (mid_1[2847:2840] > mid_1[2839:2832]) ? 1 : 0;
assign detect_max[354][13] = (mid_1[2847:2840] > mid_1[2855:2848]) ? 1 : 0;
assign detect_max[354][14] = (mid_1[2847:2840] > mid_2[2839:2832]) ? 1 : 0;
assign detect_max[354][15] = (mid_1[2847:2840] > mid_2[2847:2840]) ? 1 : 0;
assign detect_max[354][16] = (mid_1[2847:2840] > mid_2[2855:2848]) ? 1 : 0;
assign detect_max[354][17] = (mid_1[2847:2840] > btm_0[2839:2832]) ? 1 : 0;
assign detect_max[354][18] = (mid_1[2847:2840] > btm_0[2847:2840]) ? 1 : 0;
assign detect_max[354][19] = (mid_1[2847:2840] > btm_0[2855:2848]) ? 1 : 0;
assign detect_max[354][20] = (mid_1[2847:2840] > btm_1[2839:2832]) ? 1 : 0;
assign detect_max[354][21] = (mid_1[2847:2840] > btm_1[2847:2840]) ? 1 : 0;
assign detect_max[354][22] = (mid_1[2847:2840] > btm_1[2855:2848]) ? 1 : 0;
assign detect_max[354][23] = (mid_1[2847:2840] > btm_2[2839:2832]) ? 1 : 0;
assign detect_max[354][24] = (mid_1[2847:2840] > btm_2[2847:2840]) ? 1 : 0;
assign detect_max[354][25] = (mid_1[2847:2840] > btm_2[2855:2848]) ? 1 : 0;

assign detect_max[355][0] = (mid_1[2855:2848] > top_0[2847:2840]) ? 1 : 0;
assign detect_max[355][1] = (mid_1[2855:2848] > top_0[2855:2848]) ? 1 : 0;
assign detect_max[355][2] = (mid_1[2855:2848] > top_0[2863:2856]) ? 1 : 0;
assign detect_max[355][3] = (mid_1[2855:2848] > top_1[2847:2840]) ? 1 : 0;
assign detect_max[355][4] = (mid_1[2855:2848] > top_1[2855:2848]) ? 1 : 0;
assign detect_max[355][5] = (mid_1[2855:2848] > top_1[2863:2856]) ? 1 : 0;
assign detect_max[355][6] = (mid_1[2855:2848] > top_2[2847:2840]) ? 1 : 0;
assign detect_max[355][7] = (mid_1[2855:2848] > top_2[2855:2848]) ? 1 : 0;
assign detect_max[355][8] = (mid_1[2855:2848] > top_2[2863:2856]) ? 1 : 0;
assign detect_max[355][9] = (mid_1[2855:2848] > mid_0[2847:2840]) ? 1 : 0;
assign detect_max[355][10] = (mid_1[2855:2848] > mid_0[2855:2848]) ? 1 : 0;
assign detect_max[355][11] = (mid_1[2855:2848] > mid_0[2863:2856]) ? 1 : 0;
assign detect_max[355][12] = (mid_1[2855:2848] > mid_1[2847:2840]) ? 1 : 0;
assign detect_max[355][13] = (mid_1[2855:2848] > mid_1[2863:2856]) ? 1 : 0;
assign detect_max[355][14] = (mid_1[2855:2848] > mid_2[2847:2840]) ? 1 : 0;
assign detect_max[355][15] = (mid_1[2855:2848] > mid_2[2855:2848]) ? 1 : 0;
assign detect_max[355][16] = (mid_1[2855:2848] > mid_2[2863:2856]) ? 1 : 0;
assign detect_max[355][17] = (mid_1[2855:2848] > btm_0[2847:2840]) ? 1 : 0;
assign detect_max[355][18] = (mid_1[2855:2848] > btm_0[2855:2848]) ? 1 : 0;
assign detect_max[355][19] = (mid_1[2855:2848] > btm_0[2863:2856]) ? 1 : 0;
assign detect_max[355][20] = (mid_1[2855:2848] > btm_1[2847:2840]) ? 1 : 0;
assign detect_max[355][21] = (mid_1[2855:2848] > btm_1[2855:2848]) ? 1 : 0;
assign detect_max[355][22] = (mid_1[2855:2848] > btm_1[2863:2856]) ? 1 : 0;
assign detect_max[355][23] = (mid_1[2855:2848] > btm_2[2847:2840]) ? 1 : 0;
assign detect_max[355][24] = (mid_1[2855:2848] > btm_2[2855:2848]) ? 1 : 0;
assign detect_max[355][25] = (mid_1[2855:2848] > btm_2[2863:2856]) ? 1 : 0;

assign detect_max[356][0] = (mid_1[2863:2856] > top_0[2855:2848]) ? 1 : 0;
assign detect_max[356][1] = (mid_1[2863:2856] > top_0[2863:2856]) ? 1 : 0;
assign detect_max[356][2] = (mid_1[2863:2856] > top_0[2871:2864]) ? 1 : 0;
assign detect_max[356][3] = (mid_1[2863:2856] > top_1[2855:2848]) ? 1 : 0;
assign detect_max[356][4] = (mid_1[2863:2856] > top_1[2863:2856]) ? 1 : 0;
assign detect_max[356][5] = (mid_1[2863:2856] > top_1[2871:2864]) ? 1 : 0;
assign detect_max[356][6] = (mid_1[2863:2856] > top_2[2855:2848]) ? 1 : 0;
assign detect_max[356][7] = (mid_1[2863:2856] > top_2[2863:2856]) ? 1 : 0;
assign detect_max[356][8] = (mid_1[2863:2856] > top_2[2871:2864]) ? 1 : 0;
assign detect_max[356][9] = (mid_1[2863:2856] > mid_0[2855:2848]) ? 1 : 0;
assign detect_max[356][10] = (mid_1[2863:2856] > mid_0[2863:2856]) ? 1 : 0;
assign detect_max[356][11] = (mid_1[2863:2856] > mid_0[2871:2864]) ? 1 : 0;
assign detect_max[356][12] = (mid_1[2863:2856] > mid_1[2855:2848]) ? 1 : 0;
assign detect_max[356][13] = (mid_1[2863:2856] > mid_1[2871:2864]) ? 1 : 0;
assign detect_max[356][14] = (mid_1[2863:2856] > mid_2[2855:2848]) ? 1 : 0;
assign detect_max[356][15] = (mid_1[2863:2856] > mid_2[2863:2856]) ? 1 : 0;
assign detect_max[356][16] = (mid_1[2863:2856] > mid_2[2871:2864]) ? 1 : 0;
assign detect_max[356][17] = (mid_1[2863:2856] > btm_0[2855:2848]) ? 1 : 0;
assign detect_max[356][18] = (mid_1[2863:2856] > btm_0[2863:2856]) ? 1 : 0;
assign detect_max[356][19] = (mid_1[2863:2856] > btm_0[2871:2864]) ? 1 : 0;
assign detect_max[356][20] = (mid_1[2863:2856] > btm_1[2855:2848]) ? 1 : 0;
assign detect_max[356][21] = (mid_1[2863:2856] > btm_1[2863:2856]) ? 1 : 0;
assign detect_max[356][22] = (mid_1[2863:2856] > btm_1[2871:2864]) ? 1 : 0;
assign detect_max[356][23] = (mid_1[2863:2856] > btm_2[2855:2848]) ? 1 : 0;
assign detect_max[356][24] = (mid_1[2863:2856] > btm_2[2863:2856]) ? 1 : 0;
assign detect_max[356][25] = (mid_1[2863:2856] > btm_2[2871:2864]) ? 1 : 0;

assign detect_max[357][0] = (mid_1[2871:2864] > top_0[2863:2856]) ? 1 : 0;
assign detect_max[357][1] = (mid_1[2871:2864] > top_0[2871:2864]) ? 1 : 0;
assign detect_max[357][2] = (mid_1[2871:2864] > top_0[2879:2872]) ? 1 : 0;
assign detect_max[357][3] = (mid_1[2871:2864] > top_1[2863:2856]) ? 1 : 0;
assign detect_max[357][4] = (mid_1[2871:2864] > top_1[2871:2864]) ? 1 : 0;
assign detect_max[357][5] = (mid_1[2871:2864] > top_1[2879:2872]) ? 1 : 0;
assign detect_max[357][6] = (mid_1[2871:2864] > top_2[2863:2856]) ? 1 : 0;
assign detect_max[357][7] = (mid_1[2871:2864] > top_2[2871:2864]) ? 1 : 0;
assign detect_max[357][8] = (mid_1[2871:2864] > top_2[2879:2872]) ? 1 : 0;
assign detect_max[357][9] = (mid_1[2871:2864] > mid_0[2863:2856]) ? 1 : 0;
assign detect_max[357][10] = (mid_1[2871:2864] > mid_0[2871:2864]) ? 1 : 0;
assign detect_max[357][11] = (mid_1[2871:2864] > mid_0[2879:2872]) ? 1 : 0;
assign detect_max[357][12] = (mid_1[2871:2864] > mid_1[2863:2856]) ? 1 : 0;
assign detect_max[357][13] = (mid_1[2871:2864] > mid_1[2879:2872]) ? 1 : 0;
assign detect_max[357][14] = (mid_1[2871:2864] > mid_2[2863:2856]) ? 1 : 0;
assign detect_max[357][15] = (mid_1[2871:2864] > mid_2[2871:2864]) ? 1 : 0;
assign detect_max[357][16] = (mid_1[2871:2864] > mid_2[2879:2872]) ? 1 : 0;
assign detect_max[357][17] = (mid_1[2871:2864] > btm_0[2863:2856]) ? 1 : 0;
assign detect_max[357][18] = (mid_1[2871:2864] > btm_0[2871:2864]) ? 1 : 0;
assign detect_max[357][19] = (mid_1[2871:2864] > btm_0[2879:2872]) ? 1 : 0;
assign detect_max[357][20] = (mid_1[2871:2864] > btm_1[2863:2856]) ? 1 : 0;
assign detect_max[357][21] = (mid_1[2871:2864] > btm_1[2871:2864]) ? 1 : 0;
assign detect_max[357][22] = (mid_1[2871:2864] > btm_1[2879:2872]) ? 1 : 0;
assign detect_max[357][23] = (mid_1[2871:2864] > btm_2[2863:2856]) ? 1 : 0;
assign detect_max[357][24] = (mid_1[2871:2864] > btm_2[2871:2864]) ? 1 : 0;
assign detect_max[357][25] = (mid_1[2871:2864] > btm_2[2879:2872]) ? 1 : 0;

assign detect_max[358][0] = (mid_1[2879:2872] > top_0[2871:2864]) ? 1 : 0;
assign detect_max[358][1] = (mid_1[2879:2872] > top_0[2879:2872]) ? 1 : 0;
assign detect_max[358][2] = (mid_1[2879:2872] > top_0[2887:2880]) ? 1 : 0;
assign detect_max[358][3] = (mid_1[2879:2872] > top_1[2871:2864]) ? 1 : 0;
assign detect_max[358][4] = (mid_1[2879:2872] > top_1[2879:2872]) ? 1 : 0;
assign detect_max[358][5] = (mid_1[2879:2872] > top_1[2887:2880]) ? 1 : 0;
assign detect_max[358][6] = (mid_1[2879:2872] > top_2[2871:2864]) ? 1 : 0;
assign detect_max[358][7] = (mid_1[2879:2872] > top_2[2879:2872]) ? 1 : 0;
assign detect_max[358][8] = (mid_1[2879:2872] > top_2[2887:2880]) ? 1 : 0;
assign detect_max[358][9] = (mid_1[2879:2872] > mid_0[2871:2864]) ? 1 : 0;
assign detect_max[358][10] = (mid_1[2879:2872] > mid_0[2879:2872]) ? 1 : 0;
assign detect_max[358][11] = (mid_1[2879:2872] > mid_0[2887:2880]) ? 1 : 0;
assign detect_max[358][12] = (mid_1[2879:2872] > mid_1[2871:2864]) ? 1 : 0;
assign detect_max[358][13] = (mid_1[2879:2872] > mid_1[2887:2880]) ? 1 : 0;
assign detect_max[358][14] = (mid_1[2879:2872] > mid_2[2871:2864]) ? 1 : 0;
assign detect_max[358][15] = (mid_1[2879:2872] > mid_2[2879:2872]) ? 1 : 0;
assign detect_max[358][16] = (mid_1[2879:2872] > mid_2[2887:2880]) ? 1 : 0;
assign detect_max[358][17] = (mid_1[2879:2872] > btm_0[2871:2864]) ? 1 : 0;
assign detect_max[358][18] = (mid_1[2879:2872] > btm_0[2879:2872]) ? 1 : 0;
assign detect_max[358][19] = (mid_1[2879:2872] > btm_0[2887:2880]) ? 1 : 0;
assign detect_max[358][20] = (mid_1[2879:2872] > btm_1[2871:2864]) ? 1 : 0;
assign detect_max[358][21] = (mid_1[2879:2872] > btm_1[2879:2872]) ? 1 : 0;
assign detect_max[358][22] = (mid_1[2879:2872] > btm_1[2887:2880]) ? 1 : 0;
assign detect_max[358][23] = (mid_1[2879:2872] > btm_2[2871:2864]) ? 1 : 0;
assign detect_max[358][24] = (mid_1[2879:2872] > btm_2[2879:2872]) ? 1 : 0;
assign detect_max[358][25] = (mid_1[2879:2872] > btm_2[2887:2880]) ? 1 : 0;

assign detect_max[359][0] = (mid_1[2887:2880] > top_0[2879:2872]) ? 1 : 0;
assign detect_max[359][1] = (mid_1[2887:2880] > top_0[2887:2880]) ? 1 : 0;
assign detect_max[359][2] = (mid_1[2887:2880] > top_0[2895:2888]) ? 1 : 0;
assign detect_max[359][3] = (mid_1[2887:2880] > top_1[2879:2872]) ? 1 : 0;
assign detect_max[359][4] = (mid_1[2887:2880] > top_1[2887:2880]) ? 1 : 0;
assign detect_max[359][5] = (mid_1[2887:2880] > top_1[2895:2888]) ? 1 : 0;
assign detect_max[359][6] = (mid_1[2887:2880] > top_2[2879:2872]) ? 1 : 0;
assign detect_max[359][7] = (mid_1[2887:2880] > top_2[2887:2880]) ? 1 : 0;
assign detect_max[359][8] = (mid_1[2887:2880] > top_2[2895:2888]) ? 1 : 0;
assign detect_max[359][9] = (mid_1[2887:2880] > mid_0[2879:2872]) ? 1 : 0;
assign detect_max[359][10] = (mid_1[2887:2880] > mid_0[2887:2880]) ? 1 : 0;
assign detect_max[359][11] = (mid_1[2887:2880] > mid_0[2895:2888]) ? 1 : 0;
assign detect_max[359][12] = (mid_1[2887:2880] > mid_1[2879:2872]) ? 1 : 0;
assign detect_max[359][13] = (mid_1[2887:2880] > mid_1[2895:2888]) ? 1 : 0;
assign detect_max[359][14] = (mid_1[2887:2880] > mid_2[2879:2872]) ? 1 : 0;
assign detect_max[359][15] = (mid_1[2887:2880] > mid_2[2887:2880]) ? 1 : 0;
assign detect_max[359][16] = (mid_1[2887:2880] > mid_2[2895:2888]) ? 1 : 0;
assign detect_max[359][17] = (mid_1[2887:2880] > btm_0[2879:2872]) ? 1 : 0;
assign detect_max[359][18] = (mid_1[2887:2880] > btm_0[2887:2880]) ? 1 : 0;
assign detect_max[359][19] = (mid_1[2887:2880] > btm_0[2895:2888]) ? 1 : 0;
assign detect_max[359][20] = (mid_1[2887:2880] > btm_1[2879:2872]) ? 1 : 0;
assign detect_max[359][21] = (mid_1[2887:2880] > btm_1[2887:2880]) ? 1 : 0;
assign detect_max[359][22] = (mid_1[2887:2880] > btm_1[2895:2888]) ? 1 : 0;
assign detect_max[359][23] = (mid_1[2887:2880] > btm_2[2879:2872]) ? 1 : 0;
assign detect_max[359][24] = (mid_1[2887:2880] > btm_2[2887:2880]) ? 1 : 0;
assign detect_max[359][25] = (mid_1[2887:2880] > btm_2[2895:2888]) ? 1 : 0;

assign detect_max[360][0] = (mid_1[2895:2888] > top_0[2887:2880]) ? 1 : 0;
assign detect_max[360][1] = (mid_1[2895:2888] > top_0[2895:2888]) ? 1 : 0;
assign detect_max[360][2] = (mid_1[2895:2888] > top_0[2903:2896]) ? 1 : 0;
assign detect_max[360][3] = (mid_1[2895:2888] > top_1[2887:2880]) ? 1 : 0;
assign detect_max[360][4] = (mid_1[2895:2888] > top_1[2895:2888]) ? 1 : 0;
assign detect_max[360][5] = (mid_1[2895:2888] > top_1[2903:2896]) ? 1 : 0;
assign detect_max[360][6] = (mid_1[2895:2888] > top_2[2887:2880]) ? 1 : 0;
assign detect_max[360][7] = (mid_1[2895:2888] > top_2[2895:2888]) ? 1 : 0;
assign detect_max[360][8] = (mid_1[2895:2888] > top_2[2903:2896]) ? 1 : 0;
assign detect_max[360][9] = (mid_1[2895:2888] > mid_0[2887:2880]) ? 1 : 0;
assign detect_max[360][10] = (mid_1[2895:2888] > mid_0[2895:2888]) ? 1 : 0;
assign detect_max[360][11] = (mid_1[2895:2888] > mid_0[2903:2896]) ? 1 : 0;
assign detect_max[360][12] = (mid_1[2895:2888] > mid_1[2887:2880]) ? 1 : 0;
assign detect_max[360][13] = (mid_1[2895:2888] > mid_1[2903:2896]) ? 1 : 0;
assign detect_max[360][14] = (mid_1[2895:2888] > mid_2[2887:2880]) ? 1 : 0;
assign detect_max[360][15] = (mid_1[2895:2888] > mid_2[2895:2888]) ? 1 : 0;
assign detect_max[360][16] = (mid_1[2895:2888] > mid_2[2903:2896]) ? 1 : 0;
assign detect_max[360][17] = (mid_1[2895:2888] > btm_0[2887:2880]) ? 1 : 0;
assign detect_max[360][18] = (mid_1[2895:2888] > btm_0[2895:2888]) ? 1 : 0;
assign detect_max[360][19] = (mid_1[2895:2888] > btm_0[2903:2896]) ? 1 : 0;
assign detect_max[360][20] = (mid_1[2895:2888] > btm_1[2887:2880]) ? 1 : 0;
assign detect_max[360][21] = (mid_1[2895:2888] > btm_1[2895:2888]) ? 1 : 0;
assign detect_max[360][22] = (mid_1[2895:2888] > btm_1[2903:2896]) ? 1 : 0;
assign detect_max[360][23] = (mid_1[2895:2888] > btm_2[2887:2880]) ? 1 : 0;
assign detect_max[360][24] = (mid_1[2895:2888] > btm_2[2895:2888]) ? 1 : 0;
assign detect_max[360][25] = (mid_1[2895:2888] > btm_2[2903:2896]) ? 1 : 0;

assign detect_max[361][0] = (mid_1[2903:2896] > top_0[2895:2888]) ? 1 : 0;
assign detect_max[361][1] = (mid_1[2903:2896] > top_0[2903:2896]) ? 1 : 0;
assign detect_max[361][2] = (mid_1[2903:2896] > top_0[2911:2904]) ? 1 : 0;
assign detect_max[361][3] = (mid_1[2903:2896] > top_1[2895:2888]) ? 1 : 0;
assign detect_max[361][4] = (mid_1[2903:2896] > top_1[2903:2896]) ? 1 : 0;
assign detect_max[361][5] = (mid_1[2903:2896] > top_1[2911:2904]) ? 1 : 0;
assign detect_max[361][6] = (mid_1[2903:2896] > top_2[2895:2888]) ? 1 : 0;
assign detect_max[361][7] = (mid_1[2903:2896] > top_2[2903:2896]) ? 1 : 0;
assign detect_max[361][8] = (mid_1[2903:2896] > top_2[2911:2904]) ? 1 : 0;
assign detect_max[361][9] = (mid_1[2903:2896] > mid_0[2895:2888]) ? 1 : 0;
assign detect_max[361][10] = (mid_1[2903:2896] > mid_0[2903:2896]) ? 1 : 0;
assign detect_max[361][11] = (mid_1[2903:2896] > mid_0[2911:2904]) ? 1 : 0;
assign detect_max[361][12] = (mid_1[2903:2896] > mid_1[2895:2888]) ? 1 : 0;
assign detect_max[361][13] = (mid_1[2903:2896] > mid_1[2911:2904]) ? 1 : 0;
assign detect_max[361][14] = (mid_1[2903:2896] > mid_2[2895:2888]) ? 1 : 0;
assign detect_max[361][15] = (mid_1[2903:2896] > mid_2[2903:2896]) ? 1 : 0;
assign detect_max[361][16] = (mid_1[2903:2896] > mid_2[2911:2904]) ? 1 : 0;
assign detect_max[361][17] = (mid_1[2903:2896] > btm_0[2895:2888]) ? 1 : 0;
assign detect_max[361][18] = (mid_1[2903:2896] > btm_0[2903:2896]) ? 1 : 0;
assign detect_max[361][19] = (mid_1[2903:2896] > btm_0[2911:2904]) ? 1 : 0;
assign detect_max[361][20] = (mid_1[2903:2896] > btm_1[2895:2888]) ? 1 : 0;
assign detect_max[361][21] = (mid_1[2903:2896] > btm_1[2903:2896]) ? 1 : 0;
assign detect_max[361][22] = (mid_1[2903:2896] > btm_1[2911:2904]) ? 1 : 0;
assign detect_max[361][23] = (mid_1[2903:2896] > btm_2[2895:2888]) ? 1 : 0;
assign detect_max[361][24] = (mid_1[2903:2896] > btm_2[2903:2896]) ? 1 : 0;
assign detect_max[361][25] = (mid_1[2903:2896] > btm_2[2911:2904]) ? 1 : 0;

assign detect_max[362][0] = (mid_1[2911:2904] > top_0[2903:2896]) ? 1 : 0;
assign detect_max[362][1] = (mid_1[2911:2904] > top_0[2911:2904]) ? 1 : 0;
assign detect_max[362][2] = (mid_1[2911:2904] > top_0[2919:2912]) ? 1 : 0;
assign detect_max[362][3] = (mid_1[2911:2904] > top_1[2903:2896]) ? 1 : 0;
assign detect_max[362][4] = (mid_1[2911:2904] > top_1[2911:2904]) ? 1 : 0;
assign detect_max[362][5] = (mid_1[2911:2904] > top_1[2919:2912]) ? 1 : 0;
assign detect_max[362][6] = (mid_1[2911:2904] > top_2[2903:2896]) ? 1 : 0;
assign detect_max[362][7] = (mid_1[2911:2904] > top_2[2911:2904]) ? 1 : 0;
assign detect_max[362][8] = (mid_1[2911:2904] > top_2[2919:2912]) ? 1 : 0;
assign detect_max[362][9] = (mid_1[2911:2904] > mid_0[2903:2896]) ? 1 : 0;
assign detect_max[362][10] = (mid_1[2911:2904] > mid_0[2911:2904]) ? 1 : 0;
assign detect_max[362][11] = (mid_1[2911:2904] > mid_0[2919:2912]) ? 1 : 0;
assign detect_max[362][12] = (mid_1[2911:2904] > mid_1[2903:2896]) ? 1 : 0;
assign detect_max[362][13] = (mid_1[2911:2904] > mid_1[2919:2912]) ? 1 : 0;
assign detect_max[362][14] = (mid_1[2911:2904] > mid_2[2903:2896]) ? 1 : 0;
assign detect_max[362][15] = (mid_1[2911:2904] > mid_2[2911:2904]) ? 1 : 0;
assign detect_max[362][16] = (mid_1[2911:2904] > mid_2[2919:2912]) ? 1 : 0;
assign detect_max[362][17] = (mid_1[2911:2904] > btm_0[2903:2896]) ? 1 : 0;
assign detect_max[362][18] = (mid_1[2911:2904] > btm_0[2911:2904]) ? 1 : 0;
assign detect_max[362][19] = (mid_1[2911:2904] > btm_0[2919:2912]) ? 1 : 0;
assign detect_max[362][20] = (mid_1[2911:2904] > btm_1[2903:2896]) ? 1 : 0;
assign detect_max[362][21] = (mid_1[2911:2904] > btm_1[2911:2904]) ? 1 : 0;
assign detect_max[362][22] = (mid_1[2911:2904] > btm_1[2919:2912]) ? 1 : 0;
assign detect_max[362][23] = (mid_1[2911:2904] > btm_2[2903:2896]) ? 1 : 0;
assign detect_max[362][24] = (mid_1[2911:2904] > btm_2[2911:2904]) ? 1 : 0;
assign detect_max[362][25] = (mid_1[2911:2904] > btm_2[2919:2912]) ? 1 : 0;

assign detect_max[363][0] = (mid_1[2919:2912] > top_0[2911:2904]) ? 1 : 0;
assign detect_max[363][1] = (mid_1[2919:2912] > top_0[2919:2912]) ? 1 : 0;
assign detect_max[363][2] = (mid_1[2919:2912] > top_0[2927:2920]) ? 1 : 0;
assign detect_max[363][3] = (mid_1[2919:2912] > top_1[2911:2904]) ? 1 : 0;
assign detect_max[363][4] = (mid_1[2919:2912] > top_1[2919:2912]) ? 1 : 0;
assign detect_max[363][5] = (mid_1[2919:2912] > top_1[2927:2920]) ? 1 : 0;
assign detect_max[363][6] = (mid_1[2919:2912] > top_2[2911:2904]) ? 1 : 0;
assign detect_max[363][7] = (mid_1[2919:2912] > top_2[2919:2912]) ? 1 : 0;
assign detect_max[363][8] = (mid_1[2919:2912] > top_2[2927:2920]) ? 1 : 0;
assign detect_max[363][9] = (mid_1[2919:2912] > mid_0[2911:2904]) ? 1 : 0;
assign detect_max[363][10] = (mid_1[2919:2912] > mid_0[2919:2912]) ? 1 : 0;
assign detect_max[363][11] = (mid_1[2919:2912] > mid_0[2927:2920]) ? 1 : 0;
assign detect_max[363][12] = (mid_1[2919:2912] > mid_1[2911:2904]) ? 1 : 0;
assign detect_max[363][13] = (mid_1[2919:2912] > mid_1[2927:2920]) ? 1 : 0;
assign detect_max[363][14] = (mid_1[2919:2912] > mid_2[2911:2904]) ? 1 : 0;
assign detect_max[363][15] = (mid_1[2919:2912] > mid_2[2919:2912]) ? 1 : 0;
assign detect_max[363][16] = (mid_1[2919:2912] > mid_2[2927:2920]) ? 1 : 0;
assign detect_max[363][17] = (mid_1[2919:2912] > btm_0[2911:2904]) ? 1 : 0;
assign detect_max[363][18] = (mid_1[2919:2912] > btm_0[2919:2912]) ? 1 : 0;
assign detect_max[363][19] = (mid_1[2919:2912] > btm_0[2927:2920]) ? 1 : 0;
assign detect_max[363][20] = (mid_1[2919:2912] > btm_1[2911:2904]) ? 1 : 0;
assign detect_max[363][21] = (mid_1[2919:2912] > btm_1[2919:2912]) ? 1 : 0;
assign detect_max[363][22] = (mid_1[2919:2912] > btm_1[2927:2920]) ? 1 : 0;
assign detect_max[363][23] = (mid_1[2919:2912] > btm_2[2911:2904]) ? 1 : 0;
assign detect_max[363][24] = (mid_1[2919:2912] > btm_2[2919:2912]) ? 1 : 0;
assign detect_max[363][25] = (mid_1[2919:2912] > btm_2[2927:2920]) ? 1 : 0;

assign detect_max[364][0] = (mid_1[2927:2920] > top_0[2919:2912]) ? 1 : 0;
assign detect_max[364][1] = (mid_1[2927:2920] > top_0[2927:2920]) ? 1 : 0;
assign detect_max[364][2] = (mid_1[2927:2920] > top_0[2935:2928]) ? 1 : 0;
assign detect_max[364][3] = (mid_1[2927:2920] > top_1[2919:2912]) ? 1 : 0;
assign detect_max[364][4] = (mid_1[2927:2920] > top_1[2927:2920]) ? 1 : 0;
assign detect_max[364][5] = (mid_1[2927:2920] > top_1[2935:2928]) ? 1 : 0;
assign detect_max[364][6] = (mid_1[2927:2920] > top_2[2919:2912]) ? 1 : 0;
assign detect_max[364][7] = (mid_1[2927:2920] > top_2[2927:2920]) ? 1 : 0;
assign detect_max[364][8] = (mid_1[2927:2920] > top_2[2935:2928]) ? 1 : 0;
assign detect_max[364][9] = (mid_1[2927:2920] > mid_0[2919:2912]) ? 1 : 0;
assign detect_max[364][10] = (mid_1[2927:2920] > mid_0[2927:2920]) ? 1 : 0;
assign detect_max[364][11] = (mid_1[2927:2920] > mid_0[2935:2928]) ? 1 : 0;
assign detect_max[364][12] = (mid_1[2927:2920] > mid_1[2919:2912]) ? 1 : 0;
assign detect_max[364][13] = (mid_1[2927:2920] > mid_1[2935:2928]) ? 1 : 0;
assign detect_max[364][14] = (mid_1[2927:2920] > mid_2[2919:2912]) ? 1 : 0;
assign detect_max[364][15] = (mid_1[2927:2920] > mid_2[2927:2920]) ? 1 : 0;
assign detect_max[364][16] = (mid_1[2927:2920] > mid_2[2935:2928]) ? 1 : 0;
assign detect_max[364][17] = (mid_1[2927:2920] > btm_0[2919:2912]) ? 1 : 0;
assign detect_max[364][18] = (mid_1[2927:2920] > btm_0[2927:2920]) ? 1 : 0;
assign detect_max[364][19] = (mid_1[2927:2920] > btm_0[2935:2928]) ? 1 : 0;
assign detect_max[364][20] = (mid_1[2927:2920] > btm_1[2919:2912]) ? 1 : 0;
assign detect_max[364][21] = (mid_1[2927:2920] > btm_1[2927:2920]) ? 1 : 0;
assign detect_max[364][22] = (mid_1[2927:2920] > btm_1[2935:2928]) ? 1 : 0;
assign detect_max[364][23] = (mid_1[2927:2920] > btm_2[2919:2912]) ? 1 : 0;
assign detect_max[364][24] = (mid_1[2927:2920] > btm_2[2927:2920]) ? 1 : 0;
assign detect_max[364][25] = (mid_1[2927:2920] > btm_2[2935:2928]) ? 1 : 0;

assign detect_max[365][0] = (mid_1[2935:2928] > top_0[2927:2920]) ? 1 : 0;
assign detect_max[365][1] = (mid_1[2935:2928] > top_0[2935:2928]) ? 1 : 0;
assign detect_max[365][2] = (mid_1[2935:2928] > top_0[2943:2936]) ? 1 : 0;
assign detect_max[365][3] = (mid_1[2935:2928] > top_1[2927:2920]) ? 1 : 0;
assign detect_max[365][4] = (mid_1[2935:2928] > top_1[2935:2928]) ? 1 : 0;
assign detect_max[365][5] = (mid_1[2935:2928] > top_1[2943:2936]) ? 1 : 0;
assign detect_max[365][6] = (mid_1[2935:2928] > top_2[2927:2920]) ? 1 : 0;
assign detect_max[365][7] = (mid_1[2935:2928] > top_2[2935:2928]) ? 1 : 0;
assign detect_max[365][8] = (mid_1[2935:2928] > top_2[2943:2936]) ? 1 : 0;
assign detect_max[365][9] = (mid_1[2935:2928] > mid_0[2927:2920]) ? 1 : 0;
assign detect_max[365][10] = (mid_1[2935:2928] > mid_0[2935:2928]) ? 1 : 0;
assign detect_max[365][11] = (mid_1[2935:2928] > mid_0[2943:2936]) ? 1 : 0;
assign detect_max[365][12] = (mid_1[2935:2928] > mid_1[2927:2920]) ? 1 : 0;
assign detect_max[365][13] = (mid_1[2935:2928] > mid_1[2943:2936]) ? 1 : 0;
assign detect_max[365][14] = (mid_1[2935:2928] > mid_2[2927:2920]) ? 1 : 0;
assign detect_max[365][15] = (mid_1[2935:2928] > mid_2[2935:2928]) ? 1 : 0;
assign detect_max[365][16] = (mid_1[2935:2928] > mid_2[2943:2936]) ? 1 : 0;
assign detect_max[365][17] = (mid_1[2935:2928] > btm_0[2927:2920]) ? 1 : 0;
assign detect_max[365][18] = (mid_1[2935:2928] > btm_0[2935:2928]) ? 1 : 0;
assign detect_max[365][19] = (mid_1[2935:2928] > btm_0[2943:2936]) ? 1 : 0;
assign detect_max[365][20] = (mid_1[2935:2928] > btm_1[2927:2920]) ? 1 : 0;
assign detect_max[365][21] = (mid_1[2935:2928] > btm_1[2935:2928]) ? 1 : 0;
assign detect_max[365][22] = (mid_1[2935:2928] > btm_1[2943:2936]) ? 1 : 0;
assign detect_max[365][23] = (mid_1[2935:2928] > btm_2[2927:2920]) ? 1 : 0;
assign detect_max[365][24] = (mid_1[2935:2928] > btm_2[2935:2928]) ? 1 : 0;
assign detect_max[365][25] = (mid_1[2935:2928] > btm_2[2943:2936]) ? 1 : 0;

assign detect_max[366][0] = (mid_1[2943:2936] > top_0[2935:2928]) ? 1 : 0;
assign detect_max[366][1] = (mid_1[2943:2936] > top_0[2943:2936]) ? 1 : 0;
assign detect_max[366][2] = (mid_1[2943:2936] > top_0[2951:2944]) ? 1 : 0;
assign detect_max[366][3] = (mid_1[2943:2936] > top_1[2935:2928]) ? 1 : 0;
assign detect_max[366][4] = (mid_1[2943:2936] > top_1[2943:2936]) ? 1 : 0;
assign detect_max[366][5] = (mid_1[2943:2936] > top_1[2951:2944]) ? 1 : 0;
assign detect_max[366][6] = (mid_1[2943:2936] > top_2[2935:2928]) ? 1 : 0;
assign detect_max[366][7] = (mid_1[2943:2936] > top_2[2943:2936]) ? 1 : 0;
assign detect_max[366][8] = (mid_1[2943:2936] > top_2[2951:2944]) ? 1 : 0;
assign detect_max[366][9] = (mid_1[2943:2936] > mid_0[2935:2928]) ? 1 : 0;
assign detect_max[366][10] = (mid_1[2943:2936] > mid_0[2943:2936]) ? 1 : 0;
assign detect_max[366][11] = (mid_1[2943:2936] > mid_0[2951:2944]) ? 1 : 0;
assign detect_max[366][12] = (mid_1[2943:2936] > mid_1[2935:2928]) ? 1 : 0;
assign detect_max[366][13] = (mid_1[2943:2936] > mid_1[2951:2944]) ? 1 : 0;
assign detect_max[366][14] = (mid_1[2943:2936] > mid_2[2935:2928]) ? 1 : 0;
assign detect_max[366][15] = (mid_1[2943:2936] > mid_2[2943:2936]) ? 1 : 0;
assign detect_max[366][16] = (mid_1[2943:2936] > mid_2[2951:2944]) ? 1 : 0;
assign detect_max[366][17] = (mid_1[2943:2936] > btm_0[2935:2928]) ? 1 : 0;
assign detect_max[366][18] = (mid_1[2943:2936] > btm_0[2943:2936]) ? 1 : 0;
assign detect_max[366][19] = (mid_1[2943:2936] > btm_0[2951:2944]) ? 1 : 0;
assign detect_max[366][20] = (mid_1[2943:2936] > btm_1[2935:2928]) ? 1 : 0;
assign detect_max[366][21] = (mid_1[2943:2936] > btm_1[2943:2936]) ? 1 : 0;
assign detect_max[366][22] = (mid_1[2943:2936] > btm_1[2951:2944]) ? 1 : 0;
assign detect_max[366][23] = (mid_1[2943:2936] > btm_2[2935:2928]) ? 1 : 0;
assign detect_max[366][24] = (mid_1[2943:2936] > btm_2[2943:2936]) ? 1 : 0;
assign detect_max[366][25] = (mid_1[2943:2936] > btm_2[2951:2944]) ? 1 : 0;

assign detect_max[367][0] = (mid_1[2951:2944] > top_0[2943:2936]) ? 1 : 0;
assign detect_max[367][1] = (mid_1[2951:2944] > top_0[2951:2944]) ? 1 : 0;
assign detect_max[367][2] = (mid_1[2951:2944] > top_0[2959:2952]) ? 1 : 0;
assign detect_max[367][3] = (mid_1[2951:2944] > top_1[2943:2936]) ? 1 : 0;
assign detect_max[367][4] = (mid_1[2951:2944] > top_1[2951:2944]) ? 1 : 0;
assign detect_max[367][5] = (mid_1[2951:2944] > top_1[2959:2952]) ? 1 : 0;
assign detect_max[367][6] = (mid_1[2951:2944] > top_2[2943:2936]) ? 1 : 0;
assign detect_max[367][7] = (mid_1[2951:2944] > top_2[2951:2944]) ? 1 : 0;
assign detect_max[367][8] = (mid_1[2951:2944] > top_2[2959:2952]) ? 1 : 0;
assign detect_max[367][9] = (mid_1[2951:2944] > mid_0[2943:2936]) ? 1 : 0;
assign detect_max[367][10] = (mid_1[2951:2944] > mid_0[2951:2944]) ? 1 : 0;
assign detect_max[367][11] = (mid_1[2951:2944] > mid_0[2959:2952]) ? 1 : 0;
assign detect_max[367][12] = (mid_1[2951:2944] > mid_1[2943:2936]) ? 1 : 0;
assign detect_max[367][13] = (mid_1[2951:2944] > mid_1[2959:2952]) ? 1 : 0;
assign detect_max[367][14] = (mid_1[2951:2944] > mid_2[2943:2936]) ? 1 : 0;
assign detect_max[367][15] = (mid_1[2951:2944] > mid_2[2951:2944]) ? 1 : 0;
assign detect_max[367][16] = (mid_1[2951:2944] > mid_2[2959:2952]) ? 1 : 0;
assign detect_max[367][17] = (mid_1[2951:2944] > btm_0[2943:2936]) ? 1 : 0;
assign detect_max[367][18] = (mid_1[2951:2944] > btm_0[2951:2944]) ? 1 : 0;
assign detect_max[367][19] = (mid_1[2951:2944] > btm_0[2959:2952]) ? 1 : 0;
assign detect_max[367][20] = (mid_1[2951:2944] > btm_1[2943:2936]) ? 1 : 0;
assign detect_max[367][21] = (mid_1[2951:2944] > btm_1[2951:2944]) ? 1 : 0;
assign detect_max[367][22] = (mid_1[2951:2944] > btm_1[2959:2952]) ? 1 : 0;
assign detect_max[367][23] = (mid_1[2951:2944] > btm_2[2943:2936]) ? 1 : 0;
assign detect_max[367][24] = (mid_1[2951:2944] > btm_2[2951:2944]) ? 1 : 0;
assign detect_max[367][25] = (mid_1[2951:2944] > btm_2[2959:2952]) ? 1 : 0;

assign detect_max[368][0] = (mid_1[2959:2952] > top_0[2951:2944]) ? 1 : 0;
assign detect_max[368][1] = (mid_1[2959:2952] > top_0[2959:2952]) ? 1 : 0;
assign detect_max[368][2] = (mid_1[2959:2952] > top_0[2967:2960]) ? 1 : 0;
assign detect_max[368][3] = (mid_1[2959:2952] > top_1[2951:2944]) ? 1 : 0;
assign detect_max[368][4] = (mid_1[2959:2952] > top_1[2959:2952]) ? 1 : 0;
assign detect_max[368][5] = (mid_1[2959:2952] > top_1[2967:2960]) ? 1 : 0;
assign detect_max[368][6] = (mid_1[2959:2952] > top_2[2951:2944]) ? 1 : 0;
assign detect_max[368][7] = (mid_1[2959:2952] > top_2[2959:2952]) ? 1 : 0;
assign detect_max[368][8] = (mid_1[2959:2952] > top_2[2967:2960]) ? 1 : 0;
assign detect_max[368][9] = (mid_1[2959:2952] > mid_0[2951:2944]) ? 1 : 0;
assign detect_max[368][10] = (mid_1[2959:2952] > mid_0[2959:2952]) ? 1 : 0;
assign detect_max[368][11] = (mid_1[2959:2952] > mid_0[2967:2960]) ? 1 : 0;
assign detect_max[368][12] = (mid_1[2959:2952] > mid_1[2951:2944]) ? 1 : 0;
assign detect_max[368][13] = (mid_1[2959:2952] > mid_1[2967:2960]) ? 1 : 0;
assign detect_max[368][14] = (mid_1[2959:2952] > mid_2[2951:2944]) ? 1 : 0;
assign detect_max[368][15] = (mid_1[2959:2952] > mid_2[2959:2952]) ? 1 : 0;
assign detect_max[368][16] = (mid_1[2959:2952] > mid_2[2967:2960]) ? 1 : 0;
assign detect_max[368][17] = (mid_1[2959:2952] > btm_0[2951:2944]) ? 1 : 0;
assign detect_max[368][18] = (mid_1[2959:2952] > btm_0[2959:2952]) ? 1 : 0;
assign detect_max[368][19] = (mid_1[2959:2952] > btm_0[2967:2960]) ? 1 : 0;
assign detect_max[368][20] = (mid_1[2959:2952] > btm_1[2951:2944]) ? 1 : 0;
assign detect_max[368][21] = (mid_1[2959:2952] > btm_1[2959:2952]) ? 1 : 0;
assign detect_max[368][22] = (mid_1[2959:2952] > btm_1[2967:2960]) ? 1 : 0;
assign detect_max[368][23] = (mid_1[2959:2952] > btm_2[2951:2944]) ? 1 : 0;
assign detect_max[368][24] = (mid_1[2959:2952] > btm_2[2959:2952]) ? 1 : 0;
assign detect_max[368][25] = (mid_1[2959:2952] > btm_2[2967:2960]) ? 1 : 0;

assign detect_max[369][0] = (mid_1[2967:2960] > top_0[2959:2952]) ? 1 : 0;
assign detect_max[369][1] = (mid_1[2967:2960] > top_0[2967:2960]) ? 1 : 0;
assign detect_max[369][2] = (mid_1[2967:2960] > top_0[2975:2968]) ? 1 : 0;
assign detect_max[369][3] = (mid_1[2967:2960] > top_1[2959:2952]) ? 1 : 0;
assign detect_max[369][4] = (mid_1[2967:2960] > top_1[2967:2960]) ? 1 : 0;
assign detect_max[369][5] = (mid_1[2967:2960] > top_1[2975:2968]) ? 1 : 0;
assign detect_max[369][6] = (mid_1[2967:2960] > top_2[2959:2952]) ? 1 : 0;
assign detect_max[369][7] = (mid_1[2967:2960] > top_2[2967:2960]) ? 1 : 0;
assign detect_max[369][8] = (mid_1[2967:2960] > top_2[2975:2968]) ? 1 : 0;
assign detect_max[369][9] = (mid_1[2967:2960] > mid_0[2959:2952]) ? 1 : 0;
assign detect_max[369][10] = (mid_1[2967:2960] > mid_0[2967:2960]) ? 1 : 0;
assign detect_max[369][11] = (mid_1[2967:2960] > mid_0[2975:2968]) ? 1 : 0;
assign detect_max[369][12] = (mid_1[2967:2960] > mid_1[2959:2952]) ? 1 : 0;
assign detect_max[369][13] = (mid_1[2967:2960] > mid_1[2975:2968]) ? 1 : 0;
assign detect_max[369][14] = (mid_1[2967:2960] > mid_2[2959:2952]) ? 1 : 0;
assign detect_max[369][15] = (mid_1[2967:2960] > mid_2[2967:2960]) ? 1 : 0;
assign detect_max[369][16] = (mid_1[2967:2960] > mid_2[2975:2968]) ? 1 : 0;
assign detect_max[369][17] = (mid_1[2967:2960] > btm_0[2959:2952]) ? 1 : 0;
assign detect_max[369][18] = (mid_1[2967:2960] > btm_0[2967:2960]) ? 1 : 0;
assign detect_max[369][19] = (mid_1[2967:2960] > btm_0[2975:2968]) ? 1 : 0;
assign detect_max[369][20] = (mid_1[2967:2960] > btm_1[2959:2952]) ? 1 : 0;
assign detect_max[369][21] = (mid_1[2967:2960] > btm_1[2967:2960]) ? 1 : 0;
assign detect_max[369][22] = (mid_1[2967:2960] > btm_1[2975:2968]) ? 1 : 0;
assign detect_max[369][23] = (mid_1[2967:2960] > btm_2[2959:2952]) ? 1 : 0;
assign detect_max[369][24] = (mid_1[2967:2960] > btm_2[2967:2960]) ? 1 : 0;
assign detect_max[369][25] = (mid_1[2967:2960] > btm_2[2975:2968]) ? 1 : 0;

assign detect_max[370][0] = (mid_1[2975:2968] > top_0[2967:2960]) ? 1 : 0;
assign detect_max[370][1] = (mid_1[2975:2968] > top_0[2975:2968]) ? 1 : 0;
assign detect_max[370][2] = (mid_1[2975:2968] > top_0[2983:2976]) ? 1 : 0;
assign detect_max[370][3] = (mid_1[2975:2968] > top_1[2967:2960]) ? 1 : 0;
assign detect_max[370][4] = (mid_1[2975:2968] > top_1[2975:2968]) ? 1 : 0;
assign detect_max[370][5] = (mid_1[2975:2968] > top_1[2983:2976]) ? 1 : 0;
assign detect_max[370][6] = (mid_1[2975:2968] > top_2[2967:2960]) ? 1 : 0;
assign detect_max[370][7] = (mid_1[2975:2968] > top_2[2975:2968]) ? 1 : 0;
assign detect_max[370][8] = (mid_1[2975:2968] > top_2[2983:2976]) ? 1 : 0;
assign detect_max[370][9] = (mid_1[2975:2968] > mid_0[2967:2960]) ? 1 : 0;
assign detect_max[370][10] = (mid_1[2975:2968] > mid_0[2975:2968]) ? 1 : 0;
assign detect_max[370][11] = (mid_1[2975:2968] > mid_0[2983:2976]) ? 1 : 0;
assign detect_max[370][12] = (mid_1[2975:2968] > mid_1[2967:2960]) ? 1 : 0;
assign detect_max[370][13] = (mid_1[2975:2968] > mid_1[2983:2976]) ? 1 : 0;
assign detect_max[370][14] = (mid_1[2975:2968] > mid_2[2967:2960]) ? 1 : 0;
assign detect_max[370][15] = (mid_1[2975:2968] > mid_2[2975:2968]) ? 1 : 0;
assign detect_max[370][16] = (mid_1[2975:2968] > mid_2[2983:2976]) ? 1 : 0;
assign detect_max[370][17] = (mid_1[2975:2968] > btm_0[2967:2960]) ? 1 : 0;
assign detect_max[370][18] = (mid_1[2975:2968] > btm_0[2975:2968]) ? 1 : 0;
assign detect_max[370][19] = (mid_1[2975:2968] > btm_0[2983:2976]) ? 1 : 0;
assign detect_max[370][20] = (mid_1[2975:2968] > btm_1[2967:2960]) ? 1 : 0;
assign detect_max[370][21] = (mid_1[2975:2968] > btm_1[2975:2968]) ? 1 : 0;
assign detect_max[370][22] = (mid_1[2975:2968] > btm_1[2983:2976]) ? 1 : 0;
assign detect_max[370][23] = (mid_1[2975:2968] > btm_2[2967:2960]) ? 1 : 0;
assign detect_max[370][24] = (mid_1[2975:2968] > btm_2[2975:2968]) ? 1 : 0;
assign detect_max[370][25] = (mid_1[2975:2968] > btm_2[2983:2976]) ? 1 : 0;

assign detect_max[371][0] = (mid_1[2983:2976] > top_0[2975:2968]) ? 1 : 0;
assign detect_max[371][1] = (mid_1[2983:2976] > top_0[2983:2976]) ? 1 : 0;
assign detect_max[371][2] = (mid_1[2983:2976] > top_0[2991:2984]) ? 1 : 0;
assign detect_max[371][3] = (mid_1[2983:2976] > top_1[2975:2968]) ? 1 : 0;
assign detect_max[371][4] = (mid_1[2983:2976] > top_1[2983:2976]) ? 1 : 0;
assign detect_max[371][5] = (mid_1[2983:2976] > top_1[2991:2984]) ? 1 : 0;
assign detect_max[371][6] = (mid_1[2983:2976] > top_2[2975:2968]) ? 1 : 0;
assign detect_max[371][7] = (mid_1[2983:2976] > top_2[2983:2976]) ? 1 : 0;
assign detect_max[371][8] = (mid_1[2983:2976] > top_2[2991:2984]) ? 1 : 0;
assign detect_max[371][9] = (mid_1[2983:2976] > mid_0[2975:2968]) ? 1 : 0;
assign detect_max[371][10] = (mid_1[2983:2976] > mid_0[2983:2976]) ? 1 : 0;
assign detect_max[371][11] = (mid_1[2983:2976] > mid_0[2991:2984]) ? 1 : 0;
assign detect_max[371][12] = (mid_1[2983:2976] > mid_1[2975:2968]) ? 1 : 0;
assign detect_max[371][13] = (mid_1[2983:2976] > mid_1[2991:2984]) ? 1 : 0;
assign detect_max[371][14] = (mid_1[2983:2976] > mid_2[2975:2968]) ? 1 : 0;
assign detect_max[371][15] = (mid_1[2983:2976] > mid_2[2983:2976]) ? 1 : 0;
assign detect_max[371][16] = (mid_1[2983:2976] > mid_2[2991:2984]) ? 1 : 0;
assign detect_max[371][17] = (mid_1[2983:2976] > btm_0[2975:2968]) ? 1 : 0;
assign detect_max[371][18] = (mid_1[2983:2976] > btm_0[2983:2976]) ? 1 : 0;
assign detect_max[371][19] = (mid_1[2983:2976] > btm_0[2991:2984]) ? 1 : 0;
assign detect_max[371][20] = (mid_1[2983:2976] > btm_1[2975:2968]) ? 1 : 0;
assign detect_max[371][21] = (mid_1[2983:2976] > btm_1[2983:2976]) ? 1 : 0;
assign detect_max[371][22] = (mid_1[2983:2976] > btm_1[2991:2984]) ? 1 : 0;
assign detect_max[371][23] = (mid_1[2983:2976] > btm_2[2975:2968]) ? 1 : 0;
assign detect_max[371][24] = (mid_1[2983:2976] > btm_2[2983:2976]) ? 1 : 0;
assign detect_max[371][25] = (mid_1[2983:2976] > btm_2[2991:2984]) ? 1 : 0;

assign detect_max[372][0] = (mid_1[2991:2984] > top_0[2983:2976]) ? 1 : 0;
assign detect_max[372][1] = (mid_1[2991:2984] > top_0[2991:2984]) ? 1 : 0;
assign detect_max[372][2] = (mid_1[2991:2984] > top_0[2999:2992]) ? 1 : 0;
assign detect_max[372][3] = (mid_1[2991:2984] > top_1[2983:2976]) ? 1 : 0;
assign detect_max[372][4] = (mid_1[2991:2984] > top_1[2991:2984]) ? 1 : 0;
assign detect_max[372][5] = (mid_1[2991:2984] > top_1[2999:2992]) ? 1 : 0;
assign detect_max[372][6] = (mid_1[2991:2984] > top_2[2983:2976]) ? 1 : 0;
assign detect_max[372][7] = (mid_1[2991:2984] > top_2[2991:2984]) ? 1 : 0;
assign detect_max[372][8] = (mid_1[2991:2984] > top_2[2999:2992]) ? 1 : 0;
assign detect_max[372][9] = (mid_1[2991:2984] > mid_0[2983:2976]) ? 1 : 0;
assign detect_max[372][10] = (mid_1[2991:2984] > mid_0[2991:2984]) ? 1 : 0;
assign detect_max[372][11] = (mid_1[2991:2984] > mid_0[2999:2992]) ? 1 : 0;
assign detect_max[372][12] = (mid_1[2991:2984] > mid_1[2983:2976]) ? 1 : 0;
assign detect_max[372][13] = (mid_1[2991:2984] > mid_1[2999:2992]) ? 1 : 0;
assign detect_max[372][14] = (mid_1[2991:2984] > mid_2[2983:2976]) ? 1 : 0;
assign detect_max[372][15] = (mid_1[2991:2984] > mid_2[2991:2984]) ? 1 : 0;
assign detect_max[372][16] = (mid_1[2991:2984] > mid_2[2999:2992]) ? 1 : 0;
assign detect_max[372][17] = (mid_1[2991:2984] > btm_0[2983:2976]) ? 1 : 0;
assign detect_max[372][18] = (mid_1[2991:2984] > btm_0[2991:2984]) ? 1 : 0;
assign detect_max[372][19] = (mid_1[2991:2984] > btm_0[2999:2992]) ? 1 : 0;
assign detect_max[372][20] = (mid_1[2991:2984] > btm_1[2983:2976]) ? 1 : 0;
assign detect_max[372][21] = (mid_1[2991:2984] > btm_1[2991:2984]) ? 1 : 0;
assign detect_max[372][22] = (mid_1[2991:2984] > btm_1[2999:2992]) ? 1 : 0;
assign detect_max[372][23] = (mid_1[2991:2984] > btm_2[2983:2976]) ? 1 : 0;
assign detect_max[372][24] = (mid_1[2991:2984] > btm_2[2991:2984]) ? 1 : 0;
assign detect_max[372][25] = (mid_1[2991:2984] > btm_2[2999:2992]) ? 1 : 0;

assign detect_max[373][0] = (mid_1[2999:2992] > top_0[2991:2984]) ? 1 : 0;
assign detect_max[373][1] = (mid_1[2999:2992] > top_0[2999:2992]) ? 1 : 0;
assign detect_max[373][2] = (mid_1[2999:2992] > top_0[3007:3000]) ? 1 : 0;
assign detect_max[373][3] = (mid_1[2999:2992] > top_1[2991:2984]) ? 1 : 0;
assign detect_max[373][4] = (mid_1[2999:2992] > top_1[2999:2992]) ? 1 : 0;
assign detect_max[373][5] = (mid_1[2999:2992] > top_1[3007:3000]) ? 1 : 0;
assign detect_max[373][6] = (mid_1[2999:2992] > top_2[2991:2984]) ? 1 : 0;
assign detect_max[373][7] = (mid_1[2999:2992] > top_2[2999:2992]) ? 1 : 0;
assign detect_max[373][8] = (mid_1[2999:2992] > top_2[3007:3000]) ? 1 : 0;
assign detect_max[373][9] = (mid_1[2999:2992] > mid_0[2991:2984]) ? 1 : 0;
assign detect_max[373][10] = (mid_1[2999:2992] > mid_0[2999:2992]) ? 1 : 0;
assign detect_max[373][11] = (mid_1[2999:2992] > mid_0[3007:3000]) ? 1 : 0;
assign detect_max[373][12] = (mid_1[2999:2992] > mid_1[2991:2984]) ? 1 : 0;
assign detect_max[373][13] = (mid_1[2999:2992] > mid_1[3007:3000]) ? 1 : 0;
assign detect_max[373][14] = (mid_1[2999:2992] > mid_2[2991:2984]) ? 1 : 0;
assign detect_max[373][15] = (mid_1[2999:2992] > mid_2[2999:2992]) ? 1 : 0;
assign detect_max[373][16] = (mid_1[2999:2992] > mid_2[3007:3000]) ? 1 : 0;
assign detect_max[373][17] = (mid_1[2999:2992] > btm_0[2991:2984]) ? 1 : 0;
assign detect_max[373][18] = (mid_1[2999:2992] > btm_0[2999:2992]) ? 1 : 0;
assign detect_max[373][19] = (mid_1[2999:2992] > btm_0[3007:3000]) ? 1 : 0;
assign detect_max[373][20] = (mid_1[2999:2992] > btm_1[2991:2984]) ? 1 : 0;
assign detect_max[373][21] = (mid_1[2999:2992] > btm_1[2999:2992]) ? 1 : 0;
assign detect_max[373][22] = (mid_1[2999:2992] > btm_1[3007:3000]) ? 1 : 0;
assign detect_max[373][23] = (mid_1[2999:2992] > btm_2[2991:2984]) ? 1 : 0;
assign detect_max[373][24] = (mid_1[2999:2992] > btm_2[2999:2992]) ? 1 : 0;
assign detect_max[373][25] = (mid_1[2999:2992] > btm_2[3007:3000]) ? 1 : 0;

assign detect_max[374][0] = (mid_1[3007:3000] > top_0[2999:2992]) ? 1 : 0;
assign detect_max[374][1] = (mid_1[3007:3000] > top_0[3007:3000]) ? 1 : 0;
assign detect_max[374][2] = (mid_1[3007:3000] > top_0[3015:3008]) ? 1 : 0;
assign detect_max[374][3] = (mid_1[3007:3000] > top_1[2999:2992]) ? 1 : 0;
assign detect_max[374][4] = (mid_1[3007:3000] > top_1[3007:3000]) ? 1 : 0;
assign detect_max[374][5] = (mid_1[3007:3000] > top_1[3015:3008]) ? 1 : 0;
assign detect_max[374][6] = (mid_1[3007:3000] > top_2[2999:2992]) ? 1 : 0;
assign detect_max[374][7] = (mid_1[3007:3000] > top_2[3007:3000]) ? 1 : 0;
assign detect_max[374][8] = (mid_1[3007:3000] > top_2[3015:3008]) ? 1 : 0;
assign detect_max[374][9] = (mid_1[3007:3000] > mid_0[2999:2992]) ? 1 : 0;
assign detect_max[374][10] = (mid_1[3007:3000] > mid_0[3007:3000]) ? 1 : 0;
assign detect_max[374][11] = (mid_1[3007:3000] > mid_0[3015:3008]) ? 1 : 0;
assign detect_max[374][12] = (mid_1[3007:3000] > mid_1[2999:2992]) ? 1 : 0;
assign detect_max[374][13] = (mid_1[3007:3000] > mid_1[3015:3008]) ? 1 : 0;
assign detect_max[374][14] = (mid_1[3007:3000] > mid_2[2999:2992]) ? 1 : 0;
assign detect_max[374][15] = (mid_1[3007:3000] > mid_2[3007:3000]) ? 1 : 0;
assign detect_max[374][16] = (mid_1[3007:3000] > mid_2[3015:3008]) ? 1 : 0;
assign detect_max[374][17] = (mid_1[3007:3000] > btm_0[2999:2992]) ? 1 : 0;
assign detect_max[374][18] = (mid_1[3007:3000] > btm_0[3007:3000]) ? 1 : 0;
assign detect_max[374][19] = (mid_1[3007:3000] > btm_0[3015:3008]) ? 1 : 0;
assign detect_max[374][20] = (mid_1[3007:3000] > btm_1[2999:2992]) ? 1 : 0;
assign detect_max[374][21] = (mid_1[3007:3000] > btm_1[3007:3000]) ? 1 : 0;
assign detect_max[374][22] = (mid_1[3007:3000] > btm_1[3015:3008]) ? 1 : 0;
assign detect_max[374][23] = (mid_1[3007:3000] > btm_2[2999:2992]) ? 1 : 0;
assign detect_max[374][24] = (mid_1[3007:3000] > btm_2[3007:3000]) ? 1 : 0;
assign detect_max[374][25] = (mid_1[3007:3000] > btm_2[3015:3008]) ? 1 : 0;

assign detect_max[375][0] = (mid_1[3015:3008] > top_0[3007:3000]) ? 1 : 0;
assign detect_max[375][1] = (mid_1[3015:3008] > top_0[3015:3008]) ? 1 : 0;
assign detect_max[375][2] = (mid_1[3015:3008] > top_0[3023:3016]) ? 1 : 0;
assign detect_max[375][3] = (mid_1[3015:3008] > top_1[3007:3000]) ? 1 : 0;
assign detect_max[375][4] = (mid_1[3015:3008] > top_1[3015:3008]) ? 1 : 0;
assign detect_max[375][5] = (mid_1[3015:3008] > top_1[3023:3016]) ? 1 : 0;
assign detect_max[375][6] = (mid_1[3015:3008] > top_2[3007:3000]) ? 1 : 0;
assign detect_max[375][7] = (mid_1[3015:3008] > top_2[3015:3008]) ? 1 : 0;
assign detect_max[375][8] = (mid_1[3015:3008] > top_2[3023:3016]) ? 1 : 0;
assign detect_max[375][9] = (mid_1[3015:3008] > mid_0[3007:3000]) ? 1 : 0;
assign detect_max[375][10] = (mid_1[3015:3008] > mid_0[3015:3008]) ? 1 : 0;
assign detect_max[375][11] = (mid_1[3015:3008] > mid_0[3023:3016]) ? 1 : 0;
assign detect_max[375][12] = (mid_1[3015:3008] > mid_1[3007:3000]) ? 1 : 0;
assign detect_max[375][13] = (mid_1[3015:3008] > mid_1[3023:3016]) ? 1 : 0;
assign detect_max[375][14] = (mid_1[3015:3008] > mid_2[3007:3000]) ? 1 : 0;
assign detect_max[375][15] = (mid_1[3015:3008] > mid_2[3015:3008]) ? 1 : 0;
assign detect_max[375][16] = (mid_1[3015:3008] > mid_2[3023:3016]) ? 1 : 0;
assign detect_max[375][17] = (mid_1[3015:3008] > btm_0[3007:3000]) ? 1 : 0;
assign detect_max[375][18] = (mid_1[3015:3008] > btm_0[3015:3008]) ? 1 : 0;
assign detect_max[375][19] = (mid_1[3015:3008] > btm_0[3023:3016]) ? 1 : 0;
assign detect_max[375][20] = (mid_1[3015:3008] > btm_1[3007:3000]) ? 1 : 0;
assign detect_max[375][21] = (mid_1[3015:3008] > btm_1[3015:3008]) ? 1 : 0;
assign detect_max[375][22] = (mid_1[3015:3008] > btm_1[3023:3016]) ? 1 : 0;
assign detect_max[375][23] = (mid_1[3015:3008] > btm_2[3007:3000]) ? 1 : 0;
assign detect_max[375][24] = (mid_1[3015:3008] > btm_2[3015:3008]) ? 1 : 0;
assign detect_max[375][25] = (mid_1[3015:3008] > btm_2[3023:3016]) ? 1 : 0;

assign detect_max[376][0] = (mid_1[3023:3016] > top_0[3015:3008]) ? 1 : 0;
assign detect_max[376][1] = (mid_1[3023:3016] > top_0[3023:3016]) ? 1 : 0;
assign detect_max[376][2] = (mid_1[3023:3016] > top_0[3031:3024]) ? 1 : 0;
assign detect_max[376][3] = (mid_1[3023:3016] > top_1[3015:3008]) ? 1 : 0;
assign detect_max[376][4] = (mid_1[3023:3016] > top_1[3023:3016]) ? 1 : 0;
assign detect_max[376][5] = (mid_1[3023:3016] > top_1[3031:3024]) ? 1 : 0;
assign detect_max[376][6] = (mid_1[3023:3016] > top_2[3015:3008]) ? 1 : 0;
assign detect_max[376][7] = (mid_1[3023:3016] > top_2[3023:3016]) ? 1 : 0;
assign detect_max[376][8] = (mid_1[3023:3016] > top_2[3031:3024]) ? 1 : 0;
assign detect_max[376][9] = (mid_1[3023:3016] > mid_0[3015:3008]) ? 1 : 0;
assign detect_max[376][10] = (mid_1[3023:3016] > mid_0[3023:3016]) ? 1 : 0;
assign detect_max[376][11] = (mid_1[3023:3016] > mid_0[3031:3024]) ? 1 : 0;
assign detect_max[376][12] = (mid_1[3023:3016] > mid_1[3015:3008]) ? 1 : 0;
assign detect_max[376][13] = (mid_1[3023:3016] > mid_1[3031:3024]) ? 1 : 0;
assign detect_max[376][14] = (mid_1[3023:3016] > mid_2[3015:3008]) ? 1 : 0;
assign detect_max[376][15] = (mid_1[3023:3016] > mid_2[3023:3016]) ? 1 : 0;
assign detect_max[376][16] = (mid_1[3023:3016] > mid_2[3031:3024]) ? 1 : 0;
assign detect_max[376][17] = (mid_1[3023:3016] > btm_0[3015:3008]) ? 1 : 0;
assign detect_max[376][18] = (mid_1[3023:3016] > btm_0[3023:3016]) ? 1 : 0;
assign detect_max[376][19] = (mid_1[3023:3016] > btm_0[3031:3024]) ? 1 : 0;
assign detect_max[376][20] = (mid_1[3023:3016] > btm_1[3015:3008]) ? 1 : 0;
assign detect_max[376][21] = (mid_1[3023:3016] > btm_1[3023:3016]) ? 1 : 0;
assign detect_max[376][22] = (mid_1[3023:3016] > btm_1[3031:3024]) ? 1 : 0;
assign detect_max[376][23] = (mid_1[3023:3016] > btm_2[3015:3008]) ? 1 : 0;
assign detect_max[376][24] = (mid_1[3023:3016] > btm_2[3023:3016]) ? 1 : 0;
assign detect_max[376][25] = (mid_1[3023:3016] > btm_2[3031:3024]) ? 1 : 0;

assign detect_max[377][0] = (mid_1[3031:3024] > top_0[3023:3016]) ? 1 : 0;
assign detect_max[377][1] = (mid_1[3031:3024] > top_0[3031:3024]) ? 1 : 0;
assign detect_max[377][2] = (mid_1[3031:3024] > top_0[3039:3032]) ? 1 : 0;
assign detect_max[377][3] = (mid_1[3031:3024] > top_1[3023:3016]) ? 1 : 0;
assign detect_max[377][4] = (mid_1[3031:3024] > top_1[3031:3024]) ? 1 : 0;
assign detect_max[377][5] = (mid_1[3031:3024] > top_1[3039:3032]) ? 1 : 0;
assign detect_max[377][6] = (mid_1[3031:3024] > top_2[3023:3016]) ? 1 : 0;
assign detect_max[377][7] = (mid_1[3031:3024] > top_2[3031:3024]) ? 1 : 0;
assign detect_max[377][8] = (mid_1[3031:3024] > top_2[3039:3032]) ? 1 : 0;
assign detect_max[377][9] = (mid_1[3031:3024] > mid_0[3023:3016]) ? 1 : 0;
assign detect_max[377][10] = (mid_1[3031:3024] > mid_0[3031:3024]) ? 1 : 0;
assign detect_max[377][11] = (mid_1[3031:3024] > mid_0[3039:3032]) ? 1 : 0;
assign detect_max[377][12] = (mid_1[3031:3024] > mid_1[3023:3016]) ? 1 : 0;
assign detect_max[377][13] = (mid_1[3031:3024] > mid_1[3039:3032]) ? 1 : 0;
assign detect_max[377][14] = (mid_1[3031:3024] > mid_2[3023:3016]) ? 1 : 0;
assign detect_max[377][15] = (mid_1[3031:3024] > mid_2[3031:3024]) ? 1 : 0;
assign detect_max[377][16] = (mid_1[3031:3024] > mid_2[3039:3032]) ? 1 : 0;
assign detect_max[377][17] = (mid_1[3031:3024] > btm_0[3023:3016]) ? 1 : 0;
assign detect_max[377][18] = (mid_1[3031:3024] > btm_0[3031:3024]) ? 1 : 0;
assign detect_max[377][19] = (mid_1[3031:3024] > btm_0[3039:3032]) ? 1 : 0;
assign detect_max[377][20] = (mid_1[3031:3024] > btm_1[3023:3016]) ? 1 : 0;
assign detect_max[377][21] = (mid_1[3031:3024] > btm_1[3031:3024]) ? 1 : 0;
assign detect_max[377][22] = (mid_1[3031:3024] > btm_1[3039:3032]) ? 1 : 0;
assign detect_max[377][23] = (mid_1[3031:3024] > btm_2[3023:3016]) ? 1 : 0;
assign detect_max[377][24] = (mid_1[3031:3024] > btm_2[3031:3024]) ? 1 : 0;
assign detect_max[377][25] = (mid_1[3031:3024] > btm_2[3039:3032]) ? 1 : 0;

assign detect_max[378][0] = (mid_1[3039:3032] > top_0[3031:3024]) ? 1 : 0;
assign detect_max[378][1] = (mid_1[3039:3032] > top_0[3039:3032]) ? 1 : 0;
assign detect_max[378][2] = (mid_1[3039:3032] > top_0[3047:3040]) ? 1 : 0;
assign detect_max[378][3] = (mid_1[3039:3032] > top_1[3031:3024]) ? 1 : 0;
assign detect_max[378][4] = (mid_1[3039:3032] > top_1[3039:3032]) ? 1 : 0;
assign detect_max[378][5] = (mid_1[3039:3032] > top_1[3047:3040]) ? 1 : 0;
assign detect_max[378][6] = (mid_1[3039:3032] > top_2[3031:3024]) ? 1 : 0;
assign detect_max[378][7] = (mid_1[3039:3032] > top_2[3039:3032]) ? 1 : 0;
assign detect_max[378][8] = (mid_1[3039:3032] > top_2[3047:3040]) ? 1 : 0;
assign detect_max[378][9] = (mid_1[3039:3032] > mid_0[3031:3024]) ? 1 : 0;
assign detect_max[378][10] = (mid_1[3039:3032] > mid_0[3039:3032]) ? 1 : 0;
assign detect_max[378][11] = (mid_1[3039:3032] > mid_0[3047:3040]) ? 1 : 0;
assign detect_max[378][12] = (mid_1[3039:3032] > mid_1[3031:3024]) ? 1 : 0;
assign detect_max[378][13] = (mid_1[3039:3032] > mid_1[3047:3040]) ? 1 : 0;
assign detect_max[378][14] = (mid_1[3039:3032] > mid_2[3031:3024]) ? 1 : 0;
assign detect_max[378][15] = (mid_1[3039:3032] > mid_2[3039:3032]) ? 1 : 0;
assign detect_max[378][16] = (mid_1[3039:3032] > mid_2[3047:3040]) ? 1 : 0;
assign detect_max[378][17] = (mid_1[3039:3032] > btm_0[3031:3024]) ? 1 : 0;
assign detect_max[378][18] = (mid_1[3039:3032] > btm_0[3039:3032]) ? 1 : 0;
assign detect_max[378][19] = (mid_1[3039:3032] > btm_0[3047:3040]) ? 1 : 0;
assign detect_max[378][20] = (mid_1[3039:3032] > btm_1[3031:3024]) ? 1 : 0;
assign detect_max[378][21] = (mid_1[3039:3032] > btm_1[3039:3032]) ? 1 : 0;
assign detect_max[378][22] = (mid_1[3039:3032] > btm_1[3047:3040]) ? 1 : 0;
assign detect_max[378][23] = (mid_1[3039:3032] > btm_2[3031:3024]) ? 1 : 0;
assign detect_max[378][24] = (mid_1[3039:3032] > btm_2[3039:3032]) ? 1 : 0;
assign detect_max[378][25] = (mid_1[3039:3032] > btm_2[3047:3040]) ? 1 : 0;

assign detect_max[379][0] = (mid_1[3047:3040] > top_0[3039:3032]) ? 1 : 0;
assign detect_max[379][1] = (mid_1[3047:3040] > top_0[3047:3040]) ? 1 : 0;
assign detect_max[379][2] = (mid_1[3047:3040] > top_0[3055:3048]) ? 1 : 0;
assign detect_max[379][3] = (mid_1[3047:3040] > top_1[3039:3032]) ? 1 : 0;
assign detect_max[379][4] = (mid_1[3047:3040] > top_1[3047:3040]) ? 1 : 0;
assign detect_max[379][5] = (mid_1[3047:3040] > top_1[3055:3048]) ? 1 : 0;
assign detect_max[379][6] = (mid_1[3047:3040] > top_2[3039:3032]) ? 1 : 0;
assign detect_max[379][7] = (mid_1[3047:3040] > top_2[3047:3040]) ? 1 : 0;
assign detect_max[379][8] = (mid_1[3047:3040] > top_2[3055:3048]) ? 1 : 0;
assign detect_max[379][9] = (mid_1[3047:3040] > mid_0[3039:3032]) ? 1 : 0;
assign detect_max[379][10] = (mid_1[3047:3040] > mid_0[3047:3040]) ? 1 : 0;
assign detect_max[379][11] = (mid_1[3047:3040] > mid_0[3055:3048]) ? 1 : 0;
assign detect_max[379][12] = (mid_1[3047:3040] > mid_1[3039:3032]) ? 1 : 0;
assign detect_max[379][13] = (mid_1[3047:3040] > mid_1[3055:3048]) ? 1 : 0;
assign detect_max[379][14] = (mid_1[3047:3040] > mid_2[3039:3032]) ? 1 : 0;
assign detect_max[379][15] = (mid_1[3047:3040] > mid_2[3047:3040]) ? 1 : 0;
assign detect_max[379][16] = (mid_1[3047:3040] > mid_2[3055:3048]) ? 1 : 0;
assign detect_max[379][17] = (mid_1[3047:3040] > btm_0[3039:3032]) ? 1 : 0;
assign detect_max[379][18] = (mid_1[3047:3040] > btm_0[3047:3040]) ? 1 : 0;
assign detect_max[379][19] = (mid_1[3047:3040] > btm_0[3055:3048]) ? 1 : 0;
assign detect_max[379][20] = (mid_1[3047:3040] > btm_1[3039:3032]) ? 1 : 0;
assign detect_max[379][21] = (mid_1[3047:3040] > btm_1[3047:3040]) ? 1 : 0;
assign detect_max[379][22] = (mid_1[3047:3040] > btm_1[3055:3048]) ? 1 : 0;
assign detect_max[379][23] = (mid_1[3047:3040] > btm_2[3039:3032]) ? 1 : 0;
assign detect_max[379][24] = (mid_1[3047:3040] > btm_2[3047:3040]) ? 1 : 0;
assign detect_max[379][25] = (mid_1[3047:3040] > btm_2[3055:3048]) ? 1 : 0;

assign detect_max[380][0] = (mid_1[3055:3048] > top_0[3047:3040]) ? 1 : 0;
assign detect_max[380][1] = (mid_1[3055:3048] > top_0[3055:3048]) ? 1 : 0;
assign detect_max[380][2] = (mid_1[3055:3048] > top_0[3063:3056]) ? 1 : 0;
assign detect_max[380][3] = (mid_1[3055:3048] > top_1[3047:3040]) ? 1 : 0;
assign detect_max[380][4] = (mid_1[3055:3048] > top_1[3055:3048]) ? 1 : 0;
assign detect_max[380][5] = (mid_1[3055:3048] > top_1[3063:3056]) ? 1 : 0;
assign detect_max[380][6] = (mid_1[3055:3048] > top_2[3047:3040]) ? 1 : 0;
assign detect_max[380][7] = (mid_1[3055:3048] > top_2[3055:3048]) ? 1 : 0;
assign detect_max[380][8] = (mid_1[3055:3048] > top_2[3063:3056]) ? 1 : 0;
assign detect_max[380][9] = (mid_1[3055:3048] > mid_0[3047:3040]) ? 1 : 0;
assign detect_max[380][10] = (mid_1[3055:3048] > mid_0[3055:3048]) ? 1 : 0;
assign detect_max[380][11] = (mid_1[3055:3048] > mid_0[3063:3056]) ? 1 : 0;
assign detect_max[380][12] = (mid_1[3055:3048] > mid_1[3047:3040]) ? 1 : 0;
assign detect_max[380][13] = (mid_1[3055:3048] > mid_1[3063:3056]) ? 1 : 0;
assign detect_max[380][14] = (mid_1[3055:3048] > mid_2[3047:3040]) ? 1 : 0;
assign detect_max[380][15] = (mid_1[3055:3048] > mid_2[3055:3048]) ? 1 : 0;
assign detect_max[380][16] = (mid_1[3055:3048] > mid_2[3063:3056]) ? 1 : 0;
assign detect_max[380][17] = (mid_1[3055:3048] > btm_0[3047:3040]) ? 1 : 0;
assign detect_max[380][18] = (mid_1[3055:3048] > btm_0[3055:3048]) ? 1 : 0;
assign detect_max[380][19] = (mid_1[3055:3048] > btm_0[3063:3056]) ? 1 : 0;
assign detect_max[380][20] = (mid_1[3055:3048] > btm_1[3047:3040]) ? 1 : 0;
assign detect_max[380][21] = (mid_1[3055:3048] > btm_1[3055:3048]) ? 1 : 0;
assign detect_max[380][22] = (mid_1[3055:3048] > btm_1[3063:3056]) ? 1 : 0;
assign detect_max[380][23] = (mid_1[3055:3048] > btm_2[3047:3040]) ? 1 : 0;
assign detect_max[380][24] = (mid_1[3055:3048] > btm_2[3055:3048]) ? 1 : 0;
assign detect_max[380][25] = (mid_1[3055:3048] > btm_2[3063:3056]) ? 1 : 0;

assign detect_max[381][0] = (mid_1[3063:3056] > top_0[3055:3048]) ? 1 : 0;
assign detect_max[381][1] = (mid_1[3063:3056] > top_0[3063:3056]) ? 1 : 0;
assign detect_max[381][2] = (mid_1[3063:3056] > top_0[3071:3064]) ? 1 : 0;
assign detect_max[381][3] = (mid_1[3063:3056] > top_1[3055:3048]) ? 1 : 0;
assign detect_max[381][4] = (mid_1[3063:3056] > top_1[3063:3056]) ? 1 : 0;
assign detect_max[381][5] = (mid_1[3063:3056] > top_1[3071:3064]) ? 1 : 0;
assign detect_max[381][6] = (mid_1[3063:3056] > top_2[3055:3048]) ? 1 : 0;
assign detect_max[381][7] = (mid_1[3063:3056] > top_2[3063:3056]) ? 1 : 0;
assign detect_max[381][8] = (mid_1[3063:3056] > top_2[3071:3064]) ? 1 : 0;
assign detect_max[381][9] = (mid_1[3063:3056] > mid_0[3055:3048]) ? 1 : 0;
assign detect_max[381][10] = (mid_1[3063:3056] > mid_0[3063:3056]) ? 1 : 0;
assign detect_max[381][11] = (mid_1[3063:3056] > mid_0[3071:3064]) ? 1 : 0;
assign detect_max[381][12] = (mid_1[3063:3056] > mid_1[3055:3048]) ? 1 : 0;
assign detect_max[381][13] = (mid_1[3063:3056] > mid_1[3071:3064]) ? 1 : 0;
assign detect_max[381][14] = (mid_1[3063:3056] > mid_2[3055:3048]) ? 1 : 0;
assign detect_max[381][15] = (mid_1[3063:3056] > mid_2[3063:3056]) ? 1 : 0;
assign detect_max[381][16] = (mid_1[3063:3056] > mid_2[3071:3064]) ? 1 : 0;
assign detect_max[381][17] = (mid_1[3063:3056] > btm_0[3055:3048]) ? 1 : 0;
assign detect_max[381][18] = (mid_1[3063:3056] > btm_0[3063:3056]) ? 1 : 0;
assign detect_max[381][19] = (mid_1[3063:3056] > btm_0[3071:3064]) ? 1 : 0;
assign detect_max[381][20] = (mid_1[3063:3056] > btm_1[3055:3048]) ? 1 : 0;
assign detect_max[381][21] = (mid_1[3063:3056] > btm_1[3063:3056]) ? 1 : 0;
assign detect_max[381][22] = (mid_1[3063:3056] > btm_1[3071:3064]) ? 1 : 0;
assign detect_max[381][23] = (mid_1[3063:3056] > btm_2[3055:3048]) ? 1 : 0;
assign detect_max[381][24] = (mid_1[3063:3056] > btm_2[3063:3056]) ? 1 : 0;
assign detect_max[381][25] = (mid_1[3063:3056] > btm_2[3071:3064]) ? 1 : 0;

assign detect_max[382][0] = (mid_1[3071:3064] > top_0[3063:3056]) ? 1 : 0;
assign detect_max[382][1] = (mid_1[3071:3064] > top_0[3071:3064]) ? 1 : 0;
assign detect_max[382][2] = (mid_1[3071:3064] > top_0[3079:3072]) ? 1 : 0;
assign detect_max[382][3] = (mid_1[3071:3064] > top_1[3063:3056]) ? 1 : 0;
assign detect_max[382][4] = (mid_1[3071:3064] > top_1[3071:3064]) ? 1 : 0;
assign detect_max[382][5] = (mid_1[3071:3064] > top_1[3079:3072]) ? 1 : 0;
assign detect_max[382][6] = (mid_1[3071:3064] > top_2[3063:3056]) ? 1 : 0;
assign detect_max[382][7] = (mid_1[3071:3064] > top_2[3071:3064]) ? 1 : 0;
assign detect_max[382][8] = (mid_1[3071:3064] > top_2[3079:3072]) ? 1 : 0;
assign detect_max[382][9] = (mid_1[3071:3064] > mid_0[3063:3056]) ? 1 : 0;
assign detect_max[382][10] = (mid_1[3071:3064] > mid_0[3071:3064]) ? 1 : 0;
assign detect_max[382][11] = (mid_1[3071:3064] > mid_0[3079:3072]) ? 1 : 0;
assign detect_max[382][12] = (mid_1[3071:3064] > mid_1[3063:3056]) ? 1 : 0;
assign detect_max[382][13] = (mid_1[3071:3064] > mid_1[3079:3072]) ? 1 : 0;
assign detect_max[382][14] = (mid_1[3071:3064] > mid_2[3063:3056]) ? 1 : 0;
assign detect_max[382][15] = (mid_1[3071:3064] > mid_2[3071:3064]) ? 1 : 0;
assign detect_max[382][16] = (mid_1[3071:3064] > mid_2[3079:3072]) ? 1 : 0;
assign detect_max[382][17] = (mid_1[3071:3064] > btm_0[3063:3056]) ? 1 : 0;
assign detect_max[382][18] = (mid_1[3071:3064] > btm_0[3071:3064]) ? 1 : 0;
assign detect_max[382][19] = (mid_1[3071:3064] > btm_0[3079:3072]) ? 1 : 0;
assign detect_max[382][20] = (mid_1[3071:3064] > btm_1[3063:3056]) ? 1 : 0;
assign detect_max[382][21] = (mid_1[3071:3064] > btm_1[3071:3064]) ? 1 : 0;
assign detect_max[382][22] = (mid_1[3071:3064] > btm_1[3079:3072]) ? 1 : 0;
assign detect_max[382][23] = (mid_1[3071:3064] > btm_2[3063:3056]) ? 1 : 0;
assign detect_max[382][24] = (mid_1[3071:3064] > btm_2[3071:3064]) ? 1 : 0;
assign detect_max[382][25] = (mid_1[3071:3064] > btm_2[3079:3072]) ? 1 : 0;

assign detect_max[383][0] = (mid_1[3079:3072] > top_0[3071:3064]) ? 1 : 0;
assign detect_max[383][1] = (mid_1[3079:3072] > top_0[3079:3072]) ? 1 : 0;
assign detect_max[383][2] = (mid_1[3079:3072] > top_0[3087:3080]) ? 1 : 0;
assign detect_max[383][3] = (mid_1[3079:3072] > top_1[3071:3064]) ? 1 : 0;
assign detect_max[383][4] = (mid_1[3079:3072] > top_1[3079:3072]) ? 1 : 0;
assign detect_max[383][5] = (mid_1[3079:3072] > top_1[3087:3080]) ? 1 : 0;
assign detect_max[383][6] = (mid_1[3079:3072] > top_2[3071:3064]) ? 1 : 0;
assign detect_max[383][7] = (mid_1[3079:3072] > top_2[3079:3072]) ? 1 : 0;
assign detect_max[383][8] = (mid_1[3079:3072] > top_2[3087:3080]) ? 1 : 0;
assign detect_max[383][9] = (mid_1[3079:3072] > mid_0[3071:3064]) ? 1 : 0;
assign detect_max[383][10] = (mid_1[3079:3072] > mid_0[3079:3072]) ? 1 : 0;
assign detect_max[383][11] = (mid_1[3079:3072] > mid_0[3087:3080]) ? 1 : 0;
assign detect_max[383][12] = (mid_1[3079:3072] > mid_1[3071:3064]) ? 1 : 0;
assign detect_max[383][13] = (mid_1[3079:3072] > mid_1[3087:3080]) ? 1 : 0;
assign detect_max[383][14] = (mid_1[3079:3072] > mid_2[3071:3064]) ? 1 : 0;
assign detect_max[383][15] = (mid_1[3079:3072] > mid_2[3079:3072]) ? 1 : 0;
assign detect_max[383][16] = (mid_1[3079:3072] > mid_2[3087:3080]) ? 1 : 0;
assign detect_max[383][17] = (mid_1[3079:3072] > btm_0[3071:3064]) ? 1 : 0;
assign detect_max[383][18] = (mid_1[3079:3072] > btm_0[3079:3072]) ? 1 : 0;
assign detect_max[383][19] = (mid_1[3079:3072] > btm_0[3087:3080]) ? 1 : 0;
assign detect_max[383][20] = (mid_1[3079:3072] > btm_1[3071:3064]) ? 1 : 0;
assign detect_max[383][21] = (mid_1[3079:3072] > btm_1[3079:3072]) ? 1 : 0;
assign detect_max[383][22] = (mid_1[3079:3072] > btm_1[3087:3080]) ? 1 : 0;
assign detect_max[383][23] = (mid_1[3079:3072] > btm_2[3071:3064]) ? 1 : 0;
assign detect_max[383][24] = (mid_1[3079:3072] > btm_2[3079:3072]) ? 1 : 0;
assign detect_max[383][25] = (mid_1[3079:3072] > btm_2[3087:3080]) ? 1 : 0;

assign detect_max[384][0] = (mid_1[3087:3080] > top_0[3079:3072]) ? 1 : 0;
assign detect_max[384][1] = (mid_1[3087:3080] > top_0[3087:3080]) ? 1 : 0;
assign detect_max[384][2] = (mid_1[3087:3080] > top_0[3095:3088]) ? 1 : 0;
assign detect_max[384][3] = (mid_1[3087:3080] > top_1[3079:3072]) ? 1 : 0;
assign detect_max[384][4] = (mid_1[3087:3080] > top_1[3087:3080]) ? 1 : 0;
assign detect_max[384][5] = (mid_1[3087:3080] > top_1[3095:3088]) ? 1 : 0;
assign detect_max[384][6] = (mid_1[3087:3080] > top_2[3079:3072]) ? 1 : 0;
assign detect_max[384][7] = (mid_1[3087:3080] > top_2[3087:3080]) ? 1 : 0;
assign detect_max[384][8] = (mid_1[3087:3080] > top_2[3095:3088]) ? 1 : 0;
assign detect_max[384][9] = (mid_1[3087:3080] > mid_0[3079:3072]) ? 1 : 0;
assign detect_max[384][10] = (mid_1[3087:3080] > mid_0[3087:3080]) ? 1 : 0;
assign detect_max[384][11] = (mid_1[3087:3080] > mid_0[3095:3088]) ? 1 : 0;
assign detect_max[384][12] = (mid_1[3087:3080] > mid_1[3079:3072]) ? 1 : 0;
assign detect_max[384][13] = (mid_1[3087:3080] > mid_1[3095:3088]) ? 1 : 0;
assign detect_max[384][14] = (mid_1[3087:3080] > mid_2[3079:3072]) ? 1 : 0;
assign detect_max[384][15] = (mid_1[3087:3080] > mid_2[3087:3080]) ? 1 : 0;
assign detect_max[384][16] = (mid_1[3087:3080] > mid_2[3095:3088]) ? 1 : 0;
assign detect_max[384][17] = (mid_1[3087:3080] > btm_0[3079:3072]) ? 1 : 0;
assign detect_max[384][18] = (mid_1[3087:3080] > btm_0[3087:3080]) ? 1 : 0;
assign detect_max[384][19] = (mid_1[3087:3080] > btm_0[3095:3088]) ? 1 : 0;
assign detect_max[384][20] = (mid_1[3087:3080] > btm_1[3079:3072]) ? 1 : 0;
assign detect_max[384][21] = (mid_1[3087:3080] > btm_1[3087:3080]) ? 1 : 0;
assign detect_max[384][22] = (mid_1[3087:3080] > btm_1[3095:3088]) ? 1 : 0;
assign detect_max[384][23] = (mid_1[3087:3080] > btm_2[3079:3072]) ? 1 : 0;
assign detect_max[384][24] = (mid_1[3087:3080] > btm_2[3087:3080]) ? 1 : 0;
assign detect_max[384][25] = (mid_1[3087:3080] > btm_2[3095:3088]) ? 1 : 0;

assign detect_max[385][0] = (mid_1[3095:3088] > top_0[3087:3080]) ? 1 : 0;
assign detect_max[385][1] = (mid_1[3095:3088] > top_0[3095:3088]) ? 1 : 0;
assign detect_max[385][2] = (mid_1[3095:3088] > top_0[3103:3096]) ? 1 : 0;
assign detect_max[385][3] = (mid_1[3095:3088] > top_1[3087:3080]) ? 1 : 0;
assign detect_max[385][4] = (mid_1[3095:3088] > top_1[3095:3088]) ? 1 : 0;
assign detect_max[385][5] = (mid_1[3095:3088] > top_1[3103:3096]) ? 1 : 0;
assign detect_max[385][6] = (mid_1[3095:3088] > top_2[3087:3080]) ? 1 : 0;
assign detect_max[385][7] = (mid_1[3095:3088] > top_2[3095:3088]) ? 1 : 0;
assign detect_max[385][8] = (mid_1[3095:3088] > top_2[3103:3096]) ? 1 : 0;
assign detect_max[385][9] = (mid_1[3095:3088] > mid_0[3087:3080]) ? 1 : 0;
assign detect_max[385][10] = (mid_1[3095:3088] > mid_0[3095:3088]) ? 1 : 0;
assign detect_max[385][11] = (mid_1[3095:3088] > mid_0[3103:3096]) ? 1 : 0;
assign detect_max[385][12] = (mid_1[3095:3088] > mid_1[3087:3080]) ? 1 : 0;
assign detect_max[385][13] = (mid_1[3095:3088] > mid_1[3103:3096]) ? 1 : 0;
assign detect_max[385][14] = (mid_1[3095:3088] > mid_2[3087:3080]) ? 1 : 0;
assign detect_max[385][15] = (mid_1[3095:3088] > mid_2[3095:3088]) ? 1 : 0;
assign detect_max[385][16] = (mid_1[3095:3088] > mid_2[3103:3096]) ? 1 : 0;
assign detect_max[385][17] = (mid_1[3095:3088] > btm_0[3087:3080]) ? 1 : 0;
assign detect_max[385][18] = (mid_1[3095:3088] > btm_0[3095:3088]) ? 1 : 0;
assign detect_max[385][19] = (mid_1[3095:3088] > btm_0[3103:3096]) ? 1 : 0;
assign detect_max[385][20] = (mid_1[3095:3088] > btm_1[3087:3080]) ? 1 : 0;
assign detect_max[385][21] = (mid_1[3095:3088] > btm_1[3095:3088]) ? 1 : 0;
assign detect_max[385][22] = (mid_1[3095:3088] > btm_1[3103:3096]) ? 1 : 0;
assign detect_max[385][23] = (mid_1[3095:3088] > btm_2[3087:3080]) ? 1 : 0;
assign detect_max[385][24] = (mid_1[3095:3088] > btm_2[3095:3088]) ? 1 : 0;
assign detect_max[385][25] = (mid_1[3095:3088] > btm_2[3103:3096]) ? 1 : 0;

assign detect_max[386][0] = (mid_1[3103:3096] > top_0[3095:3088]) ? 1 : 0;
assign detect_max[386][1] = (mid_1[3103:3096] > top_0[3103:3096]) ? 1 : 0;
assign detect_max[386][2] = (mid_1[3103:3096] > top_0[3111:3104]) ? 1 : 0;
assign detect_max[386][3] = (mid_1[3103:3096] > top_1[3095:3088]) ? 1 : 0;
assign detect_max[386][4] = (mid_1[3103:3096] > top_1[3103:3096]) ? 1 : 0;
assign detect_max[386][5] = (mid_1[3103:3096] > top_1[3111:3104]) ? 1 : 0;
assign detect_max[386][6] = (mid_1[3103:3096] > top_2[3095:3088]) ? 1 : 0;
assign detect_max[386][7] = (mid_1[3103:3096] > top_2[3103:3096]) ? 1 : 0;
assign detect_max[386][8] = (mid_1[3103:3096] > top_2[3111:3104]) ? 1 : 0;
assign detect_max[386][9] = (mid_1[3103:3096] > mid_0[3095:3088]) ? 1 : 0;
assign detect_max[386][10] = (mid_1[3103:3096] > mid_0[3103:3096]) ? 1 : 0;
assign detect_max[386][11] = (mid_1[3103:3096] > mid_0[3111:3104]) ? 1 : 0;
assign detect_max[386][12] = (mid_1[3103:3096] > mid_1[3095:3088]) ? 1 : 0;
assign detect_max[386][13] = (mid_1[3103:3096] > mid_1[3111:3104]) ? 1 : 0;
assign detect_max[386][14] = (mid_1[3103:3096] > mid_2[3095:3088]) ? 1 : 0;
assign detect_max[386][15] = (mid_1[3103:3096] > mid_2[3103:3096]) ? 1 : 0;
assign detect_max[386][16] = (mid_1[3103:3096] > mid_2[3111:3104]) ? 1 : 0;
assign detect_max[386][17] = (mid_1[3103:3096] > btm_0[3095:3088]) ? 1 : 0;
assign detect_max[386][18] = (mid_1[3103:3096] > btm_0[3103:3096]) ? 1 : 0;
assign detect_max[386][19] = (mid_1[3103:3096] > btm_0[3111:3104]) ? 1 : 0;
assign detect_max[386][20] = (mid_1[3103:3096] > btm_1[3095:3088]) ? 1 : 0;
assign detect_max[386][21] = (mid_1[3103:3096] > btm_1[3103:3096]) ? 1 : 0;
assign detect_max[386][22] = (mid_1[3103:3096] > btm_1[3111:3104]) ? 1 : 0;
assign detect_max[386][23] = (mid_1[3103:3096] > btm_2[3095:3088]) ? 1 : 0;
assign detect_max[386][24] = (mid_1[3103:3096] > btm_2[3103:3096]) ? 1 : 0;
assign detect_max[386][25] = (mid_1[3103:3096] > btm_2[3111:3104]) ? 1 : 0;

assign detect_max[387][0] = (mid_1[3111:3104] > top_0[3103:3096]) ? 1 : 0;
assign detect_max[387][1] = (mid_1[3111:3104] > top_0[3111:3104]) ? 1 : 0;
assign detect_max[387][2] = (mid_1[3111:3104] > top_0[3119:3112]) ? 1 : 0;
assign detect_max[387][3] = (mid_1[3111:3104] > top_1[3103:3096]) ? 1 : 0;
assign detect_max[387][4] = (mid_1[3111:3104] > top_1[3111:3104]) ? 1 : 0;
assign detect_max[387][5] = (mid_1[3111:3104] > top_1[3119:3112]) ? 1 : 0;
assign detect_max[387][6] = (mid_1[3111:3104] > top_2[3103:3096]) ? 1 : 0;
assign detect_max[387][7] = (mid_1[3111:3104] > top_2[3111:3104]) ? 1 : 0;
assign detect_max[387][8] = (mid_1[3111:3104] > top_2[3119:3112]) ? 1 : 0;
assign detect_max[387][9] = (mid_1[3111:3104] > mid_0[3103:3096]) ? 1 : 0;
assign detect_max[387][10] = (mid_1[3111:3104] > mid_0[3111:3104]) ? 1 : 0;
assign detect_max[387][11] = (mid_1[3111:3104] > mid_0[3119:3112]) ? 1 : 0;
assign detect_max[387][12] = (mid_1[3111:3104] > mid_1[3103:3096]) ? 1 : 0;
assign detect_max[387][13] = (mid_1[3111:3104] > mid_1[3119:3112]) ? 1 : 0;
assign detect_max[387][14] = (mid_1[3111:3104] > mid_2[3103:3096]) ? 1 : 0;
assign detect_max[387][15] = (mid_1[3111:3104] > mid_2[3111:3104]) ? 1 : 0;
assign detect_max[387][16] = (mid_1[3111:3104] > mid_2[3119:3112]) ? 1 : 0;
assign detect_max[387][17] = (mid_1[3111:3104] > btm_0[3103:3096]) ? 1 : 0;
assign detect_max[387][18] = (mid_1[3111:3104] > btm_0[3111:3104]) ? 1 : 0;
assign detect_max[387][19] = (mid_1[3111:3104] > btm_0[3119:3112]) ? 1 : 0;
assign detect_max[387][20] = (mid_1[3111:3104] > btm_1[3103:3096]) ? 1 : 0;
assign detect_max[387][21] = (mid_1[3111:3104] > btm_1[3111:3104]) ? 1 : 0;
assign detect_max[387][22] = (mid_1[3111:3104] > btm_1[3119:3112]) ? 1 : 0;
assign detect_max[387][23] = (mid_1[3111:3104] > btm_2[3103:3096]) ? 1 : 0;
assign detect_max[387][24] = (mid_1[3111:3104] > btm_2[3111:3104]) ? 1 : 0;
assign detect_max[387][25] = (mid_1[3111:3104] > btm_2[3119:3112]) ? 1 : 0;

assign detect_max[388][0] = (mid_1[3119:3112] > top_0[3111:3104]) ? 1 : 0;
assign detect_max[388][1] = (mid_1[3119:3112] > top_0[3119:3112]) ? 1 : 0;
assign detect_max[388][2] = (mid_1[3119:3112] > top_0[3127:3120]) ? 1 : 0;
assign detect_max[388][3] = (mid_1[3119:3112] > top_1[3111:3104]) ? 1 : 0;
assign detect_max[388][4] = (mid_1[3119:3112] > top_1[3119:3112]) ? 1 : 0;
assign detect_max[388][5] = (mid_1[3119:3112] > top_1[3127:3120]) ? 1 : 0;
assign detect_max[388][6] = (mid_1[3119:3112] > top_2[3111:3104]) ? 1 : 0;
assign detect_max[388][7] = (mid_1[3119:3112] > top_2[3119:3112]) ? 1 : 0;
assign detect_max[388][8] = (mid_1[3119:3112] > top_2[3127:3120]) ? 1 : 0;
assign detect_max[388][9] = (mid_1[3119:3112] > mid_0[3111:3104]) ? 1 : 0;
assign detect_max[388][10] = (mid_1[3119:3112] > mid_0[3119:3112]) ? 1 : 0;
assign detect_max[388][11] = (mid_1[3119:3112] > mid_0[3127:3120]) ? 1 : 0;
assign detect_max[388][12] = (mid_1[3119:3112] > mid_1[3111:3104]) ? 1 : 0;
assign detect_max[388][13] = (mid_1[3119:3112] > mid_1[3127:3120]) ? 1 : 0;
assign detect_max[388][14] = (mid_1[3119:3112] > mid_2[3111:3104]) ? 1 : 0;
assign detect_max[388][15] = (mid_1[3119:3112] > mid_2[3119:3112]) ? 1 : 0;
assign detect_max[388][16] = (mid_1[3119:3112] > mid_2[3127:3120]) ? 1 : 0;
assign detect_max[388][17] = (mid_1[3119:3112] > btm_0[3111:3104]) ? 1 : 0;
assign detect_max[388][18] = (mid_1[3119:3112] > btm_0[3119:3112]) ? 1 : 0;
assign detect_max[388][19] = (mid_1[3119:3112] > btm_0[3127:3120]) ? 1 : 0;
assign detect_max[388][20] = (mid_1[3119:3112] > btm_1[3111:3104]) ? 1 : 0;
assign detect_max[388][21] = (mid_1[3119:3112] > btm_1[3119:3112]) ? 1 : 0;
assign detect_max[388][22] = (mid_1[3119:3112] > btm_1[3127:3120]) ? 1 : 0;
assign detect_max[388][23] = (mid_1[3119:3112] > btm_2[3111:3104]) ? 1 : 0;
assign detect_max[388][24] = (mid_1[3119:3112] > btm_2[3119:3112]) ? 1 : 0;
assign detect_max[388][25] = (mid_1[3119:3112] > btm_2[3127:3120]) ? 1 : 0;

assign detect_max[389][0] = (mid_1[3127:3120] > top_0[3119:3112]) ? 1 : 0;
assign detect_max[389][1] = (mid_1[3127:3120] > top_0[3127:3120]) ? 1 : 0;
assign detect_max[389][2] = (mid_1[3127:3120] > top_0[3135:3128]) ? 1 : 0;
assign detect_max[389][3] = (mid_1[3127:3120] > top_1[3119:3112]) ? 1 : 0;
assign detect_max[389][4] = (mid_1[3127:3120] > top_1[3127:3120]) ? 1 : 0;
assign detect_max[389][5] = (mid_1[3127:3120] > top_1[3135:3128]) ? 1 : 0;
assign detect_max[389][6] = (mid_1[3127:3120] > top_2[3119:3112]) ? 1 : 0;
assign detect_max[389][7] = (mid_1[3127:3120] > top_2[3127:3120]) ? 1 : 0;
assign detect_max[389][8] = (mid_1[3127:3120] > top_2[3135:3128]) ? 1 : 0;
assign detect_max[389][9] = (mid_1[3127:3120] > mid_0[3119:3112]) ? 1 : 0;
assign detect_max[389][10] = (mid_1[3127:3120] > mid_0[3127:3120]) ? 1 : 0;
assign detect_max[389][11] = (mid_1[3127:3120] > mid_0[3135:3128]) ? 1 : 0;
assign detect_max[389][12] = (mid_1[3127:3120] > mid_1[3119:3112]) ? 1 : 0;
assign detect_max[389][13] = (mid_1[3127:3120] > mid_1[3135:3128]) ? 1 : 0;
assign detect_max[389][14] = (mid_1[3127:3120] > mid_2[3119:3112]) ? 1 : 0;
assign detect_max[389][15] = (mid_1[3127:3120] > mid_2[3127:3120]) ? 1 : 0;
assign detect_max[389][16] = (mid_1[3127:3120] > mid_2[3135:3128]) ? 1 : 0;
assign detect_max[389][17] = (mid_1[3127:3120] > btm_0[3119:3112]) ? 1 : 0;
assign detect_max[389][18] = (mid_1[3127:3120] > btm_0[3127:3120]) ? 1 : 0;
assign detect_max[389][19] = (mid_1[3127:3120] > btm_0[3135:3128]) ? 1 : 0;
assign detect_max[389][20] = (mid_1[3127:3120] > btm_1[3119:3112]) ? 1 : 0;
assign detect_max[389][21] = (mid_1[3127:3120] > btm_1[3127:3120]) ? 1 : 0;
assign detect_max[389][22] = (mid_1[3127:3120] > btm_1[3135:3128]) ? 1 : 0;
assign detect_max[389][23] = (mid_1[3127:3120] > btm_2[3119:3112]) ? 1 : 0;
assign detect_max[389][24] = (mid_1[3127:3120] > btm_2[3127:3120]) ? 1 : 0;
assign detect_max[389][25] = (mid_1[3127:3120] > btm_2[3135:3128]) ? 1 : 0;

assign detect_max[390][0] = (mid_1[3135:3128] > top_0[3127:3120]) ? 1 : 0;
assign detect_max[390][1] = (mid_1[3135:3128] > top_0[3135:3128]) ? 1 : 0;
assign detect_max[390][2] = (mid_1[3135:3128] > top_0[3143:3136]) ? 1 : 0;
assign detect_max[390][3] = (mid_1[3135:3128] > top_1[3127:3120]) ? 1 : 0;
assign detect_max[390][4] = (mid_1[3135:3128] > top_1[3135:3128]) ? 1 : 0;
assign detect_max[390][5] = (mid_1[3135:3128] > top_1[3143:3136]) ? 1 : 0;
assign detect_max[390][6] = (mid_1[3135:3128] > top_2[3127:3120]) ? 1 : 0;
assign detect_max[390][7] = (mid_1[3135:3128] > top_2[3135:3128]) ? 1 : 0;
assign detect_max[390][8] = (mid_1[3135:3128] > top_2[3143:3136]) ? 1 : 0;
assign detect_max[390][9] = (mid_1[3135:3128] > mid_0[3127:3120]) ? 1 : 0;
assign detect_max[390][10] = (mid_1[3135:3128] > mid_0[3135:3128]) ? 1 : 0;
assign detect_max[390][11] = (mid_1[3135:3128] > mid_0[3143:3136]) ? 1 : 0;
assign detect_max[390][12] = (mid_1[3135:3128] > mid_1[3127:3120]) ? 1 : 0;
assign detect_max[390][13] = (mid_1[3135:3128] > mid_1[3143:3136]) ? 1 : 0;
assign detect_max[390][14] = (mid_1[3135:3128] > mid_2[3127:3120]) ? 1 : 0;
assign detect_max[390][15] = (mid_1[3135:3128] > mid_2[3135:3128]) ? 1 : 0;
assign detect_max[390][16] = (mid_1[3135:3128] > mid_2[3143:3136]) ? 1 : 0;
assign detect_max[390][17] = (mid_1[3135:3128] > btm_0[3127:3120]) ? 1 : 0;
assign detect_max[390][18] = (mid_1[3135:3128] > btm_0[3135:3128]) ? 1 : 0;
assign detect_max[390][19] = (mid_1[3135:3128] > btm_0[3143:3136]) ? 1 : 0;
assign detect_max[390][20] = (mid_1[3135:3128] > btm_1[3127:3120]) ? 1 : 0;
assign detect_max[390][21] = (mid_1[3135:3128] > btm_1[3135:3128]) ? 1 : 0;
assign detect_max[390][22] = (mid_1[3135:3128] > btm_1[3143:3136]) ? 1 : 0;
assign detect_max[390][23] = (mid_1[3135:3128] > btm_2[3127:3120]) ? 1 : 0;
assign detect_max[390][24] = (mid_1[3135:3128] > btm_2[3135:3128]) ? 1 : 0;
assign detect_max[390][25] = (mid_1[3135:3128] > btm_2[3143:3136]) ? 1 : 0;

assign detect_max[391][0] = (mid_1[3143:3136] > top_0[3135:3128]) ? 1 : 0;
assign detect_max[391][1] = (mid_1[3143:3136] > top_0[3143:3136]) ? 1 : 0;
assign detect_max[391][2] = (mid_1[3143:3136] > top_0[3151:3144]) ? 1 : 0;
assign detect_max[391][3] = (mid_1[3143:3136] > top_1[3135:3128]) ? 1 : 0;
assign detect_max[391][4] = (mid_1[3143:3136] > top_1[3143:3136]) ? 1 : 0;
assign detect_max[391][5] = (mid_1[3143:3136] > top_1[3151:3144]) ? 1 : 0;
assign detect_max[391][6] = (mid_1[3143:3136] > top_2[3135:3128]) ? 1 : 0;
assign detect_max[391][7] = (mid_1[3143:3136] > top_2[3143:3136]) ? 1 : 0;
assign detect_max[391][8] = (mid_1[3143:3136] > top_2[3151:3144]) ? 1 : 0;
assign detect_max[391][9] = (mid_1[3143:3136] > mid_0[3135:3128]) ? 1 : 0;
assign detect_max[391][10] = (mid_1[3143:3136] > mid_0[3143:3136]) ? 1 : 0;
assign detect_max[391][11] = (mid_1[3143:3136] > mid_0[3151:3144]) ? 1 : 0;
assign detect_max[391][12] = (mid_1[3143:3136] > mid_1[3135:3128]) ? 1 : 0;
assign detect_max[391][13] = (mid_1[3143:3136] > mid_1[3151:3144]) ? 1 : 0;
assign detect_max[391][14] = (mid_1[3143:3136] > mid_2[3135:3128]) ? 1 : 0;
assign detect_max[391][15] = (mid_1[3143:3136] > mid_2[3143:3136]) ? 1 : 0;
assign detect_max[391][16] = (mid_1[3143:3136] > mid_2[3151:3144]) ? 1 : 0;
assign detect_max[391][17] = (mid_1[3143:3136] > btm_0[3135:3128]) ? 1 : 0;
assign detect_max[391][18] = (mid_1[3143:3136] > btm_0[3143:3136]) ? 1 : 0;
assign detect_max[391][19] = (mid_1[3143:3136] > btm_0[3151:3144]) ? 1 : 0;
assign detect_max[391][20] = (mid_1[3143:3136] > btm_1[3135:3128]) ? 1 : 0;
assign detect_max[391][21] = (mid_1[3143:3136] > btm_1[3143:3136]) ? 1 : 0;
assign detect_max[391][22] = (mid_1[3143:3136] > btm_1[3151:3144]) ? 1 : 0;
assign detect_max[391][23] = (mid_1[3143:3136] > btm_2[3135:3128]) ? 1 : 0;
assign detect_max[391][24] = (mid_1[3143:3136] > btm_2[3143:3136]) ? 1 : 0;
assign detect_max[391][25] = (mid_1[3143:3136] > btm_2[3151:3144]) ? 1 : 0;

assign detect_max[392][0] = (mid_1[3151:3144] > top_0[3143:3136]) ? 1 : 0;
assign detect_max[392][1] = (mid_1[3151:3144] > top_0[3151:3144]) ? 1 : 0;
assign detect_max[392][2] = (mid_1[3151:3144] > top_0[3159:3152]) ? 1 : 0;
assign detect_max[392][3] = (mid_1[3151:3144] > top_1[3143:3136]) ? 1 : 0;
assign detect_max[392][4] = (mid_1[3151:3144] > top_1[3151:3144]) ? 1 : 0;
assign detect_max[392][5] = (mid_1[3151:3144] > top_1[3159:3152]) ? 1 : 0;
assign detect_max[392][6] = (mid_1[3151:3144] > top_2[3143:3136]) ? 1 : 0;
assign detect_max[392][7] = (mid_1[3151:3144] > top_2[3151:3144]) ? 1 : 0;
assign detect_max[392][8] = (mid_1[3151:3144] > top_2[3159:3152]) ? 1 : 0;
assign detect_max[392][9] = (mid_1[3151:3144] > mid_0[3143:3136]) ? 1 : 0;
assign detect_max[392][10] = (mid_1[3151:3144] > mid_0[3151:3144]) ? 1 : 0;
assign detect_max[392][11] = (mid_1[3151:3144] > mid_0[3159:3152]) ? 1 : 0;
assign detect_max[392][12] = (mid_1[3151:3144] > mid_1[3143:3136]) ? 1 : 0;
assign detect_max[392][13] = (mid_1[3151:3144] > mid_1[3159:3152]) ? 1 : 0;
assign detect_max[392][14] = (mid_1[3151:3144] > mid_2[3143:3136]) ? 1 : 0;
assign detect_max[392][15] = (mid_1[3151:3144] > mid_2[3151:3144]) ? 1 : 0;
assign detect_max[392][16] = (mid_1[3151:3144] > mid_2[3159:3152]) ? 1 : 0;
assign detect_max[392][17] = (mid_1[3151:3144] > btm_0[3143:3136]) ? 1 : 0;
assign detect_max[392][18] = (mid_1[3151:3144] > btm_0[3151:3144]) ? 1 : 0;
assign detect_max[392][19] = (mid_1[3151:3144] > btm_0[3159:3152]) ? 1 : 0;
assign detect_max[392][20] = (mid_1[3151:3144] > btm_1[3143:3136]) ? 1 : 0;
assign detect_max[392][21] = (mid_1[3151:3144] > btm_1[3151:3144]) ? 1 : 0;
assign detect_max[392][22] = (mid_1[3151:3144] > btm_1[3159:3152]) ? 1 : 0;
assign detect_max[392][23] = (mid_1[3151:3144] > btm_2[3143:3136]) ? 1 : 0;
assign detect_max[392][24] = (mid_1[3151:3144] > btm_2[3151:3144]) ? 1 : 0;
assign detect_max[392][25] = (mid_1[3151:3144] > btm_2[3159:3152]) ? 1 : 0;

assign detect_max[393][0] = (mid_1[3159:3152] > top_0[3151:3144]) ? 1 : 0;
assign detect_max[393][1] = (mid_1[3159:3152] > top_0[3159:3152]) ? 1 : 0;
assign detect_max[393][2] = (mid_1[3159:3152] > top_0[3167:3160]) ? 1 : 0;
assign detect_max[393][3] = (mid_1[3159:3152] > top_1[3151:3144]) ? 1 : 0;
assign detect_max[393][4] = (mid_1[3159:3152] > top_1[3159:3152]) ? 1 : 0;
assign detect_max[393][5] = (mid_1[3159:3152] > top_1[3167:3160]) ? 1 : 0;
assign detect_max[393][6] = (mid_1[3159:3152] > top_2[3151:3144]) ? 1 : 0;
assign detect_max[393][7] = (mid_1[3159:3152] > top_2[3159:3152]) ? 1 : 0;
assign detect_max[393][8] = (mid_1[3159:3152] > top_2[3167:3160]) ? 1 : 0;
assign detect_max[393][9] = (mid_1[3159:3152] > mid_0[3151:3144]) ? 1 : 0;
assign detect_max[393][10] = (mid_1[3159:3152] > mid_0[3159:3152]) ? 1 : 0;
assign detect_max[393][11] = (mid_1[3159:3152] > mid_0[3167:3160]) ? 1 : 0;
assign detect_max[393][12] = (mid_1[3159:3152] > mid_1[3151:3144]) ? 1 : 0;
assign detect_max[393][13] = (mid_1[3159:3152] > mid_1[3167:3160]) ? 1 : 0;
assign detect_max[393][14] = (mid_1[3159:3152] > mid_2[3151:3144]) ? 1 : 0;
assign detect_max[393][15] = (mid_1[3159:3152] > mid_2[3159:3152]) ? 1 : 0;
assign detect_max[393][16] = (mid_1[3159:3152] > mid_2[3167:3160]) ? 1 : 0;
assign detect_max[393][17] = (mid_1[3159:3152] > btm_0[3151:3144]) ? 1 : 0;
assign detect_max[393][18] = (mid_1[3159:3152] > btm_0[3159:3152]) ? 1 : 0;
assign detect_max[393][19] = (mid_1[3159:3152] > btm_0[3167:3160]) ? 1 : 0;
assign detect_max[393][20] = (mid_1[3159:3152] > btm_1[3151:3144]) ? 1 : 0;
assign detect_max[393][21] = (mid_1[3159:3152] > btm_1[3159:3152]) ? 1 : 0;
assign detect_max[393][22] = (mid_1[3159:3152] > btm_1[3167:3160]) ? 1 : 0;
assign detect_max[393][23] = (mid_1[3159:3152] > btm_2[3151:3144]) ? 1 : 0;
assign detect_max[393][24] = (mid_1[3159:3152] > btm_2[3159:3152]) ? 1 : 0;
assign detect_max[393][25] = (mid_1[3159:3152] > btm_2[3167:3160]) ? 1 : 0;

assign detect_max[394][0] = (mid_1[3167:3160] > top_0[3159:3152]) ? 1 : 0;
assign detect_max[394][1] = (mid_1[3167:3160] > top_0[3167:3160]) ? 1 : 0;
assign detect_max[394][2] = (mid_1[3167:3160] > top_0[3175:3168]) ? 1 : 0;
assign detect_max[394][3] = (mid_1[3167:3160] > top_1[3159:3152]) ? 1 : 0;
assign detect_max[394][4] = (mid_1[3167:3160] > top_1[3167:3160]) ? 1 : 0;
assign detect_max[394][5] = (mid_1[3167:3160] > top_1[3175:3168]) ? 1 : 0;
assign detect_max[394][6] = (mid_1[3167:3160] > top_2[3159:3152]) ? 1 : 0;
assign detect_max[394][7] = (mid_1[3167:3160] > top_2[3167:3160]) ? 1 : 0;
assign detect_max[394][8] = (mid_1[3167:3160] > top_2[3175:3168]) ? 1 : 0;
assign detect_max[394][9] = (mid_1[3167:3160] > mid_0[3159:3152]) ? 1 : 0;
assign detect_max[394][10] = (mid_1[3167:3160] > mid_0[3167:3160]) ? 1 : 0;
assign detect_max[394][11] = (mid_1[3167:3160] > mid_0[3175:3168]) ? 1 : 0;
assign detect_max[394][12] = (mid_1[3167:3160] > mid_1[3159:3152]) ? 1 : 0;
assign detect_max[394][13] = (mid_1[3167:3160] > mid_1[3175:3168]) ? 1 : 0;
assign detect_max[394][14] = (mid_1[3167:3160] > mid_2[3159:3152]) ? 1 : 0;
assign detect_max[394][15] = (mid_1[3167:3160] > mid_2[3167:3160]) ? 1 : 0;
assign detect_max[394][16] = (mid_1[3167:3160] > mid_2[3175:3168]) ? 1 : 0;
assign detect_max[394][17] = (mid_1[3167:3160] > btm_0[3159:3152]) ? 1 : 0;
assign detect_max[394][18] = (mid_1[3167:3160] > btm_0[3167:3160]) ? 1 : 0;
assign detect_max[394][19] = (mid_1[3167:3160] > btm_0[3175:3168]) ? 1 : 0;
assign detect_max[394][20] = (mid_1[3167:3160] > btm_1[3159:3152]) ? 1 : 0;
assign detect_max[394][21] = (mid_1[3167:3160] > btm_1[3167:3160]) ? 1 : 0;
assign detect_max[394][22] = (mid_1[3167:3160] > btm_1[3175:3168]) ? 1 : 0;
assign detect_max[394][23] = (mid_1[3167:3160] > btm_2[3159:3152]) ? 1 : 0;
assign detect_max[394][24] = (mid_1[3167:3160] > btm_2[3167:3160]) ? 1 : 0;
assign detect_max[394][25] = (mid_1[3167:3160] > btm_2[3175:3168]) ? 1 : 0;

assign detect_max[395][0] = (mid_1[3175:3168] > top_0[3167:3160]) ? 1 : 0;
assign detect_max[395][1] = (mid_1[3175:3168] > top_0[3175:3168]) ? 1 : 0;
assign detect_max[395][2] = (mid_1[3175:3168] > top_0[3183:3176]) ? 1 : 0;
assign detect_max[395][3] = (mid_1[3175:3168] > top_1[3167:3160]) ? 1 : 0;
assign detect_max[395][4] = (mid_1[3175:3168] > top_1[3175:3168]) ? 1 : 0;
assign detect_max[395][5] = (mid_1[3175:3168] > top_1[3183:3176]) ? 1 : 0;
assign detect_max[395][6] = (mid_1[3175:3168] > top_2[3167:3160]) ? 1 : 0;
assign detect_max[395][7] = (mid_1[3175:3168] > top_2[3175:3168]) ? 1 : 0;
assign detect_max[395][8] = (mid_1[3175:3168] > top_2[3183:3176]) ? 1 : 0;
assign detect_max[395][9] = (mid_1[3175:3168] > mid_0[3167:3160]) ? 1 : 0;
assign detect_max[395][10] = (mid_1[3175:3168] > mid_0[3175:3168]) ? 1 : 0;
assign detect_max[395][11] = (mid_1[3175:3168] > mid_0[3183:3176]) ? 1 : 0;
assign detect_max[395][12] = (mid_1[3175:3168] > mid_1[3167:3160]) ? 1 : 0;
assign detect_max[395][13] = (mid_1[3175:3168] > mid_1[3183:3176]) ? 1 : 0;
assign detect_max[395][14] = (mid_1[3175:3168] > mid_2[3167:3160]) ? 1 : 0;
assign detect_max[395][15] = (mid_1[3175:3168] > mid_2[3175:3168]) ? 1 : 0;
assign detect_max[395][16] = (mid_1[3175:3168] > mid_2[3183:3176]) ? 1 : 0;
assign detect_max[395][17] = (mid_1[3175:3168] > btm_0[3167:3160]) ? 1 : 0;
assign detect_max[395][18] = (mid_1[3175:3168] > btm_0[3175:3168]) ? 1 : 0;
assign detect_max[395][19] = (mid_1[3175:3168] > btm_0[3183:3176]) ? 1 : 0;
assign detect_max[395][20] = (mid_1[3175:3168] > btm_1[3167:3160]) ? 1 : 0;
assign detect_max[395][21] = (mid_1[3175:3168] > btm_1[3175:3168]) ? 1 : 0;
assign detect_max[395][22] = (mid_1[3175:3168] > btm_1[3183:3176]) ? 1 : 0;
assign detect_max[395][23] = (mid_1[3175:3168] > btm_2[3167:3160]) ? 1 : 0;
assign detect_max[395][24] = (mid_1[3175:3168] > btm_2[3175:3168]) ? 1 : 0;
assign detect_max[395][25] = (mid_1[3175:3168] > btm_2[3183:3176]) ? 1 : 0;

assign detect_max[396][0] = (mid_1[3183:3176] > top_0[3175:3168]) ? 1 : 0;
assign detect_max[396][1] = (mid_1[3183:3176] > top_0[3183:3176]) ? 1 : 0;
assign detect_max[396][2] = (mid_1[3183:3176] > top_0[3191:3184]) ? 1 : 0;
assign detect_max[396][3] = (mid_1[3183:3176] > top_1[3175:3168]) ? 1 : 0;
assign detect_max[396][4] = (mid_1[3183:3176] > top_1[3183:3176]) ? 1 : 0;
assign detect_max[396][5] = (mid_1[3183:3176] > top_1[3191:3184]) ? 1 : 0;
assign detect_max[396][6] = (mid_1[3183:3176] > top_2[3175:3168]) ? 1 : 0;
assign detect_max[396][7] = (mid_1[3183:3176] > top_2[3183:3176]) ? 1 : 0;
assign detect_max[396][8] = (mid_1[3183:3176] > top_2[3191:3184]) ? 1 : 0;
assign detect_max[396][9] = (mid_1[3183:3176] > mid_0[3175:3168]) ? 1 : 0;
assign detect_max[396][10] = (mid_1[3183:3176] > mid_0[3183:3176]) ? 1 : 0;
assign detect_max[396][11] = (mid_1[3183:3176] > mid_0[3191:3184]) ? 1 : 0;
assign detect_max[396][12] = (mid_1[3183:3176] > mid_1[3175:3168]) ? 1 : 0;
assign detect_max[396][13] = (mid_1[3183:3176] > mid_1[3191:3184]) ? 1 : 0;
assign detect_max[396][14] = (mid_1[3183:3176] > mid_2[3175:3168]) ? 1 : 0;
assign detect_max[396][15] = (mid_1[3183:3176] > mid_2[3183:3176]) ? 1 : 0;
assign detect_max[396][16] = (mid_1[3183:3176] > mid_2[3191:3184]) ? 1 : 0;
assign detect_max[396][17] = (mid_1[3183:3176] > btm_0[3175:3168]) ? 1 : 0;
assign detect_max[396][18] = (mid_1[3183:3176] > btm_0[3183:3176]) ? 1 : 0;
assign detect_max[396][19] = (mid_1[3183:3176] > btm_0[3191:3184]) ? 1 : 0;
assign detect_max[396][20] = (mid_1[3183:3176] > btm_1[3175:3168]) ? 1 : 0;
assign detect_max[396][21] = (mid_1[3183:3176] > btm_1[3183:3176]) ? 1 : 0;
assign detect_max[396][22] = (mid_1[3183:3176] > btm_1[3191:3184]) ? 1 : 0;
assign detect_max[396][23] = (mid_1[3183:3176] > btm_2[3175:3168]) ? 1 : 0;
assign detect_max[396][24] = (mid_1[3183:3176] > btm_2[3183:3176]) ? 1 : 0;
assign detect_max[396][25] = (mid_1[3183:3176] > btm_2[3191:3184]) ? 1 : 0;

assign detect_max[397][0] = (mid_1[3191:3184] > top_0[3183:3176]) ? 1 : 0;
assign detect_max[397][1] = (mid_1[3191:3184] > top_0[3191:3184]) ? 1 : 0;
assign detect_max[397][2] = (mid_1[3191:3184] > top_0[3199:3192]) ? 1 : 0;
assign detect_max[397][3] = (mid_1[3191:3184] > top_1[3183:3176]) ? 1 : 0;
assign detect_max[397][4] = (mid_1[3191:3184] > top_1[3191:3184]) ? 1 : 0;
assign detect_max[397][5] = (mid_1[3191:3184] > top_1[3199:3192]) ? 1 : 0;
assign detect_max[397][6] = (mid_1[3191:3184] > top_2[3183:3176]) ? 1 : 0;
assign detect_max[397][7] = (mid_1[3191:3184] > top_2[3191:3184]) ? 1 : 0;
assign detect_max[397][8] = (mid_1[3191:3184] > top_2[3199:3192]) ? 1 : 0;
assign detect_max[397][9] = (mid_1[3191:3184] > mid_0[3183:3176]) ? 1 : 0;
assign detect_max[397][10] = (mid_1[3191:3184] > mid_0[3191:3184]) ? 1 : 0;
assign detect_max[397][11] = (mid_1[3191:3184] > mid_0[3199:3192]) ? 1 : 0;
assign detect_max[397][12] = (mid_1[3191:3184] > mid_1[3183:3176]) ? 1 : 0;
assign detect_max[397][13] = (mid_1[3191:3184] > mid_1[3199:3192]) ? 1 : 0;
assign detect_max[397][14] = (mid_1[3191:3184] > mid_2[3183:3176]) ? 1 : 0;
assign detect_max[397][15] = (mid_1[3191:3184] > mid_2[3191:3184]) ? 1 : 0;
assign detect_max[397][16] = (mid_1[3191:3184] > mid_2[3199:3192]) ? 1 : 0;
assign detect_max[397][17] = (mid_1[3191:3184] > btm_0[3183:3176]) ? 1 : 0;
assign detect_max[397][18] = (mid_1[3191:3184] > btm_0[3191:3184]) ? 1 : 0;
assign detect_max[397][19] = (mid_1[3191:3184] > btm_0[3199:3192]) ? 1 : 0;
assign detect_max[397][20] = (mid_1[3191:3184] > btm_1[3183:3176]) ? 1 : 0;
assign detect_max[397][21] = (mid_1[3191:3184] > btm_1[3191:3184]) ? 1 : 0;
assign detect_max[397][22] = (mid_1[3191:3184] > btm_1[3199:3192]) ? 1 : 0;
assign detect_max[397][23] = (mid_1[3191:3184] > btm_2[3183:3176]) ? 1 : 0;
assign detect_max[397][24] = (mid_1[3191:3184] > btm_2[3191:3184]) ? 1 : 0;
assign detect_max[397][25] = (mid_1[3191:3184] > btm_2[3199:3192]) ? 1 : 0;

assign detect_max[398][0] = (mid_1[3199:3192] > top_0[3191:3184]) ? 1 : 0;
assign detect_max[398][1] = (mid_1[3199:3192] > top_0[3199:3192]) ? 1 : 0;
assign detect_max[398][2] = (mid_1[3199:3192] > top_0[3207:3200]) ? 1 : 0;
assign detect_max[398][3] = (mid_1[3199:3192] > top_1[3191:3184]) ? 1 : 0;
assign detect_max[398][4] = (mid_1[3199:3192] > top_1[3199:3192]) ? 1 : 0;
assign detect_max[398][5] = (mid_1[3199:3192] > top_1[3207:3200]) ? 1 : 0;
assign detect_max[398][6] = (mid_1[3199:3192] > top_2[3191:3184]) ? 1 : 0;
assign detect_max[398][7] = (mid_1[3199:3192] > top_2[3199:3192]) ? 1 : 0;
assign detect_max[398][8] = (mid_1[3199:3192] > top_2[3207:3200]) ? 1 : 0;
assign detect_max[398][9] = (mid_1[3199:3192] > mid_0[3191:3184]) ? 1 : 0;
assign detect_max[398][10] = (mid_1[3199:3192] > mid_0[3199:3192]) ? 1 : 0;
assign detect_max[398][11] = (mid_1[3199:3192] > mid_0[3207:3200]) ? 1 : 0;
assign detect_max[398][12] = (mid_1[3199:3192] > mid_1[3191:3184]) ? 1 : 0;
assign detect_max[398][13] = (mid_1[3199:3192] > mid_1[3207:3200]) ? 1 : 0;
assign detect_max[398][14] = (mid_1[3199:3192] > mid_2[3191:3184]) ? 1 : 0;
assign detect_max[398][15] = (mid_1[3199:3192] > mid_2[3199:3192]) ? 1 : 0;
assign detect_max[398][16] = (mid_1[3199:3192] > mid_2[3207:3200]) ? 1 : 0;
assign detect_max[398][17] = (mid_1[3199:3192] > btm_0[3191:3184]) ? 1 : 0;
assign detect_max[398][18] = (mid_1[3199:3192] > btm_0[3199:3192]) ? 1 : 0;
assign detect_max[398][19] = (mid_1[3199:3192] > btm_0[3207:3200]) ? 1 : 0;
assign detect_max[398][20] = (mid_1[3199:3192] > btm_1[3191:3184]) ? 1 : 0;
assign detect_max[398][21] = (mid_1[3199:3192] > btm_1[3199:3192]) ? 1 : 0;
assign detect_max[398][22] = (mid_1[3199:3192] > btm_1[3207:3200]) ? 1 : 0;
assign detect_max[398][23] = (mid_1[3199:3192] > btm_2[3191:3184]) ? 1 : 0;
assign detect_max[398][24] = (mid_1[3199:3192] > btm_2[3199:3192]) ? 1 : 0;
assign detect_max[398][25] = (mid_1[3199:3192] > btm_2[3207:3200]) ? 1 : 0;

assign detect_max[399][0] = (mid_1[3207:3200] > top_0[3199:3192]) ? 1 : 0;
assign detect_max[399][1] = (mid_1[3207:3200] > top_0[3207:3200]) ? 1 : 0;
assign detect_max[399][2] = (mid_1[3207:3200] > top_0[3215:3208]) ? 1 : 0;
assign detect_max[399][3] = (mid_1[3207:3200] > top_1[3199:3192]) ? 1 : 0;
assign detect_max[399][4] = (mid_1[3207:3200] > top_1[3207:3200]) ? 1 : 0;
assign detect_max[399][5] = (mid_1[3207:3200] > top_1[3215:3208]) ? 1 : 0;
assign detect_max[399][6] = (mid_1[3207:3200] > top_2[3199:3192]) ? 1 : 0;
assign detect_max[399][7] = (mid_1[3207:3200] > top_2[3207:3200]) ? 1 : 0;
assign detect_max[399][8] = (mid_1[3207:3200] > top_2[3215:3208]) ? 1 : 0;
assign detect_max[399][9] = (mid_1[3207:3200] > mid_0[3199:3192]) ? 1 : 0;
assign detect_max[399][10] = (mid_1[3207:3200] > mid_0[3207:3200]) ? 1 : 0;
assign detect_max[399][11] = (mid_1[3207:3200] > mid_0[3215:3208]) ? 1 : 0;
assign detect_max[399][12] = (mid_1[3207:3200] > mid_1[3199:3192]) ? 1 : 0;
assign detect_max[399][13] = (mid_1[3207:3200] > mid_1[3215:3208]) ? 1 : 0;
assign detect_max[399][14] = (mid_1[3207:3200] > mid_2[3199:3192]) ? 1 : 0;
assign detect_max[399][15] = (mid_1[3207:3200] > mid_2[3207:3200]) ? 1 : 0;
assign detect_max[399][16] = (mid_1[3207:3200] > mid_2[3215:3208]) ? 1 : 0;
assign detect_max[399][17] = (mid_1[3207:3200] > btm_0[3199:3192]) ? 1 : 0;
assign detect_max[399][18] = (mid_1[3207:3200] > btm_0[3207:3200]) ? 1 : 0;
assign detect_max[399][19] = (mid_1[3207:3200] > btm_0[3215:3208]) ? 1 : 0;
assign detect_max[399][20] = (mid_1[3207:3200] > btm_1[3199:3192]) ? 1 : 0;
assign detect_max[399][21] = (mid_1[3207:3200] > btm_1[3207:3200]) ? 1 : 0;
assign detect_max[399][22] = (mid_1[3207:3200] > btm_1[3215:3208]) ? 1 : 0;
assign detect_max[399][23] = (mid_1[3207:3200] > btm_2[3199:3192]) ? 1 : 0;
assign detect_max[399][24] = (mid_1[3207:3200] > btm_2[3207:3200]) ? 1 : 0;
assign detect_max[399][25] = (mid_1[3207:3200] > btm_2[3215:3208]) ? 1 : 0;

assign detect_max[400][0] = (mid_1[3215:3208] > top_0[3207:3200]) ? 1 : 0;
assign detect_max[400][1] = (mid_1[3215:3208] > top_0[3215:3208]) ? 1 : 0;
assign detect_max[400][2] = (mid_1[3215:3208] > top_0[3223:3216]) ? 1 : 0;
assign detect_max[400][3] = (mid_1[3215:3208] > top_1[3207:3200]) ? 1 : 0;
assign detect_max[400][4] = (mid_1[3215:3208] > top_1[3215:3208]) ? 1 : 0;
assign detect_max[400][5] = (mid_1[3215:3208] > top_1[3223:3216]) ? 1 : 0;
assign detect_max[400][6] = (mid_1[3215:3208] > top_2[3207:3200]) ? 1 : 0;
assign detect_max[400][7] = (mid_1[3215:3208] > top_2[3215:3208]) ? 1 : 0;
assign detect_max[400][8] = (mid_1[3215:3208] > top_2[3223:3216]) ? 1 : 0;
assign detect_max[400][9] = (mid_1[3215:3208] > mid_0[3207:3200]) ? 1 : 0;
assign detect_max[400][10] = (mid_1[3215:3208] > mid_0[3215:3208]) ? 1 : 0;
assign detect_max[400][11] = (mid_1[3215:3208] > mid_0[3223:3216]) ? 1 : 0;
assign detect_max[400][12] = (mid_1[3215:3208] > mid_1[3207:3200]) ? 1 : 0;
assign detect_max[400][13] = (mid_1[3215:3208] > mid_1[3223:3216]) ? 1 : 0;
assign detect_max[400][14] = (mid_1[3215:3208] > mid_2[3207:3200]) ? 1 : 0;
assign detect_max[400][15] = (mid_1[3215:3208] > mid_2[3215:3208]) ? 1 : 0;
assign detect_max[400][16] = (mid_1[3215:3208] > mid_2[3223:3216]) ? 1 : 0;
assign detect_max[400][17] = (mid_1[3215:3208] > btm_0[3207:3200]) ? 1 : 0;
assign detect_max[400][18] = (mid_1[3215:3208] > btm_0[3215:3208]) ? 1 : 0;
assign detect_max[400][19] = (mid_1[3215:3208] > btm_0[3223:3216]) ? 1 : 0;
assign detect_max[400][20] = (mid_1[3215:3208] > btm_1[3207:3200]) ? 1 : 0;
assign detect_max[400][21] = (mid_1[3215:3208] > btm_1[3215:3208]) ? 1 : 0;
assign detect_max[400][22] = (mid_1[3215:3208] > btm_1[3223:3216]) ? 1 : 0;
assign detect_max[400][23] = (mid_1[3215:3208] > btm_2[3207:3200]) ? 1 : 0;
assign detect_max[400][24] = (mid_1[3215:3208] > btm_2[3215:3208]) ? 1 : 0;
assign detect_max[400][25] = (mid_1[3215:3208] > btm_2[3223:3216]) ? 1 : 0;

assign detect_max[401][0] = (mid_1[3223:3216] > top_0[3215:3208]) ? 1 : 0;
assign detect_max[401][1] = (mid_1[3223:3216] > top_0[3223:3216]) ? 1 : 0;
assign detect_max[401][2] = (mid_1[3223:3216] > top_0[3231:3224]) ? 1 : 0;
assign detect_max[401][3] = (mid_1[3223:3216] > top_1[3215:3208]) ? 1 : 0;
assign detect_max[401][4] = (mid_1[3223:3216] > top_1[3223:3216]) ? 1 : 0;
assign detect_max[401][5] = (mid_1[3223:3216] > top_1[3231:3224]) ? 1 : 0;
assign detect_max[401][6] = (mid_1[3223:3216] > top_2[3215:3208]) ? 1 : 0;
assign detect_max[401][7] = (mid_1[3223:3216] > top_2[3223:3216]) ? 1 : 0;
assign detect_max[401][8] = (mid_1[3223:3216] > top_2[3231:3224]) ? 1 : 0;
assign detect_max[401][9] = (mid_1[3223:3216] > mid_0[3215:3208]) ? 1 : 0;
assign detect_max[401][10] = (mid_1[3223:3216] > mid_0[3223:3216]) ? 1 : 0;
assign detect_max[401][11] = (mid_1[3223:3216] > mid_0[3231:3224]) ? 1 : 0;
assign detect_max[401][12] = (mid_1[3223:3216] > mid_1[3215:3208]) ? 1 : 0;
assign detect_max[401][13] = (mid_1[3223:3216] > mid_1[3231:3224]) ? 1 : 0;
assign detect_max[401][14] = (mid_1[3223:3216] > mid_2[3215:3208]) ? 1 : 0;
assign detect_max[401][15] = (mid_1[3223:3216] > mid_2[3223:3216]) ? 1 : 0;
assign detect_max[401][16] = (mid_1[3223:3216] > mid_2[3231:3224]) ? 1 : 0;
assign detect_max[401][17] = (mid_1[3223:3216] > btm_0[3215:3208]) ? 1 : 0;
assign detect_max[401][18] = (mid_1[3223:3216] > btm_0[3223:3216]) ? 1 : 0;
assign detect_max[401][19] = (mid_1[3223:3216] > btm_0[3231:3224]) ? 1 : 0;
assign detect_max[401][20] = (mid_1[3223:3216] > btm_1[3215:3208]) ? 1 : 0;
assign detect_max[401][21] = (mid_1[3223:3216] > btm_1[3223:3216]) ? 1 : 0;
assign detect_max[401][22] = (mid_1[3223:3216] > btm_1[3231:3224]) ? 1 : 0;
assign detect_max[401][23] = (mid_1[3223:3216] > btm_2[3215:3208]) ? 1 : 0;
assign detect_max[401][24] = (mid_1[3223:3216] > btm_2[3223:3216]) ? 1 : 0;
assign detect_max[401][25] = (mid_1[3223:3216] > btm_2[3231:3224]) ? 1 : 0;

assign detect_max[402][0] = (mid_1[3231:3224] > top_0[3223:3216]) ? 1 : 0;
assign detect_max[402][1] = (mid_1[3231:3224] > top_0[3231:3224]) ? 1 : 0;
assign detect_max[402][2] = (mid_1[3231:3224] > top_0[3239:3232]) ? 1 : 0;
assign detect_max[402][3] = (mid_1[3231:3224] > top_1[3223:3216]) ? 1 : 0;
assign detect_max[402][4] = (mid_1[3231:3224] > top_1[3231:3224]) ? 1 : 0;
assign detect_max[402][5] = (mid_1[3231:3224] > top_1[3239:3232]) ? 1 : 0;
assign detect_max[402][6] = (mid_1[3231:3224] > top_2[3223:3216]) ? 1 : 0;
assign detect_max[402][7] = (mid_1[3231:3224] > top_2[3231:3224]) ? 1 : 0;
assign detect_max[402][8] = (mid_1[3231:3224] > top_2[3239:3232]) ? 1 : 0;
assign detect_max[402][9] = (mid_1[3231:3224] > mid_0[3223:3216]) ? 1 : 0;
assign detect_max[402][10] = (mid_1[3231:3224] > mid_0[3231:3224]) ? 1 : 0;
assign detect_max[402][11] = (mid_1[3231:3224] > mid_0[3239:3232]) ? 1 : 0;
assign detect_max[402][12] = (mid_1[3231:3224] > mid_1[3223:3216]) ? 1 : 0;
assign detect_max[402][13] = (mid_1[3231:3224] > mid_1[3239:3232]) ? 1 : 0;
assign detect_max[402][14] = (mid_1[3231:3224] > mid_2[3223:3216]) ? 1 : 0;
assign detect_max[402][15] = (mid_1[3231:3224] > mid_2[3231:3224]) ? 1 : 0;
assign detect_max[402][16] = (mid_1[3231:3224] > mid_2[3239:3232]) ? 1 : 0;
assign detect_max[402][17] = (mid_1[3231:3224] > btm_0[3223:3216]) ? 1 : 0;
assign detect_max[402][18] = (mid_1[3231:3224] > btm_0[3231:3224]) ? 1 : 0;
assign detect_max[402][19] = (mid_1[3231:3224] > btm_0[3239:3232]) ? 1 : 0;
assign detect_max[402][20] = (mid_1[3231:3224] > btm_1[3223:3216]) ? 1 : 0;
assign detect_max[402][21] = (mid_1[3231:3224] > btm_1[3231:3224]) ? 1 : 0;
assign detect_max[402][22] = (mid_1[3231:3224] > btm_1[3239:3232]) ? 1 : 0;
assign detect_max[402][23] = (mid_1[3231:3224] > btm_2[3223:3216]) ? 1 : 0;
assign detect_max[402][24] = (mid_1[3231:3224] > btm_2[3231:3224]) ? 1 : 0;
assign detect_max[402][25] = (mid_1[3231:3224] > btm_2[3239:3232]) ? 1 : 0;

assign detect_max[403][0] = (mid_1[3239:3232] > top_0[3231:3224]) ? 1 : 0;
assign detect_max[403][1] = (mid_1[3239:3232] > top_0[3239:3232]) ? 1 : 0;
assign detect_max[403][2] = (mid_1[3239:3232] > top_0[3247:3240]) ? 1 : 0;
assign detect_max[403][3] = (mid_1[3239:3232] > top_1[3231:3224]) ? 1 : 0;
assign detect_max[403][4] = (mid_1[3239:3232] > top_1[3239:3232]) ? 1 : 0;
assign detect_max[403][5] = (mid_1[3239:3232] > top_1[3247:3240]) ? 1 : 0;
assign detect_max[403][6] = (mid_1[3239:3232] > top_2[3231:3224]) ? 1 : 0;
assign detect_max[403][7] = (mid_1[3239:3232] > top_2[3239:3232]) ? 1 : 0;
assign detect_max[403][8] = (mid_1[3239:3232] > top_2[3247:3240]) ? 1 : 0;
assign detect_max[403][9] = (mid_1[3239:3232] > mid_0[3231:3224]) ? 1 : 0;
assign detect_max[403][10] = (mid_1[3239:3232] > mid_0[3239:3232]) ? 1 : 0;
assign detect_max[403][11] = (mid_1[3239:3232] > mid_0[3247:3240]) ? 1 : 0;
assign detect_max[403][12] = (mid_1[3239:3232] > mid_1[3231:3224]) ? 1 : 0;
assign detect_max[403][13] = (mid_1[3239:3232] > mid_1[3247:3240]) ? 1 : 0;
assign detect_max[403][14] = (mid_1[3239:3232] > mid_2[3231:3224]) ? 1 : 0;
assign detect_max[403][15] = (mid_1[3239:3232] > mid_2[3239:3232]) ? 1 : 0;
assign detect_max[403][16] = (mid_1[3239:3232] > mid_2[3247:3240]) ? 1 : 0;
assign detect_max[403][17] = (mid_1[3239:3232] > btm_0[3231:3224]) ? 1 : 0;
assign detect_max[403][18] = (mid_1[3239:3232] > btm_0[3239:3232]) ? 1 : 0;
assign detect_max[403][19] = (mid_1[3239:3232] > btm_0[3247:3240]) ? 1 : 0;
assign detect_max[403][20] = (mid_1[3239:3232] > btm_1[3231:3224]) ? 1 : 0;
assign detect_max[403][21] = (mid_1[3239:3232] > btm_1[3239:3232]) ? 1 : 0;
assign detect_max[403][22] = (mid_1[3239:3232] > btm_1[3247:3240]) ? 1 : 0;
assign detect_max[403][23] = (mid_1[3239:3232] > btm_2[3231:3224]) ? 1 : 0;
assign detect_max[403][24] = (mid_1[3239:3232] > btm_2[3239:3232]) ? 1 : 0;
assign detect_max[403][25] = (mid_1[3239:3232] > btm_2[3247:3240]) ? 1 : 0;

assign detect_max[404][0] = (mid_1[3247:3240] > top_0[3239:3232]) ? 1 : 0;
assign detect_max[404][1] = (mid_1[3247:3240] > top_0[3247:3240]) ? 1 : 0;
assign detect_max[404][2] = (mid_1[3247:3240] > top_0[3255:3248]) ? 1 : 0;
assign detect_max[404][3] = (mid_1[3247:3240] > top_1[3239:3232]) ? 1 : 0;
assign detect_max[404][4] = (mid_1[3247:3240] > top_1[3247:3240]) ? 1 : 0;
assign detect_max[404][5] = (mid_1[3247:3240] > top_1[3255:3248]) ? 1 : 0;
assign detect_max[404][6] = (mid_1[3247:3240] > top_2[3239:3232]) ? 1 : 0;
assign detect_max[404][7] = (mid_1[3247:3240] > top_2[3247:3240]) ? 1 : 0;
assign detect_max[404][8] = (mid_1[3247:3240] > top_2[3255:3248]) ? 1 : 0;
assign detect_max[404][9] = (mid_1[3247:3240] > mid_0[3239:3232]) ? 1 : 0;
assign detect_max[404][10] = (mid_1[3247:3240] > mid_0[3247:3240]) ? 1 : 0;
assign detect_max[404][11] = (mid_1[3247:3240] > mid_0[3255:3248]) ? 1 : 0;
assign detect_max[404][12] = (mid_1[3247:3240] > mid_1[3239:3232]) ? 1 : 0;
assign detect_max[404][13] = (mid_1[3247:3240] > mid_1[3255:3248]) ? 1 : 0;
assign detect_max[404][14] = (mid_1[3247:3240] > mid_2[3239:3232]) ? 1 : 0;
assign detect_max[404][15] = (mid_1[3247:3240] > mid_2[3247:3240]) ? 1 : 0;
assign detect_max[404][16] = (mid_1[3247:3240] > mid_2[3255:3248]) ? 1 : 0;
assign detect_max[404][17] = (mid_1[3247:3240] > btm_0[3239:3232]) ? 1 : 0;
assign detect_max[404][18] = (mid_1[3247:3240] > btm_0[3247:3240]) ? 1 : 0;
assign detect_max[404][19] = (mid_1[3247:3240] > btm_0[3255:3248]) ? 1 : 0;
assign detect_max[404][20] = (mid_1[3247:3240] > btm_1[3239:3232]) ? 1 : 0;
assign detect_max[404][21] = (mid_1[3247:3240] > btm_1[3247:3240]) ? 1 : 0;
assign detect_max[404][22] = (mid_1[3247:3240] > btm_1[3255:3248]) ? 1 : 0;
assign detect_max[404][23] = (mid_1[3247:3240] > btm_2[3239:3232]) ? 1 : 0;
assign detect_max[404][24] = (mid_1[3247:3240] > btm_2[3247:3240]) ? 1 : 0;
assign detect_max[404][25] = (mid_1[3247:3240] > btm_2[3255:3248]) ? 1 : 0;

assign detect_max[405][0] = (mid_1[3255:3248] > top_0[3247:3240]) ? 1 : 0;
assign detect_max[405][1] = (mid_1[3255:3248] > top_0[3255:3248]) ? 1 : 0;
assign detect_max[405][2] = (mid_1[3255:3248] > top_0[3263:3256]) ? 1 : 0;
assign detect_max[405][3] = (mid_1[3255:3248] > top_1[3247:3240]) ? 1 : 0;
assign detect_max[405][4] = (mid_1[3255:3248] > top_1[3255:3248]) ? 1 : 0;
assign detect_max[405][5] = (mid_1[3255:3248] > top_1[3263:3256]) ? 1 : 0;
assign detect_max[405][6] = (mid_1[3255:3248] > top_2[3247:3240]) ? 1 : 0;
assign detect_max[405][7] = (mid_1[3255:3248] > top_2[3255:3248]) ? 1 : 0;
assign detect_max[405][8] = (mid_1[3255:3248] > top_2[3263:3256]) ? 1 : 0;
assign detect_max[405][9] = (mid_1[3255:3248] > mid_0[3247:3240]) ? 1 : 0;
assign detect_max[405][10] = (mid_1[3255:3248] > mid_0[3255:3248]) ? 1 : 0;
assign detect_max[405][11] = (mid_1[3255:3248] > mid_0[3263:3256]) ? 1 : 0;
assign detect_max[405][12] = (mid_1[3255:3248] > mid_1[3247:3240]) ? 1 : 0;
assign detect_max[405][13] = (mid_1[3255:3248] > mid_1[3263:3256]) ? 1 : 0;
assign detect_max[405][14] = (mid_1[3255:3248] > mid_2[3247:3240]) ? 1 : 0;
assign detect_max[405][15] = (mid_1[3255:3248] > mid_2[3255:3248]) ? 1 : 0;
assign detect_max[405][16] = (mid_1[3255:3248] > mid_2[3263:3256]) ? 1 : 0;
assign detect_max[405][17] = (mid_1[3255:3248] > btm_0[3247:3240]) ? 1 : 0;
assign detect_max[405][18] = (mid_1[3255:3248] > btm_0[3255:3248]) ? 1 : 0;
assign detect_max[405][19] = (mid_1[3255:3248] > btm_0[3263:3256]) ? 1 : 0;
assign detect_max[405][20] = (mid_1[3255:3248] > btm_1[3247:3240]) ? 1 : 0;
assign detect_max[405][21] = (mid_1[3255:3248] > btm_1[3255:3248]) ? 1 : 0;
assign detect_max[405][22] = (mid_1[3255:3248] > btm_1[3263:3256]) ? 1 : 0;
assign detect_max[405][23] = (mid_1[3255:3248] > btm_2[3247:3240]) ? 1 : 0;
assign detect_max[405][24] = (mid_1[3255:3248] > btm_2[3255:3248]) ? 1 : 0;
assign detect_max[405][25] = (mid_1[3255:3248] > btm_2[3263:3256]) ? 1 : 0;

assign detect_max[406][0] = (mid_1[3263:3256] > top_0[3255:3248]) ? 1 : 0;
assign detect_max[406][1] = (mid_1[3263:3256] > top_0[3263:3256]) ? 1 : 0;
assign detect_max[406][2] = (mid_1[3263:3256] > top_0[3271:3264]) ? 1 : 0;
assign detect_max[406][3] = (mid_1[3263:3256] > top_1[3255:3248]) ? 1 : 0;
assign detect_max[406][4] = (mid_1[3263:3256] > top_1[3263:3256]) ? 1 : 0;
assign detect_max[406][5] = (mid_1[3263:3256] > top_1[3271:3264]) ? 1 : 0;
assign detect_max[406][6] = (mid_1[3263:3256] > top_2[3255:3248]) ? 1 : 0;
assign detect_max[406][7] = (mid_1[3263:3256] > top_2[3263:3256]) ? 1 : 0;
assign detect_max[406][8] = (mid_1[3263:3256] > top_2[3271:3264]) ? 1 : 0;
assign detect_max[406][9] = (mid_1[3263:3256] > mid_0[3255:3248]) ? 1 : 0;
assign detect_max[406][10] = (mid_1[3263:3256] > mid_0[3263:3256]) ? 1 : 0;
assign detect_max[406][11] = (mid_1[3263:3256] > mid_0[3271:3264]) ? 1 : 0;
assign detect_max[406][12] = (mid_1[3263:3256] > mid_1[3255:3248]) ? 1 : 0;
assign detect_max[406][13] = (mid_1[3263:3256] > mid_1[3271:3264]) ? 1 : 0;
assign detect_max[406][14] = (mid_1[3263:3256] > mid_2[3255:3248]) ? 1 : 0;
assign detect_max[406][15] = (mid_1[3263:3256] > mid_2[3263:3256]) ? 1 : 0;
assign detect_max[406][16] = (mid_1[3263:3256] > mid_2[3271:3264]) ? 1 : 0;
assign detect_max[406][17] = (mid_1[3263:3256] > btm_0[3255:3248]) ? 1 : 0;
assign detect_max[406][18] = (mid_1[3263:3256] > btm_0[3263:3256]) ? 1 : 0;
assign detect_max[406][19] = (mid_1[3263:3256] > btm_0[3271:3264]) ? 1 : 0;
assign detect_max[406][20] = (mid_1[3263:3256] > btm_1[3255:3248]) ? 1 : 0;
assign detect_max[406][21] = (mid_1[3263:3256] > btm_1[3263:3256]) ? 1 : 0;
assign detect_max[406][22] = (mid_1[3263:3256] > btm_1[3271:3264]) ? 1 : 0;
assign detect_max[406][23] = (mid_1[3263:3256] > btm_2[3255:3248]) ? 1 : 0;
assign detect_max[406][24] = (mid_1[3263:3256] > btm_2[3263:3256]) ? 1 : 0;
assign detect_max[406][25] = (mid_1[3263:3256] > btm_2[3271:3264]) ? 1 : 0;

assign detect_max[407][0] = (mid_1[3271:3264] > top_0[3263:3256]) ? 1 : 0;
assign detect_max[407][1] = (mid_1[3271:3264] > top_0[3271:3264]) ? 1 : 0;
assign detect_max[407][2] = (mid_1[3271:3264] > top_0[3279:3272]) ? 1 : 0;
assign detect_max[407][3] = (mid_1[3271:3264] > top_1[3263:3256]) ? 1 : 0;
assign detect_max[407][4] = (mid_1[3271:3264] > top_1[3271:3264]) ? 1 : 0;
assign detect_max[407][5] = (mid_1[3271:3264] > top_1[3279:3272]) ? 1 : 0;
assign detect_max[407][6] = (mid_1[3271:3264] > top_2[3263:3256]) ? 1 : 0;
assign detect_max[407][7] = (mid_1[3271:3264] > top_2[3271:3264]) ? 1 : 0;
assign detect_max[407][8] = (mid_1[3271:3264] > top_2[3279:3272]) ? 1 : 0;
assign detect_max[407][9] = (mid_1[3271:3264] > mid_0[3263:3256]) ? 1 : 0;
assign detect_max[407][10] = (mid_1[3271:3264] > mid_0[3271:3264]) ? 1 : 0;
assign detect_max[407][11] = (mid_1[3271:3264] > mid_0[3279:3272]) ? 1 : 0;
assign detect_max[407][12] = (mid_1[3271:3264] > mid_1[3263:3256]) ? 1 : 0;
assign detect_max[407][13] = (mid_1[3271:3264] > mid_1[3279:3272]) ? 1 : 0;
assign detect_max[407][14] = (mid_1[3271:3264] > mid_2[3263:3256]) ? 1 : 0;
assign detect_max[407][15] = (mid_1[3271:3264] > mid_2[3271:3264]) ? 1 : 0;
assign detect_max[407][16] = (mid_1[3271:3264] > mid_2[3279:3272]) ? 1 : 0;
assign detect_max[407][17] = (mid_1[3271:3264] > btm_0[3263:3256]) ? 1 : 0;
assign detect_max[407][18] = (mid_1[3271:3264] > btm_0[3271:3264]) ? 1 : 0;
assign detect_max[407][19] = (mid_1[3271:3264] > btm_0[3279:3272]) ? 1 : 0;
assign detect_max[407][20] = (mid_1[3271:3264] > btm_1[3263:3256]) ? 1 : 0;
assign detect_max[407][21] = (mid_1[3271:3264] > btm_1[3271:3264]) ? 1 : 0;
assign detect_max[407][22] = (mid_1[3271:3264] > btm_1[3279:3272]) ? 1 : 0;
assign detect_max[407][23] = (mid_1[3271:3264] > btm_2[3263:3256]) ? 1 : 0;
assign detect_max[407][24] = (mid_1[3271:3264] > btm_2[3271:3264]) ? 1 : 0;
assign detect_max[407][25] = (mid_1[3271:3264] > btm_2[3279:3272]) ? 1 : 0;

assign detect_max[408][0] = (mid_1[3279:3272] > top_0[3271:3264]) ? 1 : 0;
assign detect_max[408][1] = (mid_1[3279:3272] > top_0[3279:3272]) ? 1 : 0;
assign detect_max[408][2] = (mid_1[3279:3272] > top_0[3287:3280]) ? 1 : 0;
assign detect_max[408][3] = (mid_1[3279:3272] > top_1[3271:3264]) ? 1 : 0;
assign detect_max[408][4] = (mid_1[3279:3272] > top_1[3279:3272]) ? 1 : 0;
assign detect_max[408][5] = (mid_1[3279:3272] > top_1[3287:3280]) ? 1 : 0;
assign detect_max[408][6] = (mid_1[3279:3272] > top_2[3271:3264]) ? 1 : 0;
assign detect_max[408][7] = (mid_1[3279:3272] > top_2[3279:3272]) ? 1 : 0;
assign detect_max[408][8] = (mid_1[3279:3272] > top_2[3287:3280]) ? 1 : 0;
assign detect_max[408][9] = (mid_1[3279:3272] > mid_0[3271:3264]) ? 1 : 0;
assign detect_max[408][10] = (mid_1[3279:3272] > mid_0[3279:3272]) ? 1 : 0;
assign detect_max[408][11] = (mid_1[3279:3272] > mid_0[3287:3280]) ? 1 : 0;
assign detect_max[408][12] = (mid_1[3279:3272] > mid_1[3271:3264]) ? 1 : 0;
assign detect_max[408][13] = (mid_1[3279:3272] > mid_1[3287:3280]) ? 1 : 0;
assign detect_max[408][14] = (mid_1[3279:3272] > mid_2[3271:3264]) ? 1 : 0;
assign detect_max[408][15] = (mid_1[3279:3272] > mid_2[3279:3272]) ? 1 : 0;
assign detect_max[408][16] = (mid_1[3279:3272] > mid_2[3287:3280]) ? 1 : 0;
assign detect_max[408][17] = (mid_1[3279:3272] > btm_0[3271:3264]) ? 1 : 0;
assign detect_max[408][18] = (mid_1[3279:3272] > btm_0[3279:3272]) ? 1 : 0;
assign detect_max[408][19] = (mid_1[3279:3272] > btm_0[3287:3280]) ? 1 : 0;
assign detect_max[408][20] = (mid_1[3279:3272] > btm_1[3271:3264]) ? 1 : 0;
assign detect_max[408][21] = (mid_1[3279:3272] > btm_1[3279:3272]) ? 1 : 0;
assign detect_max[408][22] = (mid_1[3279:3272] > btm_1[3287:3280]) ? 1 : 0;
assign detect_max[408][23] = (mid_1[3279:3272] > btm_2[3271:3264]) ? 1 : 0;
assign detect_max[408][24] = (mid_1[3279:3272] > btm_2[3279:3272]) ? 1 : 0;
assign detect_max[408][25] = (mid_1[3279:3272] > btm_2[3287:3280]) ? 1 : 0;

assign detect_max[409][0] = (mid_1[3287:3280] > top_0[3279:3272]) ? 1 : 0;
assign detect_max[409][1] = (mid_1[3287:3280] > top_0[3287:3280]) ? 1 : 0;
assign detect_max[409][2] = (mid_1[3287:3280] > top_0[3295:3288]) ? 1 : 0;
assign detect_max[409][3] = (mid_1[3287:3280] > top_1[3279:3272]) ? 1 : 0;
assign detect_max[409][4] = (mid_1[3287:3280] > top_1[3287:3280]) ? 1 : 0;
assign detect_max[409][5] = (mid_1[3287:3280] > top_1[3295:3288]) ? 1 : 0;
assign detect_max[409][6] = (mid_1[3287:3280] > top_2[3279:3272]) ? 1 : 0;
assign detect_max[409][7] = (mid_1[3287:3280] > top_2[3287:3280]) ? 1 : 0;
assign detect_max[409][8] = (mid_1[3287:3280] > top_2[3295:3288]) ? 1 : 0;
assign detect_max[409][9] = (mid_1[3287:3280] > mid_0[3279:3272]) ? 1 : 0;
assign detect_max[409][10] = (mid_1[3287:3280] > mid_0[3287:3280]) ? 1 : 0;
assign detect_max[409][11] = (mid_1[3287:3280] > mid_0[3295:3288]) ? 1 : 0;
assign detect_max[409][12] = (mid_1[3287:3280] > mid_1[3279:3272]) ? 1 : 0;
assign detect_max[409][13] = (mid_1[3287:3280] > mid_1[3295:3288]) ? 1 : 0;
assign detect_max[409][14] = (mid_1[3287:3280] > mid_2[3279:3272]) ? 1 : 0;
assign detect_max[409][15] = (mid_1[3287:3280] > mid_2[3287:3280]) ? 1 : 0;
assign detect_max[409][16] = (mid_1[3287:3280] > mid_2[3295:3288]) ? 1 : 0;
assign detect_max[409][17] = (mid_1[3287:3280] > btm_0[3279:3272]) ? 1 : 0;
assign detect_max[409][18] = (mid_1[3287:3280] > btm_0[3287:3280]) ? 1 : 0;
assign detect_max[409][19] = (mid_1[3287:3280] > btm_0[3295:3288]) ? 1 : 0;
assign detect_max[409][20] = (mid_1[3287:3280] > btm_1[3279:3272]) ? 1 : 0;
assign detect_max[409][21] = (mid_1[3287:3280] > btm_1[3287:3280]) ? 1 : 0;
assign detect_max[409][22] = (mid_1[3287:3280] > btm_1[3295:3288]) ? 1 : 0;
assign detect_max[409][23] = (mid_1[3287:3280] > btm_2[3279:3272]) ? 1 : 0;
assign detect_max[409][24] = (mid_1[3287:3280] > btm_2[3287:3280]) ? 1 : 0;
assign detect_max[409][25] = (mid_1[3287:3280] > btm_2[3295:3288]) ? 1 : 0;

assign detect_max[410][0] = (mid_1[3295:3288] > top_0[3287:3280]) ? 1 : 0;
assign detect_max[410][1] = (mid_1[3295:3288] > top_0[3295:3288]) ? 1 : 0;
assign detect_max[410][2] = (mid_1[3295:3288] > top_0[3303:3296]) ? 1 : 0;
assign detect_max[410][3] = (mid_1[3295:3288] > top_1[3287:3280]) ? 1 : 0;
assign detect_max[410][4] = (mid_1[3295:3288] > top_1[3295:3288]) ? 1 : 0;
assign detect_max[410][5] = (mid_1[3295:3288] > top_1[3303:3296]) ? 1 : 0;
assign detect_max[410][6] = (mid_1[3295:3288] > top_2[3287:3280]) ? 1 : 0;
assign detect_max[410][7] = (mid_1[3295:3288] > top_2[3295:3288]) ? 1 : 0;
assign detect_max[410][8] = (mid_1[3295:3288] > top_2[3303:3296]) ? 1 : 0;
assign detect_max[410][9] = (mid_1[3295:3288] > mid_0[3287:3280]) ? 1 : 0;
assign detect_max[410][10] = (mid_1[3295:3288] > mid_0[3295:3288]) ? 1 : 0;
assign detect_max[410][11] = (mid_1[3295:3288] > mid_0[3303:3296]) ? 1 : 0;
assign detect_max[410][12] = (mid_1[3295:3288] > mid_1[3287:3280]) ? 1 : 0;
assign detect_max[410][13] = (mid_1[3295:3288] > mid_1[3303:3296]) ? 1 : 0;
assign detect_max[410][14] = (mid_1[3295:3288] > mid_2[3287:3280]) ? 1 : 0;
assign detect_max[410][15] = (mid_1[3295:3288] > mid_2[3295:3288]) ? 1 : 0;
assign detect_max[410][16] = (mid_1[3295:3288] > mid_2[3303:3296]) ? 1 : 0;
assign detect_max[410][17] = (mid_1[3295:3288] > btm_0[3287:3280]) ? 1 : 0;
assign detect_max[410][18] = (mid_1[3295:3288] > btm_0[3295:3288]) ? 1 : 0;
assign detect_max[410][19] = (mid_1[3295:3288] > btm_0[3303:3296]) ? 1 : 0;
assign detect_max[410][20] = (mid_1[3295:3288] > btm_1[3287:3280]) ? 1 : 0;
assign detect_max[410][21] = (mid_1[3295:3288] > btm_1[3295:3288]) ? 1 : 0;
assign detect_max[410][22] = (mid_1[3295:3288] > btm_1[3303:3296]) ? 1 : 0;
assign detect_max[410][23] = (mid_1[3295:3288] > btm_2[3287:3280]) ? 1 : 0;
assign detect_max[410][24] = (mid_1[3295:3288] > btm_2[3295:3288]) ? 1 : 0;
assign detect_max[410][25] = (mid_1[3295:3288] > btm_2[3303:3296]) ? 1 : 0;

assign detect_max[411][0] = (mid_1[3303:3296] > top_0[3295:3288]) ? 1 : 0;
assign detect_max[411][1] = (mid_1[3303:3296] > top_0[3303:3296]) ? 1 : 0;
assign detect_max[411][2] = (mid_1[3303:3296] > top_0[3311:3304]) ? 1 : 0;
assign detect_max[411][3] = (mid_1[3303:3296] > top_1[3295:3288]) ? 1 : 0;
assign detect_max[411][4] = (mid_1[3303:3296] > top_1[3303:3296]) ? 1 : 0;
assign detect_max[411][5] = (mid_1[3303:3296] > top_1[3311:3304]) ? 1 : 0;
assign detect_max[411][6] = (mid_1[3303:3296] > top_2[3295:3288]) ? 1 : 0;
assign detect_max[411][7] = (mid_1[3303:3296] > top_2[3303:3296]) ? 1 : 0;
assign detect_max[411][8] = (mid_1[3303:3296] > top_2[3311:3304]) ? 1 : 0;
assign detect_max[411][9] = (mid_1[3303:3296] > mid_0[3295:3288]) ? 1 : 0;
assign detect_max[411][10] = (mid_1[3303:3296] > mid_0[3303:3296]) ? 1 : 0;
assign detect_max[411][11] = (mid_1[3303:3296] > mid_0[3311:3304]) ? 1 : 0;
assign detect_max[411][12] = (mid_1[3303:3296] > mid_1[3295:3288]) ? 1 : 0;
assign detect_max[411][13] = (mid_1[3303:3296] > mid_1[3311:3304]) ? 1 : 0;
assign detect_max[411][14] = (mid_1[3303:3296] > mid_2[3295:3288]) ? 1 : 0;
assign detect_max[411][15] = (mid_1[3303:3296] > mid_2[3303:3296]) ? 1 : 0;
assign detect_max[411][16] = (mid_1[3303:3296] > mid_2[3311:3304]) ? 1 : 0;
assign detect_max[411][17] = (mid_1[3303:3296] > btm_0[3295:3288]) ? 1 : 0;
assign detect_max[411][18] = (mid_1[3303:3296] > btm_0[3303:3296]) ? 1 : 0;
assign detect_max[411][19] = (mid_1[3303:3296] > btm_0[3311:3304]) ? 1 : 0;
assign detect_max[411][20] = (mid_1[3303:3296] > btm_1[3295:3288]) ? 1 : 0;
assign detect_max[411][21] = (mid_1[3303:3296] > btm_1[3303:3296]) ? 1 : 0;
assign detect_max[411][22] = (mid_1[3303:3296] > btm_1[3311:3304]) ? 1 : 0;
assign detect_max[411][23] = (mid_1[3303:3296] > btm_2[3295:3288]) ? 1 : 0;
assign detect_max[411][24] = (mid_1[3303:3296] > btm_2[3303:3296]) ? 1 : 0;
assign detect_max[411][25] = (mid_1[3303:3296] > btm_2[3311:3304]) ? 1 : 0;

assign detect_max[412][0] = (mid_1[3311:3304] > top_0[3303:3296]) ? 1 : 0;
assign detect_max[412][1] = (mid_1[3311:3304] > top_0[3311:3304]) ? 1 : 0;
assign detect_max[412][2] = (mid_1[3311:3304] > top_0[3319:3312]) ? 1 : 0;
assign detect_max[412][3] = (mid_1[3311:3304] > top_1[3303:3296]) ? 1 : 0;
assign detect_max[412][4] = (mid_1[3311:3304] > top_1[3311:3304]) ? 1 : 0;
assign detect_max[412][5] = (mid_1[3311:3304] > top_1[3319:3312]) ? 1 : 0;
assign detect_max[412][6] = (mid_1[3311:3304] > top_2[3303:3296]) ? 1 : 0;
assign detect_max[412][7] = (mid_1[3311:3304] > top_2[3311:3304]) ? 1 : 0;
assign detect_max[412][8] = (mid_1[3311:3304] > top_2[3319:3312]) ? 1 : 0;
assign detect_max[412][9] = (mid_1[3311:3304] > mid_0[3303:3296]) ? 1 : 0;
assign detect_max[412][10] = (mid_1[3311:3304] > mid_0[3311:3304]) ? 1 : 0;
assign detect_max[412][11] = (mid_1[3311:3304] > mid_0[3319:3312]) ? 1 : 0;
assign detect_max[412][12] = (mid_1[3311:3304] > mid_1[3303:3296]) ? 1 : 0;
assign detect_max[412][13] = (mid_1[3311:3304] > mid_1[3319:3312]) ? 1 : 0;
assign detect_max[412][14] = (mid_1[3311:3304] > mid_2[3303:3296]) ? 1 : 0;
assign detect_max[412][15] = (mid_1[3311:3304] > mid_2[3311:3304]) ? 1 : 0;
assign detect_max[412][16] = (mid_1[3311:3304] > mid_2[3319:3312]) ? 1 : 0;
assign detect_max[412][17] = (mid_1[3311:3304] > btm_0[3303:3296]) ? 1 : 0;
assign detect_max[412][18] = (mid_1[3311:3304] > btm_0[3311:3304]) ? 1 : 0;
assign detect_max[412][19] = (mid_1[3311:3304] > btm_0[3319:3312]) ? 1 : 0;
assign detect_max[412][20] = (mid_1[3311:3304] > btm_1[3303:3296]) ? 1 : 0;
assign detect_max[412][21] = (mid_1[3311:3304] > btm_1[3311:3304]) ? 1 : 0;
assign detect_max[412][22] = (mid_1[3311:3304] > btm_1[3319:3312]) ? 1 : 0;
assign detect_max[412][23] = (mid_1[3311:3304] > btm_2[3303:3296]) ? 1 : 0;
assign detect_max[412][24] = (mid_1[3311:3304] > btm_2[3311:3304]) ? 1 : 0;
assign detect_max[412][25] = (mid_1[3311:3304] > btm_2[3319:3312]) ? 1 : 0;

assign detect_max[413][0] = (mid_1[3319:3312] > top_0[3311:3304]) ? 1 : 0;
assign detect_max[413][1] = (mid_1[3319:3312] > top_0[3319:3312]) ? 1 : 0;
assign detect_max[413][2] = (mid_1[3319:3312] > top_0[3327:3320]) ? 1 : 0;
assign detect_max[413][3] = (mid_1[3319:3312] > top_1[3311:3304]) ? 1 : 0;
assign detect_max[413][4] = (mid_1[3319:3312] > top_1[3319:3312]) ? 1 : 0;
assign detect_max[413][5] = (mid_1[3319:3312] > top_1[3327:3320]) ? 1 : 0;
assign detect_max[413][6] = (mid_1[3319:3312] > top_2[3311:3304]) ? 1 : 0;
assign detect_max[413][7] = (mid_1[3319:3312] > top_2[3319:3312]) ? 1 : 0;
assign detect_max[413][8] = (mid_1[3319:3312] > top_2[3327:3320]) ? 1 : 0;
assign detect_max[413][9] = (mid_1[3319:3312] > mid_0[3311:3304]) ? 1 : 0;
assign detect_max[413][10] = (mid_1[3319:3312] > mid_0[3319:3312]) ? 1 : 0;
assign detect_max[413][11] = (mid_1[3319:3312] > mid_0[3327:3320]) ? 1 : 0;
assign detect_max[413][12] = (mid_1[3319:3312] > mid_1[3311:3304]) ? 1 : 0;
assign detect_max[413][13] = (mid_1[3319:3312] > mid_1[3327:3320]) ? 1 : 0;
assign detect_max[413][14] = (mid_1[3319:3312] > mid_2[3311:3304]) ? 1 : 0;
assign detect_max[413][15] = (mid_1[3319:3312] > mid_2[3319:3312]) ? 1 : 0;
assign detect_max[413][16] = (mid_1[3319:3312] > mid_2[3327:3320]) ? 1 : 0;
assign detect_max[413][17] = (mid_1[3319:3312] > btm_0[3311:3304]) ? 1 : 0;
assign detect_max[413][18] = (mid_1[3319:3312] > btm_0[3319:3312]) ? 1 : 0;
assign detect_max[413][19] = (mid_1[3319:3312] > btm_0[3327:3320]) ? 1 : 0;
assign detect_max[413][20] = (mid_1[3319:3312] > btm_1[3311:3304]) ? 1 : 0;
assign detect_max[413][21] = (mid_1[3319:3312] > btm_1[3319:3312]) ? 1 : 0;
assign detect_max[413][22] = (mid_1[3319:3312] > btm_1[3327:3320]) ? 1 : 0;
assign detect_max[413][23] = (mid_1[3319:3312] > btm_2[3311:3304]) ? 1 : 0;
assign detect_max[413][24] = (mid_1[3319:3312] > btm_2[3319:3312]) ? 1 : 0;
assign detect_max[413][25] = (mid_1[3319:3312] > btm_2[3327:3320]) ? 1 : 0;

assign detect_max[414][0] = (mid_1[3327:3320] > top_0[3319:3312]) ? 1 : 0;
assign detect_max[414][1] = (mid_1[3327:3320] > top_0[3327:3320]) ? 1 : 0;
assign detect_max[414][2] = (mid_1[3327:3320] > top_0[3335:3328]) ? 1 : 0;
assign detect_max[414][3] = (mid_1[3327:3320] > top_1[3319:3312]) ? 1 : 0;
assign detect_max[414][4] = (mid_1[3327:3320] > top_1[3327:3320]) ? 1 : 0;
assign detect_max[414][5] = (mid_1[3327:3320] > top_1[3335:3328]) ? 1 : 0;
assign detect_max[414][6] = (mid_1[3327:3320] > top_2[3319:3312]) ? 1 : 0;
assign detect_max[414][7] = (mid_1[3327:3320] > top_2[3327:3320]) ? 1 : 0;
assign detect_max[414][8] = (mid_1[3327:3320] > top_2[3335:3328]) ? 1 : 0;
assign detect_max[414][9] = (mid_1[3327:3320] > mid_0[3319:3312]) ? 1 : 0;
assign detect_max[414][10] = (mid_1[3327:3320] > mid_0[3327:3320]) ? 1 : 0;
assign detect_max[414][11] = (mid_1[3327:3320] > mid_0[3335:3328]) ? 1 : 0;
assign detect_max[414][12] = (mid_1[3327:3320] > mid_1[3319:3312]) ? 1 : 0;
assign detect_max[414][13] = (mid_1[3327:3320] > mid_1[3335:3328]) ? 1 : 0;
assign detect_max[414][14] = (mid_1[3327:3320] > mid_2[3319:3312]) ? 1 : 0;
assign detect_max[414][15] = (mid_1[3327:3320] > mid_2[3327:3320]) ? 1 : 0;
assign detect_max[414][16] = (mid_1[3327:3320] > mid_2[3335:3328]) ? 1 : 0;
assign detect_max[414][17] = (mid_1[3327:3320] > btm_0[3319:3312]) ? 1 : 0;
assign detect_max[414][18] = (mid_1[3327:3320] > btm_0[3327:3320]) ? 1 : 0;
assign detect_max[414][19] = (mid_1[3327:3320] > btm_0[3335:3328]) ? 1 : 0;
assign detect_max[414][20] = (mid_1[3327:3320] > btm_1[3319:3312]) ? 1 : 0;
assign detect_max[414][21] = (mid_1[3327:3320] > btm_1[3327:3320]) ? 1 : 0;
assign detect_max[414][22] = (mid_1[3327:3320] > btm_1[3335:3328]) ? 1 : 0;
assign detect_max[414][23] = (mid_1[3327:3320] > btm_2[3319:3312]) ? 1 : 0;
assign detect_max[414][24] = (mid_1[3327:3320] > btm_2[3327:3320]) ? 1 : 0;
assign detect_max[414][25] = (mid_1[3327:3320] > btm_2[3335:3328]) ? 1 : 0;

assign detect_max[415][0] = (mid_1[3335:3328] > top_0[3327:3320]) ? 1 : 0;
assign detect_max[415][1] = (mid_1[3335:3328] > top_0[3335:3328]) ? 1 : 0;
assign detect_max[415][2] = (mid_1[3335:3328] > top_0[3343:3336]) ? 1 : 0;
assign detect_max[415][3] = (mid_1[3335:3328] > top_1[3327:3320]) ? 1 : 0;
assign detect_max[415][4] = (mid_1[3335:3328] > top_1[3335:3328]) ? 1 : 0;
assign detect_max[415][5] = (mid_1[3335:3328] > top_1[3343:3336]) ? 1 : 0;
assign detect_max[415][6] = (mid_1[3335:3328] > top_2[3327:3320]) ? 1 : 0;
assign detect_max[415][7] = (mid_1[3335:3328] > top_2[3335:3328]) ? 1 : 0;
assign detect_max[415][8] = (mid_1[3335:3328] > top_2[3343:3336]) ? 1 : 0;
assign detect_max[415][9] = (mid_1[3335:3328] > mid_0[3327:3320]) ? 1 : 0;
assign detect_max[415][10] = (mid_1[3335:3328] > mid_0[3335:3328]) ? 1 : 0;
assign detect_max[415][11] = (mid_1[3335:3328] > mid_0[3343:3336]) ? 1 : 0;
assign detect_max[415][12] = (mid_1[3335:3328] > mid_1[3327:3320]) ? 1 : 0;
assign detect_max[415][13] = (mid_1[3335:3328] > mid_1[3343:3336]) ? 1 : 0;
assign detect_max[415][14] = (mid_1[3335:3328] > mid_2[3327:3320]) ? 1 : 0;
assign detect_max[415][15] = (mid_1[3335:3328] > mid_2[3335:3328]) ? 1 : 0;
assign detect_max[415][16] = (mid_1[3335:3328] > mid_2[3343:3336]) ? 1 : 0;
assign detect_max[415][17] = (mid_1[3335:3328] > btm_0[3327:3320]) ? 1 : 0;
assign detect_max[415][18] = (mid_1[3335:3328] > btm_0[3335:3328]) ? 1 : 0;
assign detect_max[415][19] = (mid_1[3335:3328] > btm_0[3343:3336]) ? 1 : 0;
assign detect_max[415][20] = (mid_1[3335:3328] > btm_1[3327:3320]) ? 1 : 0;
assign detect_max[415][21] = (mid_1[3335:3328] > btm_1[3335:3328]) ? 1 : 0;
assign detect_max[415][22] = (mid_1[3335:3328] > btm_1[3343:3336]) ? 1 : 0;
assign detect_max[415][23] = (mid_1[3335:3328] > btm_2[3327:3320]) ? 1 : 0;
assign detect_max[415][24] = (mid_1[3335:3328] > btm_2[3335:3328]) ? 1 : 0;
assign detect_max[415][25] = (mid_1[3335:3328] > btm_2[3343:3336]) ? 1 : 0;

assign detect_max[416][0] = (mid_1[3343:3336] > top_0[3335:3328]) ? 1 : 0;
assign detect_max[416][1] = (mid_1[3343:3336] > top_0[3343:3336]) ? 1 : 0;
assign detect_max[416][2] = (mid_1[3343:3336] > top_0[3351:3344]) ? 1 : 0;
assign detect_max[416][3] = (mid_1[3343:3336] > top_1[3335:3328]) ? 1 : 0;
assign detect_max[416][4] = (mid_1[3343:3336] > top_1[3343:3336]) ? 1 : 0;
assign detect_max[416][5] = (mid_1[3343:3336] > top_1[3351:3344]) ? 1 : 0;
assign detect_max[416][6] = (mid_1[3343:3336] > top_2[3335:3328]) ? 1 : 0;
assign detect_max[416][7] = (mid_1[3343:3336] > top_2[3343:3336]) ? 1 : 0;
assign detect_max[416][8] = (mid_1[3343:3336] > top_2[3351:3344]) ? 1 : 0;
assign detect_max[416][9] = (mid_1[3343:3336] > mid_0[3335:3328]) ? 1 : 0;
assign detect_max[416][10] = (mid_1[3343:3336] > mid_0[3343:3336]) ? 1 : 0;
assign detect_max[416][11] = (mid_1[3343:3336] > mid_0[3351:3344]) ? 1 : 0;
assign detect_max[416][12] = (mid_1[3343:3336] > mid_1[3335:3328]) ? 1 : 0;
assign detect_max[416][13] = (mid_1[3343:3336] > mid_1[3351:3344]) ? 1 : 0;
assign detect_max[416][14] = (mid_1[3343:3336] > mid_2[3335:3328]) ? 1 : 0;
assign detect_max[416][15] = (mid_1[3343:3336] > mid_2[3343:3336]) ? 1 : 0;
assign detect_max[416][16] = (mid_1[3343:3336] > mid_2[3351:3344]) ? 1 : 0;
assign detect_max[416][17] = (mid_1[3343:3336] > btm_0[3335:3328]) ? 1 : 0;
assign detect_max[416][18] = (mid_1[3343:3336] > btm_0[3343:3336]) ? 1 : 0;
assign detect_max[416][19] = (mid_1[3343:3336] > btm_0[3351:3344]) ? 1 : 0;
assign detect_max[416][20] = (mid_1[3343:3336] > btm_1[3335:3328]) ? 1 : 0;
assign detect_max[416][21] = (mid_1[3343:3336] > btm_1[3343:3336]) ? 1 : 0;
assign detect_max[416][22] = (mid_1[3343:3336] > btm_1[3351:3344]) ? 1 : 0;
assign detect_max[416][23] = (mid_1[3343:3336] > btm_2[3335:3328]) ? 1 : 0;
assign detect_max[416][24] = (mid_1[3343:3336] > btm_2[3343:3336]) ? 1 : 0;
assign detect_max[416][25] = (mid_1[3343:3336] > btm_2[3351:3344]) ? 1 : 0;

assign detect_max[417][0] = (mid_1[3351:3344] > top_0[3343:3336]) ? 1 : 0;
assign detect_max[417][1] = (mid_1[3351:3344] > top_0[3351:3344]) ? 1 : 0;
assign detect_max[417][2] = (mid_1[3351:3344] > top_0[3359:3352]) ? 1 : 0;
assign detect_max[417][3] = (mid_1[3351:3344] > top_1[3343:3336]) ? 1 : 0;
assign detect_max[417][4] = (mid_1[3351:3344] > top_1[3351:3344]) ? 1 : 0;
assign detect_max[417][5] = (mid_1[3351:3344] > top_1[3359:3352]) ? 1 : 0;
assign detect_max[417][6] = (mid_1[3351:3344] > top_2[3343:3336]) ? 1 : 0;
assign detect_max[417][7] = (mid_1[3351:3344] > top_2[3351:3344]) ? 1 : 0;
assign detect_max[417][8] = (mid_1[3351:3344] > top_2[3359:3352]) ? 1 : 0;
assign detect_max[417][9] = (mid_1[3351:3344] > mid_0[3343:3336]) ? 1 : 0;
assign detect_max[417][10] = (mid_1[3351:3344] > mid_0[3351:3344]) ? 1 : 0;
assign detect_max[417][11] = (mid_1[3351:3344] > mid_0[3359:3352]) ? 1 : 0;
assign detect_max[417][12] = (mid_1[3351:3344] > mid_1[3343:3336]) ? 1 : 0;
assign detect_max[417][13] = (mid_1[3351:3344] > mid_1[3359:3352]) ? 1 : 0;
assign detect_max[417][14] = (mid_1[3351:3344] > mid_2[3343:3336]) ? 1 : 0;
assign detect_max[417][15] = (mid_1[3351:3344] > mid_2[3351:3344]) ? 1 : 0;
assign detect_max[417][16] = (mid_1[3351:3344] > mid_2[3359:3352]) ? 1 : 0;
assign detect_max[417][17] = (mid_1[3351:3344] > btm_0[3343:3336]) ? 1 : 0;
assign detect_max[417][18] = (mid_1[3351:3344] > btm_0[3351:3344]) ? 1 : 0;
assign detect_max[417][19] = (mid_1[3351:3344] > btm_0[3359:3352]) ? 1 : 0;
assign detect_max[417][20] = (mid_1[3351:3344] > btm_1[3343:3336]) ? 1 : 0;
assign detect_max[417][21] = (mid_1[3351:3344] > btm_1[3351:3344]) ? 1 : 0;
assign detect_max[417][22] = (mid_1[3351:3344] > btm_1[3359:3352]) ? 1 : 0;
assign detect_max[417][23] = (mid_1[3351:3344] > btm_2[3343:3336]) ? 1 : 0;
assign detect_max[417][24] = (mid_1[3351:3344] > btm_2[3351:3344]) ? 1 : 0;
assign detect_max[417][25] = (mid_1[3351:3344] > btm_2[3359:3352]) ? 1 : 0;

assign detect_max[418][0] = (mid_1[3359:3352] > top_0[3351:3344]) ? 1 : 0;
assign detect_max[418][1] = (mid_1[3359:3352] > top_0[3359:3352]) ? 1 : 0;
assign detect_max[418][2] = (mid_1[3359:3352] > top_0[3367:3360]) ? 1 : 0;
assign detect_max[418][3] = (mid_1[3359:3352] > top_1[3351:3344]) ? 1 : 0;
assign detect_max[418][4] = (mid_1[3359:3352] > top_1[3359:3352]) ? 1 : 0;
assign detect_max[418][5] = (mid_1[3359:3352] > top_1[3367:3360]) ? 1 : 0;
assign detect_max[418][6] = (mid_1[3359:3352] > top_2[3351:3344]) ? 1 : 0;
assign detect_max[418][7] = (mid_1[3359:3352] > top_2[3359:3352]) ? 1 : 0;
assign detect_max[418][8] = (mid_1[3359:3352] > top_2[3367:3360]) ? 1 : 0;
assign detect_max[418][9] = (mid_1[3359:3352] > mid_0[3351:3344]) ? 1 : 0;
assign detect_max[418][10] = (mid_1[3359:3352] > mid_0[3359:3352]) ? 1 : 0;
assign detect_max[418][11] = (mid_1[3359:3352] > mid_0[3367:3360]) ? 1 : 0;
assign detect_max[418][12] = (mid_1[3359:3352] > mid_1[3351:3344]) ? 1 : 0;
assign detect_max[418][13] = (mid_1[3359:3352] > mid_1[3367:3360]) ? 1 : 0;
assign detect_max[418][14] = (mid_1[3359:3352] > mid_2[3351:3344]) ? 1 : 0;
assign detect_max[418][15] = (mid_1[3359:3352] > mid_2[3359:3352]) ? 1 : 0;
assign detect_max[418][16] = (mid_1[3359:3352] > mid_2[3367:3360]) ? 1 : 0;
assign detect_max[418][17] = (mid_1[3359:3352] > btm_0[3351:3344]) ? 1 : 0;
assign detect_max[418][18] = (mid_1[3359:3352] > btm_0[3359:3352]) ? 1 : 0;
assign detect_max[418][19] = (mid_1[3359:3352] > btm_0[3367:3360]) ? 1 : 0;
assign detect_max[418][20] = (mid_1[3359:3352] > btm_1[3351:3344]) ? 1 : 0;
assign detect_max[418][21] = (mid_1[3359:3352] > btm_1[3359:3352]) ? 1 : 0;
assign detect_max[418][22] = (mid_1[3359:3352] > btm_1[3367:3360]) ? 1 : 0;
assign detect_max[418][23] = (mid_1[3359:3352] > btm_2[3351:3344]) ? 1 : 0;
assign detect_max[418][24] = (mid_1[3359:3352] > btm_2[3359:3352]) ? 1 : 0;
assign detect_max[418][25] = (mid_1[3359:3352] > btm_2[3367:3360]) ? 1 : 0;

assign detect_max[419][0] = (mid_1[3367:3360] > top_0[3359:3352]) ? 1 : 0;
assign detect_max[419][1] = (mid_1[3367:3360] > top_0[3367:3360]) ? 1 : 0;
assign detect_max[419][2] = (mid_1[3367:3360] > top_0[3375:3368]) ? 1 : 0;
assign detect_max[419][3] = (mid_1[3367:3360] > top_1[3359:3352]) ? 1 : 0;
assign detect_max[419][4] = (mid_1[3367:3360] > top_1[3367:3360]) ? 1 : 0;
assign detect_max[419][5] = (mid_1[3367:3360] > top_1[3375:3368]) ? 1 : 0;
assign detect_max[419][6] = (mid_1[3367:3360] > top_2[3359:3352]) ? 1 : 0;
assign detect_max[419][7] = (mid_1[3367:3360] > top_2[3367:3360]) ? 1 : 0;
assign detect_max[419][8] = (mid_1[3367:3360] > top_2[3375:3368]) ? 1 : 0;
assign detect_max[419][9] = (mid_1[3367:3360] > mid_0[3359:3352]) ? 1 : 0;
assign detect_max[419][10] = (mid_1[3367:3360] > mid_0[3367:3360]) ? 1 : 0;
assign detect_max[419][11] = (mid_1[3367:3360] > mid_0[3375:3368]) ? 1 : 0;
assign detect_max[419][12] = (mid_1[3367:3360] > mid_1[3359:3352]) ? 1 : 0;
assign detect_max[419][13] = (mid_1[3367:3360] > mid_1[3375:3368]) ? 1 : 0;
assign detect_max[419][14] = (mid_1[3367:3360] > mid_2[3359:3352]) ? 1 : 0;
assign detect_max[419][15] = (mid_1[3367:3360] > mid_2[3367:3360]) ? 1 : 0;
assign detect_max[419][16] = (mid_1[3367:3360] > mid_2[3375:3368]) ? 1 : 0;
assign detect_max[419][17] = (mid_1[3367:3360] > btm_0[3359:3352]) ? 1 : 0;
assign detect_max[419][18] = (mid_1[3367:3360] > btm_0[3367:3360]) ? 1 : 0;
assign detect_max[419][19] = (mid_1[3367:3360] > btm_0[3375:3368]) ? 1 : 0;
assign detect_max[419][20] = (mid_1[3367:3360] > btm_1[3359:3352]) ? 1 : 0;
assign detect_max[419][21] = (mid_1[3367:3360] > btm_1[3367:3360]) ? 1 : 0;
assign detect_max[419][22] = (mid_1[3367:3360] > btm_1[3375:3368]) ? 1 : 0;
assign detect_max[419][23] = (mid_1[3367:3360] > btm_2[3359:3352]) ? 1 : 0;
assign detect_max[419][24] = (mid_1[3367:3360] > btm_2[3367:3360]) ? 1 : 0;
assign detect_max[419][25] = (mid_1[3367:3360] > btm_2[3375:3368]) ? 1 : 0;

assign detect_max[420][0] = (mid_1[3375:3368] > top_0[3367:3360]) ? 1 : 0;
assign detect_max[420][1] = (mid_1[3375:3368] > top_0[3375:3368]) ? 1 : 0;
assign detect_max[420][2] = (mid_1[3375:3368] > top_0[3383:3376]) ? 1 : 0;
assign detect_max[420][3] = (mid_1[3375:3368] > top_1[3367:3360]) ? 1 : 0;
assign detect_max[420][4] = (mid_1[3375:3368] > top_1[3375:3368]) ? 1 : 0;
assign detect_max[420][5] = (mid_1[3375:3368] > top_1[3383:3376]) ? 1 : 0;
assign detect_max[420][6] = (mid_1[3375:3368] > top_2[3367:3360]) ? 1 : 0;
assign detect_max[420][7] = (mid_1[3375:3368] > top_2[3375:3368]) ? 1 : 0;
assign detect_max[420][8] = (mid_1[3375:3368] > top_2[3383:3376]) ? 1 : 0;
assign detect_max[420][9] = (mid_1[3375:3368] > mid_0[3367:3360]) ? 1 : 0;
assign detect_max[420][10] = (mid_1[3375:3368] > mid_0[3375:3368]) ? 1 : 0;
assign detect_max[420][11] = (mid_1[3375:3368] > mid_0[3383:3376]) ? 1 : 0;
assign detect_max[420][12] = (mid_1[3375:3368] > mid_1[3367:3360]) ? 1 : 0;
assign detect_max[420][13] = (mid_1[3375:3368] > mid_1[3383:3376]) ? 1 : 0;
assign detect_max[420][14] = (mid_1[3375:3368] > mid_2[3367:3360]) ? 1 : 0;
assign detect_max[420][15] = (mid_1[3375:3368] > mid_2[3375:3368]) ? 1 : 0;
assign detect_max[420][16] = (mid_1[3375:3368] > mid_2[3383:3376]) ? 1 : 0;
assign detect_max[420][17] = (mid_1[3375:3368] > btm_0[3367:3360]) ? 1 : 0;
assign detect_max[420][18] = (mid_1[3375:3368] > btm_0[3375:3368]) ? 1 : 0;
assign detect_max[420][19] = (mid_1[3375:3368] > btm_0[3383:3376]) ? 1 : 0;
assign detect_max[420][20] = (mid_1[3375:3368] > btm_1[3367:3360]) ? 1 : 0;
assign detect_max[420][21] = (mid_1[3375:3368] > btm_1[3375:3368]) ? 1 : 0;
assign detect_max[420][22] = (mid_1[3375:3368] > btm_1[3383:3376]) ? 1 : 0;
assign detect_max[420][23] = (mid_1[3375:3368] > btm_2[3367:3360]) ? 1 : 0;
assign detect_max[420][24] = (mid_1[3375:3368] > btm_2[3375:3368]) ? 1 : 0;
assign detect_max[420][25] = (mid_1[3375:3368] > btm_2[3383:3376]) ? 1 : 0;

assign detect_max[421][0] = (mid_1[3383:3376] > top_0[3375:3368]) ? 1 : 0;
assign detect_max[421][1] = (mid_1[3383:3376] > top_0[3383:3376]) ? 1 : 0;
assign detect_max[421][2] = (mid_1[3383:3376] > top_0[3391:3384]) ? 1 : 0;
assign detect_max[421][3] = (mid_1[3383:3376] > top_1[3375:3368]) ? 1 : 0;
assign detect_max[421][4] = (mid_1[3383:3376] > top_1[3383:3376]) ? 1 : 0;
assign detect_max[421][5] = (mid_1[3383:3376] > top_1[3391:3384]) ? 1 : 0;
assign detect_max[421][6] = (mid_1[3383:3376] > top_2[3375:3368]) ? 1 : 0;
assign detect_max[421][7] = (mid_1[3383:3376] > top_2[3383:3376]) ? 1 : 0;
assign detect_max[421][8] = (mid_1[3383:3376] > top_2[3391:3384]) ? 1 : 0;
assign detect_max[421][9] = (mid_1[3383:3376] > mid_0[3375:3368]) ? 1 : 0;
assign detect_max[421][10] = (mid_1[3383:3376] > mid_0[3383:3376]) ? 1 : 0;
assign detect_max[421][11] = (mid_1[3383:3376] > mid_0[3391:3384]) ? 1 : 0;
assign detect_max[421][12] = (mid_1[3383:3376] > mid_1[3375:3368]) ? 1 : 0;
assign detect_max[421][13] = (mid_1[3383:3376] > mid_1[3391:3384]) ? 1 : 0;
assign detect_max[421][14] = (mid_1[3383:3376] > mid_2[3375:3368]) ? 1 : 0;
assign detect_max[421][15] = (mid_1[3383:3376] > mid_2[3383:3376]) ? 1 : 0;
assign detect_max[421][16] = (mid_1[3383:3376] > mid_2[3391:3384]) ? 1 : 0;
assign detect_max[421][17] = (mid_1[3383:3376] > btm_0[3375:3368]) ? 1 : 0;
assign detect_max[421][18] = (mid_1[3383:3376] > btm_0[3383:3376]) ? 1 : 0;
assign detect_max[421][19] = (mid_1[3383:3376] > btm_0[3391:3384]) ? 1 : 0;
assign detect_max[421][20] = (mid_1[3383:3376] > btm_1[3375:3368]) ? 1 : 0;
assign detect_max[421][21] = (mid_1[3383:3376] > btm_1[3383:3376]) ? 1 : 0;
assign detect_max[421][22] = (mid_1[3383:3376] > btm_1[3391:3384]) ? 1 : 0;
assign detect_max[421][23] = (mid_1[3383:3376] > btm_2[3375:3368]) ? 1 : 0;
assign detect_max[421][24] = (mid_1[3383:3376] > btm_2[3383:3376]) ? 1 : 0;
assign detect_max[421][25] = (mid_1[3383:3376] > btm_2[3391:3384]) ? 1 : 0;

assign detect_max[422][0] = (mid_1[3391:3384] > top_0[3383:3376]) ? 1 : 0;
assign detect_max[422][1] = (mid_1[3391:3384] > top_0[3391:3384]) ? 1 : 0;
assign detect_max[422][2] = (mid_1[3391:3384] > top_0[3399:3392]) ? 1 : 0;
assign detect_max[422][3] = (mid_1[3391:3384] > top_1[3383:3376]) ? 1 : 0;
assign detect_max[422][4] = (mid_1[3391:3384] > top_1[3391:3384]) ? 1 : 0;
assign detect_max[422][5] = (mid_1[3391:3384] > top_1[3399:3392]) ? 1 : 0;
assign detect_max[422][6] = (mid_1[3391:3384] > top_2[3383:3376]) ? 1 : 0;
assign detect_max[422][7] = (mid_1[3391:3384] > top_2[3391:3384]) ? 1 : 0;
assign detect_max[422][8] = (mid_1[3391:3384] > top_2[3399:3392]) ? 1 : 0;
assign detect_max[422][9] = (mid_1[3391:3384] > mid_0[3383:3376]) ? 1 : 0;
assign detect_max[422][10] = (mid_1[3391:3384] > mid_0[3391:3384]) ? 1 : 0;
assign detect_max[422][11] = (mid_1[3391:3384] > mid_0[3399:3392]) ? 1 : 0;
assign detect_max[422][12] = (mid_1[3391:3384] > mid_1[3383:3376]) ? 1 : 0;
assign detect_max[422][13] = (mid_1[3391:3384] > mid_1[3399:3392]) ? 1 : 0;
assign detect_max[422][14] = (mid_1[3391:3384] > mid_2[3383:3376]) ? 1 : 0;
assign detect_max[422][15] = (mid_1[3391:3384] > mid_2[3391:3384]) ? 1 : 0;
assign detect_max[422][16] = (mid_1[3391:3384] > mid_2[3399:3392]) ? 1 : 0;
assign detect_max[422][17] = (mid_1[3391:3384] > btm_0[3383:3376]) ? 1 : 0;
assign detect_max[422][18] = (mid_1[3391:3384] > btm_0[3391:3384]) ? 1 : 0;
assign detect_max[422][19] = (mid_1[3391:3384] > btm_0[3399:3392]) ? 1 : 0;
assign detect_max[422][20] = (mid_1[3391:3384] > btm_1[3383:3376]) ? 1 : 0;
assign detect_max[422][21] = (mid_1[3391:3384] > btm_1[3391:3384]) ? 1 : 0;
assign detect_max[422][22] = (mid_1[3391:3384] > btm_1[3399:3392]) ? 1 : 0;
assign detect_max[422][23] = (mid_1[3391:3384] > btm_2[3383:3376]) ? 1 : 0;
assign detect_max[422][24] = (mid_1[3391:3384] > btm_2[3391:3384]) ? 1 : 0;
assign detect_max[422][25] = (mid_1[3391:3384] > btm_2[3399:3392]) ? 1 : 0;

assign detect_max[423][0] = (mid_1[3399:3392] > top_0[3391:3384]) ? 1 : 0;
assign detect_max[423][1] = (mid_1[3399:3392] > top_0[3399:3392]) ? 1 : 0;
assign detect_max[423][2] = (mid_1[3399:3392] > top_0[3407:3400]) ? 1 : 0;
assign detect_max[423][3] = (mid_1[3399:3392] > top_1[3391:3384]) ? 1 : 0;
assign detect_max[423][4] = (mid_1[3399:3392] > top_1[3399:3392]) ? 1 : 0;
assign detect_max[423][5] = (mid_1[3399:3392] > top_1[3407:3400]) ? 1 : 0;
assign detect_max[423][6] = (mid_1[3399:3392] > top_2[3391:3384]) ? 1 : 0;
assign detect_max[423][7] = (mid_1[3399:3392] > top_2[3399:3392]) ? 1 : 0;
assign detect_max[423][8] = (mid_1[3399:3392] > top_2[3407:3400]) ? 1 : 0;
assign detect_max[423][9] = (mid_1[3399:3392] > mid_0[3391:3384]) ? 1 : 0;
assign detect_max[423][10] = (mid_1[3399:3392] > mid_0[3399:3392]) ? 1 : 0;
assign detect_max[423][11] = (mid_1[3399:3392] > mid_0[3407:3400]) ? 1 : 0;
assign detect_max[423][12] = (mid_1[3399:3392] > mid_1[3391:3384]) ? 1 : 0;
assign detect_max[423][13] = (mid_1[3399:3392] > mid_1[3407:3400]) ? 1 : 0;
assign detect_max[423][14] = (mid_1[3399:3392] > mid_2[3391:3384]) ? 1 : 0;
assign detect_max[423][15] = (mid_1[3399:3392] > mid_2[3399:3392]) ? 1 : 0;
assign detect_max[423][16] = (mid_1[3399:3392] > mid_2[3407:3400]) ? 1 : 0;
assign detect_max[423][17] = (mid_1[3399:3392] > btm_0[3391:3384]) ? 1 : 0;
assign detect_max[423][18] = (mid_1[3399:3392] > btm_0[3399:3392]) ? 1 : 0;
assign detect_max[423][19] = (mid_1[3399:3392] > btm_0[3407:3400]) ? 1 : 0;
assign detect_max[423][20] = (mid_1[3399:3392] > btm_1[3391:3384]) ? 1 : 0;
assign detect_max[423][21] = (mid_1[3399:3392] > btm_1[3399:3392]) ? 1 : 0;
assign detect_max[423][22] = (mid_1[3399:3392] > btm_1[3407:3400]) ? 1 : 0;
assign detect_max[423][23] = (mid_1[3399:3392] > btm_2[3391:3384]) ? 1 : 0;
assign detect_max[423][24] = (mid_1[3399:3392] > btm_2[3399:3392]) ? 1 : 0;
assign detect_max[423][25] = (mid_1[3399:3392] > btm_2[3407:3400]) ? 1 : 0;

assign detect_max[424][0] = (mid_1[3407:3400] > top_0[3399:3392]) ? 1 : 0;
assign detect_max[424][1] = (mid_1[3407:3400] > top_0[3407:3400]) ? 1 : 0;
assign detect_max[424][2] = (mid_1[3407:3400] > top_0[3415:3408]) ? 1 : 0;
assign detect_max[424][3] = (mid_1[3407:3400] > top_1[3399:3392]) ? 1 : 0;
assign detect_max[424][4] = (mid_1[3407:3400] > top_1[3407:3400]) ? 1 : 0;
assign detect_max[424][5] = (mid_1[3407:3400] > top_1[3415:3408]) ? 1 : 0;
assign detect_max[424][6] = (mid_1[3407:3400] > top_2[3399:3392]) ? 1 : 0;
assign detect_max[424][7] = (mid_1[3407:3400] > top_2[3407:3400]) ? 1 : 0;
assign detect_max[424][8] = (mid_1[3407:3400] > top_2[3415:3408]) ? 1 : 0;
assign detect_max[424][9] = (mid_1[3407:3400] > mid_0[3399:3392]) ? 1 : 0;
assign detect_max[424][10] = (mid_1[3407:3400] > mid_0[3407:3400]) ? 1 : 0;
assign detect_max[424][11] = (mid_1[3407:3400] > mid_0[3415:3408]) ? 1 : 0;
assign detect_max[424][12] = (mid_1[3407:3400] > mid_1[3399:3392]) ? 1 : 0;
assign detect_max[424][13] = (mid_1[3407:3400] > mid_1[3415:3408]) ? 1 : 0;
assign detect_max[424][14] = (mid_1[3407:3400] > mid_2[3399:3392]) ? 1 : 0;
assign detect_max[424][15] = (mid_1[3407:3400] > mid_2[3407:3400]) ? 1 : 0;
assign detect_max[424][16] = (mid_1[3407:3400] > mid_2[3415:3408]) ? 1 : 0;
assign detect_max[424][17] = (mid_1[3407:3400] > btm_0[3399:3392]) ? 1 : 0;
assign detect_max[424][18] = (mid_1[3407:3400] > btm_0[3407:3400]) ? 1 : 0;
assign detect_max[424][19] = (mid_1[3407:3400] > btm_0[3415:3408]) ? 1 : 0;
assign detect_max[424][20] = (mid_1[3407:3400] > btm_1[3399:3392]) ? 1 : 0;
assign detect_max[424][21] = (mid_1[3407:3400] > btm_1[3407:3400]) ? 1 : 0;
assign detect_max[424][22] = (mid_1[3407:3400] > btm_1[3415:3408]) ? 1 : 0;
assign detect_max[424][23] = (mid_1[3407:3400] > btm_2[3399:3392]) ? 1 : 0;
assign detect_max[424][24] = (mid_1[3407:3400] > btm_2[3407:3400]) ? 1 : 0;
assign detect_max[424][25] = (mid_1[3407:3400] > btm_2[3415:3408]) ? 1 : 0;

assign detect_max[425][0] = (mid_1[3415:3408] > top_0[3407:3400]) ? 1 : 0;
assign detect_max[425][1] = (mid_1[3415:3408] > top_0[3415:3408]) ? 1 : 0;
assign detect_max[425][2] = (mid_1[3415:3408] > top_0[3423:3416]) ? 1 : 0;
assign detect_max[425][3] = (mid_1[3415:3408] > top_1[3407:3400]) ? 1 : 0;
assign detect_max[425][4] = (mid_1[3415:3408] > top_1[3415:3408]) ? 1 : 0;
assign detect_max[425][5] = (mid_1[3415:3408] > top_1[3423:3416]) ? 1 : 0;
assign detect_max[425][6] = (mid_1[3415:3408] > top_2[3407:3400]) ? 1 : 0;
assign detect_max[425][7] = (mid_1[3415:3408] > top_2[3415:3408]) ? 1 : 0;
assign detect_max[425][8] = (mid_1[3415:3408] > top_2[3423:3416]) ? 1 : 0;
assign detect_max[425][9] = (mid_1[3415:3408] > mid_0[3407:3400]) ? 1 : 0;
assign detect_max[425][10] = (mid_1[3415:3408] > mid_0[3415:3408]) ? 1 : 0;
assign detect_max[425][11] = (mid_1[3415:3408] > mid_0[3423:3416]) ? 1 : 0;
assign detect_max[425][12] = (mid_1[3415:3408] > mid_1[3407:3400]) ? 1 : 0;
assign detect_max[425][13] = (mid_1[3415:3408] > mid_1[3423:3416]) ? 1 : 0;
assign detect_max[425][14] = (mid_1[3415:3408] > mid_2[3407:3400]) ? 1 : 0;
assign detect_max[425][15] = (mid_1[3415:3408] > mid_2[3415:3408]) ? 1 : 0;
assign detect_max[425][16] = (mid_1[3415:3408] > mid_2[3423:3416]) ? 1 : 0;
assign detect_max[425][17] = (mid_1[3415:3408] > btm_0[3407:3400]) ? 1 : 0;
assign detect_max[425][18] = (mid_1[3415:3408] > btm_0[3415:3408]) ? 1 : 0;
assign detect_max[425][19] = (mid_1[3415:3408] > btm_0[3423:3416]) ? 1 : 0;
assign detect_max[425][20] = (mid_1[3415:3408] > btm_1[3407:3400]) ? 1 : 0;
assign detect_max[425][21] = (mid_1[3415:3408] > btm_1[3415:3408]) ? 1 : 0;
assign detect_max[425][22] = (mid_1[3415:3408] > btm_1[3423:3416]) ? 1 : 0;
assign detect_max[425][23] = (mid_1[3415:3408] > btm_2[3407:3400]) ? 1 : 0;
assign detect_max[425][24] = (mid_1[3415:3408] > btm_2[3415:3408]) ? 1 : 0;
assign detect_max[425][25] = (mid_1[3415:3408] > btm_2[3423:3416]) ? 1 : 0;

assign detect_max[426][0] = (mid_1[3423:3416] > top_0[3415:3408]) ? 1 : 0;
assign detect_max[426][1] = (mid_1[3423:3416] > top_0[3423:3416]) ? 1 : 0;
assign detect_max[426][2] = (mid_1[3423:3416] > top_0[3431:3424]) ? 1 : 0;
assign detect_max[426][3] = (mid_1[3423:3416] > top_1[3415:3408]) ? 1 : 0;
assign detect_max[426][4] = (mid_1[3423:3416] > top_1[3423:3416]) ? 1 : 0;
assign detect_max[426][5] = (mid_1[3423:3416] > top_1[3431:3424]) ? 1 : 0;
assign detect_max[426][6] = (mid_1[3423:3416] > top_2[3415:3408]) ? 1 : 0;
assign detect_max[426][7] = (mid_1[3423:3416] > top_2[3423:3416]) ? 1 : 0;
assign detect_max[426][8] = (mid_1[3423:3416] > top_2[3431:3424]) ? 1 : 0;
assign detect_max[426][9] = (mid_1[3423:3416] > mid_0[3415:3408]) ? 1 : 0;
assign detect_max[426][10] = (mid_1[3423:3416] > mid_0[3423:3416]) ? 1 : 0;
assign detect_max[426][11] = (mid_1[3423:3416] > mid_0[3431:3424]) ? 1 : 0;
assign detect_max[426][12] = (mid_1[3423:3416] > mid_1[3415:3408]) ? 1 : 0;
assign detect_max[426][13] = (mid_1[3423:3416] > mid_1[3431:3424]) ? 1 : 0;
assign detect_max[426][14] = (mid_1[3423:3416] > mid_2[3415:3408]) ? 1 : 0;
assign detect_max[426][15] = (mid_1[3423:3416] > mid_2[3423:3416]) ? 1 : 0;
assign detect_max[426][16] = (mid_1[3423:3416] > mid_2[3431:3424]) ? 1 : 0;
assign detect_max[426][17] = (mid_1[3423:3416] > btm_0[3415:3408]) ? 1 : 0;
assign detect_max[426][18] = (mid_1[3423:3416] > btm_0[3423:3416]) ? 1 : 0;
assign detect_max[426][19] = (mid_1[3423:3416] > btm_0[3431:3424]) ? 1 : 0;
assign detect_max[426][20] = (mid_1[3423:3416] > btm_1[3415:3408]) ? 1 : 0;
assign detect_max[426][21] = (mid_1[3423:3416] > btm_1[3423:3416]) ? 1 : 0;
assign detect_max[426][22] = (mid_1[3423:3416] > btm_1[3431:3424]) ? 1 : 0;
assign detect_max[426][23] = (mid_1[3423:3416] > btm_2[3415:3408]) ? 1 : 0;
assign detect_max[426][24] = (mid_1[3423:3416] > btm_2[3423:3416]) ? 1 : 0;
assign detect_max[426][25] = (mid_1[3423:3416] > btm_2[3431:3424]) ? 1 : 0;

assign detect_max[427][0] = (mid_1[3431:3424] > top_0[3423:3416]) ? 1 : 0;
assign detect_max[427][1] = (mid_1[3431:3424] > top_0[3431:3424]) ? 1 : 0;
assign detect_max[427][2] = (mid_1[3431:3424] > top_0[3439:3432]) ? 1 : 0;
assign detect_max[427][3] = (mid_1[3431:3424] > top_1[3423:3416]) ? 1 : 0;
assign detect_max[427][4] = (mid_1[3431:3424] > top_1[3431:3424]) ? 1 : 0;
assign detect_max[427][5] = (mid_1[3431:3424] > top_1[3439:3432]) ? 1 : 0;
assign detect_max[427][6] = (mid_1[3431:3424] > top_2[3423:3416]) ? 1 : 0;
assign detect_max[427][7] = (mid_1[3431:3424] > top_2[3431:3424]) ? 1 : 0;
assign detect_max[427][8] = (mid_1[3431:3424] > top_2[3439:3432]) ? 1 : 0;
assign detect_max[427][9] = (mid_1[3431:3424] > mid_0[3423:3416]) ? 1 : 0;
assign detect_max[427][10] = (mid_1[3431:3424] > mid_0[3431:3424]) ? 1 : 0;
assign detect_max[427][11] = (mid_1[3431:3424] > mid_0[3439:3432]) ? 1 : 0;
assign detect_max[427][12] = (mid_1[3431:3424] > mid_1[3423:3416]) ? 1 : 0;
assign detect_max[427][13] = (mid_1[3431:3424] > mid_1[3439:3432]) ? 1 : 0;
assign detect_max[427][14] = (mid_1[3431:3424] > mid_2[3423:3416]) ? 1 : 0;
assign detect_max[427][15] = (mid_1[3431:3424] > mid_2[3431:3424]) ? 1 : 0;
assign detect_max[427][16] = (mid_1[3431:3424] > mid_2[3439:3432]) ? 1 : 0;
assign detect_max[427][17] = (mid_1[3431:3424] > btm_0[3423:3416]) ? 1 : 0;
assign detect_max[427][18] = (mid_1[3431:3424] > btm_0[3431:3424]) ? 1 : 0;
assign detect_max[427][19] = (mid_1[3431:3424] > btm_0[3439:3432]) ? 1 : 0;
assign detect_max[427][20] = (mid_1[3431:3424] > btm_1[3423:3416]) ? 1 : 0;
assign detect_max[427][21] = (mid_1[3431:3424] > btm_1[3431:3424]) ? 1 : 0;
assign detect_max[427][22] = (mid_1[3431:3424] > btm_1[3439:3432]) ? 1 : 0;
assign detect_max[427][23] = (mid_1[3431:3424] > btm_2[3423:3416]) ? 1 : 0;
assign detect_max[427][24] = (mid_1[3431:3424] > btm_2[3431:3424]) ? 1 : 0;
assign detect_max[427][25] = (mid_1[3431:3424] > btm_2[3439:3432]) ? 1 : 0;

assign detect_max[428][0] = (mid_1[3439:3432] > top_0[3431:3424]) ? 1 : 0;
assign detect_max[428][1] = (mid_1[3439:3432] > top_0[3439:3432]) ? 1 : 0;
assign detect_max[428][2] = (mid_1[3439:3432] > top_0[3447:3440]) ? 1 : 0;
assign detect_max[428][3] = (mid_1[3439:3432] > top_1[3431:3424]) ? 1 : 0;
assign detect_max[428][4] = (mid_1[3439:3432] > top_1[3439:3432]) ? 1 : 0;
assign detect_max[428][5] = (mid_1[3439:3432] > top_1[3447:3440]) ? 1 : 0;
assign detect_max[428][6] = (mid_1[3439:3432] > top_2[3431:3424]) ? 1 : 0;
assign detect_max[428][7] = (mid_1[3439:3432] > top_2[3439:3432]) ? 1 : 0;
assign detect_max[428][8] = (mid_1[3439:3432] > top_2[3447:3440]) ? 1 : 0;
assign detect_max[428][9] = (mid_1[3439:3432] > mid_0[3431:3424]) ? 1 : 0;
assign detect_max[428][10] = (mid_1[3439:3432] > mid_0[3439:3432]) ? 1 : 0;
assign detect_max[428][11] = (mid_1[3439:3432] > mid_0[3447:3440]) ? 1 : 0;
assign detect_max[428][12] = (mid_1[3439:3432] > mid_1[3431:3424]) ? 1 : 0;
assign detect_max[428][13] = (mid_1[3439:3432] > mid_1[3447:3440]) ? 1 : 0;
assign detect_max[428][14] = (mid_1[3439:3432] > mid_2[3431:3424]) ? 1 : 0;
assign detect_max[428][15] = (mid_1[3439:3432] > mid_2[3439:3432]) ? 1 : 0;
assign detect_max[428][16] = (mid_1[3439:3432] > mid_2[3447:3440]) ? 1 : 0;
assign detect_max[428][17] = (mid_1[3439:3432] > btm_0[3431:3424]) ? 1 : 0;
assign detect_max[428][18] = (mid_1[3439:3432] > btm_0[3439:3432]) ? 1 : 0;
assign detect_max[428][19] = (mid_1[3439:3432] > btm_0[3447:3440]) ? 1 : 0;
assign detect_max[428][20] = (mid_1[3439:3432] > btm_1[3431:3424]) ? 1 : 0;
assign detect_max[428][21] = (mid_1[3439:3432] > btm_1[3439:3432]) ? 1 : 0;
assign detect_max[428][22] = (mid_1[3439:3432] > btm_1[3447:3440]) ? 1 : 0;
assign detect_max[428][23] = (mid_1[3439:3432] > btm_2[3431:3424]) ? 1 : 0;
assign detect_max[428][24] = (mid_1[3439:3432] > btm_2[3439:3432]) ? 1 : 0;
assign detect_max[428][25] = (mid_1[3439:3432] > btm_2[3447:3440]) ? 1 : 0;

assign detect_max[429][0] = (mid_1[3447:3440] > top_0[3439:3432]) ? 1 : 0;
assign detect_max[429][1] = (mid_1[3447:3440] > top_0[3447:3440]) ? 1 : 0;
assign detect_max[429][2] = (mid_1[3447:3440] > top_0[3455:3448]) ? 1 : 0;
assign detect_max[429][3] = (mid_1[3447:3440] > top_1[3439:3432]) ? 1 : 0;
assign detect_max[429][4] = (mid_1[3447:3440] > top_1[3447:3440]) ? 1 : 0;
assign detect_max[429][5] = (mid_1[3447:3440] > top_1[3455:3448]) ? 1 : 0;
assign detect_max[429][6] = (mid_1[3447:3440] > top_2[3439:3432]) ? 1 : 0;
assign detect_max[429][7] = (mid_1[3447:3440] > top_2[3447:3440]) ? 1 : 0;
assign detect_max[429][8] = (mid_1[3447:3440] > top_2[3455:3448]) ? 1 : 0;
assign detect_max[429][9] = (mid_1[3447:3440] > mid_0[3439:3432]) ? 1 : 0;
assign detect_max[429][10] = (mid_1[3447:3440] > mid_0[3447:3440]) ? 1 : 0;
assign detect_max[429][11] = (mid_1[3447:3440] > mid_0[3455:3448]) ? 1 : 0;
assign detect_max[429][12] = (mid_1[3447:3440] > mid_1[3439:3432]) ? 1 : 0;
assign detect_max[429][13] = (mid_1[3447:3440] > mid_1[3455:3448]) ? 1 : 0;
assign detect_max[429][14] = (mid_1[3447:3440] > mid_2[3439:3432]) ? 1 : 0;
assign detect_max[429][15] = (mid_1[3447:3440] > mid_2[3447:3440]) ? 1 : 0;
assign detect_max[429][16] = (mid_1[3447:3440] > mid_2[3455:3448]) ? 1 : 0;
assign detect_max[429][17] = (mid_1[3447:3440] > btm_0[3439:3432]) ? 1 : 0;
assign detect_max[429][18] = (mid_1[3447:3440] > btm_0[3447:3440]) ? 1 : 0;
assign detect_max[429][19] = (mid_1[3447:3440] > btm_0[3455:3448]) ? 1 : 0;
assign detect_max[429][20] = (mid_1[3447:3440] > btm_1[3439:3432]) ? 1 : 0;
assign detect_max[429][21] = (mid_1[3447:3440] > btm_1[3447:3440]) ? 1 : 0;
assign detect_max[429][22] = (mid_1[3447:3440] > btm_1[3455:3448]) ? 1 : 0;
assign detect_max[429][23] = (mid_1[3447:3440] > btm_2[3439:3432]) ? 1 : 0;
assign detect_max[429][24] = (mid_1[3447:3440] > btm_2[3447:3440]) ? 1 : 0;
assign detect_max[429][25] = (mid_1[3447:3440] > btm_2[3455:3448]) ? 1 : 0;

assign detect_max[430][0] = (mid_1[3455:3448] > top_0[3447:3440]) ? 1 : 0;
assign detect_max[430][1] = (mid_1[3455:3448] > top_0[3455:3448]) ? 1 : 0;
assign detect_max[430][2] = (mid_1[3455:3448] > top_0[3463:3456]) ? 1 : 0;
assign detect_max[430][3] = (mid_1[3455:3448] > top_1[3447:3440]) ? 1 : 0;
assign detect_max[430][4] = (mid_1[3455:3448] > top_1[3455:3448]) ? 1 : 0;
assign detect_max[430][5] = (mid_1[3455:3448] > top_1[3463:3456]) ? 1 : 0;
assign detect_max[430][6] = (mid_1[3455:3448] > top_2[3447:3440]) ? 1 : 0;
assign detect_max[430][7] = (mid_1[3455:3448] > top_2[3455:3448]) ? 1 : 0;
assign detect_max[430][8] = (mid_1[3455:3448] > top_2[3463:3456]) ? 1 : 0;
assign detect_max[430][9] = (mid_1[3455:3448] > mid_0[3447:3440]) ? 1 : 0;
assign detect_max[430][10] = (mid_1[3455:3448] > mid_0[3455:3448]) ? 1 : 0;
assign detect_max[430][11] = (mid_1[3455:3448] > mid_0[3463:3456]) ? 1 : 0;
assign detect_max[430][12] = (mid_1[3455:3448] > mid_1[3447:3440]) ? 1 : 0;
assign detect_max[430][13] = (mid_1[3455:3448] > mid_1[3463:3456]) ? 1 : 0;
assign detect_max[430][14] = (mid_1[3455:3448] > mid_2[3447:3440]) ? 1 : 0;
assign detect_max[430][15] = (mid_1[3455:3448] > mid_2[3455:3448]) ? 1 : 0;
assign detect_max[430][16] = (mid_1[3455:3448] > mid_2[3463:3456]) ? 1 : 0;
assign detect_max[430][17] = (mid_1[3455:3448] > btm_0[3447:3440]) ? 1 : 0;
assign detect_max[430][18] = (mid_1[3455:3448] > btm_0[3455:3448]) ? 1 : 0;
assign detect_max[430][19] = (mid_1[3455:3448] > btm_0[3463:3456]) ? 1 : 0;
assign detect_max[430][20] = (mid_1[3455:3448] > btm_1[3447:3440]) ? 1 : 0;
assign detect_max[430][21] = (mid_1[3455:3448] > btm_1[3455:3448]) ? 1 : 0;
assign detect_max[430][22] = (mid_1[3455:3448] > btm_1[3463:3456]) ? 1 : 0;
assign detect_max[430][23] = (mid_1[3455:3448] > btm_2[3447:3440]) ? 1 : 0;
assign detect_max[430][24] = (mid_1[3455:3448] > btm_2[3455:3448]) ? 1 : 0;
assign detect_max[430][25] = (mid_1[3455:3448] > btm_2[3463:3456]) ? 1 : 0;

assign detect_max[431][0] = (mid_1[3463:3456] > top_0[3455:3448]) ? 1 : 0;
assign detect_max[431][1] = (mid_1[3463:3456] > top_0[3463:3456]) ? 1 : 0;
assign detect_max[431][2] = (mid_1[3463:3456] > top_0[3471:3464]) ? 1 : 0;
assign detect_max[431][3] = (mid_1[3463:3456] > top_1[3455:3448]) ? 1 : 0;
assign detect_max[431][4] = (mid_1[3463:3456] > top_1[3463:3456]) ? 1 : 0;
assign detect_max[431][5] = (mid_1[3463:3456] > top_1[3471:3464]) ? 1 : 0;
assign detect_max[431][6] = (mid_1[3463:3456] > top_2[3455:3448]) ? 1 : 0;
assign detect_max[431][7] = (mid_1[3463:3456] > top_2[3463:3456]) ? 1 : 0;
assign detect_max[431][8] = (mid_1[3463:3456] > top_2[3471:3464]) ? 1 : 0;
assign detect_max[431][9] = (mid_1[3463:3456] > mid_0[3455:3448]) ? 1 : 0;
assign detect_max[431][10] = (mid_1[3463:3456] > mid_0[3463:3456]) ? 1 : 0;
assign detect_max[431][11] = (mid_1[3463:3456] > mid_0[3471:3464]) ? 1 : 0;
assign detect_max[431][12] = (mid_1[3463:3456] > mid_1[3455:3448]) ? 1 : 0;
assign detect_max[431][13] = (mid_1[3463:3456] > mid_1[3471:3464]) ? 1 : 0;
assign detect_max[431][14] = (mid_1[3463:3456] > mid_2[3455:3448]) ? 1 : 0;
assign detect_max[431][15] = (mid_1[3463:3456] > mid_2[3463:3456]) ? 1 : 0;
assign detect_max[431][16] = (mid_1[3463:3456] > mid_2[3471:3464]) ? 1 : 0;
assign detect_max[431][17] = (mid_1[3463:3456] > btm_0[3455:3448]) ? 1 : 0;
assign detect_max[431][18] = (mid_1[3463:3456] > btm_0[3463:3456]) ? 1 : 0;
assign detect_max[431][19] = (mid_1[3463:3456] > btm_0[3471:3464]) ? 1 : 0;
assign detect_max[431][20] = (mid_1[3463:3456] > btm_1[3455:3448]) ? 1 : 0;
assign detect_max[431][21] = (mid_1[3463:3456] > btm_1[3463:3456]) ? 1 : 0;
assign detect_max[431][22] = (mid_1[3463:3456] > btm_1[3471:3464]) ? 1 : 0;
assign detect_max[431][23] = (mid_1[3463:3456] > btm_2[3455:3448]) ? 1 : 0;
assign detect_max[431][24] = (mid_1[3463:3456] > btm_2[3463:3456]) ? 1 : 0;
assign detect_max[431][25] = (mid_1[3463:3456] > btm_2[3471:3464]) ? 1 : 0;

assign detect_max[432][0] = (mid_1[3471:3464] > top_0[3463:3456]) ? 1 : 0;
assign detect_max[432][1] = (mid_1[3471:3464] > top_0[3471:3464]) ? 1 : 0;
assign detect_max[432][2] = (mid_1[3471:3464] > top_0[3479:3472]) ? 1 : 0;
assign detect_max[432][3] = (mid_1[3471:3464] > top_1[3463:3456]) ? 1 : 0;
assign detect_max[432][4] = (mid_1[3471:3464] > top_1[3471:3464]) ? 1 : 0;
assign detect_max[432][5] = (mid_1[3471:3464] > top_1[3479:3472]) ? 1 : 0;
assign detect_max[432][6] = (mid_1[3471:3464] > top_2[3463:3456]) ? 1 : 0;
assign detect_max[432][7] = (mid_1[3471:3464] > top_2[3471:3464]) ? 1 : 0;
assign detect_max[432][8] = (mid_1[3471:3464] > top_2[3479:3472]) ? 1 : 0;
assign detect_max[432][9] = (mid_1[3471:3464] > mid_0[3463:3456]) ? 1 : 0;
assign detect_max[432][10] = (mid_1[3471:3464] > mid_0[3471:3464]) ? 1 : 0;
assign detect_max[432][11] = (mid_1[3471:3464] > mid_0[3479:3472]) ? 1 : 0;
assign detect_max[432][12] = (mid_1[3471:3464] > mid_1[3463:3456]) ? 1 : 0;
assign detect_max[432][13] = (mid_1[3471:3464] > mid_1[3479:3472]) ? 1 : 0;
assign detect_max[432][14] = (mid_1[3471:3464] > mid_2[3463:3456]) ? 1 : 0;
assign detect_max[432][15] = (mid_1[3471:3464] > mid_2[3471:3464]) ? 1 : 0;
assign detect_max[432][16] = (mid_1[3471:3464] > mid_2[3479:3472]) ? 1 : 0;
assign detect_max[432][17] = (mid_1[3471:3464] > btm_0[3463:3456]) ? 1 : 0;
assign detect_max[432][18] = (mid_1[3471:3464] > btm_0[3471:3464]) ? 1 : 0;
assign detect_max[432][19] = (mid_1[3471:3464] > btm_0[3479:3472]) ? 1 : 0;
assign detect_max[432][20] = (mid_1[3471:3464] > btm_1[3463:3456]) ? 1 : 0;
assign detect_max[432][21] = (mid_1[3471:3464] > btm_1[3471:3464]) ? 1 : 0;
assign detect_max[432][22] = (mid_1[3471:3464] > btm_1[3479:3472]) ? 1 : 0;
assign detect_max[432][23] = (mid_1[3471:3464] > btm_2[3463:3456]) ? 1 : 0;
assign detect_max[432][24] = (mid_1[3471:3464] > btm_2[3471:3464]) ? 1 : 0;
assign detect_max[432][25] = (mid_1[3471:3464] > btm_2[3479:3472]) ? 1 : 0;

assign detect_max[433][0] = (mid_1[3479:3472] > top_0[3471:3464]) ? 1 : 0;
assign detect_max[433][1] = (mid_1[3479:3472] > top_0[3479:3472]) ? 1 : 0;
assign detect_max[433][2] = (mid_1[3479:3472] > top_0[3487:3480]) ? 1 : 0;
assign detect_max[433][3] = (mid_1[3479:3472] > top_1[3471:3464]) ? 1 : 0;
assign detect_max[433][4] = (mid_1[3479:3472] > top_1[3479:3472]) ? 1 : 0;
assign detect_max[433][5] = (mid_1[3479:3472] > top_1[3487:3480]) ? 1 : 0;
assign detect_max[433][6] = (mid_1[3479:3472] > top_2[3471:3464]) ? 1 : 0;
assign detect_max[433][7] = (mid_1[3479:3472] > top_2[3479:3472]) ? 1 : 0;
assign detect_max[433][8] = (mid_1[3479:3472] > top_2[3487:3480]) ? 1 : 0;
assign detect_max[433][9] = (mid_1[3479:3472] > mid_0[3471:3464]) ? 1 : 0;
assign detect_max[433][10] = (mid_1[3479:3472] > mid_0[3479:3472]) ? 1 : 0;
assign detect_max[433][11] = (mid_1[3479:3472] > mid_0[3487:3480]) ? 1 : 0;
assign detect_max[433][12] = (mid_1[3479:3472] > mid_1[3471:3464]) ? 1 : 0;
assign detect_max[433][13] = (mid_1[3479:3472] > mid_1[3487:3480]) ? 1 : 0;
assign detect_max[433][14] = (mid_1[3479:3472] > mid_2[3471:3464]) ? 1 : 0;
assign detect_max[433][15] = (mid_1[3479:3472] > mid_2[3479:3472]) ? 1 : 0;
assign detect_max[433][16] = (mid_1[3479:3472] > mid_2[3487:3480]) ? 1 : 0;
assign detect_max[433][17] = (mid_1[3479:3472] > btm_0[3471:3464]) ? 1 : 0;
assign detect_max[433][18] = (mid_1[3479:3472] > btm_0[3479:3472]) ? 1 : 0;
assign detect_max[433][19] = (mid_1[3479:3472] > btm_0[3487:3480]) ? 1 : 0;
assign detect_max[433][20] = (mid_1[3479:3472] > btm_1[3471:3464]) ? 1 : 0;
assign detect_max[433][21] = (mid_1[3479:3472] > btm_1[3479:3472]) ? 1 : 0;
assign detect_max[433][22] = (mid_1[3479:3472] > btm_1[3487:3480]) ? 1 : 0;
assign detect_max[433][23] = (mid_1[3479:3472] > btm_2[3471:3464]) ? 1 : 0;
assign detect_max[433][24] = (mid_1[3479:3472] > btm_2[3479:3472]) ? 1 : 0;
assign detect_max[433][25] = (mid_1[3479:3472] > btm_2[3487:3480]) ? 1 : 0;

assign detect_max[434][0] = (mid_1[3487:3480] > top_0[3479:3472]) ? 1 : 0;
assign detect_max[434][1] = (mid_1[3487:3480] > top_0[3487:3480]) ? 1 : 0;
assign detect_max[434][2] = (mid_1[3487:3480] > top_0[3495:3488]) ? 1 : 0;
assign detect_max[434][3] = (mid_1[3487:3480] > top_1[3479:3472]) ? 1 : 0;
assign detect_max[434][4] = (mid_1[3487:3480] > top_1[3487:3480]) ? 1 : 0;
assign detect_max[434][5] = (mid_1[3487:3480] > top_1[3495:3488]) ? 1 : 0;
assign detect_max[434][6] = (mid_1[3487:3480] > top_2[3479:3472]) ? 1 : 0;
assign detect_max[434][7] = (mid_1[3487:3480] > top_2[3487:3480]) ? 1 : 0;
assign detect_max[434][8] = (mid_1[3487:3480] > top_2[3495:3488]) ? 1 : 0;
assign detect_max[434][9] = (mid_1[3487:3480] > mid_0[3479:3472]) ? 1 : 0;
assign detect_max[434][10] = (mid_1[3487:3480] > mid_0[3487:3480]) ? 1 : 0;
assign detect_max[434][11] = (mid_1[3487:3480] > mid_0[3495:3488]) ? 1 : 0;
assign detect_max[434][12] = (mid_1[3487:3480] > mid_1[3479:3472]) ? 1 : 0;
assign detect_max[434][13] = (mid_1[3487:3480] > mid_1[3495:3488]) ? 1 : 0;
assign detect_max[434][14] = (mid_1[3487:3480] > mid_2[3479:3472]) ? 1 : 0;
assign detect_max[434][15] = (mid_1[3487:3480] > mid_2[3487:3480]) ? 1 : 0;
assign detect_max[434][16] = (mid_1[3487:3480] > mid_2[3495:3488]) ? 1 : 0;
assign detect_max[434][17] = (mid_1[3487:3480] > btm_0[3479:3472]) ? 1 : 0;
assign detect_max[434][18] = (mid_1[3487:3480] > btm_0[3487:3480]) ? 1 : 0;
assign detect_max[434][19] = (mid_1[3487:3480] > btm_0[3495:3488]) ? 1 : 0;
assign detect_max[434][20] = (mid_1[3487:3480] > btm_1[3479:3472]) ? 1 : 0;
assign detect_max[434][21] = (mid_1[3487:3480] > btm_1[3487:3480]) ? 1 : 0;
assign detect_max[434][22] = (mid_1[3487:3480] > btm_1[3495:3488]) ? 1 : 0;
assign detect_max[434][23] = (mid_1[3487:3480] > btm_2[3479:3472]) ? 1 : 0;
assign detect_max[434][24] = (mid_1[3487:3480] > btm_2[3487:3480]) ? 1 : 0;
assign detect_max[434][25] = (mid_1[3487:3480] > btm_2[3495:3488]) ? 1 : 0;

assign detect_max[435][0] = (mid_1[3495:3488] > top_0[3487:3480]) ? 1 : 0;
assign detect_max[435][1] = (mid_1[3495:3488] > top_0[3495:3488]) ? 1 : 0;
assign detect_max[435][2] = (mid_1[3495:3488] > top_0[3503:3496]) ? 1 : 0;
assign detect_max[435][3] = (mid_1[3495:3488] > top_1[3487:3480]) ? 1 : 0;
assign detect_max[435][4] = (mid_1[3495:3488] > top_1[3495:3488]) ? 1 : 0;
assign detect_max[435][5] = (mid_1[3495:3488] > top_1[3503:3496]) ? 1 : 0;
assign detect_max[435][6] = (mid_1[3495:3488] > top_2[3487:3480]) ? 1 : 0;
assign detect_max[435][7] = (mid_1[3495:3488] > top_2[3495:3488]) ? 1 : 0;
assign detect_max[435][8] = (mid_1[3495:3488] > top_2[3503:3496]) ? 1 : 0;
assign detect_max[435][9] = (mid_1[3495:3488] > mid_0[3487:3480]) ? 1 : 0;
assign detect_max[435][10] = (mid_1[3495:3488] > mid_0[3495:3488]) ? 1 : 0;
assign detect_max[435][11] = (mid_1[3495:3488] > mid_0[3503:3496]) ? 1 : 0;
assign detect_max[435][12] = (mid_1[3495:3488] > mid_1[3487:3480]) ? 1 : 0;
assign detect_max[435][13] = (mid_1[3495:3488] > mid_1[3503:3496]) ? 1 : 0;
assign detect_max[435][14] = (mid_1[3495:3488] > mid_2[3487:3480]) ? 1 : 0;
assign detect_max[435][15] = (mid_1[3495:3488] > mid_2[3495:3488]) ? 1 : 0;
assign detect_max[435][16] = (mid_1[3495:3488] > mid_2[3503:3496]) ? 1 : 0;
assign detect_max[435][17] = (mid_1[3495:3488] > btm_0[3487:3480]) ? 1 : 0;
assign detect_max[435][18] = (mid_1[3495:3488] > btm_0[3495:3488]) ? 1 : 0;
assign detect_max[435][19] = (mid_1[3495:3488] > btm_0[3503:3496]) ? 1 : 0;
assign detect_max[435][20] = (mid_1[3495:3488] > btm_1[3487:3480]) ? 1 : 0;
assign detect_max[435][21] = (mid_1[3495:3488] > btm_1[3495:3488]) ? 1 : 0;
assign detect_max[435][22] = (mid_1[3495:3488] > btm_1[3503:3496]) ? 1 : 0;
assign detect_max[435][23] = (mid_1[3495:3488] > btm_2[3487:3480]) ? 1 : 0;
assign detect_max[435][24] = (mid_1[3495:3488] > btm_2[3495:3488]) ? 1 : 0;
assign detect_max[435][25] = (mid_1[3495:3488] > btm_2[3503:3496]) ? 1 : 0;

assign detect_max[436][0] = (mid_1[3503:3496] > top_0[3495:3488]) ? 1 : 0;
assign detect_max[436][1] = (mid_1[3503:3496] > top_0[3503:3496]) ? 1 : 0;
assign detect_max[436][2] = (mid_1[3503:3496] > top_0[3511:3504]) ? 1 : 0;
assign detect_max[436][3] = (mid_1[3503:3496] > top_1[3495:3488]) ? 1 : 0;
assign detect_max[436][4] = (mid_1[3503:3496] > top_1[3503:3496]) ? 1 : 0;
assign detect_max[436][5] = (mid_1[3503:3496] > top_1[3511:3504]) ? 1 : 0;
assign detect_max[436][6] = (mid_1[3503:3496] > top_2[3495:3488]) ? 1 : 0;
assign detect_max[436][7] = (mid_1[3503:3496] > top_2[3503:3496]) ? 1 : 0;
assign detect_max[436][8] = (mid_1[3503:3496] > top_2[3511:3504]) ? 1 : 0;
assign detect_max[436][9] = (mid_1[3503:3496] > mid_0[3495:3488]) ? 1 : 0;
assign detect_max[436][10] = (mid_1[3503:3496] > mid_0[3503:3496]) ? 1 : 0;
assign detect_max[436][11] = (mid_1[3503:3496] > mid_0[3511:3504]) ? 1 : 0;
assign detect_max[436][12] = (mid_1[3503:3496] > mid_1[3495:3488]) ? 1 : 0;
assign detect_max[436][13] = (mid_1[3503:3496] > mid_1[3511:3504]) ? 1 : 0;
assign detect_max[436][14] = (mid_1[3503:3496] > mid_2[3495:3488]) ? 1 : 0;
assign detect_max[436][15] = (mid_1[3503:3496] > mid_2[3503:3496]) ? 1 : 0;
assign detect_max[436][16] = (mid_1[3503:3496] > mid_2[3511:3504]) ? 1 : 0;
assign detect_max[436][17] = (mid_1[3503:3496] > btm_0[3495:3488]) ? 1 : 0;
assign detect_max[436][18] = (mid_1[3503:3496] > btm_0[3503:3496]) ? 1 : 0;
assign detect_max[436][19] = (mid_1[3503:3496] > btm_0[3511:3504]) ? 1 : 0;
assign detect_max[436][20] = (mid_1[3503:3496] > btm_1[3495:3488]) ? 1 : 0;
assign detect_max[436][21] = (mid_1[3503:3496] > btm_1[3503:3496]) ? 1 : 0;
assign detect_max[436][22] = (mid_1[3503:3496] > btm_1[3511:3504]) ? 1 : 0;
assign detect_max[436][23] = (mid_1[3503:3496] > btm_2[3495:3488]) ? 1 : 0;
assign detect_max[436][24] = (mid_1[3503:3496] > btm_2[3503:3496]) ? 1 : 0;
assign detect_max[436][25] = (mid_1[3503:3496] > btm_2[3511:3504]) ? 1 : 0;

assign detect_max[437][0] = (mid_1[3511:3504] > top_0[3503:3496]) ? 1 : 0;
assign detect_max[437][1] = (mid_1[3511:3504] > top_0[3511:3504]) ? 1 : 0;
assign detect_max[437][2] = (mid_1[3511:3504] > top_0[3519:3512]) ? 1 : 0;
assign detect_max[437][3] = (mid_1[3511:3504] > top_1[3503:3496]) ? 1 : 0;
assign detect_max[437][4] = (mid_1[3511:3504] > top_1[3511:3504]) ? 1 : 0;
assign detect_max[437][5] = (mid_1[3511:3504] > top_1[3519:3512]) ? 1 : 0;
assign detect_max[437][6] = (mid_1[3511:3504] > top_2[3503:3496]) ? 1 : 0;
assign detect_max[437][7] = (mid_1[3511:3504] > top_2[3511:3504]) ? 1 : 0;
assign detect_max[437][8] = (mid_1[3511:3504] > top_2[3519:3512]) ? 1 : 0;
assign detect_max[437][9] = (mid_1[3511:3504] > mid_0[3503:3496]) ? 1 : 0;
assign detect_max[437][10] = (mid_1[3511:3504] > mid_0[3511:3504]) ? 1 : 0;
assign detect_max[437][11] = (mid_1[3511:3504] > mid_0[3519:3512]) ? 1 : 0;
assign detect_max[437][12] = (mid_1[3511:3504] > mid_1[3503:3496]) ? 1 : 0;
assign detect_max[437][13] = (mid_1[3511:3504] > mid_1[3519:3512]) ? 1 : 0;
assign detect_max[437][14] = (mid_1[3511:3504] > mid_2[3503:3496]) ? 1 : 0;
assign detect_max[437][15] = (mid_1[3511:3504] > mid_2[3511:3504]) ? 1 : 0;
assign detect_max[437][16] = (mid_1[3511:3504] > mid_2[3519:3512]) ? 1 : 0;
assign detect_max[437][17] = (mid_1[3511:3504] > btm_0[3503:3496]) ? 1 : 0;
assign detect_max[437][18] = (mid_1[3511:3504] > btm_0[3511:3504]) ? 1 : 0;
assign detect_max[437][19] = (mid_1[3511:3504] > btm_0[3519:3512]) ? 1 : 0;
assign detect_max[437][20] = (mid_1[3511:3504] > btm_1[3503:3496]) ? 1 : 0;
assign detect_max[437][21] = (mid_1[3511:3504] > btm_1[3511:3504]) ? 1 : 0;
assign detect_max[437][22] = (mid_1[3511:3504] > btm_1[3519:3512]) ? 1 : 0;
assign detect_max[437][23] = (mid_1[3511:3504] > btm_2[3503:3496]) ? 1 : 0;
assign detect_max[437][24] = (mid_1[3511:3504] > btm_2[3511:3504]) ? 1 : 0;
assign detect_max[437][25] = (mid_1[3511:3504] > btm_2[3519:3512]) ? 1 : 0;

assign detect_max[438][0] = (mid_1[3519:3512] > top_0[3511:3504]) ? 1 : 0;
assign detect_max[438][1] = (mid_1[3519:3512] > top_0[3519:3512]) ? 1 : 0;
assign detect_max[438][2] = (mid_1[3519:3512] > top_0[3527:3520]) ? 1 : 0;
assign detect_max[438][3] = (mid_1[3519:3512] > top_1[3511:3504]) ? 1 : 0;
assign detect_max[438][4] = (mid_1[3519:3512] > top_1[3519:3512]) ? 1 : 0;
assign detect_max[438][5] = (mid_1[3519:3512] > top_1[3527:3520]) ? 1 : 0;
assign detect_max[438][6] = (mid_1[3519:3512] > top_2[3511:3504]) ? 1 : 0;
assign detect_max[438][7] = (mid_1[3519:3512] > top_2[3519:3512]) ? 1 : 0;
assign detect_max[438][8] = (mid_1[3519:3512] > top_2[3527:3520]) ? 1 : 0;
assign detect_max[438][9] = (mid_1[3519:3512] > mid_0[3511:3504]) ? 1 : 0;
assign detect_max[438][10] = (mid_1[3519:3512] > mid_0[3519:3512]) ? 1 : 0;
assign detect_max[438][11] = (mid_1[3519:3512] > mid_0[3527:3520]) ? 1 : 0;
assign detect_max[438][12] = (mid_1[3519:3512] > mid_1[3511:3504]) ? 1 : 0;
assign detect_max[438][13] = (mid_1[3519:3512] > mid_1[3527:3520]) ? 1 : 0;
assign detect_max[438][14] = (mid_1[3519:3512] > mid_2[3511:3504]) ? 1 : 0;
assign detect_max[438][15] = (mid_1[3519:3512] > mid_2[3519:3512]) ? 1 : 0;
assign detect_max[438][16] = (mid_1[3519:3512] > mid_2[3527:3520]) ? 1 : 0;
assign detect_max[438][17] = (mid_1[3519:3512] > btm_0[3511:3504]) ? 1 : 0;
assign detect_max[438][18] = (mid_1[3519:3512] > btm_0[3519:3512]) ? 1 : 0;
assign detect_max[438][19] = (mid_1[3519:3512] > btm_0[3527:3520]) ? 1 : 0;
assign detect_max[438][20] = (mid_1[3519:3512] > btm_1[3511:3504]) ? 1 : 0;
assign detect_max[438][21] = (mid_1[3519:3512] > btm_1[3519:3512]) ? 1 : 0;
assign detect_max[438][22] = (mid_1[3519:3512] > btm_1[3527:3520]) ? 1 : 0;
assign detect_max[438][23] = (mid_1[3519:3512] > btm_2[3511:3504]) ? 1 : 0;
assign detect_max[438][24] = (mid_1[3519:3512] > btm_2[3519:3512]) ? 1 : 0;
assign detect_max[438][25] = (mid_1[3519:3512] > btm_2[3527:3520]) ? 1 : 0;

assign detect_max[439][0] = (mid_1[3527:3520] > top_0[3519:3512]) ? 1 : 0;
assign detect_max[439][1] = (mid_1[3527:3520] > top_0[3527:3520]) ? 1 : 0;
assign detect_max[439][2] = (mid_1[3527:3520] > top_0[3535:3528]) ? 1 : 0;
assign detect_max[439][3] = (mid_1[3527:3520] > top_1[3519:3512]) ? 1 : 0;
assign detect_max[439][4] = (mid_1[3527:3520] > top_1[3527:3520]) ? 1 : 0;
assign detect_max[439][5] = (mid_1[3527:3520] > top_1[3535:3528]) ? 1 : 0;
assign detect_max[439][6] = (mid_1[3527:3520] > top_2[3519:3512]) ? 1 : 0;
assign detect_max[439][7] = (mid_1[3527:3520] > top_2[3527:3520]) ? 1 : 0;
assign detect_max[439][8] = (mid_1[3527:3520] > top_2[3535:3528]) ? 1 : 0;
assign detect_max[439][9] = (mid_1[3527:3520] > mid_0[3519:3512]) ? 1 : 0;
assign detect_max[439][10] = (mid_1[3527:3520] > mid_0[3527:3520]) ? 1 : 0;
assign detect_max[439][11] = (mid_1[3527:3520] > mid_0[3535:3528]) ? 1 : 0;
assign detect_max[439][12] = (mid_1[3527:3520] > mid_1[3519:3512]) ? 1 : 0;
assign detect_max[439][13] = (mid_1[3527:3520] > mid_1[3535:3528]) ? 1 : 0;
assign detect_max[439][14] = (mid_1[3527:3520] > mid_2[3519:3512]) ? 1 : 0;
assign detect_max[439][15] = (mid_1[3527:3520] > mid_2[3527:3520]) ? 1 : 0;
assign detect_max[439][16] = (mid_1[3527:3520] > mid_2[3535:3528]) ? 1 : 0;
assign detect_max[439][17] = (mid_1[3527:3520] > btm_0[3519:3512]) ? 1 : 0;
assign detect_max[439][18] = (mid_1[3527:3520] > btm_0[3527:3520]) ? 1 : 0;
assign detect_max[439][19] = (mid_1[3527:3520] > btm_0[3535:3528]) ? 1 : 0;
assign detect_max[439][20] = (mid_1[3527:3520] > btm_1[3519:3512]) ? 1 : 0;
assign detect_max[439][21] = (mid_1[3527:3520] > btm_1[3527:3520]) ? 1 : 0;
assign detect_max[439][22] = (mid_1[3527:3520] > btm_1[3535:3528]) ? 1 : 0;
assign detect_max[439][23] = (mid_1[3527:3520] > btm_2[3519:3512]) ? 1 : 0;
assign detect_max[439][24] = (mid_1[3527:3520] > btm_2[3527:3520]) ? 1 : 0;
assign detect_max[439][25] = (mid_1[3527:3520] > btm_2[3535:3528]) ? 1 : 0;

assign detect_max[440][0] = (mid_1[3535:3528] > top_0[3527:3520]) ? 1 : 0;
assign detect_max[440][1] = (mid_1[3535:3528] > top_0[3535:3528]) ? 1 : 0;
assign detect_max[440][2] = (mid_1[3535:3528] > top_0[3543:3536]) ? 1 : 0;
assign detect_max[440][3] = (mid_1[3535:3528] > top_1[3527:3520]) ? 1 : 0;
assign detect_max[440][4] = (mid_1[3535:3528] > top_1[3535:3528]) ? 1 : 0;
assign detect_max[440][5] = (mid_1[3535:3528] > top_1[3543:3536]) ? 1 : 0;
assign detect_max[440][6] = (mid_1[3535:3528] > top_2[3527:3520]) ? 1 : 0;
assign detect_max[440][7] = (mid_1[3535:3528] > top_2[3535:3528]) ? 1 : 0;
assign detect_max[440][8] = (mid_1[3535:3528] > top_2[3543:3536]) ? 1 : 0;
assign detect_max[440][9] = (mid_1[3535:3528] > mid_0[3527:3520]) ? 1 : 0;
assign detect_max[440][10] = (mid_1[3535:3528] > mid_0[3535:3528]) ? 1 : 0;
assign detect_max[440][11] = (mid_1[3535:3528] > mid_0[3543:3536]) ? 1 : 0;
assign detect_max[440][12] = (mid_1[3535:3528] > mid_1[3527:3520]) ? 1 : 0;
assign detect_max[440][13] = (mid_1[3535:3528] > mid_1[3543:3536]) ? 1 : 0;
assign detect_max[440][14] = (mid_1[3535:3528] > mid_2[3527:3520]) ? 1 : 0;
assign detect_max[440][15] = (mid_1[3535:3528] > mid_2[3535:3528]) ? 1 : 0;
assign detect_max[440][16] = (mid_1[3535:3528] > mid_2[3543:3536]) ? 1 : 0;
assign detect_max[440][17] = (mid_1[3535:3528] > btm_0[3527:3520]) ? 1 : 0;
assign detect_max[440][18] = (mid_1[3535:3528] > btm_0[3535:3528]) ? 1 : 0;
assign detect_max[440][19] = (mid_1[3535:3528] > btm_0[3543:3536]) ? 1 : 0;
assign detect_max[440][20] = (mid_1[3535:3528] > btm_1[3527:3520]) ? 1 : 0;
assign detect_max[440][21] = (mid_1[3535:3528] > btm_1[3535:3528]) ? 1 : 0;
assign detect_max[440][22] = (mid_1[3535:3528] > btm_1[3543:3536]) ? 1 : 0;
assign detect_max[440][23] = (mid_1[3535:3528] > btm_2[3527:3520]) ? 1 : 0;
assign detect_max[440][24] = (mid_1[3535:3528] > btm_2[3535:3528]) ? 1 : 0;
assign detect_max[440][25] = (mid_1[3535:3528] > btm_2[3543:3536]) ? 1 : 0;

assign detect_max[441][0] = (mid_1[3543:3536] > top_0[3535:3528]) ? 1 : 0;
assign detect_max[441][1] = (mid_1[3543:3536] > top_0[3543:3536]) ? 1 : 0;
assign detect_max[441][2] = (mid_1[3543:3536] > top_0[3551:3544]) ? 1 : 0;
assign detect_max[441][3] = (mid_1[3543:3536] > top_1[3535:3528]) ? 1 : 0;
assign detect_max[441][4] = (mid_1[3543:3536] > top_1[3543:3536]) ? 1 : 0;
assign detect_max[441][5] = (mid_1[3543:3536] > top_1[3551:3544]) ? 1 : 0;
assign detect_max[441][6] = (mid_1[3543:3536] > top_2[3535:3528]) ? 1 : 0;
assign detect_max[441][7] = (mid_1[3543:3536] > top_2[3543:3536]) ? 1 : 0;
assign detect_max[441][8] = (mid_1[3543:3536] > top_2[3551:3544]) ? 1 : 0;
assign detect_max[441][9] = (mid_1[3543:3536] > mid_0[3535:3528]) ? 1 : 0;
assign detect_max[441][10] = (mid_1[3543:3536] > mid_0[3543:3536]) ? 1 : 0;
assign detect_max[441][11] = (mid_1[3543:3536] > mid_0[3551:3544]) ? 1 : 0;
assign detect_max[441][12] = (mid_1[3543:3536] > mid_1[3535:3528]) ? 1 : 0;
assign detect_max[441][13] = (mid_1[3543:3536] > mid_1[3551:3544]) ? 1 : 0;
assign detect_max[441][14] = (mid_1[3543:3536] > mid_2[3535:3528]) ? 1 : 0;
assign detect_max[441][15] = (mid_1[3543:3536] > mid_2[3543:3536]) ? 1 : 0;
assign detect_max[441][16] = (mid_1[3543:3536] > mid_2[3551:3544]) ? 1 : 0;
assign detect_max[441][17] = (mid_1[3543:3536] > btm_0[3535:3528]) ? 1 : 0;
assign detect_max[441][18] = (mid_1[3543:3536] > btm_0[3543:3536]) ? 1 : 0;
assign detect_max[441][19] = (mid_1[3543:3536] > btm_0[3551:3544]) ? 1 : 0;
assign detect_max[441][20] = (mid_1[3543:3536] > btm_1[3535:3528]) ? 1 : 0;
assign detect_max[441][21] = (mid_1[3543:3536] > btm_1[3543:3536]) ? 1 : 0;
assign detect_max[441][22] = (mid_1[3543:3536] > btm_1[3551:3544]) ? 1 : 0;
assign detect_max[441][23] = (mid_1[3543:3536] > btm_2[3535:3528]) ? 1 : 0;
assign detect_max[441][24] = (mid_1[3543:3536] > btm_2[3543:3536]) ? 1 : 0;
assign detect_max[441][25] = (mid_1[3543:3536] > btm_2[3551:3544]) ? 1 : 0;

assign detect_max[442][0] = (mid_1[3551:3544] > top_0[3543:3536]) ? 1 : 0;
assign detect_max[442][1] = (mid_1[3551:3544] > top_0[3551:3544]) ? 1 : 0;
assign detect_max[442][2] = (mid_1[3551:3544] > top_0[3559:3552]) ? 1 : 0;
assign detect_max[442][3] = (mid_1[3551:3544] > top_1[3543:3536]) ? 1 : 0;
assign detect_max[442][4] = (mid_1[3551:3544] > top_1[3551:3544]) ? 1 : 0;
assign detect_max[442][5] = (mid_1[3551:3544] > top_1[3559:3552]) ? 1 : 0;
assign detect_max[442][6] = (mid_1[3551:3544] > top_2[3543:3536]) ? 1 : 0;
assign detect_max[442][7] = (mid_1[3551:3544] > top_2[3551:3544]) ? 1 : 0;
assign detect_max[442][8] = (mid_1[3551:3544] > top_2[3559:3552]) ? 1 : 0;
assign detect_max[442][9] = (mid_1[3551:3544] > mid_0[3543:3536]) ? 1 : 0;
assign detect_max[442][10] = (mid_1[3551:3544] > mid_0[3551:3544]) ? 1 : 0;
assign detect_max[442][11] = (mid_1[3551:3544] > mid_0[3559:3552]) ? 1 : 0;
assign detect_max[442][12] = (mid_1[3551:3544] > mid_1[3543:3536]) ? 1 : 0;
assign detect_max[442][13] = (mid_1[3551:3544] > mid_1[3559:3552]) ? 1 : 0;
assign detect_max[442][14] = (mid_1[3551:3544] > mid_2[3543:3536]) ? 1 : 0;
assign detect_max[442][15] = (mid_1[3551:3544] > mid_2[3551:3544]) ? 1 : 0;
assign detect_max[442][16] = (mid_1[3551:3544] > mid_2[3559:3552]) ? 1 : 0;
assign detect_max[442][17] = (mid_1[3551:3544] > btm_0[3543:3536]) ? 1 : 0;
assign detect_max[442][18] = (mid_1[3551:3544] > btm_0[3551:3544]) ? 1 : 0;
assign detect_max[442][19] = (mid_1[3551:3544] > btm_0[3559:3552]) ? 1 : 0;
assign detect_max[442][20] = (mid_1[3551:3544] > btm_1[3543:3536]) ? 1 : 0;
assign detect_max[442][21] = (mid_1[3551:3544] > btm_1[3551:3544]) ? 1 : 0;
assign detect_max[442][22] = (mid_1[3551:3544] > btm_1[3559:3552]) ? 1 : 0;
assign detect_max[442][23] = (mid_1[3551:3544] > btm_2[3543:3536]) ? 1 : 0;
assign detect_max[442][24] = (mid_1[3551:3544] > btm_2[3551:3544]) ? 1 : 0;
assign detect_max[442][25] = (mid_1[3551:3544] > btm_2[3559:3552]) ? 1 : 0;

assign detect_max[443][0] = (mid_1[3559:3552] > top_0[3551:3544]) ? 1 : 0;
assign detect_max[443][1] = (mid_1[3559:3552] > top_0[3559:3552]) ? 1 : 0;
assign detect_max[443][2] = (mid_1[3559:3552] > top_0[3567:3560]) ? 1 : 0;
assign detect_max[443][3] = (mid_1[3559:3552] > top_1[3551:3544]) ? 1 : 0;
assign detect_max[443][4] = (mid_1[3559:3552] > top_1[3559:3552]) ? 1 : 0;
assign detect_max[443][5] = (mid_1[3559:3552] > top_1[3567:3560]) ? 1 : 0;
assign detect_max[443][6] = (mid_1[3559:3552] > top_2[3551:3544]) ? 1 : 0;
assign detect_max[443][7] = (mid_1[3559:3552] > top_2[3559:3552]) ? 1 : 0;
assign detect_max[443][8] = (mid_1[3559:3552] > top_2[3567:3560]) ? 1 : 0;
assign detect_max[443][9] = (mid_1[3559:3552] > mid_0[3551:3544]) ? 1 : 0;
assign detect_max[443][10] = (mid_1[3559:3552] > mid_0[3559:3552]) ? 1 : 0;
assign detect_max[443][11] = (mid_1[3559:3552] > mid_0[3567:3560]) ? 1 : 0;
assign detect_max[443][12] = (mid_1[3559:3552] > mid_1[3551:3544]) ? 1 : 0;
assign detect_max[443][13] = (mid_1[3559:3552] > mid_1[3567:3560]) ? 1 : 0;
assign detect_max[443][14] = (mid_1[3559:3552] > mid_2[3551:3544]) ? 1 : 0;
assign detect_max[443][15] = (mid_1[3559:3552] > mid_2[3559:3552]) ? 1 : 0;
assign detect_max[443][16] = (mid_1[3559:3552] > mid_2[3567:3560]) ? 1 : 0;
assign detect_max[443][17] = (mid_1[3559:3552] > btm_0[3551:3544]) ? 1 : 0;
assign detect_max[443][18] = (mid_1[3559:3552] > btm_0[3559:3552]) ? 1 : 0;
assign detect_max[443][19] = (mid_1[3559:3552] > btm_0[3567:3560]) ? 1 : 0;
assign detect_max[443][20] = (mid_1[3559:3552] > btm_1[3551:3544]) ? 1 : 0;
assign detect_max[443][21] = (mid_1[3559:3552] > btm_1[3559:3552]) ? 1 : 0;
assign detect_max[443][22] = (mid_1[3559:3552] > btm_1[3567:3560]) ? 1 : 0;
assign detect_max[443][23] = (mid_1[3559:3552] > btm_2[3551:3544]) ? 1 : 0;
assign detect_max[443][24] = (mid_1[3559:3552] > btm_2[3559:3552]) ? 1 : 0;
assign detect_max[443][25] = (mid_1[3559:3552] > btm_2[3567:3560]) ? 1 : 0;

assign detect_max[444][0] = (mid_1[3567:3560] > top_0[3559:3552]) ? 1 : 0;
assign detect_max[444][1] = (mid_1[3567:3560] > top_0[3567:3560]) ? 1 : 0;
assign detect_max[444][2] = (mid_1[3567:3560] > top_0[3575:3568]) ? 1 : 0;
assign detect_max[444][3] = (mid_1[3567:3560] > top_1[3559:3552]) ? 1 : 0;
assign detect_max[444][4] = (mid_1[3567:3560] > top_1[3567:3560]) ? 1 : 0;
assign detect_max[444][5] = (mid_1[3567:3560] > top_1[3575:3568]) ? 1 : 0;
assign detect_max[444][6] = (mid_1[3567:3560] > top_2[3559:3552]) ? 1 : 0;
assign detect_max[444][7] = (mid_1[3567:3560] > top_2[3567:3560]) ? 1 : 0;
assign detect_max[444][8] = (mid_1[3567:3560] > top_2[3575:3568]) ? 1 : 0;
assign detect_max[444][9] = (mid_1[3567:3560] > mid_0[3559:3552]) ? 1 : 0;
assign detect_max[444][10] = (mid_1[3567:3560] > mid_0[3567:3560]) ? 1 : 0;
assign detect_max[444][11] = (mid_1[3567:3560] > mid_0[3575:3568]) ? 1 : 0;
assign detect_max[444][12] = (mid_1[3567:3560] > mid_1[3559:3552]) ? 1 : 0;
assign detect_max[444][13] = (mid_1[3567:3560] > mid_1[3575:3568]) ? 1 : 0;
assign detect_max[444][14] = (mid_1[3567:3560] > mid_2[3559:3552]) ? 1 : 0;
assign detect_max[444][15] = (mid_1[3567:3560] > mid_2[3567:3560]) ? 1 : 0;
assign detect_max[444][16] = (mid_1[3567:3560] > mid_2[3575:3568]) ? 1 : 0;
assign detect_max[444][17] = (mid_1[3567:3560] > btm_0[3559:3552]) ? 1 : 0;
assign detect_max[444][18] = (mid_1[3567:3560] > btm_0[3567:3560]) ? 1 : 0;
assign detect_max[444][19] = (mid_1[3567:3560] > btm_0[3575:3568]) ? 1 : 0;
assign detect_max[444][20] = (mid_1[3567:3560] > btm_1[3559:3552]) ? 1 : 0;
assign detect_max[444][21] = (mid_1[3567:3560] > btm_1[3567:3560]) ? 1 : 0;
assign detect_max[444][22] = (mid_1[3567:3560] > btm_1[3575:3568]) ? 1 : 0;
assign detect_max[444][23] = (mid_1[3567:3560] > btm_2[3559:3552]) ? 1 : 0;
assign detect_max[444][24] = (mid_1[3567:3560] > btm_2[3567:3560]) ? 1 : 0;
assign detect_max[444][25] = (mid_1[3567:3560] > btm_2[3575:3568]) ? 1 : 0;

assign detect_max[445][0] = (mid_1[3575:3568] > top_0[3567:3560]) ? 1 : 0;
assign detect_max[445][1] = (mid_1[3575:3568] > top_0[3575:3568]) ? 1 : 0;
assign detect_max[445][2] = (mid_1[3575:3568] > top_0[3583:3576]) ? 1 : 0;
assign detect_max[445][3] = (mid_1[3575:3568] > top_1[3567:3560]) ? 1 : 0;
assign detect_max[445][4] = (mid_1[3575:3568] > top_1[3575:3568]) ? 1 : 0;
assign detect_max[445][5] = (mid_1[3575:3568] > top_1[3583:3576]) ? 1 : 0;
assign detect_max[445][6] = (mid_1[3575:3568] > top_2[3567:3560]) ? 1 : 0;
assign detect_max[445][7] = (mid_1[3575:3568] > top_2[3575:3568]) ? 1 : 0;
assign detect_max[445][8] = (mid_1[3575:3568] > top_2[3583:3576]) ? 1 : 0;
assign detect_max[445][9] = (mid_1[3575:3568] > mid_0[3567:3560]) ? 1 : 0;
assign detect_max[445][10] = (mid_1[3575:3568] > mid_0[3575:3568]) ? 1 : 0;
assign detect_max[445][11] = (mid_1[3575:3568] > mid_0[3583:3576]) ? 1 : 0;
assign detect_max[445][12] = (mid_1[3575:3568] > mid_1[3567:3560]) ? 1 : 0;
assign detect_max[445][13] = (mid_1[3575:3568] > mid_1[3583:3576]) ? 1 : 0;
assign detect_max[445][14] = (mid_1[3575:3568] > mid_2[3567:3560]) ? 1 : 0;
assign detect_max[445][15] = (mid_1[3575:3568] > mid_2[3575:3568]) ? 1 : 0;
assign detect_max[445][16] = (mid_1[3575:3568] > mid_2[3583:3576]) ? 1 : 0;
assign detect_max[445][17] = (mid_1[3575:3568] > btm_0[3567:3560]) ? 1 : 0;
assign detect_max[445][18] = (mid_1[3575:3568] > btm_0[3575:3568]) ? 1 : 0;
assign detect_max[445][19] = (mid_1[3575:3568] > btm_0[3583:3576]) ? 1 : 0;
assign detect_max[445][20] = (mid_1[3575:3568] > btm_1[3567:3560]) ? 1 : 0;
assign detect_max[445][21] = (mid_1[3575:3568] > btm_1[3575:3568]) ? 1 : 0;
assign detect_max[445][22] = (mid_1[3575:3568] > btm_1[3583:3576]) ? 1 : 0;
assign detect_max[445][23] = (mid_1[3575:3568] > btm_2[3567:3560]) ? 1 : 0;
assign detect_max[445][24] = (mid_1[3575:3568] > btm_2[3575:3568]) ? 1 : 0;
assign detect_max[445][25] = (mid_1[3575:3568] > btm_2[3583:3576]) ? 1 : 0;

assign detect_max[446][0] = (mid_1[3583:3576] > top_0[3575:3568]) ? 1 : 0;
assign detect_max[446][1] = (mid_1[3583:3576] > top_0[3583:3576]) ? 1 : 0;
assign detect_max[446][2] = (mid_1[3583:3576] > top_0[3591:3584]) ? 1 : 0;
assign detect_max[446][3] = (mid_1[3583:3576] > top_1[3575:3568]) ? 1 : 0;
assign detect_max[446][4] = (mid_1[3583:3576] > top_1[3583:3576]) ? 1 : 0;
assign detect_max[446][5] = (mid_1[3583:3576] > top_1[3591:3584]) ? 1 : 0;
assign detect_max[446][6] = (mid_1[3583:3576] > top_2[3575:3568]) ? 1 : 0;
assign detect_max[446][7] = (mid_1[3583:3576] > top_2[3583:3576]) ? 1 : 0;
assign detect_max[446][8] = (mid_1[3583:3576] > top_2[3591:3584]) ? 1 : 0;
assign detect_max[446][9] = (mid_1[3583:3576] > mid_0[3575:3568]) ? 1 : 0;
assign detect_max[446][10] = (mid_1[3583:3576] > mid_0[3583:3576]) ? 1 : 0;
assign detect_max[446][11] = (mid_1[3583:3576] > mid_0[3591:3584]) ? 1 : 0;
assign detect_max[446][12] = (mid_1[3583:3576] > mid_1[3575:3568]) ? 1 : 0;
assign detect_max[446][13] = (mid_1[3583:3576] > mid_1[3591:3584]) ? 1 : 0;
assign detect_max[446][14] = (mid_1[3583:3576] > mid_2[3575:3568]) ? 1 : 0;
assign detect_max[446][15] = (mid_1[3583:3576] > mid_2[3583:3576]) ? 1 : 0;
assign detect_max[446][16] = (mid_1[3583:3576] > mid_2[3591:3584]) ? 1 : 0;
assign detect_max[446][17] = (mid_1[3583:3576] > btm_0[3575:3568]) ? 1 : 0;
assign detect_max[446][18] = (mid_1[3583:3576] > btm_0[3583:3576]) ? 1 : 0;
assign detect_max[446][19] = (mid_1[3583:3576] > btm_0[3591:3584]) ? 1 : 0;
assign detect_max[446][20] = (mid_1[3583:3576] > btm_1[3575:3568]) ? 1 : 0;
assign detect_max[446][21] = (mid_1[3583:3576] > btm_1[3583:3576]) ? 1 : 0;
assign detect_max[446][22] = (mid_1[3583:3576] > btm_1[3591:3584]) ? 1 : 0;
assign detect_max[446][23] = (mid_1[3583:3576] > btm_2[3575:3568]) ? 1 : 0;
assign detect_max[446][24] = (mid_1[3583:3576] > btm_2[3583:3576]) ? 1 : 0;
assign detect_max[446][25] = (mid_1[3583:3576] > btm_2[3591:3584]) ? 1 : 0;

assign detect_max[447][0] = (mid_1[3591:3584] > top_0[3583:3576]) ? 1 : 0;
assign detect_max[447][1] = (mid_1[3591:3584] > top_0[3591:3584]) ? 1 : 0;
assign detect_max[447][2] = (mid_1[3591:3584] > top_0[3599:3592]) ? 1 : 0;
assign detect_max[447][3] = (mid_1[3591:3584] > top_1[3583:3576]) ? 1 : 0;
assign detect_max[447][4] = (mid_1[3591:3584] > top_1[3591:3584]) ? 1 : 0;
assign detect_max[447][5] = (mid_1[3591:3584] > top_1[3599:3592]) ? 1 : 0;
assign detect_max[447][6] = (mid_1[3591:3584] > top_2[3583:3576]) ? 1 : 0;
assign detect_max[447][7] = (mid_1[3591:3584] > top_2[3591:3584]) ? 1 : 0;
assign detect_max[447][8] = (mid_1[3591:3584] > top_2[3599:3592]) ? 1 : 0;
assign detect_max[447][9] = (mid_1[3591:3584] > mid_0[3583:3576]) ? 1 : 0;
assign detect_max[447][10] = (mid_1[3591:3584] > mid_0[3591:3584]) ? 1 : 0;
assign detect_max[447][11] = (mid_1[3591:3584] > mid_0[3599:3592]) ? 1 : 0;
assign detect_max[447][12] = (mid_1[3591:3584] > mid_1[3583:3576]) ? 1 : 0;
assign detect_max[447][13] = (mid_1[3591:3584] > mid_1[3599:3592]) ? 1 : 0;
assign detect_max[447][14] = (mid_1[3591:3584] > mid_2[3583:3576]) ? 1 : 0;
assign detect_max[447][15] = (mid_1[3591:3584] > mid_2[3591:3584]) ? 1 : 0;
assign detect_max[447][16] = (mid_1[3591:3584] > mid_2[3599:3592]) ? 1 : 0;
assign detect_max[447][17] = (mid_1[3591:3584] > btm_0[3583:3576]) ? 1 : 0;
assign detect_max[447][18] = (mid_1[3591:3584] > btm_0[3591:3584]) ? 1 : 0;
assign detect_max[447][19] = (mid_1[3591:3584] > btm_0[3599:3592]) ? 1 : 0;
assign detect_max[447][20] = (mid_1[3591:3584] > btm_1[3583:3576]) ? 1 : 0;
assign detect_max[447][21] = (mid_1[3591:3584] > btm_1[3591:3584]) ? 1 : 0;
assign detect_max[447][22] = (mid_1[3591:3584] > btm_1[3599:3592]) ? 1 : 0;
assign detect_max[447][23] = (mid_1[3591:3584] > btm_2[3583:3576]) ? 1 : 0;
assign detect_max[447][24] = (mid_1[3591:3584] > btm_2[3591:3584]) ? 1 : 0;
assign detect_max[447][25] = (mid_1[3591:3584] > btm_2[3599:3592]) ? 1 : 0;

assign detect_max[448][0] = (mid_1[3599:3592] > top_0[3591:3584]) ? 1 : 0;
assign detect_max[448][1] = (mid_1[3599:3592] > top_0[3599:3592]) ? 1 : 0;
assign detect_max[448][2] = (mid_1[3599:3592] > top_0[3607:3600]) ? 1 : 0;
assign detect_max[448][3] = (mid_1[3599:3592] > top_1[3591:3584]) ? 1 : 0;
assign detect_max[448][4] = (mid_1[3599:3592] > top_1[3599:3592]) ? 1 : 0;
assign detect_max[448][5] = (mid_1[3599:3592] > top_1[3607:3600]) ? 1 : 0;
assign detect_max[448][6] = (mid_1[3599:3592] > top_2[3591:3584]) ? 1 : 0;
assign detect_max[448][7] = (mid_1[3599:3592] > top_2[3599:3592]) ? 1 : 0;
assign detect_max[448][8] = (mid_1[3599:3592] > top_2[3607:3600]) ? 1 : 0;
assign detect_max[448][9] = (mid_1[3599:3592] > mid_0[3591:3584]) ? 1 : 0;
assign detect_max[448][10] = (mid_1[3599:3592] > mid_0[3599:3592]) ? 1 : 0;
assign detect_max[448][11] = (mid_1[3599:3592] > mid_0[3607:3600]) ? 1 : 0;
assign detect_max[448][12] = (mid_1[3599:3592] > mid_1[3591:3584]) ? 1 : 0;
assign detect_max[448][13] = (mid_1[3599:3592] > mid_1[3607:3600]) ? 1 : 0;
assign detect_max[448][14] = (mid_1[3599:3592] > mid_2[3591:3584]) ? 1 : 0;
assign detect_max[448][15] = (mid_1[3599:3592] > mid_2[3599:3592]) ? 1 : 0;
assign detect_max[448][16] = (mid_1[3599:3592] > mid_2[3607:3600]) ? 1 : 0;
assign detect_max[448][17] = (mid_1[3599:3592] > btm_0[3591:3584]) ? 1 : 0;
assign detect_max[448][18] = (mid_1[3599:3592] > btm_0[3599:3592]) ? 1 : 0;
assign detect_max[448][19] = (mid_1[3599:3592] > btm_0[3607:3600]) ? 1 : 0;
assign detect_max[448][20] = (mid_1[3599:3592] > btm_1[3591:3584]) ? 1 : 0;
assign detect_max[448][21] = (mid_1[3599:3592] > btm_1[3599:3592]) ? 1 : 0;
assign detect_max[448][22] = (mid_1[3599:3592] > btm_1[3607:3600]) ? 1 : 0;
assign detect_max[448][23] = (mid_1[3599:3592] > btm_2[3591:3584]) ? 1 : 0;
assign detect_max[448][24] = (mid_1[3599:3592] > btm_2[3599:3592]) ? 1 : 0;
assign detect_max[448][25] = (mid_1[3599:3592] > btm_2[3607:3600]) ? 1 : 0;

assign detect_max[449][0] = (mid_1[3607:3600] > top_0[3599:3592]) ? 1 : 0;
assign detect_max[449][1] = (mid_1[3607:3600] > top_0[3607:3600]) ? 1 : 0;
assign detect_max[449][2] = (mid_1[3607:3600] > top_0[3615:3608]) ? 1 : 0;
assign detect_max[449][3] = (mid_1[3607:3600] > top_1[3599:3592]) ? 1 : 0;
assign detect_max[449][4] = (mid_1[3607:3600] > top_1[3607:3600]) ? 1 : 0;
assign detect_max[449][5] = (mid_1[3607:3600] > top_1[3615:3608]) ? 1 : 0;
assign detect_max[449][6] = (mid_1[3607:3600] > top_2[3599:3592]) ? 1 : 0;
assign detect_max[449][7] = (mid_1[3607:3600] > top_2[3607:3600]) ? 1 : 0;
assign detect_max[449][8] = (mid_1[3607:3600] > top_2[3615:3608]) ? 1 : 0;
assign detect_max[449][9] = (mid_1[3607:3600] > mid_0[3599:3592]) ? 1 : 0;
assign detect_max[449][10] = (mid_1[3607:3600] > mid_0[3607:3600]) ? 1 : 0;
assign detect_max[449][11] = (mid_1[3607:3600] > mid_0[3615:3608]) ? 1 : 0;
assign detect_max[449][12] = (mid_1[3607:3600] > mid_1[3599:3592]) ? 1 : 0;
assign detect_max[449][13] = (mid_1[3607:3600] > mid_1[3615:3608]) ? 1 : 0;
assign detect_max[449][14] = (mid_1[3607:3600] > mid_2[3599:3592]) ? 1 : 0;
assign detect_max[449][15] = (mid_1[3607:3600] > mid_2[3607:3600]) ? 1 : 0;
assign detect_max[449][16] = (mid_1[3607:3600] > mid_2[3615:3608]) ? 1 : 0;
assign detect_max[449][17] = (mid_1[3607:3600] > btm_0[3599:3592]) ? 1 : 0;
assign detect_max[449][18] = (mid_1[3607:3600] > btm_0[3607:3600]) ? 1 : 0;
assign detect_max[449][19] = (mid_1[3607:3600] > btm_0[3615:3608]) ? 1 : 0;
assign detect_max[449][20] = (mid_1[3607:3600] > btm_1[3599:3592]) ? 1 : 0;
assign detect_max[449][21] = (mid_1[3607:3600] > btm_1[3607:3600]) ? 1 : 0;
assign detect_max[449][22] = (mid_1[3607:3600] > btm_1[3615:3608]) ? 1 : 0;
assign detect_max[449][23] = (mid_1[3607:3600] > btm_2[3599:3592]) ? 1 : 0;
assign detect_max[449][24] = (mid_1[3607:3600] > btm_2[3607:3600]) ? 1 : 0;
assign detect_max[449][25] = (mid_1[3607:3600] > btm_2[3615:3608]) ? 1 : 0;

assign detect_max[450][0] = (mid_1[3615:3608] > top_0[3607:3600]) ? 1 : 0;
assign detect_max[450][1] = (mid_1[3615:3608] > top_0[3615:3608]) ? 1 : 0;
assign detect_max[450][2] = (mid_1[3615:3608] > top_0[3623:3616]) ? 1 : 0;
assign detect_max[450][3] = (mid_1[3615:3608] > top_1[3607:3600]) ? 1 : 0;
assign detect_max[450][4] = (mid_1[3615:3608] > top_1[3615:3608]) ? 1 : 0;
assign detect_max[450][5] = (mid_1[3615:3608] > top_1[3623:3616]) ? 1 : 0;
assign detect_max[450][6] = (mid_1[3615:3608] > top_2[3607:3600]) ? 1 : 0;
assign detect_max[450][7] = (mid_1[3615:3608] > top_2[3615:3608]) ? 1 : 0;
assign detect_max[450][8] = (mid_1[3615:3608] > top_2[3623:3616]) ? 1 : 0;
assign detect_max[450][9] = (mid_1[3615:3608] > mid_0[3607:3600]) ? 1 : 0;
assign detect_max[450][10] = (mid_1[3615:3608] > mid_0[3615:3608]) ? 1 : 0;
assign detect_max[450][11] = (mid_1[3615:3608] > mid_0[3623:3616]) ? 1 : 0;
assign detect_max[450][12] = (mid_1[3615:3608] > mid_1[3607:3600]) ? 1 : 0;
assign detect_max[450][13] = (mid_1[3615:3608] > mid_1[3623:3616]) ? 1 : 0;
assign detect_max[450][14] = (mid_1[3615:3608] > mid_2[3607:3600]) ? 1 : 0;
assign detect_max[450][15] = (mid_1[3615:3608] > mid_2[3615:3608]) ? 1 : 0;
assign detect_max[450][16] = (mid_1[3615:3608] > mid_2[3623:3616]) ? 1 : 0;
assign detect_max[450][17] = (mid_1[3615:3608] > btm_0[3607:3600]) ? 1 : 0;
assign detect_max[450][18] = (mid_1[3615:3608] > btm_0[3615:3608]) ? 1 : 0;
assign detect_max[450][19] = (mid_1[3615:3608] > btm_0[3623:3616]) ? 1 : 0;
assign detect_max[450][20] = (mid_1[3615:3608] > btm_1[3607:3600]) ? 1 : 0;
assign detect_max[450][21] = (mid_1[3615:3608] > btm_1[3615:3608]) ? 1 : 0;
assign detect_max[450][22] = (mid_1[3615:3608] > btm_1[3623:3616]) ? 1 : 0;
assign detect_max[450][23] = (mid_1[3615:3608] > btm_2[3607:3600]) ? 1 : 0;
assign detect_max[450][24] = (mid_1[3615:3608] > btm_2[3615:3608]) ? 1 : 0;
assign detect_max[450][25] = (mid_1[3615:3608] > btm_2[3623:3616]) ? 1 : 0;

assign detect_max[451][0] = (mid_1[3623:3616] > top_0[3615:3608]) ? 1 : 0;
assign detect_max[451][1] = (mid_1[3623:3616] > top_0[3623:3616]) ? 1 : 0;
assign detect_max[451][2] = (mid_1[3623:3616] > top_0[3631:3624]) ? 1 : 0;
assign detect_max[451][3] = (mid_1[3623:3616] > top_1[3615:3608]) ? 1 : 0;
assign detect_max[451][4] = (mid_1[3623:3616] > top_1[3623:3616]) ? 1 : 0;
assign detect_max[451][5] = (mid_1[3623:3616] > top_1[3631:3624]) ? 1 : 0;
assign detect_max[451][6] = (mid_1[3623:3616] > top_2[3615:3608]) ? 1 : 0;
assign detect_max[451][7] = (mid_1[3623:3616] > top_2[3623:3616]) ? 1 : 0;
assign detect_max[451][8] = (mid_1[3623:3616] > top_2[3631:3624]) ? 1 : 0;
assign detect_max[451][9] = (mid_1[3623:3616] > mid_0[3615:3608]) ? 1 : 0;
assign detect_max[451][10] = (mid_1[3623:3616] > mid_0[3623:3616]) ? 1 : 0;
assign detect_max[451][11] = (mid_1[3623:3616] > mid_0[3631:3624]) ? 1 : 0;
assign detect_max[451][12] = (mid_1[3623:3616] > mid_1[3615:3608]) ? 1 : 0;
assign detect_max[451][13] = (mid_1[3623:3616] > mid_1[3631:3624]) ? 1 : 0;
assign detect_max[451][14] = (mid_1[3623:3616] > mid_2[3615:3608]) ? 1 : 0;
assign detect_max[451][15] = (mid_1[3623:3616] > mid_2[3623:3616]) ? 1 : 0;
assign detect_max[451][16] = (mid_1[3623:3616] > mid_2[3631:3624]) ? 1 : 0;
assign detect_max[451][17] = (mid_1[3623:3616] > btm_0[3615:3608]) ? 1 : 0;
assign detect_max[451][18] = (mid_1[3623:3616] > btm_0[3623:3616]) ? 1 : 0;
assign detect_max[451][19] = (mid_1[3623:3616] > btm_0[3631:3624]) ? 1 : 0;
assign detect_max[451][20] = (mid_1[3623:3616] > btm_1[3615:3608]) ? 1 : 0;
assign detect_max[451][21] = (mid_1[3623:3616] > btm_1[3623:3616]) ? 1 : 0;
assign detect_max[451][22] = (mid_1[3623:3616] > btm_1[3631:3624]) ? 1 : 0;
assign detect_max[451][23] = (mid_1[3623:3616] > btm_2[3615:3608]) ? 1 : 0;
assign detect_max[451][24] = (mid_1[3623:3616] > btm_2[3623:3616]) ? 1 : 0;
assign detect_max[451][25] = (mid_1[3623:3616] > btm_2[3631:3624]) ? 1 : 0;

assign detect_max[452][0] = (mid_1[3631:3624] > top_0[3623:3616]) ? 1 : 0;
assign detect_max[452][1] = (mid_1[3631:3624] > top_0[3631:3624]) ? 1 : 0;
assign detect_max[452][2] = (mid_1[3631:3624] > top_0[3639:3632]) ? 1 : 0;
assign detect_max[452][3] = (mid_1[3631:3624] > top_1[3623:3616]) ? 1 : 0;
assign detect_max[452][4] = (mid_1[3631:3624] > top_1[3631:3624]) ? 1 : 0;
assign detect_max[452][5] = (mid_1[3631:3624] > top_1[3639:3632]) ? 1 : 0;
assign detect_max[452][6] = (mid_1[3631:3624] > top_2[3623:3616]) ? 1 : 0;
assign detect_max[452][7] = (mid_1[3631:3624] > top_2[3631:3624]) ? 1 : 0;
assign detect_max[452][8] = (mid_1[3631:3624] > top_2[3639:3632]) ? 1 : 0;
assign detect_max[452][9] = (mid_1[3631:3624] > mid_0[3623:3616]) ? 1 : 0;
assign detect_max[452][10] = (mid_1[3631:3624] > mid_0[3631:3624]) ? 1 : 0;
assign detect_max[452][11] = (mid_1[3631:3624] > mid_0[3639:3632]) ? 1 : 0;
assign detect_max[452][12] = (mid_1[3631:3624] > mid_1[3623:3616]) ? 1 : 0;
assign detect_max[452][13] = (mid_1[3631:3624] > mid_1[3639:3632]) ? 1 : 0;
assign detect_max[452][14] = (mid_1[3631:3624] > mid_2[3623:3616]) ? 1 : 0;
assign detect_max[452][15] = (mid_1[3631:3624] > mid_2[3631:3624]) ? 1 : 0;
assign detect_max[452][16] = (mid_1[3631:3624] > mid_2[3639:3632]) ? 1 : 0;
assign detect_max[452][17] = (mid_1[3631:3624] > btm_0[3623:3616]) ? 1 : 0;
assign detect_max[452][18] = (mid_1[3631:3624] > btm_0[3631:3624]) ? 1 : 0;
assign detect_max[452][19] = (mid_1[3631:3624] > btm_0[3639:3632]) ? 1 : 0;
assign detect_max[452][20] = (mid_1[3631:3624] > btm_1[3623:3616]) ? 1 : 0;
assign detect_max[452][21] = (mid_1[3631:3624] > btm_1[3631:3624]) ? 1 : 0;
assign detect_max[452][22] = (mid_1[3631:3624] > btm_1[3639:3632]) ? 1 : 0;
assign detect_max[452][23] = (mid_1[3631:3624] > btm_2[3623:3616]) ? 1 : 0;
assign detect_max[452][24] = (mid_1[3631:3624] > btm_2[3631:3624]) ? 1 : 0;
assign detect_max[452][25] = (mid_1[3631:3624] > btm_2[3639:3632]) ? 1 : 0;

assign detect_max[453][0] = (mid_1[3639:3632] > top_0[3631:3624]) ? 1 : 0;
assign detect_max[453][1] = (mid_1[3639:3632] > top_0[3639:3632]) ? 1 : 0;
assign detect_max[453][2] = (mid_1[3639:3632] > top_0[3647:3640]) ? 1 : 0;
assign detect_max[453][3] = (mid_1[3639:3632] > top_1[3631:3624]) ? 1 : 0;
assign detect_max[453][4] = (mid_1[3639:3632] > top_1[3639:3632]) ? 1 : 0;
assign detect_max[453][5] = (mid_1[3639:3632] > top_1[3647:3640]) ? 1 : 0;
assign detect_max[453][6] = (mid_1[3639:3632] > top_2[3631:3624]) ? 1 : 0;
assign detect_max[453][7] = (mid_1[3639:3632] > top_2[3639:3632]) ? 1 : 0;
assign detect_max[453][8] = (mid_1[3639:3632] > top_2[3647:3640]) ? 1 : 0;
assign detect_max[453][9] = (mid_1[3639:3632] > mid_0[3631:3624]) ? 1 : 0;
assign detect_max[453][10] = (mid_1[3639:3632] > mid_0[3639:3632]) ? 1 : 0;
assign detect_max[453][11] = (mid_1[3639:3632] > mid_0[3647:3640]) ? 1 : 0;
assign detect_max[453][12] = (mid_1[3639:3632] > mid_1[3631:3624]) ? 1 : 0;
assign detect_max[453][13] = (mid_1[3639:3632] > mid_1[3647:3640]) ? 1 : 0;
assign detect_max[453][14] = (mid_1[3639:3632] > mid_2[3631:3624]) ? 1 : 0;
assign detect_max[453][15] = (mid_1[3639:3632] > mid_2[3639:3632]) ? 1 : 0;
assign detect_max[453][16] = (mid_1[3639:3632] > mid_2[3647:3640]) ? 1 : 0;
assign detect_max[453][17] = (mid_1[3639:3632] > btm_0[3631:3624]) ? 1 : 0;
assign detect_max[453][18] = (mid_1[3639:3632] > btm_0[3639:3632]) ? 1 : 0;
assign detect_max[453][19] = (mid_1[3639:3632] > btm_0[3647:3640]) ? 1 : 0;
assign detect_max[453][20] = (mid_1[3639:3632] > btm_1[3631:3624]) ? 1 : 0;
assign detect_max[453][21] = (mid_1[3639:3632] > btm_1[3639:3632]) ? 1 : 0;
assign detect_max[453][22] = (mid_1[3639:3632] > btm_1[3647:3640]) ? 1 : 0;
assign detect_max[453][23] = (mid_1[3639:3632] > btm_2[3631:3624]) ? 1 : 0;
assign detect_max[453][24] = (mid_1[3639:3632] > btm_2[3639:3632]) ? 1 : 0;
assign detect_max[453][25] = (mid_1[3639:3632] > btm_2[3647:3640]) ? 1 : 0;

assign detect_max[454][0] = (mid_1[3647:3640] > top_0[3639:3632]) ? 1 : 0;
assign detect_max[454][1] = (mid_1[3647:3640] > top_0[3647:3640]) ? 1 : 0;
assign detect_max[454][2] = (mid_1[3647:3640] > top_0[3655:3648]) ? 1 : 0;
assign detect_max[454][3] = (mid_1[3647:3640] > top_1[3639:3632]) ? 1 : 0;
assign detect_max[454][4] = (mid_1[3647:3640] > top_1[3647:3640]) ? 1 : 0;
assign detect_max[454][5] = (mid_1[3647:3640] > top_1[3655:3648]) ? 1 : 0;
assign detect_max[454][6] = (mid_1[3647:3640] > top_2[3639:3632]) ? 1 : 0;
assign detect_max[454][7] = (mid_1[3647:3640] > top_2[3647:3640]) ? 1 : 0;
assign detect_max[454][8] = (mid_1[3647:3640] > top_2[3655:3648]) ? 1 : 0;
assign detect_max[454][9] = (mid_1[3647:3640] > mid_0[3639:3632]) ? 1 : 0;
assign detect_max[454][10] = (mid_1[3647:3640] > mid_0[3647:3640]) ? 1 : 0;
assign detect_max[454][11] = (mid_1[3647:3640] > mid_0[3655:3648]) ? 1 : 0;
assign detect_max[454][12] = (mid_1[3647:3640] > mid_1[3639:3632]) ? 1 : 0;
assign detect_max[454][13] = (mid_1[3647:3640] > mid_1[3655:3648]) ? 1 : 0;
assign detect_max[454][14] = (mid_1[3647:3640] > mid_2[3639:3632]) ? 1 : 0;
assign detect_max[454][15] = (mid_1[3647:3640] > mid_2[3647:3640]) ? 1 : 0;
assign detect_max[454][16] = (mid_1[3647:3640] > mid_2[3655:3648]) ? 1 : 0;
assign detect_max[454][17] = (mid_1[3647:3640] > btm_0[3639:3632]) ? 1 : 0;
assign detect_max[454][18] = (mid_1[3647:3640] > btm_0[3647:3640]) ? 1 : 0;
assign detect_max[454][19] = (mid_1[3647:3640] > btm_0[3655:3648]) ? 1 : 0;
assign detect_max[454][20] = (mid_1[3647:3640] > btm_1[3639:3632]) ? 1 : 0;
assign detect_max[454][21] = (mid_1[3647:3640] > btm_1[3647:3640]) ? 1 : 0;
assign detect_max[454][22] = (mid_1[3647:3640] > btm_1[3655:3648]) ? 1 : 0;
assign detect_max[454][23] = (mid_1[3647:3640] > btm_2[3639:3632]) ? 1 : 0;
assign detect_max[454][24] = (mid_1[3647:3640] > btm_2[3647:3640]) ? 1 : 0;
assign detect_max[454][25] = (mid_1[3647:3640] > btm_2[3655:3648]) ? 1 : 0;

assign detect_max[455][0] = (mid_1[3655:3648] > top_0[3647:3640]) ? 1 : 0;
assign detect_max[455][1] = (mid_1[3655:3648] > top_0[3655:3648]) ? 1 : 0;
assign detect_max[455][2] = (mid_1[3655:3648] > top_0[3663:3656]) ? 1 : 0;
assign detect_max[455][3] = (mid_1[3655:3648] > top_1[3647:3640]) ? 1 : 0;
assign detect_max[455][4] = (mid_1[3655:3648] > top_1[3655:3648]) ? 1 : 0;
assign detect_max[455][5] = (mid_1[3655:3648] > top_1[3663:3656]) ? 1 : 0;
assign detect_max[455][6] = (mid_1[3655:3648] > top_2[3647:3640]) ? 1 : 0;
assign detect_max[455][7] = (mid_1[3655:3648] > top_2[3655:3648]) ? 1 : 0;
assign detect_max[455][8] = (mid_1[3655:3648] > top_2[3663:3656]) ? 1 : 0;
assign detect_max[455][9] = (mid_1[3655:3648] > mid_0[3647:3640]) ? 1 : 0;
assign detect_max[455][10] = (mid_1[3655:3648] > mid_0[3655:3648]) ? 1 : 0;
assign detect_max[455][11] = (mid_1[3655:3648] > mid_0[3663:3656]) ? 1 : 0;
assign detect_max[455][12] = (mid_1[3655:3648] > mid_1[3647:3640]) ? 1 : 0;
assign detect_max[455][13] = (mid_1[3655:3648] > mid_1[3663:3656]) ? 1 : 0;
assign detect_max[455][14] = (mid_1[3655:3648] > mid_2[3647:3640]) ? 1 : 0;
assign detect_max[455][15] = (mid_1[3655:3648] > mid_2[3655:3648]) ? 1 : 0;
assign detect_max[455][16] = (mid_1[3655:3648] > mid_2[3663:3656]) ? 1 : 0;
assign detect_max[455][17] = (mid_1[3655:3648] > btm_0[3647:3640]) ? 1 : 0;
assign detect_max[455][18] = (mid_1[3655:3648] > btm_0[3655:3648]) ? 1 : 0;
assign detect_max[455][19] = (mid_1[3655:3648] > btm_0[3663:3656]) ? 1 : 0;
assign detect_max[455][20] = (mid_1[3655:3648] > btm_1[3647:3640]) ? 1 : 0;
assign detect_max[455][21] = (mid_1[3655:3648] > btm_1[3655:3648]) ? 1 : 0;
assign detect_max[455][22] = (mid_1[3655:3648] > btm_1[3663:3656]) ? 1 : 0;
assign detect_max[455][23] = (mid_1[3655:3648] > btm_2[3647:3640]) ? 1 : 0;
assign detect_max[455][24] = (mid_1[3655:3648] > btm_2[3655:3648]) ? 1 : 0;
assign detect_max[455][25] = (mid_1[3655:3648] > btm_2[3663:3656]) ? 1 : 0;

assign detect_max[456][0] = (mid_1[3663:3656] > top_0[3655:3648]) ? 1 : 0;
assign detect_max[456][1] = (mid_1[3663:3656] > top_0[3663:3656]) ? 1 : 0;
assign detect_max[456][2] = (mid_1[3663:3656] > top_0[3671:3664]) ? 1 : 0;
assign detect_max[456][3] = (mid_1[3663:3656] > top_1[3655:3648]) ? 1 : 0;
assign detect_max[456][4] = (mid_1[3663:3656] > top_1[3663:3656]) ? 1 : 0;
assign detect_max[456][5] = (mid_1[3663:3656] > top_1[3671:3664]) ? 1 : 0;
assign detect_max[456][6] = (mid_1[3663:3656] > top_2[3655:3648]) ? 1 : 0;
assign detect_max[456][7] = (mid_1[3663:3656] > top_2[3663:3656]) ? 1 : 0;
assign detect_max[456][8] = (mid_1[3663:3656] > top_2[3671:3664]) ? 1 : 0;
assign detect_max[456][9] = (mid_1[3663:3656] > mid_0[3655:3648]) ? 1 : 0;
assign detect_max[456][10] = (mid_1[3663:3656] > mid_0[3663:3656]) ? 1 : 0;
assign detect_max[456][11] = (mid_1[3663:3656] > mid_0[3671:3664]) ? 1 : 0;
assign detect_max[456][12] = (mid_1[3663:3656] > mid_1[3655:3648]) ? 1 : 0;
assign detect_max[456][13] = (mid_1[3663:3656] > mid_1[3671:3664]) ? 1 : 0;
assign detect_max[456][14] = (mid_1[3663:3656] > mid_2[3655:3648]) ? 1 : 0;
assign detect_max[456][15] = (mid_1[3663:3656] > mid_2[3663:3656]) ? 1 : 0;
assign detect_max[456][16] = (mid_1[3663:3656] > mid_2[3671:3664]) ? 1 : 0;
assign detect_max[456][17] = (mid_1[3663:3656] > btm_0[3655:3648]) ? 1 : 0;
assign detect_max[456][18] = (mid_1[3663:3656] > btm_0[3663:3656]) ? 1 : 0;
assign detect_max[456][19] = (mid_1[3663:3656] > btm_0[3671:3664]) ? 1 : 0;
assign detect_max[456][20] = (mid_1[3663:3656] > btm_1[3655:3648]) ? 1 : 0;
assign detect_max[456][21] = (mid_1[3663:3656] > btm_1[3663:3656]) ? 1 : 0;
assign detect_max[456][22] = (mid_1[3663:3656] > btm_1[3671:3664]) ? 1 : 0;
assign detect_max[456][23] = (mid_1[3663:3656] > btm_2[3655:3648]) ? 1 : 0;
assign detect_max[456][24] = (mid_1[3663:3656] > btm_2[3663:3656]) ? 1 : 0;
assign detect_max[456][25] = (mid_1[3663:3656] > btm_2[3671:3664]) ? 1 : 0;

assign detect_max[457][0] = (mid_1[3671:3664] > top_0[3663:3656]) ? 1 : 0;
assign detect_max[457][1] = (mid_1[3671:3664] > top_0[3671:3664]) ? 1 : 0;
assign detect_max[457][2] = (mid_1[3671:3664] > top_0[3679:3672]) ? 1 : 0;
assign detect_max[457][3] = (mid_1[3671:3664] > top_1[3663:3656]) ? 1 : 0;
assign detect_max[457][4] = (mid_1[3671:3664] > top_1[3671:3664]) ? 1 : 0;
assign detect_max[457][5] = (mid_1[3671:3664] > top_1[3679:3672]) ? 1 : 0;
assign detect_max[457][6] = (mid_1[3671:3664] > top_2[3663:3656]) ? 1 : 0;
assign detect_max[457][7] = (mid_1[3671:3664] > top_2[3671:3664]) ? 1 : 0;
assign detect_max[457][8] = (mid_1[3671:3664] > top_2[3679:3672]) ? 1 : 0;
assign detect_max[457][9] = (mid_1[3671:3664] > mid_0[3663:3656]) ? 1 : 0;
assign detect_max[457][10] = (mid_1[3671:3664] > mid_0[3671:3664]) ? 1 : 0;
assign detect_max[457][11] = (mid_1[3671:3664] > mid_0[3679:3672]) ? 1 : 0;
assign detect_max[457][12] = (mid_1[3671:3664] > mid_1[3663:3656]) ? 1 : 0;
assign detect_max[457][13] = (mid_1[3671:3664] > mid_1[3679:3672]) ? 1 : 0;
assign detect_max[457][14] = (mid_1[3671:3664] > mid_2[3663:3656]) ? 1 : 0;
assign detect_max[457][15] = (mid_1[3671:3664] > mid_2[3671:3664]) ? 1 : 0;
assign detect_max[457][16] = (mid_1[3671:3664] > mid_2[3679:3672]) ? 1 : 0;
assign detect_max[457][17] = (mid_1[3671:3664] > btm_0[3663:3656]) ? 1 : 0;
assign detect_max[457][18] = (mid_1[3671:3664] > btm_0[3671:3664]) ? 1 : 0;
assign detect_max[457][19] = (mid_1[3671:3664] > btm_0[3679:3672]) ? 1 : 0;
assign detect_max[457][20] = (mid_1[3671:3664] > btm_1[3663:3656]) ? 1 : 0;
assign detect_max[457][21] = (mid_1[3671:3664] > btm_1[3671:3664]) ? 1 : 0;
assign detect_max[457][22] = (mid_1[3671:3664] > btm_1[3679:3672]) ? 1 : 0;
assign detect_max[457][23] = (mid_1[3671:3664] > btm_2[3663:3656]) ? 1 : 0;
assign detect_max[457][24] = (mid_1[3671:3664] > btm_2[3671:3664]) ? 1 : 0;
assign detect_max[457][25] = (mid_1[3671:3664] > btm_2[3679:3672]) ? 1 : 0;

assign detect_max[458][0] = (mid_1[3679:3672] > top_0[3671:3664]) ? 1 : 0;
assign detect_max[458][1] = (mid_1[3679:3672] > top_0[3679:3672]) ? 1 : 0;
assign detect_max[458][2] = (mid_1[3679:3672] > top_0[3687:3680]) ? 1 : 0;
assign detect_max[458][3] = (mid_1[3679:3672] > top_1[3671:3664]) ? 1 : 0;
assign detect_max[458][4] = (mid_1[3679:3672] > top_1[3679:3672]) ? 1 : 0;
assign detect_max[458][5] = (mid_1[3679:3672] > top_1[3687:3680]) ? 1 : 0;
assign detect_max[458][6] = (mid_1[3679:3672] > top_2[3671:3664]) ? 1 : 0;
assign detect_max[458][7] = (mid_1[3679:3672] > top_2[3679:3672]) ? 1 : 0;
assign detect_max[458][8] = (mid_1[3679:3672] > top_2[3687:3680]) ? 1 : 0;
assign detect_max[458][9] = (mid_1[3679:3672] > mid_0[3671:3664]) ? 1 : 0;
assign detect_max[458][10] = (mid_1[3679:3672] > mid_0[3679:3672]) ? 1 : 0;
assign detect_max[458][11] = (mid_1[3679:3672] > mid_0[3687:3680]) ? 1 : 0;
assign detect_max[458][12] = (mid_1[3679:3672] > mid_1[3671:3664]) ? 1 : 0;
assign detect_max[458][13] = (mid_1[3679:3672] > mid_1[3687:3680]) ? 1 : 0;
assign detect_max[458][14] = (mid_1[3679:3672] > mid_2[3671:3664]) ? 1 : 0;
assign detect_max[458][15] = (mid_1[3679:3672] > mid_2[3679:3672]) ? 1 : 0;
assign detect_max[458][16] = (mid_1[3679:3672] > mid_2[3687:3680]) ? 1 : 0;
assign detect_max[458][17] = (mid_1[3679:3672] > btm_0[3671:3664]) ? 1 : 0;
assign detect_max[458][18] = (mid_1[3679:3672] > btm_0[3679:3672]) ? 1 : 0;
assign detect_max[458][19] = (mid_1[3679:3672] > btm_0[3687:3680]) ? 1 : 0;
assign detect_max[458][20] = (mid_1[3679:3672] > btm_1[3671:3664]) ? 1 : 0;
assign detect_max[458][21] = (mid_1[3679:3672] > btm_1[3679:3672]) ? 1 : 0;
assign detect_max[458][22] = (mid_1[3679:3672] > btm_1[3687:3680]) ? 1 : 0;
assign detect_max[458][23] = (mid_1[3679:3672] > btm_2[3671:3664]) ? 1 : 0;
assign detect_max[458][24] = (mid_1[3679:3672] > btm_2[3679:3672]) ? 1 : 0;
assign detect_max[458][25] = (mid_1[3679:3672] > btm_2[3687:3680]) ? 1 : 0;

assign detect_max[459][0] = (mid_1[3687:3680] > top_0[3679:3672]) ? 1 : 0;
assign detect_max[459][1] = (mid_1[3687:3680] > top_0[3687:3680]) ? 1 : 0;
assign detect_max[459][2] = (mid_1[3687:3680] > top_0[3695:3688]) ? 1 : 0;
assign detect_max[459][3] = (mid_1[3687:3680] > top_1[3679:3672]) ? 1 : 0;
assign detect_max[459][4] = (mid_1[3687:3680] > top_1[3687:3680]) ? 1 : 0;
assign detect_max[459][5] = (mid_1[3687:3680] > top_1[3695:3688]) ? 1 : 0;
assign detect_max[459][6] = (mid_1[3687:3680] > top_2[3679:3672]) ? 1 : 0;
assign detect_max[459][7] = (mid_1[3687:3680] > top_2[3687:3680]) ? 1 : 0;
assign detect_max[459][8] = (mid_1[3687:3680] > top_2[3695:3688]) ? 1 : 0;
assign detect_max[459][9] = (mid_1[3687:3680] > mid_0[3679:3672]) ? 1 : 0;
assign detect_max[459][10] = (mid_1[3687:3680] > mid_0[3687:3680]) ? 1 : 0;
assign detect_max[459][11] = (mid_1[3687:3680] > mid_0[3695:3688]) ? 1 : 0;
assign detect_max[459][12] = (mid_1[3687:3680] > mid_1[3679:3672]) ? 1 : 0;
assign detect_max[459][13] = (mid_1[3687:3680] > mid_1[3695:3688]) ? 1 : 0;
assign detect_max[459][14] = (mid_1[3687:3680] > mid_2[3679:3672]) ? 1 : 0;
assign detect_max[459][15] = (mid_1[3687:3680] > mid_2[3687:3680]) ? 1 : 0;
assign detect_max[459][16] = (mid_1[3687:3680] > mid_2[3695:3688]) ? 1 : 0;
assign detect_max[459][17] = (mid_1[3687:3680] > btm_0[3679:3672]) ? 1 : 0;
assign detect_max[459][18] = (mid_1[3687:3680] > btm_0[3687:3680]) ? 1 : 0;
assign detect_max[459][19] = (mid_1[3687:3680] > btm_0[3695:3688]) ? 1 : 0;
assign detect_max[459][20] = (mid_1[3687:3680] > btm_1[3679:3672]) ? 1 : 0;
assign detect_max[459][21] = (mid_1[3687:3680] > btm_1[3687:3680]) ? 1 : 0;
assign detect_max[459][22] = (mid_1[3687:3680] > btm_1[3695:3688]) ? 1 : 0;
assign detect_max[459][23] = (mid_1[3687:3680] > btm_2[3679:3672]) ? 1 : 0;
assign detect_max[459][24] = (mid_1[3687:3680] > btm_2[3687:3680]) ? 1 : 0;
assign detect_max[459][25] = (mid_1[3687:3680] > btm_2[3695:3688]) ? 1 : 0;

assign detect_max[460][0] = (mid_1[3695:3688] > top_0[3687:3680]) ? 1 : 0;
assign detect_max[460][1] = (mid_1[3695:3688] > top_0[3695:3688]) ? 1 : 0;
assign detect_max[460][2] = (mid_1[3695:3688] > top_0[3703:3696]) ? 1 : 0;
assign detect_max[460][3] = (mid_1[3695:3688] > top_1[3687:3680]) ? 1 : 0;
assign detect_max[460][4] = (mid_1[3695:3688] > top_1[3695:3688]) ? 1 : 0;
assign detect_max[460][5] = (mid_1[3695:3688] > top_1[3703:3696]) ? 1 : 0;
assign detect_max[460][6] = (mid_1[3695:3688] > top_2[3687:3680]) ? 1 : 0;
assign detect_max[460][7] = (mid_1[3695:3688] > top_2[3695:3688]) ? 1 : 0;
assign detect_max[460][8] = (mid_1[3695:3688] > top_2[3703:3696]) ? 1 : 0;
assign detect_max[460][9] = (mid_1[3695:3688] > mid_0[3687:3680]) ? 1 : 0;
assign detect_max[460][10] = (mid_1[3695:3688] > mid_0[3695:3688]) ? 1 : 0;
assign detect_max[460][11] = (mid_1[3695:3688] > mid_0[3703:3696]) ? 1 : 0;
assign detect_max[460][12] = (mid_1[3695:3688] > mid_1[3687:3680]) ? 1 : 0;
assign detect_max[460][13] = (mid_1[3695:3688] > mid_1[3703:3696]) ? 1 : 0;
assign detect_max[460][14] = (mid_1[3695:3688] > mid_2[3687:3680]) ? 1 : 0;
assign detect_max[460][15] = (mid_1[3695:3688] > mid_2[3695:3688]) ? 1 : 0;
assign detect_max[460][16] = (mid_1[3695:3688] > mid_2[3703:3696]) ? 1 : 0;
assign detect_max[460][17] = (mid_1[3695:3688] > btm_0[3687:3680]) ? 1 : 0;
assign detect_max[460][18] = (mid_1[3695:3688] > btm_0[3695:3688]) ? 1 : 0;
assign detect_max[460][19] = (mid_1[3695:3688] > btm_0[3703:3696]) ? 1 : 0;
assign detect_max[460][20] = (mid_1[3695:3688] > btm_1[3687:3680]) ? 1 : 0;
assign detect_max[460][21] = (mid_1[3695:3688] > btm_1[3695:3688]) ? 1 : 0;
assign detect_max[460][22] = (mid_1[3695:3688] > btm_1[3703:3696]) ? 1 : 0;
assign detect_max[460][23] = (mid_1[3695:3688] > btm_2[3687:3680]) ? 1 : 0;
assign detect_max[460][24] = (mid_1[3695:3688] > btm_2[3695:3688]) ? 1 : 0;
assign detect_max[460][25] = (mid_1[3695:3688] > btm_2[3703:3696]) ? 1 : 0;

assign detect_max[461][0] = (mid_1[3703:3696] > top_0[3695:3688]) ? 1 : 0;
assign detect_max[461][1] = (mid_1[3703:3696] > top_0[3703:3696]) ? 1 : 0;
assign detect_max[461][2] = (mid_1[3703:3696] > top_0[3711:3704]) ? 1 : 0;
assign detect_max[461][3] = (mid_1[3703:3696] > top_1[3695:3688]) ? 1 : 0;
assign detect_max[461][4] = (mid_1[3703:3696] > top_1[3703:3696]) ? 1 : 0;
assign detect_max[461][5] = (mid_1[3703:3696] > top_1[3711:3704]) ? 1 : 0;
assign detect_max[461][6] = (mid_1[3703:3696] > top_2[3695:3688]) ? 1 : 0;
assign detect_max[461][7] = (mid_1[3703:3696] > top_2[3703:3696]) ? 1 : 0;
assign detect_max[461][8] = (mid_1[3703:3696] > top_2[3711:3704]) ? 1 : 0;
assign detect_max[461][9] = (mid_1[3703:3696] > mid_0[3695:3688]) ? 1 : 0;
assign detect_max[461][10] = (mid_1[3703:3696] > mid_0[3703:3696]) ? 1 : 0;
assign detect_max[461][11] = (mid_1[3703:3696] > mid_0[3711:3704]) ? 1 : 0;
assign detect_max[461][12] = (mid_1[3703:3696] > mid_1[3695:3688]) ? 1 : 0;
assign detect_max[461][13] = (mid_1[3703:3696] > mid_1[3711:3704]) ? 1 : 0;
assign detect_max[461][14] = (mid_1[3703:3696] > mid_2[3695:3688]) ? 1 : 0;
assign detect_max[461][15] = (mid_1[3703:3696] > mid_2[3703:3696]) ? 1 : 0;
assign detect_max[461][16] = (mid_1[3703:3696] > mid_2[3711:3704]) ? 1 : 0;
assign detect_max[461][17] = (mid_1[3703:3696] > btm_0[3695:3688]) ? 1 : 0;
assign detect_max[461][18] = (mid_1[3703:3696] > btm_0[3703:3696]) ? 1 : 0;
assign detect_max[461][19] = (mid_1[3703:3696] > btm_0[3711:3704]) ? 1 : 0;
assign detect_max[461][20] = (mid_1[3703:3696] > btm_1[3695:3688]) ? 1 : 0;
assign detect_max[461][21] = (mid_1[3703:3696] > btm_1[3703:3696]) ? 1 : 0;
assign detect_max[461][22] = (mid_1[3703:3696] > btm_1[3711:3704]) ? 1 : 0;
assign detect_max[461][23] = (mid_1[3703:3696] > btm_2[3695:3688]) ? 1 : 0;
assign detect_max[461][24] = (mid_1[3703:3696] > btm_2[3703:3696]) ? 1 : 0;
assign detect_max[461][25] = (mid_1[3703:3696] > btm_2[3711:3704]) ? 1 : 0;

assign detect_max[462][0] = (mid_1[3711:3704] > top_0[3703:3696]) ? 1 : 0;
assign detect_max[462][1] = (mid_1[3711:3704] > top_0[3711:3704]) ? 1 : 0;
assign detect_max[462][2] = (mid_1[3711:3704] > top_0[3719:3712]) ? 1 : 0;
assign detect_max[462][3] = (mid_1[3711:3704] > top_1[3703:3696]) ? 1 : 0;
assign detect_max[462][4] = (mid_1[3711:3704] > top_1[3711:3704]) ? 1 : 0;
assign detect_max[462][5] = (mid_1[3711:3704] > top_1[3719:3712]) ? 1 : 0;
assign detect_max[462][6] = (mid_1[3711:3704] > top_2[3703:3696]) ? 1 : 0;
assign detect_max[462][7] = (mid_1[3711:3704] > top_2[3711:3704]) ? 1 : 0;
assign detect_max[462][8] = (mid_1[3711:3704] > top_2[3719:3712]) ? 1 : 0;
assign detect_max[462][9] = (mid_1[3711:3704] > mid_0[3703:3696]) ? 1 : 0;
assign detect_max[462][10] = (mid_1[3711:3704] > mid_0[3711:3704]) ? 1 : 0;
assign detect_max[462][11] = (mid_1[3711:3704] > mid_0[3719:3712]) ? 1 : 0;
assign detect_max[462][12] = (mid_1[3711:3704] > mid_1[3703:3696]) ? 1 : 0;
assign detect_max[462][13] = (mid_1[3711:3704] > mid_1[3719:3712]) ? 1 : 0;
assign detect_max[462][14] = (mid_1[3711:3704] > mid_2[3703:3696]) ? 1 : 0;
assign detect_max[462][15] = (mid_1[3711:3704] > mid_2[3711:3704]) ? 1 : 0;
assign detect_max[462][16] = (mid_1[3711:3704] > mid_2[3719:3712]) ? 1 : 0;
assign detect_max[462][17] = (mid_1[3711:3704] > btm_0[3703:3696]) ? 1 : 0;
assign detect_max[462][18] = (mid_1[3711:3704] > btm_0[3711:3704]) ? 1 : 0;
assign detect_max[462][19] = (mid_1[3711:3704] > btm_0[3719:3712]) ? 1 : 0;
assign detect_max[462][20] = (mid_1[3711:3704] > btm_1[3703:3696]) ? 1 : 0;
assign detect_max[462][21] = (mid_1[3711:3704] > btm_1[3711:3704]) ? 1 : 0;
assign detect_max[462][22] = (mid_1[3711:3704] > btm_1[3719:3712]) ? 1 : 0;
assign detect_max[462][23] = (mid_1[3711:3704] > btm_2[3703:3696]) ? 1 : 0;
assign detect_max[462][24] = (mid_1[3711:3704] > btm_2[3711:3704]) ? 1 : 0;
assign detect_max[462][25] = (mid_1[3711:3704] > btm_2[3719:3712]) ? 1 : 0;

assign detect_max[463][0] = (mid_1[3719:3712] > top_0[3711:3704]) ? 1 : 0;
assign detect_max[463][1] = (mid_1[3719:3712] > top_0[3719:3712]) ? 1 : 0;
assign detect_max[463][2] = (mid_1[3719:3712] > top_0[3727:3720]) ? 1 : 0;
assign detect_max[463][3] = (mid_1[3719:3712] > top_1[3711:3704]) ? 1 : 0;
assign detect_max[463][4] = (mid_1[3719:3712] > top_1[3719:3712]) ? 1 : 0;
assign detect_max[463][5] = (mid_1[3719:3712] > top_1[3727:3720]) ? 1 : 0;
assign detect_max[463][6] = (mid_1[3719:3712] > top_2[3711:3704]) ? 1 : 0;
assign detect_max[463][7] = (mid_1[3719:3712] > top_2[3719:3712]) ? 1 : 0;
assign detect_max[463][8] = (mid_1[3719:3712] > top_2[3727:3720]) ? 1 : 0;
assign detect_max[463][9] = (mid_1[3719:3712] > mid_0[3711:3704]) ? 1 : 0;
assign detect_max[463][10] = (mid_1[3719:3712] > mid_0[3719:3712]) ? 1 : 0;
assign detect_max[463][11] = (mid_1[3719:3712] > mid_0[3727:3720]) ? 1 : 0;
assign detect_max[463][12] = (mid_1[3719:3712] > mid_1[3711:3704]) ? 1 : 0;
assign detect_max[463][13] = (mid_1[3719:3712] > mid_1[3727:3720]) ? 1 : 0;
assign detect_max[463][14] = (mid_1[3719:3712] > mid_2[3711:3704]) ? 1 : 0;
assign detect_max[463][15] = (mid_1[3719:3712] > mid_2[3719:3712]) ? 1 : 0;
assign detect_max[463][16] = (mid_1[3719:3712] > mid_2[3727:3720]) ? 1 : 0;
assign detect_max[463][17] = (mid_1[3719:3712] > btm_0[3711:3704]) ? 1 : 0;
assign detect_max[463][18] = (mid_1[3719:3712] > btm_0[3719:3712]) ? 1 : 0;
assign detect_max[463][19] = (mid_1[3719:3712] > btm_0[3727:3720]) ? 1 : 0;
assign detect_max[463][20] = (mid_1[3719:3712] > btm_1[3711:3704]) ? 1 : 0;
assign detect_max[463][21] = (mid_1[3719:3712] > btm_1[3719:3712]) ? 1 : 0;
assign detect_max[463][22] = (mid_1[3719:3712] > btm_1[3727:3720]) ? 1 : 0;
assign detect_max[463][23] = (mid_1[3719:3712] > btm_2[3711:3704]) ? 1 : 0;
assign detect_max[463][24] = (mid_1[3719:3712] > btm_2[3719:3712]) ? 1 : 0;
assign detect_max[463][25] = (mid_1[3719:3712] > btm_2[3727:3720]) ? 1 : 0;

assign detect_max[464][0] = (mid_1[3727:3720] > top_0[3719:3712]) ? 1 : 0;
assign detect_max[464][1] = (mid_1[3727:3720] > top_0[3727:3720]) ? 1 : 0;
assign detect_max[464][2] = (mid_1[3727:3720] > top_0[3735:3728]) ? 1 : 0;
assign detect_max[464][3] = (mid_1[3727:3720] > top_1[3719:3712]) ? 1 : 0;
assign detect_max[464][4] = (mid_1[3727:3720] > top_1[3727:3720]) ? 1 : 0;
assign detect_max[464][5] = (mid_1[3727:3720] > top_1[3735:3728]) ? 1 : 0;
assign detect_max[464][6] = (mid_1[3727:3720] > top_2[3719:3712]) ? 1 : 0;
assign detect_max[464][7] = (mid_1[3727:3720] > top_2[3727:3720]) ? 1 : 0;
assign detect_max[464][8] = (mid_1[3727:3720] > top_2[3735:3728]) ? 1 : 0;
assign detect_max[464][9] = (mid_1[3727:3720] > mid_0[3719:3712]) ? 1 : 0;
assign detect_max[464][10] = (mid_1[3727:3720] > mid_0[3727:3720]) ? 1 : 0;
assign detect_max[464][11] = (mid_1[3727:3720] > mid_0[3735:3728]) ? 1 : 0;
assign detect_max[464][12] = (mid_1[3727:3720] > mid_1[3719:3712]) ? 1 : 0;
assign detect_max[464][13] = (mid_1[3727:3720] > mid_1[3735:3728]) ? 1 : 0;
assign detect_max[464][14] = (mid_1[3727:3720] > mid_2[3719:3712]) ? 1 : 0;
assign detect_max[464][15] = (mid_1[3727:3720] > mid_2[3727:3720]) ? 1 : 0;
assign detect_max[464][16] = (mid_1[3727:3720] > mid_2[3735:3728]) ? 1 : 0;
assign detect_max[464][17] = (mid_1[3727:3720] > btm_0[3719:3712]) ? 1 : 0;
assign detect_max[464][18] = (mid_1[3727:3720] > btm_0[3727:3720]) ? 1 : 0;
assign detect_max[464][19] = (mid_1[3727:3720] > btm_0[3735:3728]) ? 1 : 0;
assign detect_max[464][20] = (mid_1[3727:3720] > btm_1[3719:3712]) ? 1 : 0;
assign detect_max[464][21] = (mid_1[3727:3720] > btm_1[3727:3720]) ? 1 : 0;
assign detect_max[464][22] = (mid_1[3727:3720] > btm_1[3735:3728]) ? 1 : 0;
assign detect_max[464][23] = (mid_1[3727:3720] > btm_2[3719:3712]) ? 1 : 0;
assign detect_max[464][24] = (mid_1[3727:3720] > btm_2[3727:3720]) ? 1 : 0;
assign detect_max[464][25] = (mid_1[3727:3720] > btm_2[3735:3728]) ? 1 : 0;

assign detect_max[465][0] = (mid_1[3735:3728] > top_0[3727:3720]) ? 1 : 0;
assign detect_max[465][1] = (mid_1[3735:3728] > top_0[3735:3728]) ? 1 : 0;
assign detect_max[465][2] = (mid_1[3735:3728] > top_0[3743:3736]) ? 1 : 0;
assign detect_max[465][3] = (mid_1[3735:3728] > top_1[3727:3720]) ? 1 : 0;
assign detect_max[465][4] = (mid_1[3735:3728] > top_1[3735:3728]) ? 1 : 0;
assign detect_max[465][5] = (mid_1[3735:3728] > top_1[3743:3736]) ? 1 : 0;
assign detect_max[465][6] = (mid_1[3735:3728] > top_2[3727:3720]) ? 1 : 0;
assign detect_max[465][7] = (mid_1[3735:3728] > top_2[3735:3728]) ? 1 : 0;
assign detect_max[465][8] = (mid_1[3735:3728] > top_2[3743:3736]) ? 1 : 0;
assign detect_max[465][9] = (mid_1[3735:3728] > mid_0[3727:3720]) ? 1 : 0;
assign detect_max[465][10] = (mid_1[3735:3728] > mid_0[3735:3728]) ? 1 : 0;
assign detect_max[465][11] = (mid_1[3735:3728] > mid_0[3743:3736]) ? 1 : 0;
assign detect_max[465][12] = (mid_1[3735:3728] > mid_1[3727:3720]) ? 1 : 0;
assign detect_max[465][13] = (mid_1[3735:3728] > mid_1[3743:3736]) ? 1 : 0;
assign detect_max[465][14] = (mid_1[3735:3728] > mid_2[3727:3720]) ? 1 : 0;
assign detect_max[465][15] = (mid_1[3735:3728] > mid_2[3735:3728]) ? 1 : 0;
assign detect_max[465][16] = (mid_1[3735:3728] > mid_2[3743:3736]) ? 1 : 0;
assign detect_max[465][17] = (mid_1[3735:3728] > btm_0[3727:3720]) ? 1 : 0;
assign detect_max[465][18] = (mid_1[3735:3728] > btm_0[3735:3728]) ? 1 : 0;
assign detect_max[465][19] = (mid_1[3735:3728] > btm_0[3743:3736]) ? 1 : 0;
assign detect_max[465][20] = (mid_1[3735:3728] > btm_1[3727:3720]) ? 1 : 0;
assign detect_max[465][21] = (mid_1[3735:3728] > btm_1[3735:3728]) ? 1 : 0;
assign detect_max[465][22] = (mid_1[3735:3728] > btm_1[3743:3736]) ? 1 : 0;
assign detect_max[465][23] = (mid_1[3735:3728] > btm_2[3727:3720]) ? 1 : 0;
assign detect_max[465][24] = (mid_1[3735:3728] > btm_2[3735:3728]) ? 1 : 0;
assign detect_max[465][25] = (mid_1[3735:3728] > btm_2[3743:3736]) ? 1 : 0;

assign detect_max[466][0] = (mid_1[3743:3736] > top_0[3735:3728]) ? 1 : 0;
assign detect_max[466][1] = (mid_1[3743:3736] > top_0[3743:3736]) ? 1 : 0;
assign detect_max[466][2] = (mid_1[3743:3736] > top_0[3751:3744]) ? 1 : 0;
assign detect_max[466][3] = (mid_1[3743:3736] > top_1[3735:3728]) ? 1 : 0;
assign detect_max[466][4] = (mid_1[3743:3736] > top_1[3743:3736]) ? 1 : 0;
assign detect_max[466][5] = (mid_1[3743:3736] > top_1[3751:3744]) ? 1 : 0;
assign detect_max[466][6] = (mid_1[3743:3736] > top_2[3735:3728]) ? 1 : 0;
assign detect_max[466][7] = (mid_1[3743:3736] > top_2[3743:3736]) ? 1 : 0;
assign detect_max[466][8] = (mid_1[3743:3736] > top_2[3751:3744]) ? 1 : 0;
assign detect_max[466][9] = (mid_1[3743:3736] > mid_0[3735:3728]) ? 1 : 0;
assign detect_max[466][10] = (mid_1[3743:3736] > mid_0[3743:3736]) ? 1 : 0;
assign detect_max[466][11] = (mid_1[3743:3736] > mid_0[3751:3744]) ? 1 : 0;
assign detect_max[466][12] = (mid_1[3743:3736] > mid_1[3735:3728]) ? 1 : 0;
assign detect_max[466][13] = (mid_1[3743:3736] > mid_1[3751:3744]) ? 1 : 0;
assign detect_max[466][14] = (mid_1[3743:3736] > mid_2[3735:3728]) ? 1 : 0;
assign detect_max[466][15] = (mid_1[3743:3736] > mid_2[3743:3736]) ? 1 : 0;
assign detect_max[466][16] = (mid_1[3743:3736] > mid_2[3751:3744]) ? 1 : 0;
assign detect_max[466][17] = (mid_1[3743:3736] > btm_0[3735:3728]) ? 1 : 0;
assign detect_max[466][18] = (mid_1[3743:3736] > btm_0[3743:3736]) ? 1 : 0;
assign detect_max[466][19] = (mid_1[3743:3736] > btm_0[3751:3744]) ? 1 : 0;
assign detect_max[466][20] = (mid_1[3743:3736] > btm_1[3735:3728]) ? 1 : 0;
assign detect_max[466][21] = (mid_1[3743:3736] > btm_1[3743:3736]) ? 1 : 0;
assign detect_max[466][22] = (mid_1[3743:3736] > btm_1[3751:3744]) ? 1 : 0;
assign detect_max[466][23] = (mid_1[3743:3736] > btm_2[3735:3728]) ? 1 : 0;
assign detect_max[466][24] = (mid_1[3743:3736] > btm_2[3743:3736]) ? 1 : 0;
assign detect_max[466][25] = (mid_1[3743:3736] > btm_2[3751:3744]) ? 1 : 0;

assign detect_max[467][0] = (mid_1[3751:3744] > top_0[3743:3736]) ? 1 : 0;
assign detect_max[467][1] = (mid_1[3751:3744] > top_0[3751:3744]) ? 1 : 0;
assign detect_max[467][2] = (mid_1[3751:3744] > top_0[3759:3752]) ? 1 : 0;
assign detect_max[467][3] = (mid_1[3751:3744] > top_1[3743:3736]) ? 1 : 0;
assign detect_max[467][4] = (mid_1[3751:3744] > top_1[3751:3744]) ? 1 : 0;
assign detect_max[467][5] = (mid_1[3751:3744] > top_1[3759:3752]) ? 1 : 0;
assign detect_max[467][6] = (mid_1[3751:3744] > top_2[3743:3736]) ? 1 : 0;
assign detect_max[467][7] = (mid_1[3751:3744] > top_2[3751:3744]) ? 1 : 0;
assign detect_max[467][8] = (mid_1[3751:3744] > top_2[3759:3752]) ? 1 : 0;
assign detect_max[467][9] = (mid_1[3751:3744] > mid_0[3743:3736]) ? 1 : 0;
assign detect_max[467][10] = (mid_1[3751:3744] > mid_0[3751:3744]) ? 1 : 0;
assign detect_max[467][11] = (mid_1[3751:3744] > mid_0[3759:3752]) ? 1 : 0;
assign detect_max[467][12] = (mid_1[3751:3744] > mid_1[3743:3736]) ? 1 : 0;
assign detect_max[467][13] = (mid_1[3751:3744] > mid_1[3759:3752]) ? 1 : 0;
assign detect_max[467][14] = (mid_1[3751:3744] > mid_2[3743:3736]) ? 1 : 0;
assign detect_max[467][15] = (mid_1[3751:3744] > mid_2[3751:3744]) ? 1 : 0;
assign detect_max[467][16] = (mid_1[3751:3744] > mid_2[3759:3752]) ? 1 : 0;
assign detect_max[467][17] = (mid_1[3751:3744] > btm_0[3743:3736]) ? 1 : 0;
assign detect_max[467][18] = (mid_1[3751:3744] > btm_0[3751:3744]) ? 1 : 0;
assign detect_max[467][19] = (mid_1[3751:3744] > btm_0[3759:3752]) ? 1 : 0;
assign detect_max[467][20] = (mid_1[3751:3744] > btm_1[3743:3736]) ? 1 : 0;
assign detect_max[467][21] = (mid_1[3751:3744] > btm_1[3751:3744]) ? 1 : 0;
assign detect_max[467][22] = (mid_1[3751:3744] > btm_1[3759:3752]) ? 1 : 0;
assign detect_max[467][23] = (mid_1[3751:3744] > btm_2[3743:3736]) ? 1 : 0;
assign detect_max[467][24] = (mid_1[3751:3744] > btm_2[3751:3744]) ? 1 : 0;
assign detect_max[467][25] = (mid_1[3751:3744] > btm_2[3759:3752]) ? 1 : 0;

assign detect_max[468][0] = (mid_1[3759:3752] > top_0[3751:3744]) ? 1 : 0;
assign detect_max[468][1] = (mid_1[3759:3752] > top_0[3759:3752]) ? 1 : 0;
assign detect_max[468][2] = (mid_1[3759:3752] > top_0[3767:3760]) ? 1 : 0;
assign detect_max[468][3] = (mid_1[3759:3752] > top_1[3751:3744]) ? 1 : 0;
assign detect_max[468][4] = (mid_1[3759:3752] > top_1[3759:3752]) ? 1 : 0;
assign detect_max[468][5] = (mid_1[3759:3752] > top_1[3767:3760]) ? 1 : 0;
assign detect_max[468][6] = (mid_1[3759:3752] > top_2[3751:3744]) ? 1 : 0;
assign detect_max[468][7] = (mid_1[3759:3752] > top_2[3759:3752]) ? 1 : 0;
assign detect_max[468][8] = (mid_1[3759:3752] > top_2[3767:3760]) ? 1 : 0;
assign detect_max[468][9] = (mid_1[3759:3752] > mid_0[3751:3744]) ? 1 : 0;
assign detect_max[468][10] = (mid_1[3759:3752] > mid_0[3759:3752]) ? 1 : 0;
assign detect_max[468][11] = (mid_1[3759:3752] > mid_0[3767:3760]) ? 1 : 0;
assign detect_max[468][12] = (mid_1[3759:3752] > mid_1[3751:3744]) ? 1 : 0;
assign detect_max[468][13] = (mid_1[3759:3752] > mid_1[3767:3760]) ? 1 : 0;
assign detect_max[468][14] = (mid_1[3759:3752] > mid_2[3751:3744]) ? 1 : 0;
assign detect_max[468][15] = (mid_1[3759:3752] > mid_2[3759:3752]) ? 1 : 0;
assign detect_max[468][16] = (mid_1[3759:3752] > mid_2[3767:3760]) ? 1 : 0;
assign detect_max[468][17] = (mid_1[3759:3752] > btm_0[3751:3744]) ? 1 : 0;
assign detect_max[468][18] = (mid_1[3759:3752] > btm_0[3759:3752]) ? 1 : 0;
assign detect_max[468][19] = (mid_1[3759:3752] > btm_0[3767:3760]) ? 1 : 0;
assign detect_max[468][20] = (mid_1[3759:3752] > btm_1[3751:3744]) ? 1 : 0;
assign detect_max[468][21] = (mid_1[3759:3752] > btm_1[3759:3752]) ? 1 : 0;
assign detect_max[468][22] = (mid_1[3759:3752] > btm_1[3767:3760]) ? 1 : 0;
assign detect_max[468][23] = (mid_1[3759:3752] > btm_2[3751:3744]) ? 1 : 0;
assign detect_max[468][24] = (mid_1[3759:3752] > btm_2[3759:3752]) ? 1 : 0;
assign detect_max[468][25] = (mid_1[3759:3752] > btm_2[3767:3760]) ? 1 : 0;

assign detect_max[469][0] = (mid_1[3767:3760] > top_0[3759:3752]) ? 1 : 0;
assign detect_max[469][1] = (mid_1[3767:3760] > top_0[3767:3760]) ? 1 : 0;
assign detect_max[469][2] = (mid_1[3767:3760] > top_0[3775:3768]) ? 1 : 0;
assign detect_max[469][3] = (mid_1[3767:3760] > top_1[3759:3752]) ? 1 : 0;
assign detect_max[469][4] = (mid_1[3767:3760] > top_1[3767:3760]) ? 1 : 0;
assign detect_max[469][5] = (mid_1[3767:3760] > top_1[3775:3768]) ? 1 : 0;
assign detect_max[469][6] = (mid_1[3767:3760] > top_2[3759:3752]) ? 1 : 0;
assign detect_max[469][7] = (mid_1[3767:3760] > top_2[3767:3760]) ? 1 : 0;
assign detect_max[469][8] = (mid_1[3767:3760] > top_2[3775:3768]) ? 1 : 0;
assign detect_max[469][9] = (mid_1[3767:3760] > mid_0[3759:3752]) ? 1 : 0;
assign detect_max[469][10] = (mid_1[3767:3760] > mid_0[3767:3760]) ? 1 : 0;
assign detect_max[469][11] = (mid_1[3767:3760] > mid_0[3775:3768]) ? 1 : 0;
assign detect_max[469][12] = (mid_1[3767:3760] > mid_1[3759:3752]) ? 1 : 0;
assign detect_max[469][13] = (mid_1[3767:3760] > mid_1[3775:3768]) ? 1 : 0;
assign detect_max[469][14] = (mid_1[3767:3760] > mid_2[3759:3752]) ? 1 : 0;
assign detect_max[469][15] = (mid_1[3767:3760] > mid_2[3767:3760]) ? 1 : 0;
assign detect_max[469][16] = (mid_1[3767:3760] > mid_2[3775:3768]) ? 1 : 0;
assign detect_max[469][17] = (mid_1[3767:3760] > btm_0[3759:3752]) ? 1 : 0;
assign detect_max[469][18] = (mid_1[3767:3760] > btm_0[3767:3760]) ? 1 : 0;
assign detect_max[469][19] = (mid_1[3767:3760] > btm_0[3775:3768]) ? 1 : 0;
assign detect_max[469][20] = (mid_1[3767:3760] > btm_1[3759:3752]) ? 1 : 0;
assign detect_max[469][21] = (mid_1[3767:3760] > btm_1[3767:3760]) ? 1 : 0;
assign detect_max[469][22] = (mid_1[3767:3760] > btm_1[3775:3768]) ? 1 : 0;
assign detect_max[469][23] = (mid_1[3767:3760] > btm_2[3759:3752]) ? 1 : 0;
assign detect_max[469][24] = (mid_1[3767:3760] > btm_2[3767:3760]) ? 1 : 0;
assign detect_max[469][25] = (mid_1[3767:3760] > btm_2[3775:3768]) ? 1 : 0;

assign detect_max[470][0] = (mid_1[3775:3768] > top_0[3767:3760]) ? 1 : 0;
assign detect_max[470][1] = (mid_1[3775:3768] > top_0[3775:3768]) ? 1 : 0;
assign detect_max[470][2] = (mid_1[3775:3768] > top_0[3783:3776]) ? 1 : 0;
assign detect_max[470][3] = (mid_1[3775:3768] > top_1[3767:3760]) ? 1 : 0;
assign detect_max[470][4] = (mid_1[3775:3768] > top_1[3775:3768]) ? 1 : 0;
assign detect_max[470][5] = (mid_1[3775:3768] > top_1[3783:3776]) ? 1 : 0;
assign detect_max[470][6] = (mid_1[3775:3768] > top_2[3767:3760]) ? 1 : 0;
assign detect_max[470][7] = (mid_1[3775:3768] > top_2[3775:3768]) ? 1 : 0;
assign detect_max[470][8] = (mid_1[3775:3768] > top_2[3783:3776]) ? 1 : 0;
assign detect_max[470][9] = (mid_1[3775:3768] > mid_0[3767:3760]) ? 1 : 0;
assign detect_max[470][10] = (mid_1[3775:3768] > mid_0[3775:3768]) ? 1 : 0;
assign detect_max[470][11] = (mid_1[3775:3768] > mid_0[3783:3776]) ? 1 : 0;
assign detect_max[470][12] = (mid_1[3775:3768] > mid_1[3767:3760]) ? 1 : 0;
assign detect_max[470][13] = (mid_1[3775:3768] > mid_1[3783:3776]) ? 1 : 0;
assign detect_max[470][14] = (mid_1[3775:3768] > mid_2[3767:3760]) ? 1 : 0;
assign detect_max[470][15] = (mid_1[3775:3768] > mid_2[3775:3768]) ? 1 : 0;
assign detect_max[470][16] = (mid_1[3775:3768] > mid_2[3783:3776]) ? 1 : 0;
assign detect_max[470][17] = (mid_1[3775:3768] > btm_0[3767:3760]) ? 1 : 0;
assign detect_max[470][18] = (mid_1[3775:3768] > btm_0[3775:3768]) ? 1 : 0;
assign detect_max[470][19] = (mid_1[3775:3768] > btm_0[3783:3776]) ? 1 : 0;
assign detect_max[470][20] = (mid_1[3775:3768] > btm_1[3767:3760]) ? 1 : 0;
assign detect_max[470][21] = (mid_1[3775:3768] > btm_1[3775:3768]) ? 1 : 0;
assign detect_max[470][22] = (mid_1[3775:3768] > btm_1[3783:3776]) ? 1 : 0;
assign detect_max[470][23] = (mid_1[3775:3768] > btm_2[3767:3760]) ? 1 : 0;
assign detect_max[470][24] = (mid_1[3775:3768] > btm_2[3775:3768]) ? 1 : 0;
assign detect_max[470][25] = (mid_1[3775:3768] > btm_2[3783:3776]) ? 1 : 0;

assign detect_max[471][0] = (mid_1[3783:3776] > top_0[3775:3768]) ? 1 : 0;
assign detect_max[471][1] = (mid_1[3783:3776] > top_0[3783:3776]) ? 1 : 0;
assign detect_max[471][2] = (mid_1[3783:3776] > top_0[3791:3784]) ? 1 : 0;
assign detect_max[471][3] = (mid_1[3783:3776] > top_1[3775:3768]) ? 1 : 0;
assign detect_max[471][4] = (mid_1[3783:3776] > top_1[3783:3776]) ? 1 : 0;
assign detect_max[471][5] = (mid_1[3783:3776] > top_1[3791:3784]) ? 1 : 0;
assign detect_max[471][6] = (mid_1[3783:3776] > top_2[3775:3768]) ? 1 : 0;
assign detect_max[471][7] = (mid_1[3783:3776] > top_2[3783:3776]) ? 1 : 0;
assign detect_max[471][8] = (mid_1[3783:3776] > top_2[3791:3784]) ? 1 : 0;
assign detect_max[471][9] = (mid_1[3783:3776] > mid_0[3775:3768]) ? 1 : 0;
assign detect_max[471][10] = (mid_1[3783:3776] > mid_0[3783:3776]) ? 1 : 0;
assign detect_max[471][11] = (mid_1[3783:3776] > mid_0[3791:3784]) ? 1 : 0;
assign detect_max[471][12] = (mid_1[3783:3776] > mid_1[3775:3768]) ? 1 : 0;
assign detect_max[471][13] = (mid_1[3783:3776] > mid_1[3791:3784]) ? 1 : 0;
assign detect_max[471][14] = (mid_1[3783:3776] > mid_2[3775:3768]) ? 1 : 0;
assign detect_max[471][15] = (mid_1[3783:3776] > mid_2[3783:3776]) ? 1 : 0;
assign detect_max[471][16] = (mid_1[3783:3776] > mid_2[3791:3784]) ? 1 : 0;
assign detect_max[471][17] = (mid_1[3783:3776] > btm_0[3775:3768]) ? 1 : 0;
assign detect_max[471][18] = (mid_1[3783:3776] > btm_0[3783:3776]) ? 1 : 0;
assign detect_max[471][19] = (mid_1[3783:3776] > btm_0[3791:3784]) ? 1 : 0;
assign detect_max[471][20] = (mid_1[3783:3776] > btm_1[3775:3768]) ? 1 : 0;
assign detect_max[471][21] = (mid_1[3783:3776] > btm_1[3783:3776]) ? 1 : 0;
assign detect_max[471][22] = (mid_1[3783:3776] > btm_1[3791:3784]) ? 1 : 0;
assign detect_max[471][23] = (mid_1[3783:3776] > btm_2[3775:3768]) ? 1 : 0;
assign detect_max[471][24] = (mid_1[3783:3776] > btm_2[3783:3776]) ? 1 : 0;
assign detect_max[471][25] = (mid_1[3783:3776] > btm_2[3791:3784]) ? 1 : 0;

assign detect_max[472][0] = (mid_1[3791:3784] > top_0[3783:3776]) ? 1 : 0;
assign detect_max[472][1] = (mid_1[3791:3784] > top_0[3791:3784]) ? 1 : 0;
assign detect_max[472][2] = (mid_1[3791:3784] > top_0[3799:3792]) ? 1 : 0;
assign detect_max[472][3] = (mid_1[3791:3784] > top_1[3783:3776]) ? 1 : 0;
assign detect_max[472][4] = (mid_1[3791:3784] > top_1[3791:3784]) ? 1 : 0;
assign detect_max[472][5] = (mid_1[3791:3784] > top_1[3799:3792]) ? 1 : 0;
assign detect_max[472][6] = (mid_1[3791:3784] > top_2[3783:3776]) ? 1 : 0;
assign detect_max[472][7] = (mid_1[3791:3784] > top_2[3791:3784]) ? 1 : 0;
assign detect_max[472][8] = (mid_1[3791:3784] > top_2[3799:3792]) ? 1 : 0;
assign detect_max[472][9] = (mid_1[3791:3784] > mid_0[3783:3776]) ? 1 : 0;
assign detect_max[472][10] = (mid_1[3791:3784] > mid_0[3791:3784]) ? 1 : 0;
assign detect_max[472][11] = (mid_1[3791:3784] > mid_0[3799:3792]) ? 1 : 0;
assign detect_max[472][12] = (mid_1[3791:3784] > mid_1[3783:3776]) ? 1 : 0;
assign detect_max[472][13] = (mid_1[3791:3784] > mid_1[3799:3792]) ? 1 : 0;
assign detect_max[472][14] = (mid_1[3791:3784] > mid_2[3783:3776]) ? 1 : 0;
assign detect_max[472][15] = (mid_1[3791:3784] > mid_2[3791:3784]) ? 1 : 0;
assign detect_max[472][16] = (mid_1[3791:3784] > mid_2[3799:3792]) ? 1 : 0;
assign detect_max[472][17] = (mid_1[3791:3784] > btm_0[3783:3776]) ? 1 : 0;
assign detect_max[472][18] = (mid_1[3791:3784] > btm_0[3791:3784]) ? 1 : 0;
assign detect_max[472][19] = (mid_1[3791:3784] > btm_0[3799:3792]) ? 1 : 0;
assign detect_max[472][20] = (mid_1[3791:3784] > btm_1[3783:3776]) ? 1 : 0;
assign detect_max[472][21] = (mid_1[3791:3784] > btm_1[3791:3784]) ? 1 : 0;
assign detect_max[472][22] = (mid_1[3791:3784] > btm_1[3799:3792]) ? 1 : 0;
assign detect_max[472][23] = (mid_1[3791:3784] > btm_2[3783:3776]) ? 1 : 0;
assign detect_max[472][24] = (mid_1[3791:3784] > btm_2[3791:3784]) ? 1 : 0;
assign detect_max[472][25] = (mid_1[3791:3784] > btm_2[3799:3792]) ? 1 : 0;

assign detect_max[473][0] = (mid_1[3799:3792] > top_0[3791:3784]) ? 1 : 0;
assign detect_max[473][1] = (mid_1[3799:3792] > top_0[3799:3792]) ? 1 : 0;
assign detect_max[473][2] = (mid_1[3799:3792] > top_0[3807:3800]) ? 1 : 0;
assign detect_max[473][3] = (mid_1[3799:3792] > top_1[3791:3784]) ? 1 : 0;
assign detect_max[473][4] = (mid_1[3799:3792] > top_1[3799:3792]) ? 1 : 0;
assign detect_max[473][5] = (mid_1[3799:3792] > top_1[3807:3800]) ? 1 : 0;
assign detect_max[473][6] = (mid_1[3799:3792] > top_2[3791:3784]) ? 1 : 0;
assign detect_max[473][7] = (mid_1[3799:3792] > top_2[3799:3792]) ? 1 : 0;
assign detect_max[473][8] = (mid_1[3799:3792] > top_2[3807:3800]) ? 1 : 0;
assign detect_max[473][9] = (mid_1[3799:3792] > mid_0[3791:3784]) ? 1 : 0;
assign detect_max[473][10] = (mid_1[3799:3792] > mid_0[3799:3792]) ? 1 : 0;
assign detect_max[473][11] = (mid_1[3799:3792] > mid_0[3807:3800]) ? 1 : 0;
assign detect_max[473][12] = (mid_1[3799:3792] > mid_1[3791:3784]) ? 1 : 0;
assign detect_max[473][13] = (mid_1[3799:3792] > mid_1[3807:3800]) ? 1 : 0;
assign detect_max[473][14] = (mid_1[3799:3792] > mid_2[3791:3784]) ? 1 : 0;
assign detect_max[473][15] = (mid_1[3799:3792] > mid_2[3799:3792]) ? 1 : 0;
assign detect_max[473][16] = (mid_1[3799:3792] > mid_2[3807:3800]) ? 1 : 0;
assign detect_max[473][17] = (mid_1[3799:3792] > btm_0[3791:3784]) ? 1 : 0;
assign detect_max[473][18] = (mid_1[3799:3792] > btm_0[3799:3792]) ? 1 : 0;
assign detect_max[473][19] = (mid_1[3799:3792] > btm_0[3807:3800]) ? 1 : 0;
assign detect_max[473][20] = (mid_1[3799:3792] > btm_1[3791:3784]) ? 1 : 0;
assign detect_max[473][21] = (mid_1[3799:3792] > btm_1[3799:3792]) ? 1 : 0;
assign detect_max[473][22] = (mid_1[3799:3792] > btm_1[3807:3800]) ? 1 : 0;
assign detect_max[473][23] = (mid_1[3799:3792] > btm_2[3791:3784]) ? 1 : 0;
assign detect_max[473][24] = (mid_1[3799:3792] > btm_2[3799:3792]) ? 1 : 0;
assign detect_max[473][25] = (mid_1[3799:3792] > btm_2[3807:3800]) ? 1 : 0;

assign detect_max[474][0] = (mid_1[3807:3800] > top_0[3799:3792]) ? 1 : 0;
assign detect_max[474][1] = (mid_1[3807:3800] > top_0[3807:3800]) ? 1 : 0;
assign detect_max[474][2] = (mid_1[3807:3800] > top_0[3815:3808]) ? 1 : 0;
assign detect_max[474][3] = (mid_1[3807:3800] > top_1[3799:3792]) ? 1 : 0;
assign detect_max[474][4] = (mid_1[3807:3800] > top_1[3807:3800]) ? 1 : 0;
assign detect_max[474][5] = (mid_1[3807:3800] > top_1[3815:3808]) ? 1 : 0;
assign detect_max[474][6] = (mid_1[3807:3800] > top_2[3799:3792]) ? 1 : 0;
assign detect_max[474][7] = (mid_1[3807:3800] > top_2[3807:3800]) ? 1 : 0;
assign detect_max[474][8] = (mid_1[3807:3800] > top_2[3815:3808]) ? 1 : 0;
assign detect_max[474][9] = (mid_1[3807:3800] > mid_0[3799:3792]) ? 1 : 0;
assign detect_max[474][10] = (mid_1[3807:3800] > mid_0[3807:3800]) ? 1 : 0;
assign detect_max[474][11] = (mid_1[3807:3800] > mid_0[3815:3808]) ? 1 : 0;
assign detect_max[474][12] = (mid_1[3807:3800] > mid_1[3799:3792]) ? 1 : 0;
assign detect_max[474][13] = (mid_1[3807:3800] > mid_1[3815:3808]) ? 1 : 0;
assign detect_max[474][14] = (mid_1[3807:3800] > mid_2[3799:3792]) ? 1 : 0;
assign detect_max[474][15] = (mid_1[3807:3800] > mid_2[3807:3800]) ? 1 : 0;
assign detect_max[474][16] = (mid_1[3807:3800] > mid_2[3815:3808]) ? 1 : 0;
assign detect_max[474][17] = (mid_1[3807:3800] > btm_0[3799:3792]) ? 1 : 0;
assign detect_max[474][18] = (mid_1[3807:3800] > btm_0[3807:3800]) ? 1 : 0;
assign detect_max[474][19] = (mid_1[3807:3800] > btm_0[3815:3808]) ? 1 : 0;
assign detect_max[474][20] = (mid_1[3807:3800] > btm_1[3799:3792]) ? 1 : 0;
assign detect_max[474][21] = (mid_1[3807:3800] > btm_1[3807:3800]) ? 1 : 0;
assign detect_max[474][22] = (mid_1[3807:3800] > btm_1[3815:3808]) ? 1 : 0;
assign detect_max[474][23] = (mid_1[3807:3800] > btm_2[3799:3792]) ? 1 : 0;
assign detect_max[474][24] = (mid_1[3807:3800] > btm_2[3807:3800]) ? 1 : 0;
assign detect_max[474][25] = (mid_1[3807:3800] > btm_2[3815:3808]) ? 1 : 0;

assign detect_max[475][0] = (mid_1[3815:3808] > top_0[3807:3800]) ? 1 : 0;
assign detect_max[475][1] = (mid_1[3815:3808] > top_0[3815:3808]) ? 1 : 0;
assign detect_max[475][2] = (mid_1[3815:3808] > top_0[3823:3816]) ? 1 : 0;
assign detect_max[475][3] = (mid_1[3815:3808] > top_1[3807:3800]) ? 1 : 0;
assign detect_max[475][4] = (mid_1[3815:3808] > top_1[3815:3808]) ? 1 : 0;
assign detect_max[475][5] = (mid_1[3815:3808] > top_1[3823:3816]) ? 1 : 0;
assign detect_max[475][6] = (mid_1[3815:3808] > top_2[3807:3800]) ? 1 : 0;
assign detect_max[475][7] = (mid_1[3815:3808] > top_2[3815:3808]) ? 1 : 0;
assign detect_max[475][8] = (mid_1[3815:3808] > top_2[3823:3816]) ? 1 : 0;
assign detect_max[475][9] = (mid_1[3815:3808] > mid_0[3807:3800]) ? 1 : 0;
assign detect_max[475][10] = (mid_1[3815:3808] > mid_0[3815:3808]) ? 1 : 0;
assign detect_max[475][11] = (mid_1[3815:3808] > mid_0[3823:3816]) ? 1 : 0;
assign detect_max[475][12] = (mid_1[3815:3808] > mid_1[3807:3800]) ? 1 : 0;
assign detect_max[475][13] = (mid_1[3815:3808] > mid_1[3823:3816]) ? 1 : 0;
assign detect_max[475][14] = (mid_1[3815:3808] > mid_2[3807:3800]) ? 1 : 0;
assign detect_max[475][15] = (mid_1[3815:3808] > mid_2[3815:3808]) ? 1 : 0;
assign detect_max[475][16] = (mid_1[3815:3808] > mid_2[3823:3816]) ? 1 : 0;
assign detect_max[475][17] = (mid_1[3815:3808] > btm_0[3807:3800]) ? 1 : 0;
assign detect_max[475][18] = (mid_1[3815:3808] > btm_0[3815:3808]) ? 1 : 0;
assign detect_max[475][19] = (mid_1[3815:3808] > btm_0[3823:3816]) ? 1 : 0;
assign detect_max[475][20] = (mid_1[3815:3808] > btm_1[3807:3800]) ? 1 : 0;
assign detect_max[475][21] = (mid_1[3815:3808] > btm_1[3815:3808]) ? 1 : 0;
assign detect_max[475][22] = (mid_1[3815:3808] > btm_1[3823:3816]) ? 1 : 0;
assign detect_max[475][23] = (mid_1[3815:3808] > btm_2[3807:3800]) ? 1 : 0;
assign detect_max[475][24] = (mid_1[3815:3808] > btm_2[3815:3808]) ? 1 : 0;
assign detect_max[475][25] = (mid_1[3815:3808] > btm_2[3823:3816]) ? 1 : 0;

assign detect_max[476][0] = (mid_1[3823:3816] > top_0[3815:3808]) ? 1 : 0;
assign detect_max[476][1] = (mid_1[3823:3816] > top_0[3823:3816]) ? 1 : 0;
assign detect_max[476][2] = (mid_1[3823:3816] > top_0[3831:3824]) ? 1 : 0;
assign detect_max[476][3] = (mid_1[3823:3816] > top_1[3815:3808]) ? 1 : 0;
assign detect_max[476][4] = (mid_1[3823:3816] > top_1[3823:3816]) ? 1 : 0;
assign detect_max[476][5] = (mid_1[3823:3816] > top_1[3831:3824]) ? 1 : 0;
assign detect_max[476][6] = (mid_1[3823:3816] > top_2[3815:3808]) ? 1 : 0;
assign detect_max[476][7] = (mid_1[3823:3816] > top_2[3823:3816]) ? 1 : 0;
assign detect_max[476][8] = (mid_1[3823:3816] > top_2[3831:3824]) ? 1 : 0;
assign detect_max[476][9] = (mid_1[3823:3816] > mid_0[3815:3808]) ? 1 : 0;
assign detect_max[476][10] = (mid_1[3823:3816] > mid_0[3823:3816]) ? 1 : 0;
assign detect_max[476][11] = (mid_1[3823:3816] > mid_0[3831:3824]) ? 1 : 0;
assign detect_max[476][12] = (mid_1[3823:3816] > mid_1[3815:3808]) ? 1 : 0;
assign detect_max[476][13] = (mid_1[3823:3816] > mid_1[3831:3824]) ? 1 : 0;
assign detect_max[476][14] = (mid_1[3823:3816] > mid_2[3815:3808]) ? 1 : 0;
assign detect_max[476][15] = (mid_1[3823:3816] > mid_2[3823:3816]) ? 1 : 0;
assign detect_max[476][16] = (mid_1[3823:3816] > mid_2[3831:3824]) ? 1 : 0;
assign detect_max[476][17] = (mid_1[3823:3816] > btm_0[3815:3808]) ? 1 : 0;
assign detect_max[476][18] = (mid_1[3823:3816] > btm_0[3823:3816]) ? 1 : 0;
assign detect_max[476][19] = (mid_1[3823:3816] > btm_0[3831:3824]) ? 1 : 0;
assign detect_max[476][20] = (mid_1[3823:3816] > btm_1[3815:3808]) ? 1 : 0;
assign detect_max[476][21] = (mid_1[3823:3816] > btm_1[3823:3816]) ? 1 : 0;
assign detect_max[476][22] = (mid_1[3823:3816] > btm_1[3831:3824]) ? 1 : 0;
assign detect_max[476][23] = (mid_1[3823:3816] > btm_2[3815:3808]) ? 1 : 0;
assign detect_max[476][24] = (mid_1[3823:3816] > btm_2[3823:3816]) ? 1 : 0;
assign detect_max[476][25] = (mid_1[3823:3816] > btm_2[3831:3824]) ? 1 : 0;

assign detect_max[477][0] = (mid_1[3831:3824] > top_0[3823:3816]) ? 1 : 0;
assign detect_max[477][1] = (mid_1[3831:3824] > top_0[3831:3824]) ? 1 : 0;
assign detect_max[477][2] = (mid_1[3831:3824] > top_0[3839:3832]) ? 1 : 0;
assign detect_max[477][3] = (mid_1[3831:3824] > top_1[3823:3816]) ? 1 : 0;
assign detect_max[477][4] = (mid_1[3831:3824] > top_1[3831:3824]) ? 1 : 0;
assign detect_max[477][5] = (mid_1[3831:3824] > top_1[3839:3832]) ? 1 : 0;
assign detect_max[477][6] = (mid_1[3831:3824] > top_2[3823:3816]) ? 1 : 0;
assign detect_max[477][7] = (mid_1[3831:3824] > top_2[3831:3824]) ? 1 : 0;
assign detect_max[477][8] = (mid_1[3831:3824] > top_2[3839:3832]) ? 1 : 0;
assign detect_max[477][9] = (mid_1[3831:3824] > mid_0[3823:3816]) ? 1 : 0;
assign detect_max[477][10] = (mid_1[3831:3824] > mid_0[3831:3824]) ? 1 : 0;
assign detect_max[477][11] = (mid_1[3831:3824] > mid_0[3839:3832]) ? 1 : 0;
assign detect_max[477][12] = (mid_1[3831:3824] > mid_1[3823:3816]) ? 1 : 0;
assign detect_max[477][13] = (mid_1[3831:3824] > mid_1[3839:3832]) ? 1 : 0;
assign detect_max[477][14] = (mid_1[3831:3824] > mid_2[3823:3816]) ? 1 : 0;
assign detect_max[477][15] = (mid_1[3831:3824] > mid_2[3831:3824]) ? 1 : 0;
assign detect_max[477][16] = (mid_1[3831:3824] > mid_2[3839:3832]) ? 1 : 0;
assign detect_max[477][17] = (mid_1[3831:3824] > btm_0[3823:3816]) ? 1 : 0;
assign detect_max[477][18] = (mid_1[3831:3824] > btm_0[3831:3824]) ? 1 : 0;
assign detect_max[477][19] = (mid_1[3831:3824] > btm_0[3839:3832]) ? 1 : 0;
assign detect_max[477][20] = (mid_1[3831:3824] > btm_1[3823:3816]) ? 1 : 0;
assign detect_max[477][21] = (mid_1[3831:3824] > btm_1[3831:3824]) ? 1 : 0;
assign detect_max[477][22] = (mid_1[3831:3824] > btm_1[3839:3832]) ? 1 : 0;
assign detect_max[477][23] = (mid_1[3831:3824] > btm_2[3823:3816]) ? 1 : 0;
assign detect_max[477][24] = (mid_1[3831:3824] > btm_2[3831:3824]) ? 1 : 0;
assign detect_max[477][25] = (mid_1[3831:3824] > btm_2[3839:3832]) ? 1 : 0;

assign detect_max[478][0] = (mid_1[3839:3832] > top_0[3831:3824]) ? 1 : 0;
assign detect_max[478][1] = (mid_1[3839:3832] > top_0[3839:3832]) ? 1 : 0;
assign detect_max[478][2] = (mid_1[3839:3832] > top_0[3847:3840]) ? 1 : 0;
assign detect_max[478][3] = (mid_1[3839:3832] > top_1[3831:3824]) ? 1 : 0;
assign detect_max[478][4] = (mid_1[3839:3832] > top_1[3839:3832]) ? 1 : 0;
assign detect_max[478][5] = (mid_1[3839:3832] > top_1[3847:3840]) ? 1 : 0;
assign detect_max[478][6] = (mid_1[3839:3832] > top_2[3831:3824]) ? 1 : 0;
assign detect_max[478][7] = (mid_1[3839:3832] > top_2[3839:3832]) ? 1 : 0;
assign detect_max[478][8] = (mid_1[3839:3832] > top_2[3847:3840]) ? 1 : 0;
assign detect_max[478][9] = (mid_1[3839:3832] > mid_0[3831:3824]) ? 1 : 0;
assign detect_max[478][10] = (mid_1[3839:3832] > mid_0[3839:3832]) ? 1 : 0;
assign detect_max[478][11] = (mid_1[3839:3832] > mid_0[3847:3840]) ? 1 : 0;
assign detect_max[478][12] = (mid_1[3839:3832] > mid_1[3831:3824]) ? 1 : 0;
assign detect_max[478][13] = (mid_1[3839:3832] > mid_1[3847:3840]) ? 1 : 0;
assign detect_max[478][14] = (mid_1[3839:3832] > mid_2[3831:3824]) ? 1 : 0;
assign detect_max[478][15] = (mid_1[3839:3832] > mid_2[3839:3832]) ? 1 : 0;
assign detect_max[478][16] = (mid_1[3839:3832] > mid_2[3847:3840]) ? 1 : 0;
assign detect_max[478][17] = (mid_1[3839:3832] > btm_0[3831:3824]) ? 1 : 0;
assign detect_max[478][18] = (mid_1[3839:3832] > btm_0[3839:3832]) ? 1 : 0;
assign detect_max[478][19] = (mid_1[3839:3832] > btm_0[3847:3840]) ? 1 : 0;
assign detect_max[478][20] = (mid_1[3839:3832] > btm_1[3831:3824]) ? 1 : 0;
assign detect_max[478][21] = (mid_1[3839:3832] > btm_1[3839:3832]) ? 1 : 0;
assign detect_max[478][22] = (mid_1[3839:3832] > btm_1[3847:3840]) ? 1 : 0;
assign detect_max[478][23] = (mid_1[3839:3832] > btm_2[3831:3824]) ? 1 : 0;
assign detect_max[478][24] = (mid_1[3839:3832] > btm_2[3839:3832]) ? 1 : 0;
assign detect_max[478][25] = (mid_1[3839:3832] > btm_2[3847:3840]) ? 1 : 0;

assign detect_max[479][0] = (mid_1[3847:3840] > top_0[3839:3832]) ? 1 : 0;
assign detect_max[479][1] = (mid_1[3847:3840] > top_0[3847:3840]) ? 1 : 0;
assign detect_max[479][2] = (mid_1[3847:3840] > top_0[3855:3848]) ? 1 : 0;
assign detect_max[479][3] = (mid_1[3847:3840] > top_1[3839:3832]) ? 1 : 0;
assign detect_max[479][4] = (mid_1[3847:3840] > top_1[3847:3840]) ? 1 : 0;
assign detect_max[479][5] = (mid_1[3847:3840] > top_1[3855:3848]) ? 1 : 0;
assign detect_max[479][6] = (mid_1[3847:3840] > top_2[3839:3832]) ? 1 : 0;
assign detect_max[479][7] = (mid_1[3847:3840] > top_2[3847:3840]) ? 1 : 0;
assign detect_max[479][8] = (mid_1[3847:3840] > top_2[3855:3848]) ? 1 : 0;
assign detect_max[479][9] = (mid_1[3847:3840] > mid_0[3839:3832]) ? 1 : 0;
assign detect_max[479][10] = (mid_1[3847:3840] > mid_0[3847:3840]) ? 1 : 0;
assign detect_max[479][11] = (mid_1[3847:3840] > mid_0[3855:3848]) ? 1 : 0;
assign detect_max[479][12] = (mid_1[3847:3840] > mid_1[3839:3832]) ? 1 : 0;
assign detect_max[479][13] = (mid_1[3847:3840] > mid_1[3855:3848]) ? 1 : 0;
assign detect_max[479][14] = (mid_1[3847:3840] > mid_2[3839:3832]) ? 1 : 0;
assign detect_max[479][15] = (mid_1[3847:3840] > mid_2[3847:3840]) ? 1 : 0;
assign detect_max[479][16] = (mid_1[3847:3840] > mid_2[3855:3848]) ? 1 : 0;
assign detect_max[479][17] = (mid_1[3847:3840] > btm_0[3839:3832]) ? 1 : 0;
assign detect_max[479][18] = (mid_1[3847:3840] > btm_0[3847:3840]) ? 1 : 0;
assign detect_max[479][19] = (mid_1[3847:3840] > btm_0[3855:3848]) ? 1 : 0;
assign detect_max[479][20] = (mid_1[3847:3840] > btm_1[3839:3832]) ? 1 : 0;
assign detect_max[479][21] = (mid_1[3847:3840] > btm_1[3847:3840]) ? 1 : 0;
assign detect_max[479][22] = (mid_1[3847:3840] > btm_1[3855:3848]) ? 1 : 0;
assign detect_max[479][23] = (mid_1[3847:3840] > btm_2[3839:3832]) ? 1 : 0;
assign detect_max[479][24] = (mid_1[3847:3840] > btm_2[3847:3840]) ? 1 : 0;
assign detect_max[479][25] = (mid_1[3847:3840] > btm_2[3855:3848]) ? 1 : 0;

assign detect_max[480][0] = (mid_1[3855:3848] > top_0[3847:3840]) ? 1 : 0;
assign detect_max[480][1] = (mid_1[3855:3848] > top_0[3855:3848]) ? 1 : 0;
assign detect_max[480][2] = (mid_1[3855:3848] > top_0[3863:3856]) ? 1 : 0;
assign detect_max[480][3] = (mid_1[3855:3848] > top_1[3847:3840]) ? 1 : 0;
assign detect_max[480][4] = (mid_1[3855:3848] > top_1[3855:3848]) ? 1 : 0;
assign detect_max[480][5] = (mid_1[3855:3848] > top_1[3863:3856]) ? 1 : 0;
assign detect_max[480][6] = (mid_1[3855:3848] > top_2[3847:3840]) ? 1 : 0;
assign detect_max[480][7] = (mid_1[3855:3848] > top_2[3855:3848]) ? 1 : 0;
assign detect_max[480][8] = (mid_1[3855:3848] > top_2[3863:3856]) ? 1 : 0;
assign detect_max[480][9] = (mid_1[3855:3848] > mid_0[3847:3840]) ? 1 : 0;
assign detect_max[480][10] = (mid_1[3855:3848] > mid_0[3855:3848]) ? 1 : 0;
assign detect_max[480][11] = (mid_1[3855:3848] > mid_0[3863:3856]) ? 1 : 0;
assign detect_max[480][12] = (mid_1[3855:3848] > mid_1[3847:3840]) ? 1 : 0;
assign detect_max[480][13] = (mid_1[3855:3848] > mid_1[3863:3856]) ? 1 : 0;
assign detect_max[480][14] = (mid_1[3855:3848] > mid_2[3847:3840]) ? 1 : 0;
assign detect_max[480][15] = (mid_1[3855:3848] > mid_2[3855:3848]) ? 1 : 0;
assign detect_max[480][16] = (mid_1[3855:3848] > mid_2[3863:3856]) ? 1 : 0;
assign detect_max[480][17] = (mid_1[3855:3848] > btm_0[3847:3840]) ? 1 : 0;
assign detect_max[480][18] = (mid_1[3855:3848] > btm_0[3855:3848]) ? 1 : 0;
assign detect_max[480][19] = (mid_1[3855:3848] > btm_0[3863:3856]) ? 1 : 0;
assign detect_max[480][20] = (mid_1[3855:3848] > btm_1[3847:3840]) ? 1 : 0;
assign detect_max[480][21] = (mid_1[3855:3848] > btm_1[3855:3848]) ? 1 : 0;
assign detect_max[480][22] = (mid_1[3855:3848] > btm_1[3863:3856]) ? 1 : 0;
assign detect_max[480][23] = (mid_1[3855:3848] > btm_2[3847:3840]) ? 1 : 0;
assign detect_max[480][24] = (mid_1[3855:3848] > btm_2[3855:3848]) ? 1 : 0;
assign detect_max[480][25] = (mid_1[3855:3848] > btm_2[3863:3856]) ? 1 : 0;

assign detect_max[481][0] = (mid_1[3863:3856] > top_0[3855:3848]) ? 1 : 0;
assign detect_max[481][1] = (mid_1[3863:3856] > top_0[3863:3856]) ? 1 : 0;
assign detect_max[481][2] = (mid_1[3863:3856] > top_0[3871:3864]) ? 1 : 0;
assign detect_max[481][3] = (mid_1[3863:3856] > top_1[3855:3848]) ? 1 : 0;
assign detect_max[481][4] = (mid_1[3863:3856] > top_1[3863:3856]) ? 1 : 0;
assign detect_max[481][5] = (mid_1[3863:3856] > top_1[3871:3864]) ? 1 : 0;
assign detect_max[481][6] = (mid_1[3863:3856] > top_2[3855:3848]) ? 1 : 0;
assign detect_max[481][7] = (mid_1[3863:3856] > top_2[3863:3856]) ? 1 : 0;
assign detect_max[481][8] = (mid_1[3863:3856] > top_2[3871:3864]) ? 1 : 0;
assign detect_max[481][9] = (mid_1[3863:3856] > mid_0[3855:3848]) ? 1 : 0;
assign detect_max[481][10] = (mid_1[3863:3856] > mid_0[3863:3856]) ? 1 : 0;
assign detect_max[481][11] = (mid_1[3863:3856] > mid_0[3871:3864]) ? 1 : 0;
assign detect_max[481][12] = (mid_1[3863:3856] > mid_1[3855:3848]) ? 1 : 0;
assign detect_max[481][13] = (mid_1[3863:3856] > mid_1[3871:3864]) ? 1 : 0;
assign detect_max[481][14] = (mid_1[3863:3856] > mid_2[3855:3848]) ? 1 : 0;
assign detect_max[481][15] = (mid_1[3863:3856] > mid_2[3863:3856]) ? 1 : 0;
assign detect_max[481][16] = (mid_1[3863:3856] > mid_2[3871:3864]) ? 1 : 0;
assign detect_max[481][17] = (mid_1[3863:3856] > btm_0[3855:3848]) ? 1 : 0;
assign detect_max[481][18] = (mid_1[3863:3856] > btm_0[3863:3856]) ? 1 : 0;
assign detect_max[481][19] = (mid_1[3863:3856] > btm_0[3871:3864]) ? 1 : 0;
assign detect_max[481][20] = (mid_1[3863:3856] > btm_1[3855:3848]) ? 1 : 0;
assign detect_max[481][21] = (mid_1[3863:3856] > btm_1[3863:3856]) ? 1 : 0;
assign detect_max[481][22] = (mid_1[3863:3856] > btm_1[3871:3864]) ? 1 : 0;
assign detect_max[481][23] = (mid_1[3863:3856] > btm_2[3855:3848]) ? 1 : 0;
assign detect_max[481][24] = (mid_1[3863:3856] > btm_2[3863:3856]) ? 1 : 0;
assign detect_max[481][25] = (mid_1[3863:3856] > btm_2[3871:3864]) ? 1 : 0;

assign detect_max[482][0] = (mid_1[3871:3864] > top_0[3863:3856]) ? 1 : 0;
assign detect_max[482][1] = (mid_1[3871:3864] > top_0[3871:3864]) ? 1 : 0;
assign detect_max[482][2] = (mid_1[3871:3864] > top_0[3879:3872]) ? 1 : 0;
assign detect_max[482][3] = (mid_1[3871:3864] > top_1[3863:3856]) ? 1 : 0;
assign detect_max[482][4] = (mid_1[3871:3864] > top_1[3871:3864]) ? 1 : 0;
assign detect_max[482][5] = (mid_1[3871:3864] > top_1[3879:3872]) ? 1 : 0;
assign detect_max[482][6] = (mid_1[3871:3864] > top_2[3863:3856]) ? 1 : 0;
assign detect_max[482][7] = (mid_1[3871:3864] > top_2[3871:3864]) ? 1 : 0;
assign detect_max[482][8] = (mid_1[3871:3864] > top_2[3879:3872]) ? 1 : 0;
assign detect_max[482][9] = (mid_1[3871:3864] > mid_0[3863:3856]) ? 1 : 0;
assign detect_max[482][10] = (mid_1[3871:3864] > mid_0[3871:3864]) ? 1 : 0;
assign detect_max[482][11] = (mid_1[3871:3864] > mid_0[3879:3872]) ? 1 : 0;
assign detect_max[482][12] = (mid_1[3871:3864] > mid_1[3863:3856]) ? 1 : 0;
assign detect_max[482][13] = (mid_1[3871:3864] > mid_1[3879:3872]) ? 1 : 0;
assign detect_max[482][14] = (mid_1[3871:3864] > mid_2[3863:3856]) ? 1 : 0;
assign detect_max[482][15] = (mid_1[3871:3864] > mid_2[3871:3864]) ? 1 : 0;
assign detect_max[482][16] = (mid_1[3871:3864] > mid_2[3879:3872]) ? 1 : 0;
assign detect_max[482][17] = (mid_1[3871:3864] > btm_0[3863:3856]) ? 1 : 0;
assign detect_max[482][18] = (mid_1[3871:3864] > btm_0[3871:3864]) ? 1 : 0;
assign detect_max[482][19] = (mid_1[3871:3864] > btm_0[3879:3872]) ? 1 : 0;
assign detect_max[482][20] = (mid_1[3871:3864] > btm_1[3863:3856]) ? 1 : 0;
assign detect_max[482][21] = (mid_1[3871:3864] > btm_1[3871:3864]) ? 1 : 0;
assign detect_max[482][22] = (mid_1[3871:3864] > btm_1[3879:3872]) ? 1 : 0;
assign detect_max[482][23] = (mid_1[3871:3864] > btm_2[3863:3856]) ? 1 : 0;
assign detect_max[482][24] = (mid_1[3871:3864] > btm_2[3871:3864]) ? 1 : 0;
assign detect_max[482][25] = (mid_1[3871:3864] > btm_2[3879:3872]) ? 1 : 0;

assign detect_max[483][0] = (mid_1[3879:3872] > top_0[3871:3864]) ? 1 : 0;
assign detect_max[483][1] = (mid_1[3879:3872] > top_0[3879:3872]) ? 1 : 0;
assign detect_max[483][2] = (mid_1[3879:3872] > top_0[3887:3880]) ? 1 : 0;
assign detect_max[483][3] = (mid_1[3879:3872] > top_1[3871:3864]) ? 1 : 0;
assign detect_max[483][4] = (mid_1[3879:3872] > top_1[3879:3872]) ? 1 : 0;
assign detect_max[483][5] = (mid_1[3879:3872] > top_1[3887:3880]) ? 1 : 0;
assign detect_max[483][6] = (mid_1[3879:3872] > top_2[3871:3864]) ? 1 : 0;
assign detect_max[483][7] = (mid_1[3879:3872] > top_2[3879:3872]) ? 1 : 0;
assign detect_max[483][8] = (mid_1[3879:3872] > top_2[3887:3880]) ? 1 : 0;
assign detect_max[483][9] = (mid_1[3879:3872] > mid_0[3871:3864]) ? 1 : 0;
assign detect_max[483][10] = (mid_1[3879:3872] > mid_0[3879:3872]) ? 1 : 0;
assign detect_max[483][11] = (mid_1[3879:3872] > mid_0[3887:3880]) ? 1 : 0;
assign detect_max[483][12] = (mid_1[3879:3872] > mid_1[3871:3864]) ? 1 : 0;
assign detect_max[483][13] = (mid_1[3879:3872] > mid_1[3887:3880]) ? 1 : 0;
assign detect_max[483][14] = (mid_1[3879:3872] > mid_2[3871:3864]) ? 1 : 0;
assign detect_max[483][15] = (mid_1[3879:3872] > mid_2[3879:3872]) ? 1 : 0;
assign detect_max[483][16] = (mid_1[3879:3872] > mid_2[3887:3880]) ? 1 : 0;
assign detect_max[483][17] = (mid_1[3879:3872] > btm_0[3871:3864]) ? 1 : 0;
assign detect_max[483][18] = (mid_1[3879:3872] > btm_0[3879:3872]) ? 1 : 0;
assign detect_max[483][19] = (mid_1[3879:3872] > btm_0[3887:3880]) ? 1 : 0;
assign detect_max[483][20] = (mid_1[3879:3872] > btm_1[3871:3864]) ? 1 : 0;
assign detect_max[483][21] = (mid_1[3879:3872] > btm_1[3879:3872]) ? 1 : 0;
assign detect_max[483][22] = (mid_1[3879:3872] > btm_1[3887:3880]) ? 1 : 0;
assign detect_max[483][23] = (mid_1[3879:3872] > btm_2[3871:3864]) ? 1 : 0;
assign detect_max[483][24] = (mid_1[3879:3872] > btm_2[3879:3872]) ? 1 : 0;
assign detect_max[483][25] = (mid_1[3879:3872] > btm_2[3887:3880]) ? 1 : 0;

assign detect_max[484][0] = (mid_1[3887:3880] > top_0[3879:3872]) ? 1 : 0;
assign detect_max[484][1] = (mid_1[3887:3880] > top_0[3887:3880]) ? 1 : 0;
assign detect_max[484][2] = (mid_1[3887:3880] > top_0[3895:3888]) ? 1 : 0;
assign detect_max[484][3] = (mid_1[3887:3880] > top_1[3879:3872]) ? 1 : 0;
assign detect_max[484][4] = (mid_1[3887:3880] > top_1[3887:3880]) ? 1 : 0;
assign detect_max[484][5] = (mid_1[3887:3880] > top_1[3895:3888]) ? 1 : 0;
assign detect_max[484][6] = (mid_1[3887:3880] > top_2[3879:3872]) ? 1 : 0;
assign detect_max[484][7] = (mid_1[3887:3880] > top_2[3887:3880]) ? 1 : 0;
assign detect_max[484][8] = (mid_1[3887:3880] > top_2[3895:3888]) ? 1 : 0;
assign detect_max[484][9] = (mid_1[3887:3880] > mid_0[3879:3872]) ? 1 : 0;
assign detect_max[484][10] = (mid_1[3887:3880] > mid_0[3887:3880]) ? 1 : 0;
assign detect_max[484][11] = (mid_1[3887:3880] > mid_0[3895:3888]) ? 1 : 0;
assign detect_max[484][12] = (mid_1[3887:3880] > mid_1[3879:3872]) ? 1 : 0;
assign detect_max[484][13] = (mid_1[3887:3880] > mid_1[3895:3888]) ? 1 : 0;
assign detect_max[484][14] = (mid_1[3887:3880] > mid_2[3879:3872]) ? 1 : 0;
assign detect_max[484][15] = (mid_1[3887:3880] > mid_2[3887:3880]) ? 1 : 0;
assign detect_max[484][16] = (mid_1[3887:3880] > mid_2[3895:3888]) ? 1 : 0;
assign detect_max[484][17] = (mid_1[3887:3880] > btm_0[3879:3872]) ? 1 : 0;
assign detect_max[484][18] = (mid_1[3887:3880] > btm_0[3887:3880]) ? 1 : 0;
assign detect_max[484][19] = (mid_1[3887:3880] > btm_0[3895:3888]) ? 1 : 0;
assign detect_max[484][20] = (mid_1[3887:3880] > btm_1[3879:3872]) ? 1 : 0;
assign detect_max[484][21] = (mid_1[3887:3880] > btm_1[3887:3880]) ? 1 : 0;
assign detect_max[484][22] = (mid_1[3887:3880] > btm_1[3895:3888]) ? 1 : 0;
assign detect_max[484][23] = (mid_1[3887:3880] > btm_2[3879:3872]) ? 1 : 0;
assign detect_max[484][24] = (mid_1[3887:3880] > btm_2[3887:3880]) ? 1 : 0;
assign detect_max[484][25] = (mid_1[3887:3880] > btm_2[3895:3888]) ? 1 : 0;

assign detect_max[485][0] = (mid_1[3895:3888] > top_0[3887:3880]) ? 1 : 0;
assign detect_max[485][1] = (mid_1[3895:3888] > top_0[3895:3888]) ? 1 : 0;
assign detect_max[485][2] = (mid_1[3895:3888] > top_0[3903:3896]) ? 1 : 0;
assign detect_max[485][3] = (mid_1[3895:3888] > top_1[3887:3880]) ? 1 : 0;
assign detect_max[485][4] = (mid_1[3895:3888] > top_1[3895:3888]) ? 1 : 0;
assign detect_max[485][5] = (mid_1[3895:3888] > top_1[3903:3896]) ? 1 : 0;
assign detect_max[485][6] = (mid_1[3895:3888] > top_2[3887:3880]) ? 1 : 0;
assign detect_max[485][7] = (mid_1[3895:3888] > top_2[3895:3888]) ? 1 : 0;
assign detect_max[485][8] = (mid_1[3895:3888] > top_2[3903:3896]) ? 1 : 0;
assign detect_max[485][9] = (mid_1[3895:3888] > mid_0[3887:3880]) ? 1 : 0;
assign detect_max[485][10] = (mid_1[3895:3888] > mid_0[3895:3888]) ? 1 : 0;
assign detect_max[485][11] = (mid_1[3895:3888] > mid_0[3903:3896]) ? 1 : 0;
assign detect_max[485][12] = (mid_1[3895:3888] > mid_1[3887:3880]) ? 1 : 0;
assign detect_max[485][13] = (mid_1[3895:3888] > mid_1[3903:3896]) ? 1 : 0;
assign detect_max[485][14] = (mid_1[3895:3888] > mid_2[3887:3880]) ? 1 : 0;
assign detect_max[485][15] = (mid_1[3895:3888] > mid_2[3895:3888]) ? 1 : 0;
assign detect_max[485][16] = (mid_1[3895:3888] > mid_2[3903:3896]) ? 1 : 0;
assign detect_max[485][17] = (mid_1[3895:3888] > btm_0[3887:3880]) ? 1 : 0;
assign detect_max[485][18] = (mid_1[3895:3888] > btm_0[3895:3888]) ? 1 : 0;
assign detect_max[485][19] = (mid_1[3895:3888] > btm_0[3903:3896]) ? 1 : 0;
assign detect_max[485][20] = (mid_1[3895:3888] > btm_1[3887:3880]) ? 1 : 0;
assign detect_max[485][21] = (mid_1[3895:3888] > btm_1[3895:3888]) ? 1 : 0;
assign detect_max[485][22] = (mid_1[3895:3888] > btm_1[3903:3896]) ? 1 : 0;
assign detect_max[485][23] = (mid_1[3895:3888] > btm_2[3887:3880]) ? 1 : 0;
assign detect_max[485][24] = (mid_1[3895:3888] > btm_2[3895:3888]) ? 1 : 0;
assign detect_max[485][25] = (mid_1[3895:3888] > btm_2[3903:3896]) ? 1 : 0;

assign detect_max[486][0] = (mid_1[3903:3896] > top_0[3895:3888]) ? 1 : 0;
assign detect_max[486][1] = (mid_1[3903:3896] > top_0[3903:3896]) ? 1 : 0;
assign detect_max[486][2] = (mid_1[3903:3896] > top_0[3911:3904]) ? 1 : 0;
assign detect_max[486][3] = (mid_1[3903:3896] > top_1[3895:3888]) ? 1 : 0;
assign detect_max[486][4] = (mid_1[3903:3896] > top_1[3903:3896]) ? 1 : 0;
assign detect_max[486][5] = (mid_1[3903:3896] > top_1[3911:3904]) ? 1 : 0;
assign detect_max[486][6] = (mid_1[3903:3896] > top_2[3895:3888]) ? 1 : 0;
assign detect_max[486][7] = (mid_1[3903:3896] > top_2[3903:3896]) ? 1 : 0;
assign detect_max[486][8] = (mid_1[3903:3896] > top_2[3911:3904]) ? 1 : 0;
assign detect_max[486][9] = (mid_1[3903:3896] > mid_0[3895:3888]) ? 1 : 0;
assign detect_max[486][10] = (mid_1[3903:3896] > mid_0[3903:3896]) ? 1 : 0;
assign detect_max[486][11] = (mid_1[3903:3896] > mid_0[3911:3904]) ? 1 : 0;
assign detect_max[486][12] = (mid_1[3903:3896] > mid_1[3895:3888]) ? 1 : 0;
assign detect_max[486][13] = (mid_1[3903:3896] > mid_1[3911:3904]) ? 1 : 0;
assign detect_max[486][14] = (mid_1[3903:3896] > mid_2[3895:3888]) ? 1 : 0;
assign detect_max[486][15] = (mid_1[3903:3896] > mid_2[3903:3896]) ? 1 : 0;
assign detect_max[486][16] = (mid_1[3903:3896] > mid_2[3911:3904]) ? 1 : 0;
assign detect_max[486][17] = (mid_1[3903:3896] > btm_0[3895:3888]) ? 1 : 0;
assign detect_max[486][18] = (mid_1[3903:3896] > btm_0[3903:3896]) ? 1 : 0;
assign detect_max[486][19] = (mid_1[3903:3896] > btm_0[3911:3904]) ? 1 : 0;
assign detect_max[486][20] = (mid_1[3903:3896] > btm_1[3895:3888]) ? 1 : 0;
assign detect_max[486][21] = (mid_1[3903:3896] > btm_1[3903:3896]) ? 1 : 0;
assign detect_max[486][22] = (mid_1[3903:3896] > btm_1[3911:3904]) ? 1 : 0;
assign detect_max[486][23] = (mid_1[3903:3896] > btm_2[3895:3888]) ? 1 : 0;
assign detect_max[486][24] = (mid_1[3903:3896] > btm_2[3903:3896]) ? 1 : 0;
assign detect_max[486][25] = (mid_1[3903:3896] > btm_2[3911:3904]) ? 1 : 0;

assign detect_max[487][0] = (mid_1[3911:3904] > top_0[3903:3896]) ? 1 : 0;
assign detect_max[487][1] = (mid_1[3911:3904] > top_0[3911:3904]) ? 1 : 0;
assign detect_max[487][2] = (mid_1[3911:3904] > top_0[3919:3912]) ? 1 : 0;
assign detect_max[487][3] = (mid_1[3911:3904] > top_1[3903:3896]) ? 1 : 0;
assign detect_max[487][4] = (mid_1[3911:3904] > top_1[3911:3904]) ? 1 : 0;
assign detect_max[487][5] = (mid_1[3911:3904] > top_1[3919:3912]) ? 1 : 0;
assign detect_max[487][6] = (mid_1[3911:3904] > top_2[3903:3896]) ? 1 : 0;
assign detect_max[487][7] = (mid_1[3911:3904] > top_2[3911:3904]) ? 1 : 0;
assign detect_max[487][8] = (mid_1[3911:3904] > top_2[3919:3912]) ? 1 : 0;
assign detect_max[487][9] = (mid_1[3911:3904] > mid_0[3903:3896]) ? 1 : 0;
assign detect_max[487][10] = (mid_1[3911:3904] > mid_0[3911:3904]) ? 1 : 0;
assign detect_max[487][11] = (mid_1[3911:3904] > mid_0[3919:3912]) ? 1 : 0;
assign detect_max[487][12] = (mid_1[3911:3904] > mid_1[3903:3896]) ? 1 : 0;
assign detect_max[487][13] = (mid_1[3911:3904] > mid_1[3919:3912]) ? 1 : 0;
assign detect_max[487][14] = (mid_1[3911:3904] > mid_2[3903:3896]) ? 1 : 0;
assign detect_max[487][15] = (mid_1[3911:3904] > mid_2[3911:3904]) ? 1 : 0;
assign detect_max[487][16] = (mid_1[3911:3904] > mid_2[3919:3912]) ? 1 : 0;
assign detect_max[487][17] = (mid_1[3911:3904] > btm_0[3903:3896]) ? 1 : 0;
assign detect_max[487][18] = (mid_1[3911:3904] > btm_0[3911:3904]) ? 1 : 0;
assign detect_max[487][19] = (mid_1[3911:3904] > btm_0[3919:3912]) ? 1 : 0;
assign detect_max[487][20] = (mid_1[3911:3904] > btm_1[3903:3896]) ? 1 : 0;
assign detect_max[487][21] = (mid_1[3911:3904] > btm_1[3911:3904]) ? 1 : 0;
assign detect_max[487][22] = (mid_1[3911:3904] > btm_1[3919:3912]) ? 1 : 0;
assign detect_max[487][23] = (mid_1[3911:3904] > btm_2[3903:3896]) ? 1 : 0;
assign detect_max[487][24] = (mid_1[3911:3904] > btm_2[3911:3904]) ? 1 : 0;
assign detect_max[487][25] = (mid_1[3911:3904] > btm_2[3919:3912]) ? 1 : 0;

assign detect_max[488][0] = (mid_1[3919:3912] > top_0[3911:3904]) ? 1 : 0;
assign detect_max[488][1] = (mid_1[3919:3912] > top_0[3919:3912]) ? 1 : 0;
assign detect_max[488][2] = (mid_1[3919:3912] > top_0[3927:3920]) ? 1 : 0;
assign detect_max[488][3] = (mid_1[3919:3912] > top_1[3911:3904]) ? 1 : 0;
assign detect_max[488][4] = (mid_1[3919:3912] > top_1[3919:3912]) ? 1 : 0;
assign detect_max[488][5] = (mid_1[3919:3912] > top_1[3927:3920]) ? 1 : 0;
assign detect_max[488][6] = (mid_1[3919:3912] > top_2[3911:3904]) ? 1 : 0;
assign detect_max[488][7] = (mid_1[3919:3912] > top_2[3919:3912]) ? 1 : 0;
assign detect_max[488][8] = (mid_1[3919:3912] > top_2[3927:3920]) ? 1 : 0;
assign detect_max[488][9] = (mid_1[3919:3912] > mid_0[3911:3904]) ? 1 : 0;
assign detect_max[488][10] = (mid_1[3919:3912] > mid_0[3919:3912]) ? 1 : 0;
assign detect_max[488][11] = (mid_1[3919:3912] > mid_0[3927:3920]) ? 1 : 0;
assign detect_max[488][12] = (mid_1[3919:3912] > mid_1[3911:3904]) ? 1 : 0;
assign detect_max[488][13] = (mid_1[3919:3912] > mid_1[3927:3920]) ? 1 : 0;
assign detect_max[488][14] = (mid_1[3919:3912] > mid_2[3911:3904]) ? 1 : 0;
assign detect_max[488][15] = (mid_1[3919:3912] > mid_2[3919:3912]) ? 1 : 0;
assign detect_max[488][16] = (mid_1[3919:3912] > mid_2[3927:3920]) ? 1 : 0;
assign detect_max[488][17] = (mid_1[3919:3912] > btm_0[3911:3904]) ? 1 : 0;
assign detect_max[488][18] = (mid_1[3919:3912] > btm_0[3919:3912]) ? 1 : 0;
assign detect_max[488][19] = (mid_1[3919:3912] > btm_0[3927:3920]) ? 1 : 0;
assign detect_max[488][20] = (mid_1[3919:3912] > btm_1[3911:3904]) ? 1 : 0;
assign detect_max[488][21] = (mid_1[3919:3912] > btm_1[3919:3912]) ? 1 : 0;
assign detect_max[488][22] = (mid_1[3919:3912] > btm_1[3927:3920]) ? 1 : 0;
assign detect_max[488][23] = (mid_1[3919:3912] > btm_2[3911:3904]) ? 1 : 0;
assign detect_max[488][24] = (mid_1[3919:3912] > btm_2[3919:3912]) ? 1 : 0;
assign detect_max[488][25] = (mid_1[3919:3912] > btm_2[3927:3920]) ? 1 : 0;

assign detect_max[489][0] = (mid_1[3927:3920] > top_0[3919:3912]) ? 1 : 0;
assign detect_max[489][1] = (mid_1[3927:3920] > top_0[3927:3920]) ? 1 : 0;
assign detect_max[489][2] = (mid_1[3927:3920] > top_0[3935:3928]) ? 1 : 0;
assign detect_max[489][3] = (mid_1[3927:3920] > top_1[3919:3912]) ? 1 : 0;
assign detect_max[489][4] = (mid_1[3927:3920] > top_1[3927:3920]) ? 1 : 0;
assign detect_max[489][5] = (mid_1[3927:3920] > top_1[3935:3928]) ? 1 : 0;
assign detect_max[489][6] = (mid_1[3927:3920] > top_2[3919:3912]) ? 1 : 0;
assign detect_max[489][7] = (mid_1[3927:3920] > top_2[3927:3920]) ? 1 : 0;
assign detect_max[489][8] = (mid_1[3927:3920] > top_2[3935:3928]) ? 1 : 0;
assign detect_max[489][9] = (mid_1[3927:3920] > mid_0[3919:3912]) ? 1 : 0;
assign detect_max[489][10] = (mid_1[3927:3920] > mid_0[3927:3920]) ? 1 : 0;
assign detect_max[489][11] = (mid_1[3927:3920] > mid_0[3935:3928]) ? 1 : 0;
assign detect_max[489][12] = (mid_1[3927:3920] > mid_1[3919:3912]) ? 1 : 0;
assign detect_max[489][13] = (mid_1[3927:3920] > mid_1[3935:3928]) ? 1 : 0;
assign detect_max[489][14] = (mid_1[3927:3920] > mid_2[3919:3912]) ? 1 : 0;
assign detect_max[489][15] = (mid_1[3927:3920] > mid_2[3927:3920]) ? 1 : 0;
assign detect_max[489][16] = (mid_1[3927:3920] > mid_2[3935:3928]) ? 1 : 0;
assign detect_max[489][17] = (mid_1[3927:3920] > btm_0[3919:3912]) ? 1 : 0;
assign detect_max[489][18] = (mid_1[3927:3920] > btm_0[3927:3920]) ? 1 : 0;
assign detect_max[489][19] = (mid_1[3927:3920] > btm_0[3935:3928]) ? 1 : 0;
assign detect_max[489][20] = (mid_1[3927:3920] > btm_1[3919:3912]) ? 1 : 0;
assign detect_max[489][21] = (mid_1[3927:3920] > btm_1[3927:3920]) ? 1 : 0;
assign detect_max[489][22] = (mid_1[3927:3920] > btm_1[3935:3928]) ? 1 : 0;
assign detect_max[489][23] = (mid_1[3927:3920] > btm_2[3919:3912]) ? 1 : 0;
assign detect_max[489][24] = (mid_1[3927:3920] > btm_2[3927:3920]) ? 1 : 0;
assign detect_max[489][25] = (mid_1[3927:3920] > btm_2[3935:3928]) ? 1 : 0;

assign detect_max[490][0] = (mid_1[3935:3928] > top_0[3927:3920]) ? 1 : 0;
assign detect_max[490][1] = (mid_1[3935:3928] > top_0[3935:3928]) ? 1 : 0;
assign detect_max[490][2] = (mid_1[3935:3928] > top_0[3943:3936]) ? 1 : 0;
assign detect_max[490][3] = (mid_1[3935:3928] > top_1[3927:3920]) ? 1 : 0;
assign detect_max[490][4] = (mid_1[3935:3928] > top_1[3935:3928]) ? 1 : 0;
assign detect_max[490][5] = (mid_1[3935:3928] > top_1[3943:3936]) ? 1 : 0;
assign detect_max[490][6] = (mid_1[3935:3928] > top_2[3927:3920]) ? 1 : 0;
assign detect_max[490][7] = (mid_1[3935:3928] > top_2[3935:3928]) ? 1 : 0;
assign detect_max[490][8] = (mid_1[3935:3928] > top_2[3943:3936]) ? 1 : 0;
assign detect_max[490][9] = (mid_1[3935:3928] > mid_0[3927:3920]) ? 1 : 0;
assign detect_max[490][10] = (mid_1[3935:3928] > mid_0[3935:3928]) ? 1 : 0;
assign detect_max[490][11] = (mid_1[3935:3928] > mid_0[3943:3936]) ? 1 : 0;
assign detect_max[490][12] = (mid_1[3935:3928] > mid_1[3927:3920]) ? 1 : 0;
assign detect_max[490][13] = (mid_1[3935:3928] > mid_1[3943:3936]) ? 1 : 0;
assign detect_max[490][14] = (mid_1[3935:3928] > mid_2[3927:3920]) ? 1 : 0;
assign detect_max[490][15] = (mid_1[3935:3928] > mid_2[3935:3928]) ? 1 : 0;
assign detect_max[490][16] = (mid_1[3935:3928] > mid_2[3943:3936]) ? 1 : 0;
assign detect_max[490][17] = (mid_1[3935:3928] > btm_0[3927:3920]) ? 1 : 0;
assign detect_max[490][18] = (mid_1[3935:3928] > btm_0[3935:3928]) ? 1 : 0;
assign detect_max[490][19] = (mid_1[3935:3928] > btm_0[3943:3936]) ? 1 : 0;
assign detect_max[490][20] = (mid_1[3935:3928] > btm_1[3927:3920]) ? 1 : 0;
assign detect_max[490][21] = (mid_1[3935:3928] > btm_1[3935:3928]) ? 1 : 0;
assign detect_max[490][22] = (mid_1[3935:3928] > btm_1[3943:3936]) ? 1 : 0;
assign detect_max[490][23] = (mid_1[3935:3928] > btm_2[3927:3920]) ? 1 : 0;
assign detect_max[490][24] = (mid_1[3935:3928] > btm_2[3935:3928]) ? 1 : 0;
assign detect_max[490][25] = (mid_1[3935:3928] > btm_2[3943:3936]) ? 1 : 0;

assign detect_max[491][0] = (mid_1[3943:3936] > top_0[3935:3928]) ? 1 : 0;
assign detect_max[491][1] = (mid_1[3943:3936] > top_0[3943:3936]) ? 1 : 0;
assign detect_max[491][2] = (mid_1[3943:3936] > top_0[3951:3944]) ? 1 : 0;
assign detect_max[491][3] = (mid_1[3943:3936] > top_1[3935:3928]) ? 1 : 0;
assign detect_max[491][4] = (mid_1[3943:3936] > top_1[3943:3936]) ? 1 : 0;
assign detect_max[491][5] = (mid_1[3943:3936] > top_1[3951:3944]) ? 1 : 0;
assign detect_max[491][6] = (mid_1[3943:3936] > top_2[3935:3928]) ? 1 : 0;
assign detect_max[491][7] = (mid_1[3943:3936] > top_2[3943:3936]) ? 1 : 0;
assign detect_max[491][8] = (mid_1[3943:3936] > top_2[3951:3944]) ? 1 : 0;
assign detect_max[491][9] = (mid_1[3943:3936] > mid_0[3935:3928]) ? 1 : 0;
assign detect_max[491][10] = (mid_1[3943:3936] > mid_0[3943:3936]) ? 1 : 0;
assign detect_max[491][11] = (mid_1[3943:3936] > mid_0[3951:3944]) ? 1 : 0;
assign detect_max[491][12] = (mid_1[3943:3936] > mid_1[3935:3928]) ? 1 : 0;
assign detect_max[491][13] = (mid_1[3943:3936] > mid_1[3951:3944]) ? 1 : 0;
assign detect_max[491][14] = (mid_1[3943:3936] > mid_2[3935:3928]) ? 1 : 0;
assign detect_max[491][15] = (mid_1[3943:3936] > mid_2[3943:3936]) ? 1 : 0;
assign detect_max[491][16] = (mid_1[3943:3936] > mid_2[3951:3944]) ? 1 : 0;
assign detect_max[491][17] = (mid_1[3943:3936] > btm_0[3935:3928]) ? 1 : 0;
assign detect_max[491][18] = (mid_1[3943:3936] > btm_0[3943:3936]) ? 1 : 0;
assign detect_max[491][19] = (mid_1[3943:3936] > btm_0[3951:3944]) ? 1 : 0;
assign detect_max[491][20] = (mid_1[3943:3936] > btm_1[3935:3928]) ? 1 : 0;
assign detect_max[491][21] = (mid_1[3943:3936] > btm_1[3943:3936]) ? 1 : 0;
assign detect_max[491][22] = (mid_1[3943:3936] > btm_1[3951:3944]) ? 1 : 0;
assign detect_max[491][23] = (mid_1[3943:3936] > btm_2[3935:3928]) ? 1 : 0;
assign detect_max[491][24] = (mid_1[3943:3936] > btm_2[3943:3936]) ? 1 : 0;
assign detect_max[491][25] = (mid_1[3943:3936] > btm_2[3951:3944]) ? 1 : 0;

assign detect_max[492][0] = (mid_1[3951:3944] > top_0[3943:3936]) ? 1 : 0;
assign detect_max[492][1] = (mid_1[3951:3944] > top_0[3951:3944]) ? 1 : 0;
assign detect_max[492][2] = (mid_1[3951:3944] > top_0[3959:3952]) ? 1 : 0;
assign detect_max[492][3] = (mid_1[3951:3944] > top_1[3943:3936]) ? 1 : 0;
assign detect_max[492][4] = (mid_1[3951:3944] > top_1[3951:3944]) ? 1 : 0;
assign detect_max[492][5] = (mid_1[3951:3944] > top_1[3959:3952]) ? 1 : 0;
assign detect_max[492][6] = (mid_1[3951:3944] > top_2[3943:3936]) ? 1 : 0;
assign detect_max[492][7] = (mid_1[3951:3944] > top_2[3951:3944]) ? 1 : 0;
assign detect_max[492][8] = (mid_1[3951:3944] > top_2[3959:3952]) ? 1 : 0;
assign detect_max[492][9] = (mid_1[3951:3944] > mid_0[3943:3936]) ? 1 : 0;
assign detect_max[492][10] = (mid_1[3951:3944] > mid_0[3951:3944]) ? 1 : 0;
assign detect_max[492][11] = (mid_1[3951:3944] > mid_0[3959:3952]) ? 1 : 0;
assign detect_max[492][12] = (mid_1[3951:3944] > mid_1[3943:3936]) ? 1 : 0;
assign detect_max[492][13] = (mid_1[3951:3944] > mid_1[3959:3952]) ? 1 : 0;
assign detect_max[492][14] = (mid_1[3951:3944] > mid_2[3943:3936]) ? 1 : 0;
assign detect_max[492][15] = (mid_1[3951:3944] > mid_2[3951:3944]) ? 1 : 0;
assign detect_max[492][16] = (mid_1[3951:3944] > mid_2[3959:3952]) ? 1 : 0;
assign detect_max[492][17] = (mid_1[3951:3944] > btm_0[3943:3936]) ? 1 : 0;
assign detect_max[492][18] = (mid_1[3951:3944] > btm_0[3951:3944]) ? 1 : 0;
assign detect_max[492][19] = (mid_1[3951:3944] > btm_0[3959:3952]) ? 1 : 0;
assign detect_max[492][20] = (mid_1[3951:3944] > btm_1[3943:3936]) ? 1 : 0;
assign detect_max[492][21] = (mid_1[3951:3944] > btm_1[3951:3944]) ? 1 : 0;
assign detect_max[492][22] = (mid_1[3951:3944] > btm_1[3959:3952]) ? 1 : 0;
assign detect_max[492][23] = (mid_1[3951:3944] > btm_2[3943:3936]) ? 1 : 0;
assign detect_max[492][24] = (mid_1[3951:3944] > btm_2[3951:3944]) ? 1 : 0;
assign detect_max[492][25] = (mid_1[3951:3944] > btm_2[3959:3952]) ? 1 : 0;

assign detect_max[493][0] = (mid_1[3959:3952] > top_0[3951:3944]) ? 1 : 0;
assign detect_max[493][1] = (mid_1[3959:3952] > top_0[3959:3952]) ? 1 : 0;
assign detect_max[493][2] = (mid_1[3959:3952] > top_0[3967:3960]) ? 1 : 0;
assign detect_max[493][3] = (mid_1[3959:3952] > top_1[3951:3944]) ? 1 : 0;
assign detect_max[493][4] = (mid_1[3959:3952] > top_1[3959:3952]) ? 1 : 0;
assign detect_max[493][5] = (mid_1[3959:3952] > top_1[3967:3960]) ? 1 : 0;
assign detect_max[493][6] = (mid_1[3959:3952] > top_2[3951:3944]) ? 1 : 0;
assign detect_max[493][7] = (mid_1[3959:3952] > top_2[3959:3952]) ? 1 : 0;
assign detect_max[493][8] = (mid_1[3959:3952] > top_2[3967:3960]) ? 1 : 0;
assign detect_max[493][9] = (mid_1[3959:3952] > mid_0[3951:3944]) ? 1 : 0;
assign detect_max[493][10] = (mid_1[3959:3952] > mid_0[3959:3952]) ? 1 : 0;
assign detect_max[493][11] = (mid_1[3959:3952] > mid_0[3967:3960]) ? 1 : 0;
assign detect_max[493][12] = (mid_1[3959:3952] > mid_1[3951:3944]) ? 1 : 0;
assign detect_max[493][13] = (mid_1[3959:3952] > mid_1[3967:3960]) ? 1 : 0;
assign detect_max[493][14] = (mid_1[3959:3952] > mid_2[3951:3944]) ? 1 : 0;
assign detect_max[493][15] = (mid_1[3959:3952] > mid_2[3959:3952]) ? 1 : 0;
assign detect_max[493][16] = (mid_1[3959:3952] > mid_2[3967:3960]) ? 1 : 0;
assign detect_max[493][17] = (mid_1[3959:3952] > btm_0[3951:3944]) ? 1 : 0;
assign detect_max[493][18] = (mid_1[3959:3952] > btm_0[3959:3952]) ? 1 : 0;
assign detect_max[493][19] = (mid_1[3959:3952] > btm_0[3967:3960]) ? 1 : 0;
assign detect_max[493][20] = (mid_1[3959:3952] > btm_1[3951:3944]) ? 1 : 0;
assign detect_max[493][21] = (mid_1[3959:3952] > btm_1[3959:3952]) ? 1 : 0;
assign detect_max[493][22] = (mid_1[3959:3952] > btm_1[3967:3960]) ? 1 : 0;
assign detect_max[493][23] = (mid_1[3959:3952] > btm_2[3951:3944]) ? 1 : 0;
assign detect_max[493][24] = (mid_1[3959:3952] > btm_2[3959:3952]) ? 1 : 0;
assign detect_max[493][25] = (mid_1[3959:3952] > btm_2[3967:3960]) ? 1 : 0;

assign detect_max[494][0] = (mid_1[3967:3960] > top_0[3959:3952]) ? 1 : 0;
assign detect_max[494][1] = (mid_1[3967:3960] > top_0[3967:3960]) ? 1 : 0;
assign detect_max[494][2] = (mid_1[3967:3960] > top_0[3975:3968]) ? 1 : 0;
assign detect_max[494][3] = (mid_1[3967:3960] > top_1[3959:3952]) ? 1 : 0;
assign detect_max[494][4] = (mid_1[3967:3960] > top_1[3967:3960]) ? 1 : 0;
assign detect_max[494][5] = (mid_1[3967:3960] > top_1[3975:3968]) ? 1 : 0;
assign detect_max[494][6] = (mid_1[3967:3960] > top_2[3959:3952]) ? 1 : 0;
assign detect_max[494][7] = (mid_1[3967:3960] > top_2[3967:3960]) ? 1 : 0;
assign detect_max[494][8] = (mid_1[3967:3960] > top_2[3975:3968]) ? 1 : 0;
assign detect_max[494][9] = (mid_1[3967:3960] > mid_0[3959:3952]) ? 1 : 0;
assign detect_max[494][10] = (mid_1[3967:3960] > mid_0[3967:3960]) ? 1 : 0;
assign detect_max[494][11] = (mid_1[3967:3960] > mid_0[3975:3968]) ? 1 : 0;
assign detect_max[494][12] = (mid_1[3967:3960] > mid_1[3959:3952]) ? 1 : 0;
assign detect_max[494][13] = (mid_1[3967:3960] > mid_1[3975:3968]) ? 1 : 0;
assign detect_max[494][14] = (mid_1[3967:3960] > mid_2[3959:3952]) ? 1 : 0;
assign detect_max[494][15] = (mid_1[3967:3960] > mid_2[3967:3960]) ? 1 : 0;
assign detect_max[494][16] = (mid_1[3967:3960] > mid_2[3975:3968]) ? 1 : 0;
assign detect_max[494][17] = (mid_1[3967:3960] > btm_0[3959:3952]) ? 1 : 0;
assign detect_max[494][18] = (mid_1[3967:3960] > btm_0[3967:3960]) ? 1 : 0;
assign detect_max[494][19] = (mid_1[3967:3960] > btm_0[3975:3968]) ? 1 : 0;
assign detect_max[494][20] = (mid_1[3967:3960] > btm_1[3959:3952]) ? 1 : 0;
assign detect_max[494][21] = (mid_1[3967:3960] > btm_1[3967:3960]) ? 1 : 0;
assign detect_max[494][22] = (mid_1[3967:3960] > btm_1[3975:3968]) ? 1 : 0;
assign detect_max[494][23] = (mid_1[3967:3960] > btm_2[3959:3952]) ? 1 : 0;
assign detect_max[494][24] = (mid_1[3967:3960] > btm_2[3967:3960]) ? 1 : 0;
assign detect_max[494][25] = (mid_1[3967:3960] > btm_2[3975:3968]) ? 1 : 0;

assign detect_max[495][0] = (mid_1[3975:3968] > top_0[3967:3960]) ? 1 : 0;
assign detect_max[495][1] = (mid_1[3975:3968] > top_0[3975:3968]) ? 1 : 0;
assign detect_max[495][2] = (mid_1[3975:3968] > top_0[3983:3976]) ? 1 : 0;
assign detect_max[495][3] = (mid_1[3975:3968] > top_1[3967:3960]) ? 1 : 0;
assign detect_max[495][4] = (mid_1[3975:3968] > top_1[3975:3968]) ? 1 : 0;
assign detect_max[495][5] = (mid_1[3975:3968] > top_1[3983:3976]) ? 1 : 0;
assign detect_max[495][6] = (mid_1[3975:3968] > top_2[3967:3960]) ? 1 : 0;
assign detect_max[495][7] = (mid_1[3975:3968] > top_2[3975:3968]) ? 1 : 0;
assign detect_max[495][8] = (mid_1[3975:3968] > top_2[3983:3976]) ? 1 : 0;
assign detect_max[495][9] = (mid_1[3975:3968] > mid_0[3967:3960]) ? 1 : 0;
assign detect_max[495][10] = (mid_1[3975:3968] > mid_0[3975:3968]) ? 1 : 0;
assign detect_max[495][11] = (mid_1[3975:3968] > mid_0[3983:3976]) ? 1 : 0;
assign detect_max[495][12] = (mid_1[3975:3968] > mid_1[3967:3960]) ? 1 : 0;
assign detect_max[495][13] = (mid_1[3975:3968] > mid_1[3983:3976]) ? 1 : 0;
assign detect_max[495][14] = (mid_1[3975:3968] > mid_2[3967:3960]) ? 1 : 0;
assign detect_max[495][15] = (mid_1[3975:3968] > mid_2[3975:3968]) ? 1 : 0;
assign detect_max[495][16] = (mid_1[3975:3968] > mid_2[3983:3976]) ? 1 : 0;
assign detect_max[495][17] = (mid_1[3975:3968] > btm_0[3967:3960]) ? 1 : 0;
assign detect_max[495][18] = (mid_1[3975:3968] > btm_0[3975:3968]) ? 1 : 0;
assign detect_max[495][19] = (mid_1[3975:3968] > btm_0[3983:3976]) ? 1 : 0;
assign detect_max[495][20] = (mid_1[3975:3968] > btm_1[3967:3960]) ? 1 : 0;
assign detect_max[495][21] = (mid_1[3975:3968] > btm_1[3975:3968]) ? 1 : 0;
assign detect_max[495][22] = (mid_1[3975:3968] > btm_1[3983:3976]) ? 1 : 0;
assign detect_max[495][23] = (mid_1[3975:3968] > btm_2[3967:3960]) ? 1 : 0;
assign detect_max[495][24] = (mid_1[3975:3968] > btm_2[3975:3968]) ? 1 : 0;
assign detect_max[495][25] = (mid_1[3975:3968] > btm_2[3983:3976]) ? 1 : 0;

assign detect_max[496][0] = (mid_1[3983:3976] > top_0[3975:3968]) ? 1 : 0;
assign detect_max[496][1] = (mid_1[3983:3976] > top_0[3983:3976]) ? 1 : 0;
assign detect_max[496][2] = (mid_1[3983:3976] > top_0[3991:3984]) ? 1 : 0;
assign detect_max[496][3] = (mid_1[3983:3976] > top_1[3975:3968]) ? 1 : 0;
assign detect_max[496][4] = (mid_1[3983:3976] > top_1[3983:3976]) ? 1 : 0;
assign detect_max[496][5] = (mid_1[3983:3976] > top_1[3991:3984]) ? 1 : 0;
assign detect_max[496][6] = (mid_1[3983:3976] > top_2[3975:3968]) ? 1 : 0;
assign detect_max[496][7] = (mid_1[3983:3976] > top_2[3983:3976]) ? 1 : 0;
assign detect_max[496][8] = (mid_1[3983:3976] > top_2[3991:3984]) ? 1 : 0;
assign detect_max[496][9] = (mid_1[3983:3976] > mid_0[3975:3968]) ? 1 : 0;
assign detect_max[496][10] = (mid_1[3983:3976] > mid_0[3983:3976]) ? 1 : 0;
assign detect_max[496][11] = (mid_1[3983:3976] > mid_0[3991:3984]) ? 1 : 0;
assign detect_max[496][12] = (mid_1[3983:3976] > mid_1[3975:3968]) ? 1 : 0;
assign detect_max[496][13] = (mid_1[3983:3976] > mid_1[3991:3984]) ? 1 : 0;
assign detect_max[496][14] = (mid_1[3983:3976] > mid_2[3975:3968]) ? 1 : 0;
assign detect_max[496][15] = (mid_1[3983:3976] > mid_2[3983:3976]) ? 1 : 0;
assign detect_max[496][16] = (mid_1[3983:3976] > mid_2[3991:3984]) ? 1 : 0;
assign detect_max[496][17] = (mid_1[3983:3976] > btm_0[3975:3968]) ? 1 : 0;
assign detect_max[496][18] = (mid_1[3983:3976] > btm_0[3983:3976]) ? 1 : 0;
assign detect_max[496][19] = (mid_1[3983:3976] > btm_0[3991:3984]) ? 1 : 0;
assign detect_max[496][20] = (mid_1[3983:3976] > btm_1[3975:3968]) ? 1 : 0;
assign detect_max[496][21] = (mid_1[3983:3976] > btm_1[3983:3976]) ? 1 : 0;
assign detect_max[496][22] = (mid_1[3983:3976] > btm_1[3991:3984]) ? 1 : 0;
assign detect_max[496][23] = (mid_1[3983:3976] > btm_2[3975:3968]) ? 1 : 0;
assign detect_max[496][24] = (mid_1[3983:3976] > btm_2[3983:3976]) ? 1 : 0;
assign detect_max[496][25] = (mid_1[3983:3976] > btm_2[3991:3984]) ? 1 : 0;

assign detect_max[497][0] = (mid_1[3991:3984] > top_0[3983:3976]) ? 1 : 0;
assign detect_max[497][1] = (mid_1[3991:3984] > top_0[3991:3984]) ? 1 : 0;
assign detect_max[497][2] = (mid_1[3991:3984] > top_0[3999:3992]) ? 1 : 0;
assign detect_max[497][3] = (mid_1[3991:3984] > top_1[3983:3976]) ? 1 : 0;
assign detect_max[497][4] = (mid_1[3991:3984] > top_1[3991:3984]) ? 1 : 0;
assign detect_max[497][5] = (mid_1[3991:3984] > top_1[3999:3992]) ? 1 : 0;
assign detect_max[497][6] = (mid_1[3991:3984] > top_2[3983:3976]) ? 1 : 0;
assign detect_max[497][7] = (mid_1[3991:3984] > top_2[3991:3984]) ? 1 : 0;
assign detect_max[497][8] = (mid_1[3991:3984] > top_2[3999:3992]) ? 1 : 0;
assign detect_max[497][9] = (mid_1[3991:3984] > mid_0[3983:3976]) ? 1 : 0;
assign detect_max[497][10] = (mid_1[3991:3984] > mid_0[3991:3984]) ? 1 : 0;
assign detect_max[497][11] = (mid_1[3991:3984] > mid_0[3999:3992]) ? 1 : 0;
assign detect_max[497][12] = (mid_1[3991:3984] > mid_1[3983:3976]) ? 1 : 0;
assign detect_max[497][13] = (mid_1[3991:3984] > mid_1[3999:3992]) ? 1 : 0;
assign detect_max[497][14] = (mid_1[3991:3984] > mid_2[3983:3976]) ? 1 : 0;
assign detect_max[497][15] = (mid_1[3991:3984] > mid_2[3991:3984]) ? 1 : 0;
assign detect_max[497][16] = (mid_1[3991:3984] > mid_2[3999:3992]) ? 1 : 0;
assign detect_max[497][17] = (mid_1[3991:3984] > btm_0[3983:3976]) ? 1 : 0;
assign detect_max[497][18] = (mid_1[3991:3984] > btm_0[3991:3984]) ? 1 : 0;
assign detect_max[497][19] = (mid_1[3991:3984] > btm_0[3999:3992]) ? 1 : 0;
assign detect_max[497][20] = (mid_1[3991:3984] > btm_1[3983:3976]) ? 1 : 0;
assign detect_max[497][21] = (mid_1[3991:3984] > btm_1[3991:3984]) ? 1 : 0;
assign detect_max[497][22] = (mid_1[3991:3984] > btm_1[3999:3992]) ? 1 : 0;
assign detect_max[497][23] = (mid_1[3991:3984] > btm_2[3983:3976]) ? 1 : 0;
assign detect_max[497][24] = (mid_1[3991:3984] > btm_2[3991:3984]) ? 1 : 0;
assign detect_max[497][25] = (mid_1[3991:3984] > btm_2[3999:3992]) ? 1 : 0;

assign detect_max[498][0] = (mid_1[3999:3992] > top_0[3991:3984]) ? 1 : 0;
assign detect_max[498][1] = (mid_1[3999:3992] > top_0[3999:3992]) ? 1 : 0;
assign detect_max[498][2] = (mid_1[3999:3992] > top_0[4007:4000]) ? 1 : 0;
assign detect_max[498][3] = (mid_1[3999:3992] > top_1[3991:3984]) ? 1 : 0;
assign detect_max[498][4] = (mid_1[3999:3992] > top_1[3999:3992]) ? 1 : 0;
assign detect_max[498][5] = (mid_1[3999:3992] > top_1[4007:4000]) ? 1 : 0;
assign detect_max[498][6] = (mid_1[3999:3992] > top_2[3991:3984]) ? 1 : 0;
assign detect_max[498][7] = (mid_1[3999:3992] > top_2[3999:3992]) ? 1 : 0;
assign detect_max[498][8] = (mid_1[3999:3992] > top_2[4007:4000]) ? 1 : 0;
assign detect_max[498][9] = (mid_1[3999:3992] > mid_0[3991:3984]) ? 1 : 0;
assign detect_max[498][10] = (mid_1[3999:3992] > mid_0[3999:3992]) ? 1 : 0;
assign detect_max[498][11] = (mid_1[3999:3992] > mid_0[4007:4000]) ? 1 : 0;
assign detect_max[498][12] = (mid_1[3999:3992] > mid_1[3991:3984]) ? 1 : 0;
assign detect_max[498][13] = (mid_1[3999:3992] > mid_1[4007:4000]) ? 1 : 0;
assign detect_max[498][14] = (mid_1[3999:3992] > mid_2[3991:3984]) ? 1 : 0;
assign detect_max[498][15] = (mid_1[3999:3992] > mid_2[3999:3992]) ? 1 : 0;
assign detect_max[498][16] = (mid_1[3999:3992] > mid_2[4007:4000]) ? 1 : 0;
assign detect_max[498][17] = (mid_1[3999:3992] > btm_0[3991:3984]) ? 1 : 0;
assign detect_max[498][18] = (mid_1[3999:3992] > btm_0[3999:3992]) ? 1 : 0;
assign detect_max[498][19] = (mid_1[3999:3992] > btm_0[4007:4000]) ? 1 : 0;
assign detect_max[498][20] = (mid_1[3999:3992] > btm_1[3991:3984]) ? 1 : 0;
assign detect_max[498][21] = (mid_1[3999:3992] > btm_1[3999:3992]) ? 1 : 0;
assign detect_max[498][22] = (mid_1[3999:3992] > btm_1[4007:4000]) ? 1 : 0;
assign detect_max[498][23] = (mid_1[3999:3992] > btm_2[3991:3984]) ? 1 : 0;
assign detect_max[498][24] = (mid_1[3999:3992] > btm_2[3999:3992]) ? 1 : 0;
assign detect_max[498][25] = (mid_1[3999:3992] > btm_2[4007:4000]) ? 1 : 0;

assign detect_max[499][0] = (mid_1[4007:4000] > top_0[3999:3992]) ? 1 : 0;
assign detect_max[499][1] = (mid_1[4007:4000] > top_0[4007:4000]) ? 1 : 0;
assign detect_max[499][2] = (mid_1[4007:4000] > top_0[4015:4008]) ? 1 : 0;
assign detect_max[499][3] = (mid_1[4007:4000] > top_1[3999:3992]) ? 1 : 0;
assign detect_max[499][4] = (mid_1[4007:4000] > top_1[4007:4000]) ? 1 : 0;
assign detect_max[499][5] = (mid_1[4007:4000] > top_1[4015:4008]) ? 1 : 0;
assign detect_max[499][6] = (mid_1[4007:4000] > top_2[3999:3992]) ? 1 : 0;
assign detect_max[499][7] = (mid_1[4007:4000] > top_2[4007:4000]) ? 1 : 0;
assign detect_max[499][8] = (mid_1[4007:4000] > top_2[4015:4008]) ? 1 : 0;
assign detect_max[499][9] = (mid_1[4007:4000] > mid_0[3999:3992]) ? 1 : 0;
assign detect_max[499][10] = (mid_1[4007:4000] > mid_0[4007:4000]) ? 1 : 0;
assign detect_max[499][11] = (mid_1[4007:4000] > mid_0[4015:4008]) ? 1 : 0;
assign detect_max[499][12] = (mid_1[4007:4000] > mid_1[3999:3992]) ? 1 : 0;
assign detect_max[499][13] = (mid_1[4007:4000] > mid_1[4015:4008]) ? 1 : 0;
assign detect_max[499][14] = (mid_1[4007:4000] > mid_2[3999:3992]) ? 1 : 0;
assign detect_max[499][15] = (mid_1[4007:4000] > mid_2[4007:4000]) ? 1 : 0;
assign detect_max[499][16] = (mid_1[4007:4000] > mid_2[4015:4008]) ? 1 : 0;
assign detect_max[499][17] = (mid_1[4007:4000] > btm_0[3999:3992]) ? 1 : 0;
assign detect_max[499][18] = (mid_1[4007:4000] > btm_0[4007:4000]) ? 1 : 0;
assign detect_max[499][19] = (mid_1[4007:4000] > btm_0[4015:4008]) ? 1 : 0;
assign detect_max[499][20] = (mid_1[4007:4000] > btm_1[3999:3992]) ? 1 : 0;
assign detect_max[499][21] = (mid_1[4007:4000] > btm_1[4007:4000]) ? 1 : 0;
assign detect_max[499][22] = (mid_1[4007:4000] > btm_1[4015:4008]) ? 1 : 0;
assign detect_max[499][23] = (mid_1[4007:4000] > btm_2[3999:3992]) ? 1 : 0;
assign detect_max[499][24] = (mid_1[4007:4000] > btm_2[4007:4000]) ? 1 : 0;
assign detect_max[499][25] = (mid_1[4007:4000] > btm_2[4015:4008]) ? 1 : 0;

assign detect_max[500][0] = (mid_1[4015:4008] > top_0[4007:4000]) ? 1 : 0;
assign detect_max[500][1] = (mid_1[4015:4008] > top_0[4015:4008]) ? 1 : 0;
assign detect_max[500][2] = (mid_1[4015:4008] > top_0[4023:4016]) ? 1 : 0;
assign detect_max[500][3] = (mid_1[4015:4008] > top_1[4007:4000]) ? 1 : 0;
assign detect_max[500][4] = (mid_1[4015:4008] > top_1[4015:4008]) ? 1 : 0;
assign detect_max[500][5] = (mid_1[4015:4008] > top_1[4023:4016]) ? 1 : 0;
assign detect_max[500][6] = (mid_1[4015:4008] > top_2[4007:4000]) ? 1 : 0;
assign detect_max[500][7] = (mid_1[4015:4008] > top_2[4015:4008]) ? 1 : 0;
assign detect_max[500][8] = (mid_1[4015:4008] > top_2[4023:4016]) ? 1 : 0;
assign detect_max[500][9] = (mid_1[4015:4008] > mid_0[4007:4000]) ? 1 : 0;
assign detect_max[500][10] = (mid_1[4015:4008] > mid_0[4015:4008]) ? 1 : 0;
assign detect_max[500][11] = (mid_1[4015:4008] > mid_0[4023:4016]) ? 1 : 0;
assign detect_max[500][12] = (mid_1[4015:4008] > mid_1[4007:4000]) ? 1 : 0;
assign detect_max[500][13] = (mid_1[4015:4008] > mid_1[4023:4016]) ? 1 : 0;
assign detect_max[500][14] = (mid_1[4015:4008] > mid_2[4007:4000]) ? 1 : 0;
assign detect_max[500][15] = (mid_1[4015:4008] > mid_2[4015:4008]) ? 1 : 0;
assign detect_max[500][16] = (mid_1[4015:4008] > mid_2[4023:4016]) ? 1 : 0;
assign detect_max[500][17] = (mid_1[4015:4008] > btm_0[4007:4000]) ? 1 : 0;
assign detect_max[500][18] = (mid_1[4015:4008] > btm_0[4015:4008]) ? 1 : 0;
assign detect_max[500][19] = (mid_1[4015:4008] > btm_0[4023:4016]) ? 1 : 0;
assign detect_max[500][20] = (mid_1[4015:4008] > btm_1[4007:4000]) ? 1 : 0;
assign detect_max[500][21] = (mid_1[4015:4008] > btm_1[4015:4008]) ? 1 : 0;
assign detect_max[500][22] = (mid_1[4015:4008] > btm_1[4023:4016]) ? 1 : 0;
assign detect_max[500][23] = (mid_1[4015:4008] > btm_2[4007:4000]) ? 1 : 0;
assign detect_max[500][24] = (mid_1[4015:4008] > btm_2[4015:4008]) ? 1 : 0;
assign detect_max[500][25] = (mid_1[4015:4008] > btm_2[4023:4016]) ? 1 : 0;

assign detect_max[501][0] = (mid_1[4023:4016] > top_0[4015:4008]) ? 1 : 0;
assign detect_max[501][1] = (mid_1[4023:4016] > top_0[4023:4016]) ? 1 : 0;
assign detect_max[501][2] = (mid_1[4023:4016] > top_0[4031:4024]) ? 1 : 0;
assign detect_max[501][3] = (mid_1[4023:4016] > top_1[4015:4008]) ? 1 : 0;
assign detect_max[501][4] = (mid_1[4023:4016] > top_1[4023:4016]) ? 1 : 0;
assign detect_max[501][5] = (mid_1[4023:4016] > top_1[4031:4024]) ? 1 : 0;
assign detect_max[501][6] = (mid_1[4023:4016] > top_2[4015:4008]) ? 1 : 0;
assign detect_max[501][7] = (mid_1[4023:4016] > top_2[4023:4016]) ? 1 : 0;
assign detect_max[501][8] = (mid_1[4023:4016] > top_2[4031:4024]) ? 1 : 0;
assign detect_max[501][9] = (mid_1[4023:4016] > mid_0[4015:4008]) ? 1 : 0;
assign detect_max[501][10] = (mid_1[4023:4016] > mid_0[4023:4016]) ? 1 : 0;
assign detect_max[501][11] = (mid_1[4023:4016] > mid_0[4031:4024]) ? 1 : 0;
assign detect_max[501][12] = (mid_1[4023:4016] > mid_1[4015:4008]) ? 1 : 0;
assign detect_max[501][13] = (mid_1[4023:4016] > mid_1[4031:4024]) ? 1 : 0;
assign detect_max[501][14] = (mid_1[4023:4016] > mid_2[4015:4008]) ? 1 : 0;
assign detect_max[501][15] = (mid_1[4023:4016] > mid_2[4023:4016]) ? 1 : 0;
assign detect_max[501][16] = (mid_1[4023:4016] > mid_2[4031:4024]) ? 1 : 0;
assign detect_max[501][17] = (mid_1[4023:4016] > btm_0[4015:4008]) ? 1 : 0;
assign detect_max[501][18] = (mid_1[4023:4016] > btm_0[4023:4016]) ? 1 : 0;
assign detect_max[501][19] = (mid_1[4023:4016] > btm_0[4031:4024]) ? 1 : 0;
assign detect_max[501][20] = (mid_1[4023:4016] > btm_1[4015:4008]) ? 1 : 0;
assign detect_max[501][21] = (mid_1[4023:4016] > btm_1[4023:4016]) ? 1 : 0;
assign detect_max[501][22] = (mid_1[4023:4016] > btm_1[4031:4024]) ? 1 : 0;
assign detect_max[501][23] = (mid_1[4023:4016] > btm_2[4015:4008]) ? 1 : 0;
assign detect_max[501][24] = (mid_1[4023:4016] > btm_2[4023:4016]) ? 1 : 0;
assign detect_max[501][25] = (mid_1[4023:4016] > btm_2[4031:4024]) ? 1 : 0;

assign detect_max[502][0] = (mid_1[4031:4024] > top_0[4023:4016]) ? 1 : 0;
assign detect_max[502][1] = (mid_1[4031:4024] > top_0[4031:4024]) ? 1 : 0;
assign detect_max[502][2] = (mid_1[4031:4024] > top_0[4039:4032]) ? 1 : 0;
assign detect_max[502][3] = (mid_1[4031:4024] > top_1[4023:4016]) ? 1 : 0;
assign detect_max[502][4] = (mid_1[4031:4024] > top_1[4031:4024]) ? 1 : 0;
assign detect_max[502][5] = (mid_1[4031:4024] > top_1[4039:4032]) ? 1 : 0;
assign detect_max[502][6] = (mid_1[4031:4024] > top_2[4023:4016]) ? 1 : 0;
assign detect_max[502][7] = (mid_1[4031:4024] > top_2[4031:4024]) ? 1 : 0;
assign detect_max[502][8] = (mid_1[4031:4024] > top_2[4039:4032]) ? 1 : 0;
assign detect_max[502][9] = (mid_1[4031:4024] > mid_0[4023:4016]) ? 1 : 0;
assign detect_max[502][10] = (mid_1[4031:4024] > mid_0[4031:4024]) ? 1 : 0;
assign detect_max[502][11] = (mid_1[4031:4024] > mid_0[4039:4032]) ? 1 : 0;
assign detect_max[502][12] = (mid_1[4031:4024] > mid_1[4023:4016]) ? 1 : 0;
assign detect_max[502][13] = (mid_1[4031:4024] > mid_1[4039:4032]) ? 1 : 0;
assign detect_max[502][14] = (mid_1[4031:4024] > mid_2[4023:4016]) ? 1 : 0;
assign detect_max[502][15] = (mid_1[4031:4024] > mid_2[4031:4024]) ? 1 : 0;
assign detect_max[502][16] = (mid_1[4031:4024] > mid_2[4039:4032]) ? 1 : 0;
assign detect_max[502][17] = (mid_1[4031:4024] > btm_0[4023:4016]) ? 1 : 0;
assign detect_max[502][18] = (mid_1[4031:4024] > btm_0[4031:4024]) ? 1 : 0;
assign detect_max[502][19] = (mid_1[4031:4024] > btm_0[4039:4032]) ? 1 : 0;
assign detect_max[502][20] = (mid_1[4031:4024] > btm_1[4023:4016]) ? 1 : 0;
assign detect_max[502][21] = (mid_1[4031:4024] > btm_1[4031:4024]) ? 1 : 0;
assign detect_max[502][22] = (mid_1[4031:4024] > btm_1[4039:4032]) ? 1 : 0;
assign detect_max[502][23] = (mid_1[4031:4024] > btm_2[4023:4016]) ? 1 : 0;
assign detect_max[502][24] = (mid_1[4031:4024] > btm_2[4031:4024]) ? 1 : 0;
assign detect_max[502][25] = (mid_1[4031:4024] > btm_2[4039:4032]) ? 1 : 0;

assign detect_max[503][0] = (mid_1[4039:4032] > top_0[4031:4024]) ? 1 : 0;
assign detect_max[503][1] = (mid_1[4039:4032] > top_0[4039:4032]) ? 1 : 0;
assign detect_max[503][2] = (mid_1[4039:4032] > top_0[4047:4040]) ? 1 : 0;
assign detect_max[503][3] = (mid_1[4039:4032] > top_1[4031:4024]) ? 1 : 0;
assign detect_max[503][4] = (mid_1[4039:4032] > top_1[4039:4032]) ? 1 : 0;
assign detect_max[503][5] = (mid_1[4039:4032] > top_1[4047:4040]) ? 1 : 0;
assign detect_max[503][6] = (mid_1[4039:4032] > top_2[4031:4024]) ? 1 : 0;
assign detect_max[503][7] = (mid_1[4039:4032] > top_2[4039:4032]) ? 1 : 0;
assign detect_max[503][8] = (mid_1[4039:4032] > top_2[4047:4040]) ? 1 : 0;
assign detect_max[503][9] = (mid_1[4039:4032] > mid_0[4031:4024]) ? 1 : 0;
assign detect_max[503][10] = (mid_1[4039:4032] > mid_0[4039:4032]) ? 1 : 0;
assign detect_max[503][11] = (mid_1[4039:4032] > mid_0[4047:4040]) ? 1 : 0;
assign detect_max[503][12] = (mid_1[4039:4032] > mid_1[4031:4024]) ? 1 : 0;
assign detect_max[503][13] = (mid_1[4039:4032] > mid_1[4047:4040]) ? 1 : 0;
assign detect_max[503][14] = (mid_1[4039:4032] > mid_2[4031:4024]) ? 1 : 0;
assign detect_max[503][15] = (mid_1[4039:4032] > mid_2[4039:4032]) ? 1 : 0;
assign detect_max[503][16] = (mid_1[4039:4032] > mid_2[4047:4040]) ? 1 : 0;
assign detect_max[503][17] = (mid_1[4039:4032] > btm_0[4031:4024]) ? 1 : 0;
assign detect_max[503][18] = (mid_1[4039:4032] > btm_0[4039:4032]) ? 1 : 0;
assign detect_max[503][19] = (mid_1[4039:4032] > btm_0[4047:4040]) ? 1 : 0;
assign detect_max[503][20] = (mid_1[4039:4032] > btm_1[4031:4024]) ? 1 : 0;
assign detect_max[503][21] = (mid_1[4039:4032] > btm_1[4039:4032]) ? 1 : 0;
assign detect_max[503][22] = (mid_1[4039:4032] > btm_1[4047:4040]) ? 1 : 0;
assign detect_max[503][23] = (mid_1[4039:4032] > btm_2[4031:4024]) ? 1 : 0;
assign detect_max[503][24] = (mid_1[4039:4032] > btm_2[4039:4032]) ? 1 : 0;
assign detect_max[503][25] = (mid_1[4039:4032] > btm_2[4047:4040]) ? 1 : 0;

assign detect_max[504][0] = (mid_1[4047:4040] > top_0[4039:4032]) ? 1 : 0;
assign detect_max[504][1] = (mid_1[4047:4040] > top_0[4047:4040]) ? 1 : 0;
assign detect_max[504][2] = (mid_1[4047:4040] > top_0[4055:4048]) ? 1 : 0;
assign detect_max[504][3] = (mid_1[4047:4040] > top_1[4039:4032]) ? 1 : 0;
assign detect_max[504][4] = (mid_1[4047:4040] > top_1[4047:4040]) ? 1 : 0;
assign detect_max[504][5] = (mid_1[4047:4040] > top_1[4055:4048]) ? 1 : 0;
assign detect_max[504][6] = (mid_1[4047:4040] > top_2[4039:4032]) ? 1 : 0;
assign detect_max[504][7] = (mid_1[4047:4040] > top_2[4047:4040]) ? 1 : 0;
assign detect_max[504][8] = (mid_1[4047:4040] > top_2[4055:4048]) ? 1 : 0;
assign detect_max[504][9] = (mid_1[4047:4040] > mid_0[4039:4032]) ? 1 : 0;
assign detect_max[504][10] = (mid_1[4047:4040] > mid_0[4047:4040]) ? 1 : 0;
assign detect_max[504][11] = (mid_1[4047:4040] > mid_0[4055:4048]) ? 1 : 0;
assign detect_max[504][12] = (mid_1[4047:4040] > mid_1[4039:4032]) ? 1 : 0;
assign detect_max[504][13] = (mid_1[4047:4040] > mid_1[4055:4048]) ? 1 : 0;
assign detect_max[504][14] = (mid_1[4047:4040] > mid_2[4039:4032]) ? 1 : 0;
assign detect_max[504][15] = (mid_1[4047:4040] > mid_2[4047:4040]) ? 1 : 0;
assign detect_max[504][16] = (mid_1[4047:4040] > mid_2[4055:4048]) ? 1 : 0;
assign detect_max[504][17] = (mid_1[4047:4040] > btm_0[4039:4032]) ? 1 : 0;
assign detect_max[504][18] = (mid_1[4047:4040] > btm_0[4047:4040]) ? 1 : 0;
assign detect_max[504][19] = (mid_1[4047:4040] > btm_0[4055:4048]) ? 1 : 0;
assign detect_max[504][20] = (mid_1[4047:4040] > btm_1[4039:4032]) ? 1 : 0;
assign detect_max[504][21] = (mid_1[4047:4040] > btm_1[4047:4040]) ? 1 : 0;
assign detect_max[504][22] = (mid_1[4047:4040] > btm_1[4055:4048]) ? 1 : 0;
assign detect_max[504][23] = (mid_1[4047:4040] > btm_2[4039:4032]) ? 1 : 0;
assign detect_max[504][24] = (mid_1[4047:4040] > btm_2[4047:4040]) ? 1 : 0;
assign detect_max[504][25] = (mid_1[4047:4040] > btm_2[4055:4048]) ? 1 : 0;

assign detect_max[505][0] = (mid_1[4055:4048] > top_0[4047:4040]) ? 1 : 0;
assign detect_max[505][1] = (mid_1[4055:4048] > top_0[4055:4048]) ? 1 : 0;
assign detect_max[505][2] = (mid_1[4055:4048] > top_0[4063:4056]) ? 1 : 0;
assign detect_max[505][3] = (mid_1[4055:4048] > top_1[4047:4040]) ? 1 : 0;
assign detect_max[505][4] = (mid_1[4055:4048] > top_1[4055:4048]) ? 1 : 0;
assign detect_max[505][5] = (mid_1[4055:4048] > top_1[4063:4056]) ? 1 : 0;
assign detect_max[505][6] = (mid_1[4055:4048] > top_2[4047:4040]) ? 1 : 0;
assign detect_max[505][7] = (mid_1[4055:4048] > top_2[4055:4048]) ? 1 : 0;
assign detect_max[505][8] = (mid_1[4055:4048] > top_2[4063:4056]) ? 1 : 0;
assign detect_max[505][9] = (mid_1[4055:4048] > mid_0[4047:4040]) ? 1 : 0;
assign detect_max[505][10] = (mid_1[4055:4048] > mid_0[4055:4048]) ? 1 : 0;
assign detect_max[505][11] = (mid_1[4055:4048] > mid_0[4063:4056]) ? 1 : 0;
assign detect_max[505][12] = (mid_1[4055:4048] > mid_1[4047:4040]) ? 1 : 0;
assign detect_max[505][13] = (mid_1[4055:4048] > mid_1[4063:4056]) ? 1 : 0;
assign detect_max[505][14] = (mid_1[4055:4048] > mid_2[4047:4040]) ? 1 : 0;
assign detect_max[505][15] = (mid_1[4055:4048] > mid_2[4055:4048]) ? 1 : 0;
assign detect_max[505][16] = (mid_1[4055:4048] > mid_2[4063:4056]) ? 1 : 0;
assign detect_max[505][17] = (mid_1[4055:4048] > btm_0[4047:4040]) ? 1 : 0;
assign detect_max[505][18] = (mid_1[4055:4048] > btm_0[4055:4048]) ? 1 : 0;
assign detect_max[505][19] = (mid_1[4055:4048] > btm_0[4063:4056]) ? 1 : 0;
assign detect_max[505][20] = (mid_1[4055:4048] > btm_1[4047:4040]) ? 1 : 0;
assign detect_max[505][21] = (mid_1[4055:4048] > btm_1[4055:4048]) ? 1 : 0;
assign detect_max[505][22] = (mid_1[4055:4048] > btm_1[4063:4056]) ? 1 : 0;
assign detect_max[505][23] = (mid_1[4055:4048] > btm_2[4047:4040]) ? 1 : 0;
assign detect_max[505][24] = (mid_1[4055:4048] > btm_2[4055:4048]) ? 1 : 0;
assign detect_max[505][25] = (mid_1[4055:4048] > btm_2[4063:4056]) ? 1 : 0;

assign detect_max[506][0] = (mid_1[4063:4056] > top_0[4055:4048]) ? 1 : 0;
assign detect_max[506][1] = (mid_1[4063:4056] > top_0[4063:4056]) ? 1 : 0;
assign detect_max[506][2] = (mid_1[4063:4056] > top_0[4071:4064]) ? 1 : 0;
assign detect_max[506][3] = (mid_1[4063:4056] > top_1[4055:4048]) ? 1 : 0;
assign detect_max[506][4] = (mid_1[4063:4056] > top_1[4063:4056]) ? 1 : 0;
assign detect_max[506][5] = (mid_1[4063:4056] > top_1[4071:4064]) ? 1 : 0;
assign detect_max[506][6] = (mid_1[4063:4056] > top_2[4055:4048]) ? 1 : 0;
assign detect_max[506][7] = (mid_1[4063:4056] > top_2[4063:4056]) ? 1 : 0;
assign detect_max[506][8] = (mid_1[4063:4056] > top_2[4071:4064]) ? 1 : 0;
assign detect_max[506][9] = (mid_1[4063:4056] > mid_0[4055:4048]) ? 1 : 0;
assign detect_max[506][10] = (mid_1[4063:4056] > mid_0[4063:4056]) ? 1 : 0;
assign detect_max[506][11] = (mid_1[4063:4056] > mid_0[4071:4064]) ? 1 : 0;
assign detect_max[506][12] = (mid_1[4063:4056] > mid_1[4055:4048]) ? 1 : 0;
assign detect_max[506][13] = (mid_1[4063:4056] > mid_1[4071:4064]) ? 1 : 0;
assign detect_max[506][14] = (mid_1[4063:4056] > mid_2[4055:4048]) ? 1 : 0;
assign detect_max[506][15] = (mid_1[4063:4056] > mid_2[4063:4056]) ? 1 : 0;
assign detect_max[506][16] = (mid_1[4063:4056] > mid_2[4071:4064]) ? 1 : 0;
assign detect_max[506][17] = (mid_1[4063:4056] > btm_0[4055:4048]) ? 1 : 0;
assign detect_max[506][18] = (mid_1[4063:4056] > btm_0[4063:4056]) ? 1 : 0;
assign detect_max[506][19] = (mid_1[4063:4056] > btm_0[4071:4064]) ? 1 : 0;
assign detect_max[506][20] = (mid_1[4063:4056] > btm_1[4055:4048]) ? 1 : 0;
assign detect_max[506][21] = (mid_1[4063:4056] > btm_1[4063:4056]) ? 1 : 0;
assign detect_max[506][22] = (mid_1[4063:4056] > btm_1[4071:4064]) ? 1 : 0;
assign detect_max[506][23] = (mid_1[4063:4056] > btm_2[4055:4048]) ? 1 : 0;
assign detect_max[506][24] = (mid_1[4063:4056] > btm_2[4063:4056]) ? 1 : 0;
assign detect_max[506][25] = (mid_1[4063:4056] > btm_2[4071:4064]) ? 1 : 0;

assign detect_max[507][0] = (mid_1[4071:4064] > top_0[4063:4056]) ? 1 : 0;
assign detect_max[507][1] = (mid_1[4071:4064] > top_0[4071:4064]) ? 1 : 0;
assign detect_max[507][2] = (mid_1[4071:4064] > top_0[4079:4072]) ? 1 : 0;
assign detect_max[507][3] = (mid_1[4071:4064] > top_1[4063:4056]) ? 1 : 0;
assign detect_max[507][4] = (mid_1[4071:4064] > top_1[4071:4064]) ? 1 : 0;
assign detect_max[507][5] = (mid_1[4071:4064] > top_1[4079:4072]) ? 1 : 0;
assign detect_max[507][6] = (mid_1[4071:4064] > top_2[4063:4056]) ? 1 : 0;
assign detect_max[507][7] = (mid_1[4071:4064] > top_2[4071:4064]) ? 1 : 0;
assign detect_max[507][8] = (mid_1[4071:4064] > top_2[4079:4072]) ? 1 : 0;
assign detect_max[507][9] = (mid_1[4071:4064] > mid_0[4063:4056]) ? 1 : 0;
assign detect_max[507][10] = (mid_1[4071:4064] > mid_0[4071:4064]) ? 1 : 0;
assign detect_max[507][11] = (mid_1[4071:4064] > mid_0[4079:4072]) ? 1 : 0;
assign detect_max[507][12] = (mid_1[4071:4064] > mid_1[4063:4056]) ? 1 : 0;
assign detect_max[507][13] = (mid_1[4071:4064] > mid_1[4079:4072]) ? 1 : 0;
assign detect_max[507][14] = (mid_1[4071:4064] > mid_2[4063:4056]) ? 1 : 0;
assign detect_max[507][15] = (mid_1[4071:4064] > mid_2[4071:4064]) ? 1 : 0;
assign detect_max[507][16] = (mid_1[4071:4064] > mid_2[4079:4072]) ? 1 : 0;
assign detect_max[507][17] = (mid_1[4071:4064] > btm_0[4063:4056]) ? 1 : 0;
assign detect_max[507][18] = (mid_1[4071:4064] > btm_0[4071:4064]) ? 1 : 0;
assign detect_max[507][19] = (mid_1[4071:4064] > btm_0[4079:4072]) ? 1 : 0;
assign detect_max[507][20] = (mid_1[4071:4064] > btm_1[4063:4056]) ? 1 : 0;
assign detect_max[507][21] = (mid_1[4071:4064] > btm_1[4071:4064]) ? 1 : 0;
assign detect_max[507][22] = (mid_1[4071:4064] > btm_1[4079:4072]) ? 1 : 0;
assign detect_max[507][23] = (mid_1[4071:4064] > btm_2[4063:4056]) ? 1 : 0;
assign detect_max[507][24] = (mid_1[4071:4064] > btm_2[4071:4064]) ? 1 : 0;
assign detect_max[507][25] = (mid_1[4071:4064] > btm_2[4079:4072]) ? 1 : 0;

assign detect_max[508][0] = (mid_1[4079:4072] > top_0[4071:4064]) ? 1 : 0;
assign detect_max[508][1] = (mid_1[4079:4072] > top_0[4079:4072]) ? 1 : 0;
assign detect_max[508][2] = (mid_1[4079:4072] > top_0[4087:4080]) ? 1 : 0;
assign detect_max[508][3] = (mid_1[4079:4072] > top_1[4071:4064]) ? 1 : 0;
assign detect_max[508][4] = (mid_1[4079:4072] > top_1[4079:4072]) ? 1 : 0;
assign detect_max[508][5] = (mid_1[4079:4072] > top_1[4087:4080]) ? 1 : 0;
assign detect_max[508][6] = (mid_1[4079:4072] > top_2[4071:4064]) ? 1 : 0;
assign detect_max[508][7] = (mid_1[4079:4072] > top_2[4079:4072]) ? 1 : 0;
assign detect_max[508][8] = (mid_1[4079:4072] > top_2[4087:4080]) ? 1 : 0;
assign detect_max[508][9] = (mid_1[4079:4072] > mid_0[4071:4064]) ? 1 : 0;
assign detect_max[508][10] = (mid_1[4079:4072] > mid_0[4079:4072]) ? 1 : 0;
assign detect_max[508][11] = (mid_1[4079:4072] > mid_0[4087:4080]) ? 1 : 0;
assign detect_max[508][12] = (mid_1[4079:4072] > mid_1[4071:4064]) ? 1 : 0;
assign detect_max[508][13] = (mid_1[4079:4072] > mid_1[4087:4080]) ? 1 : 0;
assign detect_max[508][14] = (mid_1[4079:4072] > mid_2[4071:4064]) ? 1 : 0;
assign detect_max[508][15] = (mid_1[4079:4072] > mid_2[4079:4072]) ? 1 : 0;
assign detect_max[508][16] = (mid_1[4079:4072] > mid_2[4087:4080]) ? 1 : 0;
assign detect_max[508][17] = (mid_1[4079:4072] > btm_0[4071:4064]) ? 1 : 0;
assign detect_max[508][18] = (mid_1[4079:4072] > btm_0[4079:4072]) ? 1 : 0;
assign detect_max[508][19] = (mid_1[4079:4072] > btm_0[4087:4080]) ? 1 : 0;
assign detect_max[508][20] = (mid_1[4079:4072] > btm_1[4071:4064]) ? 1 : 0;
assign detect_max[508][21] = (mid_1[4079:4072] > btm_1[4079:4072]) ? 1 : 0;
assign detect_max[508][22] = (mid_1[4079:4072] > btm_1[4087:4080]) ? 1 : 0;
assign detect_max[508][23] = (mid_1[4079:4072] > btm_2[4071:4064]) ? 1 : 0;
assign detect_max[508][24] = (mid_1[4079:4072] > btm_2[4079:4072]) ? 1 : 0;
assign detect_max[508][25] = (mid_1[4079:4072] > btm_2[4087:4080]) ? 1 : 0;

assign detect_max[509][0] = (mid_1[4087:4080] > top_0[4079:4072]) ? 1 : 0;
assign detect_max[509][1] = (mid_1[4087:4080] > top_0[4087:4080]) ? 1 : 0;
assign detect_max[509][2] = (mid_1[4087:4080] > top_0[4095:4088]) ? 1 : 0;
assign detect_max[509][3] = (mid_1[4087:4080] > top_1[4079:4072]) ? 1 : 0;
assign detect_max[509][4] = (mid_1[4087:4080] > top_1[4087:4080]) ? 1 : 0;
assign detect_max[509][5] = (mid_1[4087:4080] > top_1[4095:4088]) ? 1 : 0;
assign detect_max[509][6] = (mid_1[4087:4080] > top_2[4079:4072]) ? 1 : 0;
assign detect_max[509][7] = (mid_1[4087:4080] > top_2[4087:4080]) ? 1 : 0;
assign detect_max[509][8] = (mid_1[4087:4080] > top_2[4095:4088]) ? 1 : 0;
assign detect_max[509][9] = (mid_1[4087:4080] > mid_0[4079:4072]) ? 1 : 0;
assign detect_max[509][10] = (mid_1[4087:4080] > mid_0[4087:4080]) ? 1 : 0;
assign detect_max[509][11] = (mid_1[4087:4080] > mid_0[4095:4088]) ? 1 : 0;
assign detect_max[509][12] = (mid_1[4087:4080] > mid_1[4079:4072]) ? 1 : 0;
assign detect_max[509][13] = (mid_1[4087:4080] > mid_1[4095:4088]) ? 1 : 0;
assign detect_max[509][14] = (mid_1[4087:4080] > mid_2[4079:4072]) ? 1 : 0;
assign detect_max[509][15] = (mid_1[4087:4080] > mid_2[4087:4080]) ? 1 : 0;
assign detect_max[509][16] = (mid_1[4087:4080] > mid_2[4095:4088]) ? 1 : 0;
assign detect_max[509][17] = (mid_1[4087:4080] > btm_0[4079:4072]) ? 1 : 0;
assign detect_max[509][18] = (mid_1[4087:4080] > btm_0[4087:4080]) ? 1 : 0;
assign detect_max[509][19] = (mid_1[4087:4080] > btm_0[4095:4088]) ? 1 : 0;
assign detect_max[509][20] = (mid_1[4087:4080] > btm_1[4079:4072]) ? 1 : 0;
assign detect_max[509][21] = (mid_1[4087:4080] > btm_1[4087:4080]) ? 1 : 0;
assign detect_max[509][22] = (mid_1[4087:4080] > btm_1[4095:4088]) ? 1 : 0;
assign detect_max[509][23] = (mid_1[4087:4080] > btm_2[4079:4072]) ? 1 : 0;
assign detect_max[509][24] = (mid_1[4087:4080] > btm_2[4087:4080]) ? 1 : 0;
assign detect_max[509][25] = (mid_1[4087:4080] > btm_2[4095:4088]) ? 1 : 0;

assign detect_max[510][0] = (mid_1[4095:4088] > top_0[4087:4080]) ? 1 : 0;
assign detect_max[510][1] = (mid_1[4095:4088] > top_0[4095:4088]) ? 1 : 0;
assign detect_max[510][2] = (mid_1[4095:4088] > top_0[4103:4096]) ? 1 : 0;
assign detect_max[510][3] = (mid_1[4095:4088] > top_1[4087:4080]) ? 1 : 0;
assign detect_max[510][4] = (mid_1[4095:4088] > top_1[4095:4088]) ? 1 : 0;
assign detect_max[510][5] = (mid_1[4095:4088] > top_1[4103:4096]) ? 1 : 0;
assign detect_max[510][6] = (mid_1[4095:4088] > top_2[4087:4080]) ? 1 : 0;
assign detect_max[510][7] = (mid_1[4095:4088] > top_2[4095:4088]) ? 1 : 0;
assign detect_max[510][8] = (mid_1[4095:4088] > top_2[4103:4096]) ? 1 : 0;
assign detect_max[510][9] = (mid_1[4095:4088] > mid_0[4087:4080]) ? 1 : 0;
assign detect_max[510][10] = (mid_1[4095:4088] > mid_0[4095:4088]) ? 1 : 0;
assign detect_max[510][11] = (mid_1[4095:4088] > mid_0[4103:4096]) ? 1 : 0;
assign detect_max[510][12] = (mid_1[4095:4088] > mid_1[4087:4080]) ? 1 : 0;
assign detect_max[510][13] = (mid_1[4095:4088] > mid_1[4103:4096]) ? 1 : 0;
assign detect_max[510][14] = (mid_1[4095:4088] > mid_2[4087:4080]) ? 1 : 0;
assign detect_max[510][15] = (mid_1[4095:4088] > mid_2[4095:4088]) ? 1 : 0;
assign detect_max[510][16] = (mid_1[4095:4088] > mid_2[4103:4096]) ? 1 : 0;
assign detect_max[510][17] = (mid_1[4095:4088] > btm_0[4087:4080]) ? 1 : 0;
assign detect_max[510][18] = (mid_1[4095:4088] > btm_0[4095:4088]) ? 1 : 0;
assign detect_max[510][19] = (mid_1[4095:4088] > btm_0[4103:4096]) ? 1 : 0;
assign detect_max[510][20] = (mid_1[4095:4088] > btm_1[4087:4080]) ? 1 : 0;
assign detect_max[510][21] = (mid_1[4095:4088] > btm_1[4095:4088]) ? 1 : 0;
assign detect_max[510][22] = (mid_1[4095:4088] > btm_1[4103:4096]) ? 1 : 0;
assign detect_max[510][23] = (mid_1[4095:4088] > btm_2[4087:4080]) ? 1 : 0;
assign detect_max[510][24] = (mid_1[4095:4088] > btm_2[4095:4088]) ? 1 : 0;
assign detect_max[510][25] = (mid_1[4095:4088] > btm_2[4103:4096]) ? 1 : 0;

assign detect_max[511][0] = (mid_1[4103:4096] > top_0[4095:4088]) ? 1 : 0;
assign detect_max[511][1] = (mid_1[4103:4096] > top_0[4103:4096]) ? 1 : 0;
assign detect_max[511][2] = (mid_1[4103:4096] > top_0[4111:4104]) ? 1 : 0;
assign detect_max[511][3] = (mid_1[4103:4096] > top_1[4095:4088]) ? 1 : 0;
assign detect_max[511][4] = (mid_1[4103:4096] > top_1[4103:4096]) ? 1 : 0;
assign detect_max[511][5] = (mid_1[4103:4096] > top_1[4111:4104]) ? 1 : 0;
assign detect_max[511][6] = (mid_1[4103:4096] > top_2[4095:4088]) ? 1 : 0;
assign detect_max[511][7] = (mid_1[4103:4096] > top_2[4103:4096]) ? 1 : 0;
assign detect_max[511][8] = (mid_1[4103:4096] > top_2[4111:4104]) ? 1 : 0;
assign detect_max[511][9] = (mid_1[4103:4096] > mid_0[4095:4088]) ? 1 : 0;
assign detect_max[511][10] = (mid_1[4103:4096] > mid_0[4103:4096]) ? 1 : 0;
assign detect_max[511][11] = (mid_1[4103:4096] > mid_0[4111:4104]) ? 1 : 0;
assign detect_max[511][12] = (mid_1[4103:4096] > mid_1[4095:4088]) ? 1 : 0;
assign detect_max[511][13] = (mid_1[4103:4096] > mid_1[4111:4104]) ? 1 : 0;
assign detect_max[511][14] = (mid_1[4103:4096] > mid_2[4095:4088]) ? 1 : 0;
assign detect_max[511][15] = (mid_1[4103:4096] > mid_2[4103:4096]) ? 1 : 0;
assign detect_max[511][16] = (mid_1[4103:4096] > mid_2[4111:4104]) ? 1 : 0;
assign detect_max[511][17] = (mid_1[4103:4096] > btm_0[4095:4088]) ? 1 : 0;
assign detect_max[511][18] = (mid_1[4103:4096] > btm_0[4103:4096]) ? 1 : 0;
assign detect_max[511][19] = (mid_1[4103:4096] > btm_0[4111:4104]) ? 1 : 0;
assign detect_max[511][20] = (mid_1[4103:4096] > btm_1[4095:4088]) ? 1 : 0;
assign detect_max[511][21] = (mid_1[4103:4096] > btm_1[4103:4096]) ? 1 : 0;
assign detect_max[511][22] = (mid_1[4103:4096] > btm_1[4111:4104]) ? 1 : 0;
assign detect_max[511][23] = (mid_1[4103:4096] > btm_2[4095:4088]) ? 1 : 0;
assign detect_max[511][24] = (mid_1[4103:4096] > btm_2[4103:4096]) ? 1 : 0;
assign detect_max[511][25] = (mid_1[4103:4096] > btm_2[4111:4104]) ? 1 : 0;

assign detect_max[512][0] = (mid_1[4111:4104] > top_0[4103:4096]) ? 1 : 0;
assign detect_max[512][1] = (mid_1[4111:4104] > top_0[4111:4104]) ? 1 : 0;
assign detect_max[512][2] = (mid_1[4111:4104] > top_0[4119:4112]) ? 1 : 0;
assign detect_max[512][3] = (mid_1[4111:4104] > top_1[4103:4096]) ? 1 : 0;
assign detect_max[512][4] = (mid_1[4111:4104] > top_1[4111:4104]) ? 1 : 0;
assign detect_max[512][5] = (mid_1[4111:4104] > top_1[4119:4112]) ? 1 : 0;
assign detect_max[512][6] = (mid_1[4111:4104] > top_2[4103:4096]) ? 1 : 0;
assign detect_max[512][7] = (mid_1[4111:4104] > top_2[4111:4104]) ? 1 : 0;
assign detect_max[512][8] = (mid_1[4111:4104] > top_2[4119:4112]) ? 1 : 0;
assign detect_max[512][9] = (mid_1[4111:4104] > mid_0[4103:4096]) ? 1 : 0;
assign detect_max[512][10] = (mid_1[4111:4104] > mid_0[4111:4104]) ? 1 : 0;
assign detect_max[512][11] = (mid_1[4111:4104] > mid_0[4119:4112]) ? 1 : 0;
assign detect_max[512][12] = (mid_1[4111:4104] > mid_1[4103:4096]) ? 1 : 0;
assign detect_max[512][13] = (mid_1[4111:4104] > mid_1[4119:4112]) ? 1 : 0;
assign detect_max[512][14] = (mid_1[4111:4104] > mid_2[4103:4096]) ? 1 : 0;
assign detect_max[512][15] = (mid_1[4111:4104] > mid_2[4111:4104]) ? 1 : 0;
assign detect_max[512][16] = (mid_1[4111:4104] > mid_2[4119:4112]) ? 1 : 0;
assign detect_max[512][17] = (mid_1[4111:4104] > btm_0[4103:4096]) ? 1 : 0;
assign detect_max[512][18] = (mid_1[4111:4104] > btm_0[4111:4104]) ? 1 : 0;
assign detect_max[512][19] = (mid_1[4111:4104] > btm_0[4119:4112]) ? 1 : 0;
assign detect_max[512][20] = (mid_1[4111:4104] > btm_1[4103:4096]) ? 1 : 0;
assign detect_max[512][21] = (mid_1[4111:4104] > btm_1[4111:4104]) ? 1 : 0;
assign detect_max[512][22] = (mid_1[4111:4104] > btm_1[4119:4112]) ? 1 : 0;
assign detect_max[512][23] = (mid_1[4111:4104] > btm_2[4103:4096]) ? 1 : 0;
assign detect_max[512][24] = (mid_1[4111:4104] > btm_2[4111:4104]) ? 1 : 0;
assign detect_max[512][25] = (mid_1[4111:4104] > btm_2[4119:4112]) ? 1 : 0;

assign detect_max[513][0] = (mid_1[4119:4112] > top_0[4111:4104]) ? 1 : 0;
assign detect_max[513][1] = (mid_1[4119:4112] > top_0[4119:4112]) ? 1 : 0;
assign detect_max[513][2] = (mid_1[4119:4112] > top_0[4127:4120]) ? 1 : 0;
assign detect_max[513][3] = (mid_1[4119:4112] > top_1[4111:4104]) ? 1 : 0;
assign detect_max[513][4] = (mid_1[4119:4112] > top_1[4119:4112]) ? 1 : 0;
assign detect_max[513][5] = (mid_1[4119:4112] > top_1[4127:4120]) ? 1 : 0;
assign detect_max[513][6] = (mid_1[4119:4112] > top_2[4111:4104]) ? 1 : 0;
assign detect_max[513][7] = (mid_1[4119:4112] > top_2[4119:4112]) ? 1 : 0;
assign detect_max[513][8] = (mid_1[4119:4112] > top_2[4127:4120]) ? 1 : 0;
assign detect_max[513][9] = (mid_1[4119:4112] > mid_0[4111:4104]) ? 1 : 0;
assign detect_max[513][10] = (mid_1[4119:4112] > mid_0[4119:4112]) ? 1 : 0;
assign detect_max[513][11] = (mid_1[4119:4112] > mid_0[4127:4120]) ? 1 : 0;
assign detect_max[513][12] = (mid_1[4119:4112] > mid_1[4111:4104]) ? 1 : 0;
assign detect_max[513][13] = (mid_1[4119:4112] > mid_1[4127:4120]) ? 1 : 0;
assign detect_max[513][14] = (mid_1[4119:4112] > mid_2[4111:4104]) ? 1 : 0;
assign detect_max[513][15] = (mid_1[4119:4112] > mid_2[4119:4112]) ? 1 : 0;
assign detect_max[513][16] = (mid_1[4119:4112] > mid_2[4127:4120]) ? 1 : 0;
assign detect_max[513][17] = (mid_1[4119:4112] > btm_0[4111:4104]) ? 1 : 0;
assign detect_max[513][18] = (mid_1[4119:4112] > btm_0[4119:4112]) ? 1 : 0;
assign detect_max[513][19] = (mid_1[4119:4112] > btm_0[4127:4120]) ? 1 : 0;
assign detect_max[513][20] = (mid_1[4119:4112] > btm_1[4111:4104]) ? 1 : 0;
assign detect_max[513][21] = (mid_1[4119:4112] > btm_1[4119:4112]) ? 1 : 0;
assign detect_max[513][22] = (mid_1[4119:4112] > btm_1[4127:4120]) ? 1 : 0;
assign detect_max[513][23] = (mid_1[4119:4112] > btm_2[4111:4104]) ? 1 : 0;
assign detect_max[513][24] = (mid_1[4119:4112] > btm_2[4119:4112]) ? 1 : 0;
assign detect_max[513][25] = (mid_1[4119:4112] > btm_2[4127:4120]) ? 1 : 0;

assign detect_max[514][0] = (mid_1[4127:4120] > top_0[4119:4112]) ? 1 : 0;
assign detect_max[514][1] = (mid_1[4127:4120] > top_0[4127:4120]) ? 1 : 0;
assign detect_max[514][2] = (mid_1[4127:4120] > top_0[4135:4128]) ? 1 : 0;
assign detect_max[514][3] = (mid_1[4127:4120] > top_1[4119:4112]) ? 1 : 0;
assign detect_max[514][4] = (mid_1[4127:4120] > top_1[4127:4120]) ? 1 : 0;
assign detect_max[514][5] = (mid_1[4127:4120] > top_1[4135:4128]) ? 1 : 0;
assign detect_max[514][6] = (mid_1[4127:4120] > top_2[4119:4112]) ? 1 : 0;
assign detect_max[514][7] = (mid_1[4127:4120] > top_2[4127:4120]) ? 1 : 0;
assign detect_max[514][8] = (mid_1[4127:4120] > top_2[4135:4128]) ? 1 : 0;
assign detect_max[514][9] = (mid_1[4127:4120] > mid_0[4119:4112]) ? 1 : 0;
assign detect_max[514][10] = (mid_1[4127:4120] > mid_0[4127:4120]) ? 1 : 0;
assign detect_max[514][11] = (mid_1[4127:4120] > mid_0[4135:4128]) ? 1 : 0;
assign detect_max[514][12] = (mid_1[4127:4120] > mid_1[4119:4112]) ? 1 : 0;
assign detect_max[514][13] = (mid_1[4127:4120] > mid_1[4135:4128]) ? 1 : 0;
assign detect_max[514][14] = (mid_1[4127:4120] > mid_2[4119:4112]) ? 1 : 0;
assign detect_max[514][15] = (mid_1[4127:4120] > mid_2[4127:4120]) ? 1 : 0;
assign detect_max[514][16] = (mid_1[4127:4120] > mid_2[4135:4128]) ? 1 : 0;
assign detect_max[514][17] = (mid_1[4127:4120] > btm_0[4119:4112]) ? 1 : 0;
assign detect_max[514][18] = (mid_1[4127:4120] > btm_0[4127:4120]) ? 1 : 0;
assign detect_max[514][19] = (mid_1[4127:4120] > btm_0[4135:4128]) ? 1 : 0;
assign detect_max[514][20] = (mid_1[4127:4120] > btm_1[4119:4112]) ? 1 : 0;
assign detect_max[514][21] = (mid_1[4127:4120] > btm_1[4127:4120]) ? 1 : 0;
assign detect_max[514][22] = (mid_1[4127:4120] > btm_1[4135:4128]) ? 1 : 0;
assign detect_max[514][23] = (mid_1[4127:4120] > btm_2[4119:4112]) ? 1 : 0;
assign detect_max[514][24] = (mid_1[4127:4120] > btm_2[4127:4120]) ? 1 : 0;
assign detect_max[514][25] = (mid_1[4127:4120] > btm_2[4135:4128]) ? 1 : 0;

assign detect_max[515][0] = (mid_1[4135:4128] > top_0[4127:4120]) ? 1 : 0;
assign detect_max[515][1] = (mid_1[4135:4128] > top_0[4135:4128]) ? 1 : 0;
assign detect_max[515][2] = (mid_1[4135:4128] > top_0[4143:4136]) ? 1 : 0;
assign detect_max[515][3] = (mid_1[4135:4128] > top_1[4127:4120]) ? 1 : 0;
assign detect_max[515][4] = (mid_1[4135:4128] > top_1[4135:4128]) ? 1 : 0;
assign detect_max[515][5] = (mid_1[4135:4128] > top_1[4143:4136]) ? 1 : 0;
assign detect_max[515][6] = (mid_1[4135:4128] > top_2[4127:4120]) ? 1 : 0;
assign detect_max[515][7] = (mid_1[4135:4128] > top_2[4135:4128]) ? 1 : 0;
assign detect_max[515][8] = (mid_1[4135:4128] > top_2[4143:4136]) ? 1 : 0;
assign detect_max[515][9] = (mid_1[4135:4128] > mid_0[4127:4120]) ? 1 : 0;
assign detect_max[515][10] = (mid_1[4135:4128] > mid_0[4135:4128]) ? 1 : 0;
assign detect_max[515][11] = (mid_1[4135:4128] > mid_0[4143:4136]) ? 1 : 0;
assign detect_max[515][12] = (mid_1[4135:4128] > mid_1[4127:4120]) ? 1 : 0;
assign detect_max[515][13] = (mid_1[4135:4128] > mid_1[4143:4136]) ? 1 : 0;
assign detect_max[515][14] = (mid_1[4135:4128] > mid_2[4127:4120]) ? 1 : 0;
assign detect_max[515][15] = (mid_1[4135:4128] > mid_2[4135:4128]) ? 1 : 0;
assign detect_max[515][16] = (mid_1[4135:4128] > mid_2[4143:4136]) ? 1 : 0;
assign detect_max[515][17] = (mid_1[4135:4128] > btm_0[4127:4120]) ? 1 : 0;
assign detect_max[515][18] = (mid_1[4135:4128] > btm_0[4135:4128]) ? 1 : 0;
assign detect_max[515][19] = (mid_1[4135:4128] > btm_0[4143:4136]) ? 1 : 0;
assign detect_max[515][20] = (mid_1[4135:4128] > btm_1[4127:4120]) ? 1 : 0;
assign detect_max[515][21] = (mid_1[4135:4128] > btm_1[4135:4128]) ? 1 : 0;
assign detect_max[515][22] = (mid_1[4135:4128] > btm_1[4143:4136]) ? 1 : 0;
assign detect_max[515][23] = (mid_1[4135:4128] > btm_2[4127:4120]) ? 1 : 0;
assign detect_max[515][24] = (mid_1[4135:4128] > btm_2[4135:4128]) ? 1 : 0;
assign detect_max[515][25] = (mid_1[4135:4128] > btm_2[4143:4136]) ? 1 : 0;

assign detect_max[516][0] = (mid_1[4143:4136] > top_0[4135:4128]) ? 1 : 0;
assign detect_max[516][1] = (mid_1[4143:4136] > top_0[4143:4136]) ? 1 : 0;
assign detect_max[516][2] = (mid_1[4143:4136] > top_0[4151:4144]) ? 1 : 0;
assign detect_max[516][3] = (mid_1[4143:4136] > top_1[4135:4128]) ? 1 : 0;
assign detect_max[516][4] = (mid_1[4143:4136] > top_1[4143:4136]) ? 1 : 0;
assign detect_max[516][5] = (mid_1[4143:4136] > top_1[4151:4144]) ? 1 : 0;
assign detect_max[516][6] = (mid_1[4143:4136] > top_2[4135:4128]) ? 1 : 0;
assign detect_max[516][7] = (mid_1[4143:4136] > top_2[4143:4136]) ? 1 : 0;
assign detect_max[516][8] = (mid_1[4143:4136] > top_2[4151:4144]) ? 1 : 0;
assign detect_max[516][9] = (mid_1[4143:4136] > mid_0[4135:4128]) ? 1 : 0;
assign detect_max[516][10] = (mid_1[4143:4136] > mid_0[4143:4136]) ? 1 : 0;
assign detect_max[516][11] = (mid_1[4143:4136] > mid_0[4151:4144]) ? 1 : 0;
assign detect_max[516][12] = (mid_1[4143:4136] > mid_1[4135:4128]) ? 1 : 0;
assign detect_max[516][13] = (mid_1[4143:4136] > mid_1[4151:4144]) ? 1 : 0;
assign detect_max[516][14] = (mid_1[4143:4136] > mid_2[4135:4128]) ? 1 : 0;
assign detect_max[516][15] = (mid_1[4143:4136] > mid_2[4143:4136]) ? 1 : 0;
assign detect_max[516][16] = (mid_1[4143:4136] > mid_2[4151:4144]) ? 1 : 0;
assign detect_max[516][17] = (mid_1[4143:4136] > btm_0[4135:4128]) ? 1 : 0;
assign detect_max[516][18] = (mid_1[4143:4136] > btm_0[4143:4136]) ? 1 : 0;
assign detect_max[516][19] = (mid_1[4143:4136] > btm_0[4151:4144]) ? 1 : 0;
assign detect_max[516][20] = (mid_1[4143:4136] > btm_1[4135:4128]) ? 1 : 0;
assign detect_max[516][21] = (mid_1[4143:4136] > btm_1[4143:4136]) ? 1 : 0;
assign detect_max[516][22] = (mid_1[4143:4136] > btm_1[4151:4144]) ? 1 : 0;
assign detect_max[516][23] = (mid_1[4143:4136] > btm_2[4135:4128]) ? 1 : 0;
assign detect_max[516][24] = (mid_1[4143:4136] > btm_2[4143:4136]) ? 1 : 0;
assign detect_max[516][25] = (mid_1[4143:4136] > btm_2[4151:4144]) ? 1 : 0;

assign detect_max[517][0] = (mid_1[4151:4144] > top_0[4143:4136]) ? 1 : 0;
assign detect_max[517][1] = (mid_1[4151:4144] > top_0[4151:4144]) ? 1 : 0;
assign detect_max[517][2] = (mid_1[4151:4144] > top_0[4159:4152]) ? 1 : 0;
assign detect_max[517][3] = (mid_1[4151:4144] > top_1[4143:4136]) ? 1 : 0;
assign detect_max[517][4] = (mid_1[4151:4144] > top_1[4151:4144]) ? 1 : 0;
assign detect_max[517][5] = (mid_1[4151:4144] > top_1[4159:4152]) ? 1 : 0;
assign detect_max[517][6] = (mid_1[4151:4144] > top_2[4143:4136]) ? 1 : 0;
assign detect_max[517][7] = (mid_1[4151:4144] > top_2[4151:4144]) ? 1 : 0;
assign detect_max[517][8] = (mid_1[4151:4144] > top_2[4159:4152]) ? 1 : 0;
assign detect_max[517][9] = (mid_1[4151:4144] > mid_0[4143:4136]) ? 1 : 0;
assign detect_max[517][10] = (mid_1[4151:4144] > mid_0[4151:4144]) ? 1 : 0;
assign detect_max[517][11] = (mid_1[4151:4144] > mid_0[4159:4152]) ? 1 : 0;
assign detect_max[517][12] = (mid_1[4151:4144] > mid_1[4143:4136]) ? 1 : 0;
assign detect_max[517][13] = (mid_1[4151:4144] > mid_1[4159:4152]) ? 1 : 0;
assign detect_max[517][14] = (mid_1[4151:4144] > mid_2[4143:4136]) ? 1 : 0;
assign detect_max[517][15] = (mid_1[4151:4144] > mid_2[4151:4144]) ? 1 : 0;
assign detect_max[517][16] = (mid_1[4151:4144] > mid_2[4159:4152]) ? 1 : 0;
assign detect_max[517][17] = (mid_1[4151:4144] > btm_0[4143:4136]) ? 1 : 0;
assign detect_max[517][18] = (mid_1[4151:4144] > btm_0[4151:4144]) ? 1 : 0;
assign detect_max[517][19] = (mid_1[4151:4144] > btm_0[4159:4152]) ? 1 : 0;
assign detect_max[517][20] = (mid_1[4151:4144] > btm_1[4143:4136]) ? 1 : 0;
assign detect_max[517][21] = (mid_1[4151:4144] > btm_1[4151:4144]) ? 1 : 0;
assign detect_max[517][22] = (mid_1[4151:4144] > btm_1[4159:4152]) ? 1 : 0;
assign detect_max[517][23] = (mid_1[4151:4144] > btm_2[4143:4136]) ? 1 : 0;
assign detect_max[517][24] = (mid_1[4151:4144] > btm_2[4151:4144]) ? 1 : 0;
assign detect_max[517][25] = (mid_1[4151:4144] > btm_2[4159:4152]) ? 1 : 0;

assign detect_max[518][0] = (mid_1[4159:4152] > top_0[4151:4144]) ? 1 : 0;
assign detect_max[518][1] = (mid_1[4159:4152] > top_0[4159:4152]) ? 1 : 0;
assign detect_max[518][2] = (mid_1[4159:4152] > top_0[4167:4160]) ? 1 : 0;
assign detect_max[518][3] = (mid_1[4159:4152] > top_1[4151:4144]) ? 1 : 0;
assign detect_max[518][4] = (mid_1[4159:4152] > top_1[4159:4152]) ? 1 : 0;
assign detect_max[518][5] = (mid_1[4159:4152] > top_1[4167:4160]) ? 1 : 0;
assign detect_max[518][6] = (mid_1[4159:4152] > top_2[4151:4144]) ? 1 : 0;
assign detect_max[518][7] = (mid_1[4159:4152] > top_2[4159:4152]) ? 1 : 0;
assign detect_max[518][8] = (mid_1[4159:4152] > top_2[4167:4160]) ? 1 : 0;
assign detect_max[518][9] = (mid_1[4159:4152] > mid_0[4151:4144]) ? 1 : 0;
assign detect_max[518][10] = (mid_1[4159:4152] > mid_0[4159:4152]) ? 1 : 0;
assign detect_max[518][11] = (mid_1[4159:4152] > mid_0[4167:4160]) ? 1 : 0;
assign detect_max[518][12] = (mid_1[4159:4152] > mid_1[4151:4144]) ? 1 : 0;
assign detect_max[518][13] = (mid_1[4159:4152] > mid_1[4167:4160]) ? 1 : 0;
assign detect_max[518][14] = (mid_1[4159:4152] > mid_2[4151:4144]) ? 1 : 0;
assign detect_max[518][15] = (mid_1[4159:4152] > mid_2[4159:4152]) ? 1 : 0;
assign detect_max[518][16] = (mid_1[4159:4152] > mid_2[4167:4160]) ? 1 : 0;
assign detect_max[518][17] = (mid_1[4159:4152] > btm_0[4151:4144]) ? 1 : 0;
assign detect_max[518][18] = (mid_1[4159:4152] > btm_0[4159:4152]) ? 1 : 0;
assign detect_max[518][19] = (mid_1[4159:4152] > btm_0[4167:4160]) ? 1 : 0;
assign detect_max[518][20] = (mid_1[4159:4152] > btm_1[4151:4144]) ? 1 : 0;
assign detect_max[518][21] = (mid_1[4159:4152] > btm_1[4159:4152]) ? 1 : 0;
assign detect_max[518][22] = (mid_1[4159:4152] > btm_1[4167:4160]) ? 1 : 0;
assign detect_max[518][23] = (mid_1[4159:4152] > btm_2[4151:4144]) ? 1 : 0;
assign detect_max[518][24] = (mid_1[4159:4152] > btm_2[4159:4152]) ? 1 : 0;
assign detect_max[518][25] = (mid_1[4159:4152] > btm_2[4167:4160]) ? 1 : 0;

assign detect_max[519][0] = (mid_1[4167:4160] > top_0[4159:4152]) ? 1 : 0;
assign detect_max[519][1] = (mid_1[4167:4160] > top_0[4167:4160]) ? 1 : 0;
assign detect_max[519][2] = (mid_1[4167:4160] > top_0[4175:4168]) ? 1 : 0;
assign detect_max[519][3] = (mid_1[4167:4160] > top_1[4159:4152]) ? 1 : 0;
assign detect_max[519][4] = (mid_1[4167:4160] > top_1[4167:4160]) ? 1 : 0;
assign detect_max[519][5] = (mid_1[4167:4160] > top_1[4175:4168]) ? 1 : 0;
assign detect_max[519][6] = (mid_1[4167:4160] > top_2[4159:4152]) ? 1 : 0;
assign detect_max[519][7] = (mid_1[4167:4160] > top_2[4167:4160]) ? 1 : 0;
assign detect_max[519][8] = (mid_1[4167:4160] > top_2[4175:4168]) ? 1 : 0;
assign detect_max[519][9] = (mid_1[4167:4160] > mid_0[4159:4152]) ? 1 : 0;
assign detect_max[519][10] = (mid_1[4167:4160] > mid_0[4167:4160]) ? 1 : 0;
assign detect_max[519][11] = (mid_1[4167:4160] > mid_0[4175:4168]) ? 1 : 0;
assign detect_max[519][12] = (mid_1[4167:4160] > mid_1[4159:4152]) ? 1 : 0;
assign detect_max[519][13] = (mid_1[4167:4160] > mid_1[4175:4168]) ? 1 : 0;
assign detect_max[519][14] = (mid_1[4167:4160] > mid_2[4159:4152]) ? 1 : 0;
assign detect_max[519][15] = (mid_1[4167:4160] > mid_2[4167:4160]) ? 1 : 0;
assign detect_max[519][16] = (mid_1[4167:4160] > mid_2[4175:4168]) ? 1 : 0;
assign detect_max[519][17] = (mid_1[4167:4160] > btm_0[4159:4152]) ? 1 : 0;
assign detect_max[519][18] = (mid_1[4167:4160] > btm_0[4167:4160]) ? 1 : 0;
assign detect_max[519][19] = (mid_1[4167:4160] > btm_0[4175:4168]) ? 1 : 0;
assign detect_max[519][20] = (mid_1[4167:4160] > btm_1[4159:4152]) ? 1 : 0;
assign detect_max[519][21] = (mid_1[4167:4160] > btm_1[4167:4160]) ? 1 : 0;
assign detect_max[519][22] = (mid_1[4167:4160] > btm_1[4175:4168]) ? 1 : 0;
assign detect_max[519][23] = (mid_1[4167:4160] > btm_2[4159:4152]) ? 1 : 0;
assign detect_max[519][24] = (mid_1[4167:4160] > btm_2[4167:4160]) ? 1 : 0;
assign detect_max[519][25] = (mid_1[4167:4160] > btm_2[4175:4168]) ? 1 : 0;

assign detect_max[520][0] = (mid_1[4175:4168] > top_0[4167:4160]) ? 1 : 0;
assign detect_max[520][1] = (mid_1[4175:4168] > top_0[4175:4168]) ? 1 : 0;
assign detect_max[520][2] = (mid_1[4175:4168] > top_0[4183:4176]) ? 1 : 0;
assign detect_max[520][3] = (mid_1[4175:4168] > top_1[4167:4160]) ? 1 : 0;
assign detect_max[520][4] = (mid_1[4175:4168] > top_1[4175:4168]) ? 1 : 0;
assign detect_max[520][5] = (mid_1[4175:4168] > top_1[4183:4176]) ? 1 : 0;
assign detect_max[520][6] = (mid_1[4175:4168] > top_2[4167:4160]) ? 1 : 0;
assign detect_max[520][7] = (mid_1[4175:4168] > top_2[4175:4168]) ? 1 : 0;
assign detect_max[520][8] = (mid_1[4175:4168] > top_2[4183:4176]) ? 1 : 0;
assign detect_max[520][9] = (mid_1[4175:4168] > mid_0[4167:4160]) ? 1 : 0;
assign detect_max[520][10] = (mid_1[4175:4168] > mid_0[4175:4168]) ? 1 : 0;
assign detect_max[520][11] = (mid_1[4175:4168] > mid_0[4183:4176]) ? 1 : 0;
assign detect_max[520][12] = (mid_1[4175:4168] > mid_1[4167:4160]) ? 1 : 0;
assign detect_max[520][13] = (mid_1[4175:4168] > mid_1[4183:4176]) ? 1 : 0;
assign detect_max[520][14] = (mid_1[4175:4168] > mid_2[4167:4160]) ? 1 : 0;
assign detect_max[520][15] = (mid_1[4175:4168] > mid_2[4175:4168]) ? 1 : 0;
assign detect_max[520][16] = (mid_1[4175:4168] > mid_2[4183:4176]) ? 1 : 0;
assign detect_max[520][17] = (mid_1[4175:4168] > btm_0[4167:4160]) ? 1 : 0;
assign detect_max[520][18] = (mid_1[4175:4168] > btm_0[4175:4168]) ? 1 : 0;
assign detect_max[520][19] = (mid_1[4175:4168] > btm_0[4183:4176]) ? 1 : 0;
assign detect_max[520][20] = (mid_1[4175:4168] > btm_1[4167:4160]) ? 1 : 0;
assign detect_max[520][21] = (mid_1[4175:4168] > btm_1[4175:4168]) ? 1 : 0;
assign detect_max[520][22] = (mid_1[4175:4168] > btm_1[4183:4176]) ? 1 : 0;
assign detect_max[520][23] = (mid_1[4175:4168] > btm_2[4167:4160]) ? 1 : 0;
assign detect_max[520][24] = (mid_1[4175:4168] > btm_2[4175:4168]) ? 1 : 0;
assign detect_max[520][25] = (mid_1[4175:4168] > btm_2[4183:4176]) ? 1 : 0;

assign detect_max[521][0] = (mid_1[4183:4176] > top_0[4175:4168]) ? 1 : 0;
assign detect_max[521][1] = (mid_1[4183:4176] > top_0[4183:4176]) ? 1 : 0;
assign detect_max[521][2] = (mid_1[4183:4176] > top_0[4191:4184]) ? 1 : 0;
assign detect_max[521][3] = (mid_1[4183:4176] > top_1[4175:4168]) ? 1 : 0;
assign detect_max[521][4] = (mid_1[4183:4176] > top_1[4183:4176]) ? 1 : 0;
assign detect_max[521][5] = (mid_1[4183:4176] > top_1[4191:4184]) ? 1 : 0;
assign detect_max[521][6] = (mid_1[4183:4176] > top_2[4175:4168]) ? 1 : 0;
assign detect_max[521][7] = (mid_1[4183:4176] > top_2[4183:4176]) ? 1 : 0;
assign detect_max[521][8] = (mid_1[4183:4176] > top_2[4191:4184]) ? 1 : 0;
assign detect_max[521][9] = (mid_1[4183:4176] > mid_0[4175:4168]) ? 1 : 0;
assign detect_max[521][10] = (mid_1[4183:4176] > mid_0[4183:4176]) ? 1 : 0;
assign detect_max[521][11] = (mid_1[4183:4176] > mid_0[4191:4184]) ? 1 : 0;
assign detect_max[521][12] = (mid_1[4183:4176] > mid_1[4175:4168]) ? 1 : 0;
assign detect_max[521][13] = (mid_1[4183:4176] > mid_1[4191:4184]) ? 1 : 0;
assign detect_max[521][14] = (mid_1[4183:4176] > mid_2[4175:4168]) ? 1 : 0;
assign detect_max[521][15] = (mid_1[4183:4176] > mid_2[4183:4176]) ? 1 : 0;
assign detect_max[521][16] = (mid_1[4183:4176] > mid_2[4191:4184]) ? 1 : 0;
assign detect_max[521][17] = (mid_1[4183:4176] > btm_0[4175:4168]) ? 1 : 0;
assign detect_max[521][18] = (mid_1[4183:4176] > btm_0[4183:4176]) ? 1 : 0;
assign detect_max[521][19] = (mid_1[4183:4176] > btm_0[4191:4184]) ? 1 : 0;
assign detect_max[521][20] = (mid_1[4183:4176] > btm_1[4175:4168]) ? 1 : 0;
assign detect_max[521][21] = (mid_1[4183:4176] > btm_1[4183:4176]) ? 1 : 0;
assign detect_max[521][22] = (mid_1[4183:4176] > btm_1[4191:4184]) ? 1 : 0;
assign detect_max[521][23] = (mid_1[4183:4176] > btm_2[4175:4168]) ? 1 : 0;
assign detect_max[521][24] = (mid_1[4183:4176] > btm_2[4183:4176]) ? 1 : 0;
assign detect_max[521][25] = (mid_1[4183:4176] > btm_2[4191:4184]) ? 1 : 0;

assign detect_max[522][0] = (mid_1[4191:4184] > top_0[4183:4176]) ? 1 : 0;
assign detect_max[522][1] = (mid_1[4191:4184] > top_0[4191:4184]) ? 1 : 0;
assign detect_max[522][2] = (mid_1[4191:4184] > top_0[4199:4192]) ? 1 : 0;
assign detect_max[522][3] = (mid_1[4191:4184] > top_1[4183:4176]) ? 1 : 0;
assign detect_max[522][4] = (mid_1[4191:4184] > top_1[4191:4184]) ? 1 : 0;
assign detect_max[522][5] = (mid_1[4191:4184] > top_1[4199:4192]) ? 1 : 0;
assign detect_max[522][6] = (mid_1[4191:4184] > top_2[4183:4176]) ? 1 : 0;
assign detect_max[522][7] = (mid_1[4191:4184] > top_2[4191:4184]) ? 1 : 0;
assign detect_max[522][8] = (mid_1[4191:4184] > top_2[4199:4192]) ? 1 : 0;
assign detect_max[522][9] = (mid_1[4191:4184] > mid_0[4183:4176]) ? 1 : 0;
assign detect_max[522][10] = (mid_1[4191:4184] > mid_0[4191:4184]) ? 1 : 0;
assign detect_max[522][11] = (mid_1[4191:4184] > mid_0[4199:4192]) ? 1 : 0;
assign detect_max[522][12] = (mid_1[4191:4184] > mid_1[4183:4176]) ? 1 : 0;
assign detect_max[522][13] = (mid_1[4191:4184] > mid_1[4199:4192]) ? 1 : 0;
assign detect_max[522][14] = (mid_1[4191:4184] > mid_2[4183:4176]) ? 1 : 0;
assign detect_max[522][15] = (mid_1[4191:4184] > mid_2[4191:4184]) ? 1 : 0;
assign detect_max[522][16] = (mid_1[4191:4184] > mid_2[4199:4192]) ? 1 : 0;
assign detect_max[522][17] = (mid_1[4191:4184] > btm_0[4183:4176]) ? 1 : 0;
assign detect_max[522][18] = (mid_1[4191:4184] > btm_0[4191:4184]) ? 1 : 0;
assign detect_max[522][19] = (mid_1[4191:4184] > btm_0[4199:4192]) ? 1 : 0;
assign detect_max[522][20] = (mid_1[4191:4184] > btm_1[4183:4176]) ? 1 : 0;
assign detect_max[522][21] = (mid_1[4191:4184] > btm_1[4191:4184]) ? 1 : 0;
assign detect_max[522][22] = (mid_1[4191:4184] > btm_1[4199:4192]) ? 1 : 0;
assign detect_max[522][23] = (mid_1[4191:4184] > btm_2[4183:4176]) ? 1 : 0;
assign detect_max[522][24] = (mid_1[4191:4184] > btm_2[4191:4184]) ? 1 : 0;
assign detect_max[522][25] = (mid_1[4191:4184] > btm_2[4199:4192]) ? 1 : 0;

assign detect_max[523][0] = (mid_1[4199:4192] > top_0[4191:4184]) ? 1 : 0;
assign detect_max[523][1] = (mid_1[4199:4192] > top_0[4199:4192]) ? 1 : 0;
assign detect_max[523][2] = (mid_1[4199:4192] > top_0[4207:4200]) ? 1 : 0;
assign detect_max[523][3] = (mid_1[4199:4192] > top_1[4191:4184]) ? 1 : 0;
assign detect_max[523][4] = (mid_1[4199:4192] > top_1[4199:4192]) ? 1 : 0;
assign detect_max[523][5] = (mid_1[4199:4192] > top_1[4207:4200]) ? 1 : 0;
assign detect_max[523][6] = (mid_1[4199:4192] > top_2[4191:4184]) ? 1 : 0;
assign detect_max[523][7] = (mid_1[4199:4192] > top_2[4199:4192]) ? 1 : 0;
assign detect_max[523][8] = (mid_1[4199:4192] > top_2[4207:4200]) ? 1 : 0;
assign detect_max[523][9] = (mid_1[4199:4192] > mid_0[4191:4184]) ? 1 : 0;
assign detect_max[523][10] = (mid_1[4199:4192] > mid_0[4199:4192]) ? 1 : 0;
assign detect_max[523][11] = (mid_1[4199:4192] > mid_0[4207:4200]) ? 1 : 0;
assign detect_max[523][12] = (mid_1[4199:4192] > mid_1[4191:4184]) ? 1 : 0;
assign detect_max[523][13] = (mid_1[4199:4192] > mid_1[4207:4200]) ? 1 : 0;
assign detect_max[523][14] = (mid_1[4199:4192] > mid_2[4191:4184]) ? 1 : 0;
assign detect_max[523][15] = (mid_1[4199:4192] > mid_2[4199:4192]) ? 1 : 0;
assign detect_max[523][16] = (mid_1[4199:4192] > mid_2[4207:4200]) ? 1 : 0;
assign detect_max[523][17] = (mid_1[4199:4192] > btm_0[4191:4184]) ? 1 : 0;
assign detect_max[523][18] = (mid_1[4199:4192] > btm_0[4199:4192]) ? 1 : 0;
assign detect_max[523][19] = (mid_1[4199:4192] > btm_0[4207:4200]) ? 1 : 0;
assign detect_max[523][20] = (mid_1[4199:4192] > btm_1[4191:4184]) ? 1 : 0;
assign detect_max[523][21] = (mid_1[4199:4192] > btm_1[4199:4192]) ? 1 : 0;
assign detect_max[523][22] = (mid_1[4199:4192] > btm_1[4207:4200]) ? 1 : 0;
assign detect_max[523][23] = (mid_1[4199:4192] > btm_2[4191:4184]) ? 1 : 0;
assign detect_max[523][24] = (mid_1[4199:4192] > btm_2[4199:4192]) ? 1 : 0;
assign detect_max[523][25] = (mid_1[4199:4192] > btm_2[4207:4200]) ? 1 : 0;

assign detect_max[524][0] = (mid_1[4207:4200] > top_0[4199:4192]) ? 1 : 0;
assign detect_max[524][1] = (mid_1[4207:4200] > top_0[4207:4200]) ? 1 : 0;
assign detect_max[524][2] = (mid_1[4207:4200] > top_0[4215:4208]) ? 1 : 0;
assign detect_max[524][3] = (mid_1[4207:4200] > top_1[4199:4192]) ? 1 : 0;
assign detect_max[524][4] = (mid_1[4207:4200] > top_1[4207:4200]) ? 1 : 0;
assign detect_max[524][5] = (mid_1[4207:4200] > top_1[4215:4208]) ? 1 : 0;
assign detect_max[524][6] = (mid_1[4207:4200] > top_2[4199:4192]) ? 1 : 0;
assign detect_max[524][7] = (mid_1[4207:4200] > top_2[4207:4200]) ? 1 : 0;
assign detect_max[524][8] = (mid_1[4207:4200] > top_2[4215:4208]) ? 1 : 0;
assign detect_max[524][9] = (mid_1[4207:4200] > mid_0[4199:4192]) ? 1 : 0;
assign detect_max[524][10] = (mid_1[4207:4200] > mid_0[4207:4200]) ? 1 : 0;
assign detect_max[524][11] = (mid_1[4207:4200] > mid_0[4215:4208]) ? 1 : 0;
assign detect_max[524][12] = (mid_1[4207:4200] > mid_1[4199:4192]) ? 1 : 0;
assign detect_max[524][13] = (mid_1[4207:4200] > mid_1[4215:4208]) ? 1 : 0;
assign detect_max[524][14] = (mid_1[4207:4200] > mid_2[4199:4192]) ? 1 : 0;
assign detect_max[524][15] = (mid_1[4207:4200] > mid_2[4207:4200]) ? 1 : 0;
assign detect_max[524][16] = (mid_1[4207:4200] > mid_2[4215:4208]) ? 1 : 0;
assign detect_max[524][17] = (mid_1[4207:4200] > btm_0[4199:4192]) ? 1 : 0;
assign detect_max[524][18] = (mid_1[4207:4200] > btm_0[4207:4200]) ? 1 : 0;
assign detect_max[524][19] = (mid_1[4207:4200] > btm_0[4215:4208]) ? 1 : 0;
assign detect_max[524][20] = (mid_1[4207:4200] > btm_1[4199:4192]) ? 1 : 0;
assign detect_max[524][21] = (mid_1[4207:4200] > btm_1[4207:4200]) ? 1 : 0;
assign detect_max[524][22] = (mid_1[4207:4200] > btm_1[4215:4208]) ? 1 : 0;
assign detect_max[524][23] = (mid_1[4207:4200] > btm_2[4199:4192]) ? 1 : 0;
assign detect_max[524][24] = (mid_1[4207:4200] > btm_2[4207:4200]) ? 1 : 0;
assign detect_max[524][25] = (mid_1[4207:4200] > btm_2[4215:4208]) ? 1 : 0;

assign detect_max[525][0] = (mid_1[4215:4208] > top_0[4207:4200]) ? 1 : 0;
assign detect_max[525][1] = (mid_1[4215:4208] > top_0[4215:4208]) ? 1 : 0;
assign detect_max[525][2] = (mid_1[4215:4208] > top_0[4223:4216]) ? 1 : 0;
assign detect_max[525][3] = (mid_1[4215:4208] > top_1[4207:4200]) ? 1 : 0;
assign detect_max[525][4] = (mid_1[4215:4208] > top_1[4215:4208]) ? 1 : 0;
assign detect_max[525][5] = (mid_1[4215:4208] > top_1[4223:4216]) ? 1 : 0;
assign detect_max[525][6] = (mid_1[4215:4208] > top_2[4207:4200]) ? 1 : 0;
assign detect_max[525][7] = (mid_1[4215:4208] > top_2[4215:4208]) ? 1 : 0;
assign detect_max[525][8] = (mid_1[4215:4208] > top_2[4223:4216]) ? 1 : 0;
assign detect_max[525][9] = (mid_1[4215:4208] > mid_0[4207:4200]) ? 1 : 0;
assign detect_max[525][10] = (mid_1[4215:4208] > mid_0[4215:4208]) ? 1 : 0;
assign detect_max[525][11] = (mid_1[4215:4208] > mid_0[4223:4216]) ? 1 : 0;
assign detect_max[525][12] = (mid_1[4215:4208] > mid_1[4207:4200]) ? 1 : 0;
assign detect_max[525][13] = (mid_1[4215:4208] > mid_1[4223:4216]) ? 1 : 0;
assign detect_max[525][14] = (mid_1[4215:4208] > mid_2[4207:4200]) ? 1 : 0;
assign detect_max[525][15] = (mid_1[4215:4208] > mid_2[4215:4208]) ? 1 : 0;
assign detect_max[525][16] = (mid_1[4215:4208] > mid_2[4223:4216]) ? 1 : 0;
assign detect_max[525][17] = (mid_1[4215:4208] > btm_0[4207:4200]) ? 1 : 0;
assign detect_max[525][18] = (mid_1[4215:4208] > btm_0[4215:4208]) ? 1 : 0;
assign detect_max[525][19] = (mid_1[4215:4208] > btm_0[4223:4216]) ? 1 : 0;
assign detect_max[525][20] = (mid_1[4215:4208] > btm_1[4207:4200]) ? 1 : 0;
assign detect_max[525][21] = (mid_1[4215:4208] > btm_1[4215:4208]) ? 1 : 0;
assign detect_max[525][22] = (mid_1[4215:4208] > btm_1[4223:4216]) ? 1 : 0;
assign detect_max[525][23] = (mid_1[4215:4208] > btm_2[4207:4200]) ? 1 : 0;
assign detect_max[525][24] = (mid_1[4215:4208] > btm_2[4215:4208]) ? 1 : 0;
assign detect_max[525][25] = (mid_1[4215:4208] > btm_2[4223:4216]) ? 1 : 0;

assign detect_max[526][0] = (mid_1[4223:4216] > top_0[4215:4208]) ? 1 : 0;
assign detect_max[526][1] = (mid_1[4223:4216] > top_0[4223:4216]) ? 1 : 0;
assign detect_max[526][2] = (mid_1[4223:4216] > top_0[4231:4224]) ? 1 : 0;
assign detect_max[526][3] = (mid_1[4223:4216] > top_1[4215:4208]) ? 1 : 0;
assign detect_max[526][4] = (mid_1[4223:4216] > top_1[4223:4216]) ? 1 : 0;
assign detect_max[526][5] = (mid_1[4223:4216] > top_1[4231:4224]) ? 1 : 0;
assign detect_max[526][6] = (mid_1[4223:4216] > top_2[4215:4208]) ? 1 : 0;
assign detect_max[526][7] = (mid_1[4223:4216] > top_2[4223:4216]) ? 1 : 0;
assign detect_max[526][8] = (mid_1[4223:4216] > top_2[4231:4224]) ? 1 : 0;
assign detect_max[526][9] = (mid_1[4223:4216] > mid_0[4215:4208]) ? 1 : 0;
assign detect_max[526][10] = (mid_1[4223:4216] > mid_0[4223:4216]) ? 1 : 0;
assign detect_max[526][11] = (mid_1[4223:4216] > mid_0[4231:4224]) ? 1 : 0;
assign detect_max[526][12] = (mid_1[4223:4216] > mid_1[4215:4208]) ? 1 : 0;
assign detect_max[526][13] = (mid_1[4223:4216] > mid_1[4231:4224]) ? 1 : 0;
assign detect_max[526][14] = (mid_1[4223:4216] > mid_2[4215:4208]) ? 1 : 0;
assign detect_max[526][15] = (mid_1[4223:4216] > mid_2[4223:4216]) ? 1 : 0;
assign detect_max[526][16] = (mid_1[4223:4216] > mid_2[4231:4224]) ? 1 : 0;
assign detect_max[526][17] = (mid_1[4223:4216] > btm_0[4215:4208]) ? 1 : 0;
assign detect_max[526][18] = (mid_1[4223:4216] > btm_0[4223:4216]) ? 1 : 0;
assign detect_max[526][19] = (mid_1[4223:4216] > btm_0[4231:4224]) ? 1 : 0;
assign detect_max[526][20] = (mid_1[4223:4216] > btm_1[4215:4208]) ? 1 : 0;
assign detect_max[526][21] = (mid_1[4223:4216] > btm_1[4223:4216]) ? 1 : 0;
assign detect_max[526][22] = (mid_1[4223:4216] > btm_1[4231:4224]) ? 1 : 0;
assign detect_max[526][23] = (mid_1[4223:4216] > btm_2[4215:4208]) ? 1 : 0;
assign detect_max[526][24] = (mid_1[4223:4216] > btm_2[4223:4216]) ? 1 : 0;
assign detect_max[526][25] = (mid_1[4223:4216] > btm_2[4231:4224]) ? 1 : 0;

assign detect_max[527][0] = (mid_1[4231:4224] > top_0[4223:4216]) ? 1 : 0;
assign detect_max[527][1] = (mid_1[4231:4224] > top_0[4231:4224]) ? 1 : 0;
assign detect_max[527][2] = (mid_1[4231:4224] > top_0[4239:4232]) ? 1 : 0;
assign detect_max[527][3] = (mid_1[4231:4224] > top_1[4223:4216]) ? 1 : 0;
assign detect_max[527][4] = (mid_1[4231:4224] > top_1[4231:4224]) ? 1 : 0;
assign detect_max[527][5] = (mid_1[4231:4224] > top_1[4239:4232]) ? 1 : 0;
assign detect_max[527][6] = (mid_1[4231:4224] > top_2[4223:4216]) ? 1 : 0;
assign detect_max[527][7] = (mid_1[4231:4224] > top_2[4231:4224]) ? 1 : 0;
assign detect_max[527][8] = (mid_1[4231:4224] > top_2[4239:4232]) ? 1 : 0;
assign detect_max[527][9] = (mid_1[4231:4224] > mid_0[4223:4216]) ? 1 : 0;
assign detect_max[527][10] = (mid_1[4231:4224] > mid_0[4231:4224]) ? 1 : 0;
assign detect_max[527][11] = (mid_1[4231:4224] > mid_0[4239:4232]) ? 1 : 0;
assign detect_max[527][12] = (mid_1[4231:4224] > mid_1[4223:4216]) ? 1 : 0;
assign detect_max[527][13] = (mid_1[4231:4224] > mid_1[4239:4232]) ? 1 : 0;
assign detect_max[527][14] = (mid_1[4231:4224] > mid_2[4223:4216]) ? 1 : 0;
assign detect_max[527][15] = (mid_1[4231:4224] > mid_2[4231:4224]) ? 1 : 0;
assign detect_max[527][16] = (mid_1[4231:4224] > mid_2[4239:4232]) ? 1 : 0;
assign detect_max[527][17] = (mid_1[4231:4224] > btm_0[4223:4216]) ? 1 : 0;
assign detect_max[527][18] = (mid_1[4231:4224] > btm_0[4231:4224]) ? 1 : 0;
assign detect_max[527][19] = (mid_1[4231:4224] > btm_0[4239:4232]) ? 1 : 0;
assign detect_max[527][20] = (mid_1[4231:4224] > btm_1[4223:4216]) ? 1 : 0;
assign detect_max[527][21] = (mid_1[4231:4224] > btm_1[4231:4224]) ? 1 : 0;
assign detect_max[527][22] = (mid_1[4231:4224] > btm_1[4239:4232]) ? 1 : 0;
assign detect_max[527][23] = (mid_1[4231:4224] > btm_2[4223:4216]) ? 1 : 0;
assign detect_max[527][24] = (mid_1[4231:4224] > btm_2[4231:4224]) ? 1 : 0;
assign detect_max[527][25] = (mid_1[4231:4224] > btm_2[4239:4232]) ? 1 : 0;

assign detect_max[528][0] = (mid_1[4239:4232] > top_0[4231:4224]) ? 1 : 0;
assign detect_max[528][1] = (mid_1[4239:4232] > top_0[4239:4232]) ? 1 : 0;
assign detect_max[528][2] = (mid_1[4239:4232] > top_0[4247:4240]) ? 1 : 0;
assign detect_max[528][3] = (mid_1[4239:4232] > top_1[4231:4224]) ? 1 : 0;
assign detect_max[528][4] = (mid_1[4239:4232] > top_1[4239:4232]) ? 1 : 0;
assign detect_max[528][5] = (mid_1[4239:4232] > top_1[4247:4240]) ? 1 : 0;
assign detect_max[528][6] = (mid_1[4239:4232] > top_2[4231:4224]) ? 1 : 0;
assign detect_max[528][7] = (mid_1[4239:4232] > top_2[4239:4232]) ? 1 : 0;
assign detect_max[528][8] = (mid_1[4239:4232] > top_2[4247:4240]) ? 1 : 0;
assign detect_max[528][9] = (mid_1[4239:4232] > mid_0[4231:4224]) ? 1 : 0;
assign detect_max[528][10] = (mid_1[4239:4232] > mid_0[4239:4232]) ? 1 : 0;
assign detect_max[528][11] = (mid_1[4239:4232] > mid_0[4247:4240]) ? 1 : 0;
assign detect_max[528][12] = (mid_1[4239:4232] > mid_1[4231:4224]) ? 1 : 0;
assign detect_max[528][13] = (mid_1[4239:4232] > mid_1[4247:4240]) ? 1 : 0;
assign detect_max[528][14] = (mid_1[4239:4232] > mid_2[4231:4224]) ? 1 : 0;
assign detect_max[528][15] = (mid_1[4239:4232] > mid_2[4239:4232]) ? 1 : 0;
assign detect_max[528][16] = (mid_1[4239:4232] > mid_2[4247:4240]) ? 1 : 0;
assign detect_max[528][17] = (mid_1[4239:4232] > btm_0[4231:4224]) ? 1 : 0;
assign detect_max[528][18] = (mid_1[4239:4232] > btm_0[4239:4232]) ? 1 : 0;
assign detect_max[528][19] = (mid_1[4239:4232] > btm_0[4247:4240]) ? 1 : 0;
assign detect_max[528][20] = (mid_1[4239:4232] > btm_1[4231:4224]) ? 1 : 0;
assign detect_max[528][21] = (mid_1[4239:4232] > btm_1[4239:4232]) ? 1 : 0;
assign detect_max[528][22] = (mid_1[4239:4232] > btm_1[4247:4240]) ? 1 : 0;
assign detect_max[528][23] = (mid_1[4239:4232] > btm_2[4231:4224]) ? 1 : 0;
assign detect_max[528][24] = (mid_1[4239:4232] > btm_2[4239:4232]) ? 1 : 0;
assign detect_max[528][25] = (mid_1[4239:4232] > btm_2[4247:4240]) ? 1 : 0;

assign detect_max[529][0] = (mid_1[4247:4240] > top_0[4239:4232]) ? 1 : 0;
assign detect_max[529][1] = (mid_1[4247:4240] > top_0[4247:4240]) ? 1 : 0;
assign detect_max[529][2] = (mid_1[4247:4240] > top_0[4255:4248]) ? 1 : 0;
assign detect_max[529][3] = (mid_1[4247:4240] > top_1[4239:4232]) ? 1 : 0;
assign detect_max[529][4] = (mid_1[4247:4240] > top_1[4247:4240]) ? 1 : 0;
assign detect_max[529][5] = (mid_1[4247:4240] > top_1[4255:4248]) ? 1 : 0;
assign detect_max[529][6] = (mid_1[4247:4240] > top_2[4239:4232]) ? 1 : 0;
assign detect_max[529][7] = (mid_1[4247:4240] > top_2[4247:4240]) ? 1 : 0;
assign detect_max[529][8] = (mid_1[4247:4240] > top_2[4255:4248]) ? 1 : 0;
assign detect_max[529][9] = (mid_1[4247:4240] > mid_0[4239:4232]) ? 1 : 0;
assign detect_max[529][10] = (mid_1[4247:4240] > mid_0[4247:4240]) ? 1 : 0;
assign detect_max[529][11] = (mid_1[4247:4240] > mid_0[4255:4248]) ? 1 : 0;
assign detect_max[529][12] = (mid_1[4247:4240] > mid_1[4239:4232]) ? 1 : 0;
assign detect_max[529][13] = (mid_1[4247:4240] > mid_1[4255:4248]) ? 1 : 0;
assign detect_max[529][14] = (mid_1[4247:4240] > mid_2[4239:4232]) ? 1 : 0;
assign detect_max[529][15] = (mid_1[4247:4240] > mid_2[4247:4240]) ? 1 : 0;
assign detect_max[529][16] = (mid_1[4247:4240] > mid_2[4255:4248]) ? 1 : 0;
assign detect_max[529][17] = (mid_1[4247:4240] > btm_0[4239:4232]) ? 1 : 0;
assign detect_max[529][18] = (mid_1[4247:4240] > btm_0[4247:4240]) ? 1 : 0;
assign detect_max[529][19] = (mid_1[4247:4240] > btm_0[4255:4248]) ? 1 : 0;
assign detect_max[529][20] = (mid_1[4247:4240] > btm_1[4239:4232]) ? 1 : 0;
assign detect_max[529][21] = (mid_1[4247:4240] > btm_1[4247:4240]) ? 1 : 0;
assign detect_max[529][22] = (mid_1[4247:4240] > btm_1[4255:4248]) ? 1 : 0;
assign detect_max[529][23] = (mid_1[4247:4240] > btm_2[4239:4232]) ? 1 : 0;
assign detect_max[529][24] = (mid_1[4247:4240] > btm_2[4247:4240]) ? 1 : 0;
assign detect_max[529][25] = (mid_1[4247:4240] > btm_2[4255:4248]) ? 1 : 0;

assign detect_max[530][0] = (mid_1[4255:4248] > top_0[4247:4240]) ? 1 : 0;
assign detect_max[530][1] = (mid_1[4255:4248] > top_0[4255:4248]) ? 1 : 0;
assign detect_max[530][2] = (mid_1[4255:4248] > top_0[4263:4256]) ? 1 : 0;
assign detect_max[530][3] = (mid_1[4255:4248] > top_1[4247:4240]) ? 1 : 0;
assign detect_max[530][4] = (mid_1[4255:4248] > top_1[4255:4248]) ? 1 : 0;
assign detect_max[530][5] = (mid_1[4255:4248] > top_1[4263:4256]) ? 1 : 0;
assign detect_max[530][6] = (mid_1[4255:4248] > top_2[4247:4240]) ? 1 : 0;
assign detect_max[530][7] = (mid_1[4255:4248] > top_2[4255:4248]) ? 1 : 0;
assign detect_max[530][8] = (mid_1[4255:4248] > top_2[4263:4256]) ? 1 : 0;
assign detect_max[530][9] = (mid_1[4255:4248] > mid_0[4247:4240]) ? 1 : 0;
assign detect_max[530][10] = (mid_1[4255:4248] > mid_0[4255:4248]) ? 1 : 0;
assign detect_max[530][11] = (mid_1[4255:4248] > mid_0[4263:4256]) ? 1 : 0;
assign detect_max[530][12] = (mid_1[4255:4248] > mid_1[4247:4240]) ? 1 : 0;
assign detect_max[530][13] = (mid_1[4255:4248] > mid_1[4263:4256]) ? 1 : 0;
assign detect_max[530][14] = (mid_1[4255:4248] > mid_2[4247:4240]) ? 1 : 0;
assign detect_max[530][15] = (mid_1[4255:4248] > mid_2[4255:4248]) ? 1 : 0;
assign detect_max[530][16] = (mid_1[4255:4248] > mid_2[4263:4256]) ? 1 : 0;
assign detect_max[530][17] = (mid_1[4255:4248] > btm_0[4247:4240]) ? 1 : 0;
assign detect_max[530][18] = (mid_1[4255:4248] > btm_0[4255:4248]) ? 1 : 0;
assign detect_max[530][19] = (mid_1[4255:4248] > btm_0[4263:4256]) ? 1 : 0;
assign detect_max[530][20] = (mid_1[4255:4248] > btm_1[4247:4240]) ? 1 : 0;
assign detect_max[530][21] = (mid_1[4255:4248] > btm_1[4255:4248]) ? 1 : 0;
assign detect_max[530][22] = (mid_1[4255:4248] > btm_1[4263:4256]) ? 1 : 0;
assign detect_max[530][23] = (mid_1[4255:4248] > btm_2[4247:4240]) ? 1 : 0;
assign detect_max[530][24] = (mid_1[4255:4248] > btm_2[4255:4248]) ? 1 : 0;
assign detect_max[530][25] = (mid_1[4255:4248] > btm_2[4263:4256]) ? 1 : 0;

assign detect_max[531][0] = (mid_1[4263:4256] > top_0[4255:4248]) ? 1 : 0;
assign detect_max[531][1] = (mid_1[4263:4256] > top_0[4263:4256]) ? 1 : 0;
assign detect_max[531][2] = (mid_1[4263:4256] > top_0[4271:4264]) ? 1 : 0;
assign detect_max[531][3] = (mid_1[4263:4256] > top_1[4255:4248]) ? 1 : 0;
assign detect_max[531][4] = (mid_1[4263:4256] > top_1[4263:4256]) ? 1 : 0;
assign detect_max[531][5] = (mid_1[4263:4256] > top_1[4271:4264]) ? 1 : 0;
assign detect_max[531][6] = (mid_1[4263:4256] > top_2[4255:4248]) ? 1 : 0;
assign detect_max[531][7] = (mid_1[4263:4256] > top_2[4263:4256]) ? 1 : 0;
assign detect_max[531][8] = (mid_1[4263:4256] > top_2[4271:4264]) ? 1 : 0;
assign detect_max[531][9] = (mid_1[4263:4256] > mid_0[4255:4248]) ? 1 : 0;
assign detect_max[531][10] = (mid_1[4263:4256] > mid_0[4263:4256]) ? 1 : 0;
assign detect_max[531][11] = (mid_1[4263:4256] > mid_0[4271:4264]) ? 1 : 0;
assign detect_max[531][12] = (mid_1[4263:4256] > mid_1[4255:4248]) ? 1 : 0;
assign detect_max[531][13] = (mid_1[4263:4256] > mid_1[4271:4264]) ? 1 : 0;
assign detect_max[531][14] = (mid_1[4263:4256] > mid_2[4255:4248]) ? 1 : 0;
assign detect_max[531][15] = (mid_1[4263:4256] > mid_2[4263:4256]) ? 1 : 0;
assign detect_max[531][16] = (mid_1[4263:4256] > mid_2[4271:4264]) ? 1 : 0;
assign detect_max[531][17] = (mid_1[4263:4256] > btm_0[4255:4248]) ? 1 : 0;
assign detect_max[531][18] = (mid_1[4263:4256] > btm_0[4263:4256]) ? 1 : 0;
assign detect_max[531][19] = (mid_1[4263:4256] > btm_0[4271:4264]) ? 1 : 0;
assign detect_max[531][20] = (mid_1[4263:4256] > btm_1[4255:4248]) ? 1 : 0;
assign detect_max[531][21] = (mid_1[4263:4256] > btm_1[4263:4256]) ? 1 : 0;
assign detect_max[531][22] = (mid_1[4263:4256] > btm_1[4271:4264]) ? 1 : 0;
assign detect_max[531][23] = (mid_1[4263:4256] > btm_2[4255:4248]) ? 1 : 0;
assign detect_max[531][24] = (mid_1[4263:4256] > btm_2[4263:4256]) ? 1 : 0;
assign detect_max[531][25] = (mid_1[4263:4256] > btm_2[4271:4264]) ? 1 : 0;

assign detect_max[532][0] = (mid_1[4271:4264] > top_0[4263:4256]) ? 1 : 0;
assign detect_max[532][1] = (mid_1[4271:4264] > top_0[4271:4264]) ? 1 : 0;
assign detect_max[532][2] = (mid_1[4271:4264] > top_0[4279:4272]) ? 1 : 0;
assign detect_max[532][3] = (mid_1[4271:4264] > top_1[4263:4256]) ? 1 : 0;
assign detect_max[532][4] = (mid_1[4271:4264] > top_1[4271:4264]) ? 1 : 0;
assign detect_max[532][5] = (mid_1[4271:4264] > top_1[4279:4272]) ? 1 : 0;
assign detect_max[532][6] = (mid_1[4271:4264] > top_2[4263:4256]) ? 1 : 0;
assign detect_max[532][7] = (mid_1[4271:4264] > top_2[4271:4264]) ? 1 : 0;
assign detect_max[532][8] = (mid_1[4271:4264] > top_2[4279:4272]) ? 1 : 0;
assign detect_max[532][9] = (mid_1[4271:4264] > mid_0[4263:4256]) ? 1 : 0;
assign detect_max[532][10] = (mid_1[4271:4264] > mid_0[4271:4264]) ? 1 : 0;
assign detect_max[532][11] = (mid_1[4271:4264] > mid_0[4279:4272]) ? 1 : 0;
assign detect_max[532][12] = (mid_1[4271:4264] > mid_1[4263:4256]) ? 1 : 0;
assign detect_max[532][13] = (mid_1[4271:4264] > mid_1[4279:4272]) ? 1 : 0;
assign detect_max[532][14] = (mid_1[4271:4264] > mid_2[4263:4256]) ? 1 : 0;
assign detect_max[532][15] = (mid_1[4271:4264] > mid_2[4271:4264]) ? 1 : 0;
assign detect_max[532][16] = (mid_1[4271:4264] > mid_2[4279:4272]) ? 1 : 0;
assign detect_max[532][17] = (mid_1[4271:4264] > btm_0[4263:4256]) ? 1 : 0;
assign detect_max[532][18] = (mid_1[4271:4264] > btm_0[4271:4264]) ? 1 : 0;
assign detect_max[532][19] = (mid_1[4271:4264] > btm_0[4279:4272]) ? 1 : 0;
assign detect_max[532][20] = (mid_1[4271:4264] > btm_1[4263:4256]) ? 1 : 0;
assign detect_max[532][21] = (mid_1[4271:4264] > btm_1[4271:4264]) ? 1 : 0;
assign detect_max[532][22] = (mid_1[4271:4264] > btm_1[4279:4272]) ? 1 : 0;
assign detect_max[532][23] = (mid_1[4271:4264] > btm_2[4263:4256]) ? 1 : 0;
assign detect_max[532][24] = (mid_1[4271:4264] > btm_2[4271:4264]) ? 1 : 0;
assign detect_max[532][25] = (mid_1[4271:4264] > btm_2[4279:4272]) ? 1 : 0;

assign detect_max[533][0] = (mid_1[4279:4272] > top_0[4271:4264]) ? 1 : 0;
assign detect_max[533][1] = (mid_1[4279:4272] > top_0[4279:4272]) ? 1 : 0;
assign detect_max[533][2] = (mid_1[4279:4272] > top_0[4287:4280]) ? 1 : 0;
assign detect_max[533][3] = (mid_1[4279:4272] > top_1[4271:4264]) ? 1 : 0;
assign detect_max[533][4] = (mid_1[4279:4272] > top_1[4279:4272]) ? 1 : 0;
assign detect_max[533][5] = (mid_1[4279:4272] > top_1[4287:4280]) ? 1 : 0;
assign detect_max[533][6] = (mid_1[4279:4272] > top_2[4271:4264]) ? 1 : 0;
assign detect_max[533][7] = (mid_1[4279:4272] > top_2[4279:4272]) ? 1 : 0;
assign detect_max[533][8] = (mid_1[4279:4272] > top_2[4287:4280]) ? 1 : 0;
assign detect_max[533][9] = (mid_1[4279:4272] > mid_0[4271:4264]) ? 1 : 0;
assign detect_max[533][10] = (mid_1[4279:4272] > mid_0[4279:4272]) ? 1 : 0;
assign detect_max[533][11] = (mid_1[4279:4272] > mid_0[4287:4280]) ? 1 : 0;
assign detect_max[533][12] = (mid_1[4279:4272] > mid_1[4271:4264]) ? 1 : 0;
assign detect_max[533][13] = (mid_1[4279:4272] > mid_1[4287:4280]) ? 1 : 0;
assign detect_max[533][14] = (mid_1[4279:4272] > mid_2[4271:4264]) ? 1 : 0;
assign detect_max[533][15] = (mid_1[4279:4272] > mid_2[4279:4272]) ? 1 : 0;
assign detect_max[533][16] = (mid_1[4279:4272] > mid_2[4287:4280]) ? 1 : 0;
assign detect_max[533][17] = (mid_1[4279:4272] > btm_0[4271:4264]) ? 1 : 0;
assign detect_max[533][18] = (mid_1[4279:4272] > btm_0[4279:4272]) ? 1 : 0;
assign detect_max[533][19] = (mid_1[4279:4272] > btm_0[4287:4280]) ? 1 : 0;
assign detect_max[533][20] = (mid_1[4279:4272] > btm_1[4271:4264]) ? 1 : 0;
assign detect_max[533][21] = (mid_1[4279:4272] > btm_1[4279:4272]) ? 1 : 0;
assign detect_max[533][22] = (mid_1[4279:4272] > btm_1[4287:4280]) ? 1 : 0;
assign detect_max[533][23] = (mid_1[4279:4272] > btm_2[4271:4264]) ? 1 : 0;
assign detect_max[533][24] = (mid_1[4279:4272] > btm_2[4279:4272]) ? 1 : 0;
assign detect_max[533][25] = (mid_1[4279:4272] > btm_2[4287:4280]) ? 1 : 0;

assign detect_max[534][0] = (mid_1[4287:4280] > top_0[4279:4272]) ? 1 : 0;
assign detect_max[534][1] = (mid_1[4287:4280] > top_0[4287:4280]) ? 1 : 0;
assign detect_max[534][2] = (mid_1[4287:4280] > top_0[4295:4288]) ? 1 : 0;
assign detect_max[534][3] = (mid_1[4287:4280] > top_1[4279:4272]) ? 1 : 0;
assign detect_max[534][4] = (mid_1[4287:4280] > top_1[4287:4280]) ? 1 : 0;
assign detect_max[534][5] = (mid_1[4287:4280] > top_1[4295:4288]) ? 1 : 0;
assign detect_max[534][6] = (mid_1[4287:4280] > top_2[4279:4272]) ? 1 : 0;
assign detect_max[534][7] = (mid_1[4287:4280] > top_2[4287:4280]) ? 1 : 0;
assign detect_max[534][8] = (mid_1[4287:4280] > top_2[4295:4288]) ? 1 : 0;
assign detect_max[534][9] = (mid_1[4287:4280] > mid_0[4279:4272]) ? 1 : 0;
assign detect_max[534][10] = (mid_1[4287:4280] > mid_0[4287:4280]) ? 1 : 0;
assign detect_max[534][11] = (mid_1[4287:4280] > mid_0[4295:4288]) ? 1 : 0;
assign detect_max[534][12] = (mid_1[4287:4280] > mid_1[4279:4272]) ? 1 : 0;
assign detect_max[534][13] = (mid_1[4287:4280] > mid_1[4295:4288]) ? 1 : 0;
assign detect_max[534][14] = (mid_1[4287:4280] > mid_2[4279:4272]) ? 1 : 0;
assign detect_max[534][15] = (mid_1[4287:4280] > mid_2[4287:4280]) ? 1 : 0;
assign detect_max[534][16] = (mid_1[4287:4280] > mid_2[4295:4288]) ? 1 : 0;
assign detect_max[534][17] = (mid_1[4287:4280] > btm_0[4279:4272]) ? 1 : 0;
assign detect_max[534][18] = (mid_1[4287:4280] > btm_0[4287:4280]) ? 1 : 0;
assign detect_max[534][19] = (mid_1[4287:4280] > btm_0[4295:4288]) ? 1 : 0;
assign detect_max[534][20] = (mid_1[4287:4280] > btm_1[4279:4272]) ? 1 : 0;
assign detect_max[534][21] = (mid_1[4287:4280] > btm_1[4287:4280]) ? 1 : 0;
assign detect_max[534][22] = (mid_1[4287:4280] > btm_1[4295:4288]) ? 1 : 0;
assign detect_max[534][23] = (mid_1[4287:4280] > btm_2[4279:4272]) ? 1 : 0;
assign detect_max[534][24] = (mid_1[4287:4280] > btm_2[4287:4280]) ? 1 : 0;
assign detect_max[534][25] = (mid_1[4287:4280] > btm_2[4295:4288]) ? 1 : 0;

assign detect_max[535][0] = (mid_1[4295:4288] > top_0[4287:4280]) ? 1 : 0;
assign detect_max[535][1] = (mid_1[4295:4288] > top_0[4295:4288]) ? 1 : 0;
assign detect_max[535][2] = (mid_1[4295:4288] > top_0[4303:4296]) ? 1 : 0;
assign detect_max[535][3] = (mid_1[4295:4288] > top_1[4287:4280]) ? 1 : 0;
assign detect_max[535][4] = (mid_1[4295:4288] > top_1[4295:4288]) ? 1 : 0;
assign detect_max[535][5] = (mid_1[4295:4288] > top_1[4303:4296]) ? 1 : 0;
assign detect_max[535][6] = (mid_1[4295:4288] > top_2[4287:4280]) ? 1 : 0;
assign detect_max[535][7] = (mid_1[4295:4288] > top_2[4295:4288]) ? 1 : 0;
assign detect_max[535][8] = (mid_1[4295:4288] > top_2[4303:4296]) ? 1 : 0;
assign detect_max[535][9] = (mid_1[4295:4288] > mid_0[4287:4280]) ? 1 : 0;
assign detect_max[535][10] = (mid_1[4295:4288] > mid_0[4295:4288]) ? 1 : 0;
assign detect_max[535][11] = (mid_1[4295:4288] > mid_0[4303:4296]) ? 1 : 0;
assign detect_max[535][12] = (mid_1[4295:4288] > mid_1[4287:4280]) ? 1 : 0;
assign detect_max[535][13] = (mid_1[4295:4288] > mid_1[4303:4296]) ? 1 : 0;
assign detect_max[535][14] = (mid_1[4295:4288] > mid_2[4287:4280]) ? 1 : 0;
assign detect_max[535][15] = (mid_1[4295:4288] > mid_2[4295:4288]) ? 1 : 0;
assign detect_max[535][16] = (mid_1[4295:4288] > mid_2[4303:4296]) ? 1 : 0;
assign detect_max[535][17] = (mid_1[4295:4288] > btm_0[4287:4280]) ? 1 : 0;
assign detect_max[535][18] = (mid_1[4295:4288] > btm_0[4295:4288]) ? 1 : 0;
assign detect_max[535][19] = (mid_1[4295:4288] > btm_0[4303:4296]) ? 1 : 0;
assign detect_max[535][20] = (mid_1[4295:4288] > btm_1[4287:4280]) ? 1 : 0;
assign detect_max[535][21] = (mid_1[4295:4288] > btm_1[4295:4288]) ? 1 : 0;
assign detect_max[535][22] = (mid_1[4295:4288] > btm_1[4303:4296]) ? 1 : 0;
assign detect_max[535][23] = (mid_1[4295:4288] > btm_2[4287:4280]) ? 1 : 0;
assign detect_max[535][24] = (mid_1[4295:4288] > btm_2[4295:4288]) ? 1 : 0;
assign detect_max[535][25] = (mid_1[4295:4288] > btm_2[4303:4296]) ? 1 : 0;

assign detect_max[536][0] = (mid_1[4303:4296] > top_0[4295:4288]) ? 1 : 0;
assign detect_max[536][1] = (mid_1[4303:4296] > top_0[4303:4296]) ? 1 : 0;
assign detect_max[536][2] = (mid_1[4303:4296] > top_0[4311:4304]) ? 1 : 0;
assign detect_max[536][3] = (mid_1[4303:4296] > top_1[4295:4288]) ? 1 : 0;
assign detect_max[536][4] = (mid_1[4303:4296] > top_1[4303:4296]) ? 1 : 0;
assign detect_max[536][5] = (mid_1[4303:4296] > top_1[4311:4304]) ? 1 : 0;
assign detect_max[536][6] = (mid_1[4303:4296] > top_2[4295:4288]) ? 1 : 0;
assign detect_max[536][7] = (mid_1[4303:4296] > top_2[4303:4296]) ? 1 : 0;
assign detect_max[536][8] = (mid_1[4303:4296] > top_2[4311:4304]) ? 1 : 0;
assign detect_max[536][9] = (mid_1[4303:4296] > mid_0[4295:4288]) ? 1 : 0;
assign detect_max[536][10] = (mid_1[4303:4296] > mid_0[4303:4296]) ? 1 : 0;
assign detect_max[536][11] = (mid_1[4303:4296] > mid_0[4311:4304]) ? 1 : 0;
assign detect_max[536][12] = (mid_1[4303:4296] > mid_1[4295:4288]) ? 1 : 0;
assign detect_max[536][13] = (mid_1[4303:4296] > mid_1[4311:4304]) ? 1 : 0;
assign detect_max[536][14] = (mid_1[4303:4296] > mid_2[4295:4288]) ? 1 : 0;
assign detect_max[536][15] = (mid_1[4303:4296] > mid_2[4303:4296]) ? 1 : 0;
assign detect_max[536][16] = (mid_1[4303:4296] > mid_2[4311:4304]) ? 1 : 0;
assign detect_max[536][17] = (mid_1[4303:4296] > btm_0[4295:4288]) ? 1 : 0;
assign detect_max[536][18] = (mid_1[4303:4296] > btm_0[4303:4296]) ? 1 : 0;
assign detect_max[536][19] = (mid_1[4303:4296] > btm_0[4311:4304]) ? 1 : 0;
assign detect_max[536][20] = (mid_1[4303:4296] > btm_1[4295:4288]) ? 1 : 0;
assign detect_max[536][21] = (mid_1[4303:4296] > btm_1[4303:4296]) ? 1 : 0;
assign detect_max[536][22] = (mid_1[4303:4296] > btm_1[4311:4304]) ? 1 : 0;
assign detect_max[536][23] = (mid_1[4303:4296] > btm_2[4295:4288]) ? 1 : 0;
assign detect_max[536][24] = (mid_1[4303:4296] > btm_2[4303:4296]) ? 1 : 0;
assign detect_max[536][25] = (mid_1[4303:4296] > btm_2[4311:4304]) ? 1 : 0;

assign detect_max[537][0] = (mid_1[4311:4304] > top_0[4303:4296]) ? 1 : 0;
assign detect_max[537][1] = (mid_1[4311:4304] > top_0[4311:4304]) ? 1 : 0;
assign detect_max[537][2] = (mid_1[4311:4304] > top_0[4319:4312]) ? 1 : 0;
assign detect_max[537][3] = (mid_1[4311:4304] > top_1[4303:4296]) ? 1 : 0;
assign detect_max[537][4] = (mid_1[4311:4304] > top_1[4311:4304]) ? 1 : 0;
assign detect_max[537][5] = (mid_1[4311:4304] > top_1[4319:4312]) ? 1 : 0;
assign detect_max[537][6] = (mid_1[4311:4304] > top_2[4303:4296]) ? 1 : 0;
assign detect_max[537][7] = (mid_1[4311:4304] > top_2[4311:4304]) ? 1 : 0;
assign detect_max[537][8] = (mid_1[4311:4304] > top_2[4319:4312]) ? 1 : 0;
assign detect_max[537][9] = (mid_1[4311:4304] > mid_0[4303:4296]) ? 1 : 0;
assign detect_max[537][10] = (mid_1[4311:4304] > mid_0[4311:4304]) ? 1 : 0;
assign detect_max[537][11] = (mid_1[4311:4304] > mid_0[4319:4312]) ? 1 : 0;
assign detect_max[537][12] = (mid_1[4311:4304] > mid_1[4303:4296]) ? 1 : 0;
assign detect_max[537][13] = (mid_1[4311:4304] > mid_1[4319:4312]) ? 1 : 0;
assign detect_max[537][14] = (mid_1[4311:4304] > mid_2[4303:4296]) ? 1 : 0;
assign detect_max[537][15] = (mid_1[4311:4304] > mid_2[4311:4304]) ? 1 : 0;
assign detect_max[537][16] = (mid_1[4311:4304] > mid_2[4319:4312]) ? 1 : 0;
assign detect_max[537][17] = (mid_1[4311:4304] > btm_0[4303:4296]) ? 1 : 0;
assign detect_max[537][18] = (mid_1[4311:4304] > btm_0[4311:4304]) ? 1 : 0;
assign detect_max[537][19] = (mid_1[4311:4304] > btm_0[4319:4312]) ? 1 : 0;
assign detect_max[537][20] = (mid_1[4311:4304] > btm_1[4303:4296]) ? 1 : 0;
assign detect_max[537][21] = (mid_1[4311:4304] > btm_1[4311:4304]) ? 1 : 0;
assign detect_max[537][22] = (mid_1[4311:4304] > btm_1[4319:4312]) ? 1 : 0;
assign detect_max[537][23] = (mid_1[4311:4304] > btm_2[4303:4296]) ? 1 : 0;
assign detect_max[537][24] = (mid_1[4311:4304] > btm_2[4311:4304]) ? 1 : 0;
assign detect_max[537][25] = (mid_1[4311:4304] > btm_2[4319:4312]) ? 1 : 0;

assign detect_max[538][0] = (mid_1[4319:4312] > top_0[4311:4304]) ? 1 : 0;
assign detect_max[538][1] = (mid_1[4319:4312] > top_0[4319:4312]) ? 1 : 0;
assign detect_max[538][2] = (mid_1[4319:4312] > top_0[4327:4320]) ? 1 : 0;
assign detect_max[538][3] = (mid_1[4319:4312] > top_1[4311:4304]) ? 1 : 0;
assign detect_max[538][4] = (mid_1[4319:4312] > top_1[4319:4312]) ? 1 : 0;
assign detect_max[538][5] = (mid_1[4319:4312] > top_1[4327:4320]) ? 1 : 0;
assign detect_max[538][6] = (mid_1[4319:4312] > top_2[4311:4304]) ? 1 : 0;
assign detect_max[538][7] = (mid_1[4319:4312] > top_2[4319:4312]) ? 1 : 0;
assign detect_max[538][8] = (mid_1[4319:4312] > top_2[4327:4320]) ? 1 : 0;
assign detect_max[538][9] = (mid_1[4319:4312] > mid_0[4311:4304]) ? 1 : 0;
assign detect_max[538][10] = (mid_1[4319:4312] > mid_0[4319:4312]) ? 1 : 0;
assign detect_max[538][11] = (mid_1[4319:4312] > mid_0[4327:4320]) ? 1 : 0;
assign detect_max[538][12] = (mid_1[4319:4312] > mid_1[4311:4304]) ? 1 : 0;
assign detect_max[538][13] = (mid_1[4319:4312] > mid_1[4327:4320]) ? 1 : 0;
assign detect_max[538][14] = (mid_1[4319:4312] > mid_2[4311:4304]) ? 1 : 0;
assign detect_max[538][15] = (mid_1[4319:4312] > mid_2[4319:4312]) ? 1 : 0;
assign detect_max[538][16] = (mid_1[4319:4312] > mid_2[4327:4320]) ? 1 : 0;
assign detect_max[538][17] = (mid_1[4319:4312] > btm_0[4311:4304]) ? 1 : 0;
assign detect_max[538][18] = (mid_1[4319:4312] > btm_0[4319:4312]) ? 1 : 0;
assign detect_max[538][19] = (mid_1[4319:4312] > btm_0[4327:4320]) ? 1 : 0;
assign detect_max[538][20] = (mid_1[4319:4312] > btm_1[4311:4304]) ? 1 : 0;
assign detect_max[538][21] = (mid_1[4319:4312] > btm_1[4319:4312]) ? 1 : 0;
assign detect_max[538][22] = (mid_1[4319:4312] > btm_1[4327:4320]) ? 1 : 0;
assign detect_max[538][23] = (mid_1[4319:4312] > btm_2[4311:4304]) ? 1 : 0;
assign detect_max[538][24] = (mid_1[4319:4312] > btm_2[4319:4312]) ? 1 : 0;
assign detect_max[538][25] = (mid_1[4319:4312] > btm_2[4327:4320]) ? 1 : 0;

assign detect_max[539][0] = (mid_1[4327:4320] > top_0[4319:4312]) ? 1 : 0;
assign detect_max[539][1] = (mid_1[4327:4320] > top_0[4327:4320]) ? 1 : 0;
assign detect_max[539][2] = (mid_1[4327:4320] > top_0[4335:4328]) ? 1 : 0;
assign detect_max[539][3] = (mid_1[4327:4320] > top_1[4319:4312]) ? 1 : 0;
assign detect_max[539][4] = (mid_1[4327:4320] > top_1[4327:4320]) ? 1 : 0;
assign detect_max[539][5] = (mid_1[4327:4320] > top_1[4335:4328]) ? 1 : 0;
assign detect_max[539][6] = (mid_1[4327:4320] > top_2[4319:4312]) ? 1 : 0;
assign detect_max[539][7] = (mid_1[4327:4320] > top_2[4327:4320]) ? 1 : 0;
assign detect_max[539][8] = (mid_1[4327:4320] > top_2[4335:4328]) ? 1 : 0;
assign detect_max[539][9] = (mid_1[4327:4320] > mid_0[4319:4312]) ? 1 : 0;
assign detect_max[539][10] = (mid_1[4327:4320] > mid_0[4327:4320]) ? 1 : 0;
assign detect_max[539][11] = (mid_1[4327:4320] > mid_0[4335:4328]) ? 1 : 0;
assign detect_max[539][12] = (mid_1[4327:4320] > mid_1[4319:4312]) ? 1 : 0;
assign detect_max[539][13] = (mid_1[4327:4320] > mid_1[4335:4328]) ? 1 : 0;
assign detect_max[539][14] = (mid_1[4327:4320] > mid_2[4319:4312]) ? 1 : 0;
assign detect_max[539][15] = (mid_1[4327:4320] > mid_2[4327:4320]) ? 1 : 0;
assign detect_max[539][16] = (mid_1[4327:4320] > mid_2[4335:4328]) ? 1 : 0;
assign detect_max[539][17] = (mid_1[4327:4320] > btm_0[4319:4312]) ? 1 : 0;
assign detect_max[539][18] = (mid_1[4327:4320] > btm_0[4327:4320]) ? 1 : 0;
assign detect_max[539][19] = (mid_1[4327:4320] > btm_0[4335:4328]) ? 1 : 0;
assign detect_max[539][20] = (mid_1[4327:4320] > btm_1[4319:4312]) ? 1 : 0;
assign detect_max[539][21] = (mid_1[4327:4320] > btm_1[4327:4320]) ? 1 : 0;
assign detect_max[539][22] = (mid_1[4327:4320] > btm_1[4335:4328]) ? 1 : 0;
assign detect_max[539][23] = (mid_1[4327:4320] > btm_2[4319:4312]) ? 1 : 0;
assign detect_max[539][24] = (mid_1[4327:4320] > btm_2[4327:4320]) ? 1 : 0;
assign detect_max[539][25] = (mid_1[4327:4320] > btm_2[4335:4328]) ? 1 : 0;

assign detect_max[540][0] = (mid_1[4335:4328] > top_0[4327:4320]) ? 1 : 0;
assign detect_max[540][1] = (mid_1[4335:4328] > top_0[4335:4328]) ? 1 : 0;
assign detect_max[540][2] = (mid_1[4335:4328] > top_0[4343:4336]) ? 1 : 0;
assign detect_max[540][3] = (mid_1[4335:4328] > top_1[4327:4320]) ? 1 : 0;
assign detect_max[540][4] = (mid_1[4335:4328] > top_1[4335:4328]) ? 1 : 0;
assign detect_max[540][5] = (mid_1[4335:4328] > top_1[4343:4336]) ? 1 : 0;
assign detect_max[540][6] = (mid_1[4335:4328] > top_2[4327:4320]) ? 1 : 0;
assign detect_max[540][7] = (mid_1[4335:4328] > top_2[4335:4328]) ? 1 : 0;
assign detect_max[540][8] = (mid_1[4335:4328] > top_2[4343:4336]) ? 1 : 0;
assign detect_max[540][9] = (mid_1[4335:4328] > mid_0[4327:4320]) ? 1 : 0;
assign detect_max[540][10] = (mid_1[4335:4328] > mid_0[4335:4328]) ? 1 : 0;
assign detect_max[540][11] = (mid_1[4335:4328] > mid_0[4343:4336]) ? 1 : 0;
assign detect_max[540][12] = (mid_1[4335:4328] > mid_1[4327:4320]) ? 1 : 0;
assign detect_max[540][13] = (mid_1[4335:4328] > mid_1[4343:4336]) ? 1 : 0;
assign detect_max[540][14] = (mid_1[4335:4328] > mid_2[4327:4320]) ? 1 : 0;
assign detect_max[540][15] = (mid_1[4335:4328] > mid_2[4335:4328]) ? 1 : 0;
assign detect_max[540][16] = (mid_1[4335:4328] > mid_2[4343:4336]) ? 1 : 0;
assign detect_max[540][17] = (mid_1[4335:4328] > btm_0[4327:4320]) ? 1 : 0;
assign detect_max[540][18] = (mid_1[4335:4328] > btm_0[4335:4328]) ? 1 : 0;
assign detect_max[540][19] = (mid_1[4335:4328] > btm_0[4343:4336]) ? 1 : 0;
assign detect_max[540][20] = (mid_1[4335:4328] > btm_1[4327:4320]) ? 1 : 0;
assign detect_max[540][21] = (mid_1[4335:4328] > btm_1[4335:4328]) ? 1 : 0;
assign detect_max[540][22] = (mid_1[4335:4328] > btm_1[4343:4336]) ? 1 : 0;
assign detect_max[540][23] = (mid_1[4335:4328] > btm_2[4327:4320]) ? 1 : 0;
assign detect_max[540][24] = (mid_1[4335:4328] > btm_2[4335:4328]) ? 1 : 0;
assign detect_max[540][25] = (mid_1[4335:4328] > btm_2[4343:4336]) ? 1 : 0;

assign detect_max[541][0] = (mid_1[4343:4336] > top_0[4335:4328]) ? 1 : 0;
assign detect_max[541][1] = (mid_1[4343:4336] > top_0[4343:4336]) ? 1 : 0;
assign detect_max[541][2] = (mid_1[4343:4336] > top_0[4351:4344]) ? 1 : 0;
assign detect_max[541][3] = (mid_1[4343:4336] > top_1[4335:4328]) ? 1 : 0;
assign detect_max[541][4] = (mid_1[4343:4336] > top_1[4343:4336]) ? 1 : 0;
assign detect_max[541][5] = (mid_1[4343:4336] > top_1[4351:4344]) ? 1 : 0;
assign detect_max[541][6] = (mid_1[4343:4336] > top_2[4335:4328]) ? 1 : 0;
assign detect_max[541][7] = (mid_1[4343:4336] > top_2[4343:4336]) ? 1 : 0;
assign detect_max[541][8] = (mid_1[4343:4336] > top_2[4351:4344]) ? 1 : 0;
assign detect_max[541][9] = (mid_1[4343:4336] > mid_0[4335:4328]) ? 1 : 0;
assign detect_max[541][10] = (mid_1[4343:4336] > mid_0[4343:4336]) ? 1 : 0;
assign detect_max[541][11] = (mid_1[4343:4336] > mid_0[4351:4344]) ? 1 : 0;
assign detect_max[541][12] = (mid_1[4343:4336] > mid_1[4335:4328]) ? 1 : 0;
assign detect_max[541][13] = (mid_1[4343:4336] > mid_1[4351:4344]) ? 1 : 0;
assign detect_max[541][14] = (mid_1[4343:4336] > mid_2[4335:4328]) ? 1 : 0;
assign detect_max[541][15] = (mid_1[4343:4336] > mid_2[4343:4336]) ? 1 : 0;
assign detect_max[541][16] = (mid_1[4343:4336] > mid_2[4351:4344]) ? 1 : 0;
assign detect_max[541][17] = (mid_1[4343:4336] > btm_0[4335:4328]) ? 1 : 0;
assign detect_max[541][18] = (mid_1[4343:4336] > btm_0[4343:4336]) ? 1 : 0;
assign detect_max[541][19] = (mid_1[4343:4336] > btm_0[4351:4344]) ? 1 : 0;
assign detect_max[541][20] = (mid_1[4343:4336] > btm_1[4335:4328]) ? 1 : 0;
assign detect_max[541][21] = (mid_1[4343:4336] > btm_1[4343:4336]) ? 1 : 0;
assign detect_max[541][22] = (mid_1[4343:4336] > btm_1[4351:4344]) ? 1 : 0;
assign detect_max[541][23] = (mid_1[4343:4336] > btm_2[4335:4328]) ? 1 : 0;
assign detect_max[541][24] = (mid_1[4343:4336] > btm_2[4343:4336]) ? 1 : 0;
assign detect_max[541][25] = (mid_1[4343:4336] > btm_2[4351:4344]) ? 1 : 0;

assign detect_max[542][0] = (mid_1[4351:4344] > top_0[4343:4336]) ? 1 : 0;
assign detect_max[542][1] = (mid_1[4351:4344] > top_0[4351:4344]) ? 1 : 0;
assign detect_max[542][2] = (mid_1[4351:4344] > top_0[4359:4352]) ? 1 : 0;
assign detect_max[542][3] = (mid_1[4351:4344] > top_1[4343:4336]) ? 1 : 0;
assign detect_max[542][4] = (mid_1[4351:4344] > top_1[4351:4344]) ? 1 : 0;
assign detect_max[542][5] = (mid_1[4351:4344] > top_1[4359:4352]) ? 1 : 0;
assign detect_max[542][6] = (mid_1[4351:4344] > top_2[4343:4336]) ? 1 : 0;
assign detect_max[542][7] = (mid_1[4351:4344] > top_2[4351:4344]) ? 1 : 0;
assign detect_max[542][8] = (mid_1[4351:4344] > top_2[4359:4352]) ? 1 : 0;
assign detect_max[542][9] = (mid_1[4351:4344] > mid_0[4343:4336]) ? 1 : 0;
assign detect_max[542][10] = (mid_1[4351:4344] > mid_0[4351:4344]) ? 1 : 0;
assign detect_max[542][11] = (mid_1[4351:4344] > mid_0[4359:4352]) ? 1 : 0;
assign detect_max[542][12] = (mid_1[4351:4344] > mid_1[4343:4336]) ? 1 : 0;
assign detect_max[542][13] = (mid_1[4351:4344] > mid_1[4359:4352]) ? 1 : 0;
assign detect_max[542][14] = (mid_1[4351:4344] > mid_2[4343:4336]) ? 1 : 0;
assign detect_max[542][15] = (mid_1[4351:4344] > mid_2[4351:4344]) ? 1 : 0;
assign detect_max[542][16] = (mid_1[4351:4344] > mid_2[4359:4352]) ? 1 : 0;
assign detect_max[542][17] = (mid_1[4351:4344] > btm_0[4343:4336]) ? 1 : 0;
assign detect_max[542][18] = (mid_1[4351:4344] > btm_0[4351:4344]) ? 1 : 0;
assign detect_max[542][19] = (mid_1[4351:4344] > btm_0[4359:4352]) ? 1 : 0;
assign detect_max[542][20] = (mid_1[4351:4344] > btm_1[4343:4336]) ? 1 : 0;
assign detect_max[542][21] = (mid_1[4351:4344] > btm_1[4351:4344]) ? 1 : 0;
assign detect_max[542][22] = (mid_1[4351:4344] > btm_1[4359:4352]) ? 1 : 0;
assign detect_max[542][23] = (mid_1[4351:4344] > btm_2[4343:4336]) ? 1 : 0;
assign detect_max[542][24] = (mid_1[4351:4344] > btm_2[4351:4344]) ? 1 : 0;
assign detect_max[542][25] = (mid_1[4351:4344] > btm_2[4359:4352]) ? 1 : 0;

assign detect_max[543][0] = (mid_1[4359:4352] > top_0[4351:4344]) ? 1 : 0;
assign detect_max[543][1] = (mid_1[4359:4352] > top_0[4359:4352]) ? 1 : 0;
assign detect_max[543][2] = (mid_1[4359:4352] > top_0[4367:4360]) ? 1 : 0;
assign detect_max[543][3] = (mid_1[4359:4352] > top_1[4351:4344]) ? 1 : 0;
assign detect_max[543][4] = (mid_1[4359:4352] > top_1[4359:4352]) ? 1 : 0;
assign detect_max[543][5] = (mid_1[4359:4352] > top_1[4367:4360]) ? 1 : 0;
assign detect_max[543][6] = (mid_1[4359:4352] > top_2[4351:4344]) ? 1 : 0;
assign detect_max[543][7] = (mid_1[4359:4352] > top_2[4359:4352]) ? 1 : 0;
assign detect_max[543][8] = (mid_1[4359:4352] > top_2[4367:4360]) ? 1 : 0;
assign detect_max[543][9] = (mid_1[4359:4352] > mid_0[4351:4344]) ? 1 : 0;
assign detect_max[543][10] = (mid_1[4359:4352] > mid_0[4359:4352]) ? 1 : 0;
assign detect_max[543][11] = (mid_1[4359:4352] > mid_0[4367:4360]) ? 1 : 0;
assign detect_max[543][12] = (mid_1[4359:4352] > mid_1[4351:4344]) ? 1 : 0;
assign detect_max[543][13] = (mid_1[4359:4352] > mid_1[4367:4360]) ? 1 : 0;
assign detect_max[543][14] = (mid_1[4359:4352] > mid_2[4351:4344]) ? 1 : 0;
assign detect_max[543][15] = (mid_1[4359:4352] > mid_2[4359:4352]) ? 1 : 0;
assign detect_max[543][16] = (mid_1[4359:4352] > mid_2[4367:4360]) ? 1 : 0;
assign detect_max[543][17] = (mid_1[4359:4352] > btm_0[4351:4344]) ? 1 : 0;
assign detect_max[543][18] = (mid_1[4359:4352] > btm_0[4359:4352]) ? 1 : 0;
assign detect_max[543][19] = (mid_1[4359:4352] > btm_0[4367:4360]) ? 1 : 0;
assign detect_max[543][20] = (mid_1[4359:4352] > btm_1[4351:4344]) ? 1 : 0;
assign detect_max[543][21] = (mid_1[4359:4352] > btm_1[4359:4352]) ? 1 : 0;
assign detect_max[543][22] = (mid_1[4359:4352] > btm_1[4367:4360]) ? 1 : 0;
assign detect_max[543][23] = (mid_1[4359:4352] > btm_2[4351:4344]) ? 1 : 0;
assign detect_max[543][24] = (mid_1[4359:4352] > btm_2[4359:4352]) ? 1 : 0;
assign detect_max[543][25] = (mid_1[4359:4352] > btm_2[4367:4360]) ? 1 : 0;

assign detect_max[544][0] = (mid_1[4367:4360] > top_0[4359:4352]) ? 1 : 0;
assign detect_max[544][1] = (mid_1[4367:4360] > top_0[4367:4360]) ? 1 : 0;
assign detect_max[544][2] = (mid_1[4367:4360] > top_0[4375:4368]) ? 1 : 0;
assign detect_max[544][3] = (mid_1[4367:4360] > top_1[4359:4352]) ? 1 : 0;
assign detect_max[544][4] = (mid_1[4367:4360] > top_1[4367:4360]) ? 1 : 0;
assign detect_max[544][5] = (mid_1[4367:4360] > top_1[4375:4368]) ? 1 : 0;
assign detect_max[544][6] = (mid_1[4367:4360] > top_2[4359:4352]) ? 1 : 0;
assign detect_max[544][7] = (mid_1[4367:4360] > top_2[4367:4360]) ? 1 : 0;
assign detect_max[544][8] = (mid_1[4367:4360] > top_2[4375:4368]) ? 1 : 0;
assign detect_max[544][9] = (mid_1[4367:4360] > mid_0[4359:4352]) ? 1 : 0;
assign detect_max[544][10] = (mid_1[4367:4360] > mid_0[4367:4360]) ? 1 : 0;
assign detect_max[544][11] = (mid_1[4367:4360] > mid_0[4375:4368]) ? 1 : 0;
assign detect_max[544][12] = (mid_1[4367:4360] > mid_1[4359:4352]) ? 1 : 0;
assign detect_max[544][13] = (mid_1[4367:4360] > mid_1[4375:4368]) ? 1 : 0;
assign detect_max[544][14] = (mid_1[4367:4360] > mid_2[4359:4352]) ? 1 : 0;
assign detect_max[544][15] = (mid_1[4367:4360] > mid_2[4367:4360]) ? 1 : 0;
assign detect_max[544][16] = (mid_1[4367:4360] > mid_2[4375:4368]) ? 1 : 0;
assign detect_max[544][17] = (mid_1[4367:4360] > btm_0[4359:4352]) ? 1 : 0;
assign detect_max[544][18] = (mid_1[4367:4360] > btm_0[4367:4360]) ? 1 : 0;
assign detect_max[544][19] = (mid_1[4367:4360] > btm_0[4375:4368]) ? 1 : 0;
assign detect_max[544][20] = (mid_1[4367:4360] > btm_1[4359:4352]) ? 1 : 0;
assign detect_max[544][21] = (mid_1[4367:4360] > btm_1[4367:4360]) ? 1 : 0;
assign detect_max[544][22] = (mid_1[4367:4360] > btm_1[4375:4368]) ? 1 : 0;
assign detect_max[544][23] = (mid_1[4367:4360] > btm_2[4359:4352]) ? 1 : 0;
assign detect_max[544][24] = (mid_1[4367:4360] > btm_2[4367:4360]) ? 1 : 0;
assign detect_max[544][25] = (mid_1[4367:4360] > btm_2[4375:4368]) ? 1 : 0;

assign detect_max[545][0] = (mid_1[4375:4368] > top_0[4367:4360]) ? 1 : 0;
assign detect_max[545][1] = (mid_1[4375:4368] > top_0[4375:4368]) ? 1 : 0;
assign detect_max[545][2] = (mid_1[4375:4368] > top_0[4383:4376]) ? 1 : 0;
assign detect_max[545][3] = (mid_1[4375:4368] > top_1[4367:4360]) ? 1 : 0;
assign detect_max[545][4] = (mid_1[4375:4368] > top_1[4375:4368]) ? 1 : 0;
assign detect_max[545][5] = (mid_1[4375:4368] > top_1[4383:4376]) ? 1 : 0;
assign detect_max[545][6] = (mid_1[4375:4368] > top_2[4367:4360]) ? 1 : 0;
assign detect_max[545][7] = (mid_1[4375:4368] > top_2[4375:4368]) ? 1 : 0;
assign detect_max[545][8] = (mid_1[4375:4368] > top_2[4383:4376]) ? 1 : 0;
assign detect_max[545][9] = (mid_1[4375:4368] > mid_0[4367:4360]) ? 1 : 0;
assign detect_max[545][10] = (mid_1[4375:4368] > mid_0[4375:4368]) ? 1 : 0;
assign detect_max[545][11] = (mid_1[4375:4368] > mid_0[4383:4376]) ? 1 : 0;
assign detect_max[545][12] = (mid_1[4375:4368] > mid_1[4367:4360]) ? 1 : 0;
assign detect_max[545][13] = (mid_1[4375:4368] > mid_1[4383:4376]) ? 1 : 0;
assign detect_max[545][14] = (mid_1[4375:4368] > mid_2[4367:4360]) ? 1 : 0;
assign detect_max[545][15] = (mid_1[4375:4368] > mid_2[4375:4368]) ? 1 : 0;
assign detect_max[545][16] = (mid_1[4375:4368] > mid_2[4383:4376]) ? 1 : 0;
assign detect_max[545][17] = (mid_1[4375:4368] > btm_0[4367:4360]) ? 1 : 0;
assign detect_max[545][18] = (mid_1[4375:4368] > btm_0[4375:4368]) ? 1 : 0;
assign detect_max[545][19] = (mid_1[4375:4368] > btm_0[4383:4376]) ? 1 : 0;
assign detect_max[545][20] = (mid_1[4375:4368] > btm_1[4367:4360]) ? 1 : 0;
assign detect_max[545][21] = (mid_1[4375:4368] > btm_1[4375:4368]) ? 1 : 0;
assign detect_max[545][22] = (mid_1[4375:4368] > btm_1[4383:4376]) ? 1 : 0;
assign detect_max[545][23] = (mid_1[4375:4368] > btm_2[4367:4360]) ? 1 : 0;
assign detect_max[545][24] = (mid_1[4375:4368] > btm_2[4375:4368]) ? 1 : 0;
assign detect_max[545][25] = (mid_1[4375:4368] > btm_2[4383:4376]) ? 1 : 0;

assign detect_max[546][0] = (mid_1[4383:4376] > top_0[4375:4368]) ? 1 : 0;
assign detect_max[546][1] = (mid_1[4383:4376] > top_0[4383:4376]) ? 1 : 0;
assign detect_max[546][2] = (mid_1[4383:4376] > top_0[4391:4384]) ? 1 : 0;
assign detect_max[546][3] = (mid_1[4383:4376] > top_1[4375:4368]) ? 1 : 0;
assign detect_max[546][4] = (mid_1[4383:4376] > top_1[4383:4376]) ? 1 : 0;
assign detect_max[546][5] = (mid_1[4383:4376] > top_1[4391:4384]) ? 1 : 0;
assign detect_max[546][6] = (mid_1[4383:4376] > top_2[4375:4368]) ? 1 : 0;
assign detect_max[546][7] = (mid_1[4383:4376] > top_2[4383:4376]) ? 1 : 0;
assign detect_max[546][8] = (mid_1[4383:4376] > top_2[4391:4384]) ? 1 : 0;
assign detect_max[546][9] = (mid_1[4383:4376] > mid_0[4375:4368]) ? 1 : 0;
assign detect_max[546][10] = (mid_1[4383:4376] > mid_0[4383:4376]) ? 1 : 0;
assign detect_max[546][11] = (mid_1[4383:4376] > mid_0[4391:4384]) ? 1 : 0;
assign detect_max[546][12] = (mid_1[4383:4376] > mid_1[4375:4368]) ? 1 : 0;
assign detect_max[546][13] = (mid_1[4383:4376] > mid_1[4391:4384]) ? 1 : 0;
assign detect_max[546][14] = (mid_1[4383:4376] > mid_2[4375:4368]) ? 1 : 0;
assign detect_max[546][15] = (mid_1[4383:4376] > mid_2[4383:4376]) ? 1 : 0;
assign detect_max[546][16] = (mid_1[4383:4376] > mid_2[4391:4384]) ? 1 : 0;
assign detect_max[546][17] = (mid_1[4383:4376] > btm_0[4375:4368]) ? 1 : 0;
assign detect_max[546][18] = (mid_1[4383:4376] > btm_0[4383:4376]) ? 1 : 0;
assign detect_max[546][19] = (mid_1[4383:4376] > btm_0[4391:4384]) ? 1 : 0;
assign detect_max[546][20] = (mid_1[4383:4376] > btm_1[4375:4368]) ? 1 : 0;
assign detect_max[546][21] = (mid_1[4383:4376] > btm_1[4383:4376]) ? 1 : 0;
assign detect_max[546][22] = (mid_1[4383:4376] > btm_1[4391:4384]) ? 1 : 0;
assign detect_max[546][23] = (mid_1[4383:4376] > btm_2[4375:4368]) ? 1 : 0;
assign detect_max[546][24] = (mid_1[4383:4376] > btm_2[4383:4376]) ? 1 : 0;
assign detect_max[546][25] = (mid_1[4383:4376] > btm_2[4391:4384]) ? 1 : 0;

assign detect_max[547][0] = (mid_1[4391:4384] > top_0[4383:4376]) ? 1 : 0;
assign detect_max[547][1] = (mid_1[4391:4384] > top_0[4391:4384]) ? 1 : 0;
assign detect_max[547][2] = (mid_1[4391:4384] > top_0[4399:4392]) ? 1 : 0;
assign detect_max[547][3] = (mid_1[4391:4384] > top_1[4383:4376]) ? 1 : 0;
assign detect_max[547][4] = (mid_1[4391:4384] > top_1[4391:4384]) ? 1 : 0;
assign detect_max[547][5] = (mid_1[4391:4384] > top_1[4399:4392]) ? 1 : 0;
assign detect_max[547][6] = (mid_1[4391:4384] > top_2[4383:4376]) ? 1 : 0;
assign detect_max[547][7] = (mid_1[4391:4384] > top_2[4391:4384]) ? 1 : 0;
assign detect_max[547][8] = (mid_1[4391:4384] > top_2[4399:4392]) ? 1 : 0;
assign detect_max[547][9] = (mid_1[4391:4384] > mid_0[4383:4376]) ? 1 : 0;
assign detect_max[547][10] = (mid_1[4391:4384] > mid_0[4391:4384]) ? 1 : 0;
assign detect_max[547][11] = (mid_1[4391:4384] > mid_0[4399:4392]) ? 1 : 0;
assign detect_max[547][12] = (mid_1[4391:4384] > mid_1[4383:4376]) ? 1 : 0;
assign detect_max[547][13] = (mid_1[4391:4384] > mid_1[4399:4392]) ? 1 : 0;
assign detect_max[547][14] = (mid_1[4391:4384] > mid_2[4383:4376]) ? 1 : 0;
assign detect_max[547][15] = (mid_1[4391:4384] > mid_2[4391:4384]) ? 1 : 0;
assign detect_max[547][16] = (mid_1[4391:4384] > mid_2[4399:4392]) ? 1 : 0;
assign detect_max[547][17] = (mid_1[4391:4384] > btm_0[4383:4376]) ? 1 : 0;
assign detect_max[547][18] = (mid_1[4391:4384] > btm_0[4391:4384]) ? 1 : 0;
assign detect_max[547][19] = (mid_1[4391:4384] > btm_0[4399:4392]) ? 1 : 0;
assign detect_max[547][20] = (mid_1[4391:4384] > btm_1[4383:4376]) ? 1 : 0;
assign detect_max[547][21] = (mid_1[4391:4384] > btm_1[4391:4384]) ? 1 : 0;
assign detect_max[547][22] = (mid_1[4391:4384] > btm_1[4399:4392]) ? 1 : 0;
assign detect_max[547][23] = (mid_1[4391:4384] > btm_2[4383:4376]) ? 1 : 0;
assign detect_max[547][24] = (mid_1[4391:4384] > btm_2[4391:4384]) ? 1 : 0;
assign detect_max[547][25] = (mid_1[4391:4384] > btm_2[4399:4392]) ? 1 : 0;

assign detect_max[548][0] = (mid_1[4399:4392] > top_0[4391:4384]) ? 1 : 0;
assign detect_max[548][1] = (mid_1[4399:4392] > top_0[4399:4392]) ? 1 : 0;
assign detect_max[548][2] = (mid_1[4399:4392] > top_0[4407:4400]) ? 1 : 0;
assign detect_max[548][3] = (mid_1[4399:4392] > top_1[4391:4384]) ? 1 : 0;
assign detect_max[548][4] = (mid_1[4399:4392] > top_1[4399:4392]) ? 1 : 0;
assign detect_max[548][5] = (mid_1[4399:4392] > top_1[4407:4400]) ? 1 : 0;
assign detect_max[548][6] = (mid_1[4399:4392] > top_2[4391:4384]) ? 1 : 0;
assign detect_max[548][7] = (mid_1[4399:4392] > top_2[4399:4392]) ? 1 : 0;
assign detect_max[548][8] = (mid_1[4399:4392] > top_2[4407:4400]) ? 1 : 0;
assign detect_max[548][9] = (mid_1[4399:4392] > mid_0[4391:4384]) ? 1 : 0;
assign detect_max[548][10] = (mid_1[4399:4392] > mid_0[4399:4392]) ? 1 : 0;
assign detect_max[548][11] = (mid_1[4399:4392] > mid_0[4407:4400]) ? 1 : 0;
assign detect_max[548][12] = (mid_1[4399:4392] > mid_1[4391:4384]) ? 1 : 0;
assign detect_max[548][13] = (mid_1[4399:4392] > mid_1[4407:4400]) ? 1 : 0;
assign detect_max[548][14] = (mid_1[4399:4392] > mid_2[4391:4384]) ? 1 : 0;
assign detect_max[548][15] = (mid_1[4399:4392] > mid_2[4399:4392]) ? 1 : 0;
assign detect_max[548][16] = (mid_1[4399:4392] > mid_2[4407:4400]) ? 1 : 0;
assign detect_max[548][17] = (mid_1[4399:4392] > btm_0[4391:4384]) ? 1 : 0;
assign detect_max[548][18] = (mid_1[4399:4392] > btm_0[4399:4392]) ? 1 : 0;
assign detect_max[548][19] = (mid_1[4399:4392] > btm_0[4407:4400]) ? 1 : 0;
assign detect_max[548][20] = (mid_1[4399:4392] > btm_1[4391:4384]) ? 1 : 0;
assign detect_max[548][21] = (mid_1[4399:4392] > btm_1[4399:4392]) ? 1 : 0;
assign detect_max[548][22] = (mid_1[4399:4392] > btm_1[4407:4400]) ? 1 : 0;
assign detect_max[548][23] = (mid_1[4399:4392] > btm_2[4391:4384]) ? 1 : 0;
assign detect_max[548][24] = (mid_1[4399:4392] > btm_2[4399:4392]) ? 1 : 0;
assign detect_max[548][25] = (mid_1[4399:4392] > btm_2[4407:4400]) ? 1 : 0;

assign detect_max[549][0] = (mid_1[4407:4400] > top_0[4399:4392]) ? 1 : 0;
assign detect_max[549][1] = (mid_1[4407:4400] > top_0[4407:4400]) ? 1 : 0;
assign detect_max[549][2] = (mid_1[4407:4400] > top_0[4415:4408]) ? 1 : 0;
assign detect_max[549][3] = (mid_1[4407:4400] > top_1[4399:4392]) ? 1 : 0;
assign detect_max[549][4] = (mid_1[4407:4400] > top_1[4407:4400]) ? 1 : 0;
assign detect_max[549][5] = (mid_1[4407:4400] > top_1[4415:4408]) ? 1 : 0;
assign detect_max[549][6] = (mid_1[4407:4400] > top_2[4399:4392]) ? 1 : 0;
assign detect_max[549][7] = (mid_1[4407:4400] > top_2[4407:4400]) ? 1 : 0;
assign detect_max[549][8] = (mid_1[4407:4400] > top_2[4415:4408]) ? 1 : 0;
assign detect_max[549][9] = (mid_1[4407:4400] > mid_0[4399:4392]) ? 1 : 0;
assign detect_max[549][10] = (mid_1[4407:4400] > mid_0[4407:4400]) ? 1 : 0;
assign detect_max[549][11] = (mid_1[4407:4400] > mid_0[4415:4408]) ? 1 : 0;
assign detect_max[549][12] = (mid_1[4407:4400] > mid_1[4399:4392]) ? 1 : 0;
assign detect_max[549][13] = (mid_1[4407:4400] > mid_1[4415:4408]) ? 1 : 0;
assign detect_max[549][14] = (mid_1[4407:4400] > mid_2[4399:4392]) ? 1 : 0;
assign detect_max[549][15] = (mid_1[4407:4400] > mid_2[4407:4400]) ? 1 : 0;
assign detect_max[549][16] = (mid_1[4407:4400] > mid_2[4415:4408]) ? 1 : 0;
assign detect_max[549][17] = (mid_1[4407:4400] > btm_0[4399:4392]) ? 1 : 0;
assign detect_max[549][18] = (mid_1[4407:4400] > btm_0[4407:4400]) ? 1 : 0;
assign detect_max[549][19] = (mid_1[4407:4400] > btm_0[4415:4408]) ? 1 : 0;
assign detect_max[549][20] = (mid_1[4407:4400] > btm_1[4399:4392]) ? 1 : 0;
assign detect_max[549][21] = (mid_1[4407:4400] > btm_1[4407:4400]) ? 1 : 0;
assign detect_max[549][22] = (mid_1[4407:4400] > btm_1[4415:4408]) ? 1 : 0;
assign detect_max[549][23] = (mid_1[4407:4400] > btm_2[4399:4392]) ? 1 : 0;
assign detect_max[549][24] = (mid_1[4407:4400] > btm_2[4407:4400]) ? 1 : 0;
assign detect_max[549][25] = (mid_1[4407:4400] > btm_2[4415:4408]) ? 1 : 0;

assign detect_max[550][0] = (mid_1[4415:4408] > top_0[4407:4400]) ? 1 : 0;
assign detect_max[550][1] = (mid_1[4415:4408] > top_0[4415:4408]) ? 1 : 0;
assign detect_max[550][2] = (mid_1[4415:4408] > top_0[4423:4416]) ? 1 : 0;
assign detect_max[550][3] = (mid_1[4415:4408] > top_1[4407:4400]) ? 1 : 0;
assign detect_max[550][4] = (mid_1[4415:4408] > top_1[4415:4408]) ? 1 : 0;
assign detect_max[550][5] = (mid_1[4415:4408] > top_1[4423:4416]) ? 1 : 0;
assign detect_max[550][6] = (mid_1[4415:4408] > top_2[4407:4400]) ? 1 : 0;
assign detect_max[550][7] = (mid_1[4415:4408] > top_2[4415:4408]) ? 1 : 0;
assign detect_max[550][8] = (mid_1[4415:4408] > top_2[4423:4416]) ? 1 : 0;
assign detect_max[550][9] = (mid_1[4415:4408] > mid_0[4407:4400]) ? 1 : 0;
assign detect_max[550][10] = (mid_1[4415:4408] > mid_0[4415:4408]) ? 1 : 0;
assign detect_max[550][11] = (mid_1[4415:4408] > mid_0[4423:4416]) ? 1 : 0;
assign detect_max[550][12] = (mid_1[4415:4408] > mid_1[4407:4400]) ? 1 : 0;
assign detect_max[550][13] = (mid_1[4415:4408] > mid_1[4423:4416]) ? 1 : 0;
assign detect_max[550][14] = (mid_1[4415:4408] > mid_2[4407:4400]) ? 1 : 0;
assign detect_max[550][15] = (mid_1[4415:4408] > mid_2[4415:4408]) ? 1 : 0;
assign detect_max[550][16] = (mid_1[4415:4408] > mid_2[4423:4416]) ? 1 : 0;
assign detect_max[550][17] = (mid_1[4415:4408] > btm_0[4407:4400]) ? 1 : 0;
assign detect_max[550][18] = (mid_1[4415:4408] > btm_0[4415:4408]) ? 1 : 0;
assign detect_max[550][19] = (mid_1[4415:4408] > btm_0[4423:4416]) ? 1 : 0;
assign detect_max[550][20] = (mid_1[4415:4408] > btm_1[4407:4400]) ? 1 : 0;
assign detect_max[550][21] = (mid_1[4415:4408] > btm_1[4415:4408]) ? 1 : 0;
assign detect_max[550][22] = (mid_1[4415:4408] > btm_1[4423:4416]) ? 1 : 0;
assign detect_max[550][23] = (mid_1[4415:4408] > btm_2[4407:4400]) ? 1 : 0;
assign detect_max[550][24] = (mid_1[4415:4408] > btm_2[4415:4408]) ? 1 : 0;
assign detect_max[550][25] = (mid_1[4415:4408] > btm_2[4423:4416]) ? 1 : 0;

assign detect_max[551][0] = (mid_1[4423:4416] > top_0[4415:4408]) ? 1 : 0;
assign detect_max[551][1] = (mid_1[4423:4416] > top_0[4423:4416]) ? 1 : 0;
assign detect_max[551][2] = (mid_1[4423:4416] > top_0[4431:4424]) ? 1 : 0;
assign detect_max[551][3] = (mid_1[4423:4416] > top_1[4415:4408]) ? 1 : 0;
assign detect_max[551][4] = (mid_1[4423:4416] > top_1[4423:4416]) ? 1 : 0;
assign detect_max[551][5] = (mid_1[4423:4416] > top_1[4431:4424]) ? 1 : 0;
assign detect_max[551][6] = (mid_1[4423:4416] > top_2[4415:4408]) ? 1 : 0;
assign detect_max[551][7] = (mid_1[4423:4416] > top_2[4423:4416]) ? 1 : 0;
assign detect_max[551][8] = (mid_1[4423:4416] > top_2[4431:4424]) ? 1 : 0;
assign detect_max[551][9] = (mid_1[4423:4416] > mid_0[4415:4408]) ? 1 : 0;
assign detect_max[551][10] = (mid_1[4423:4416] > mid_0[4423:4416]) ? 1 : 0;
assign detect_max[551][11] = (mid_1[4423:4416] > mid_0[4431:4424]) ? 1 : 0;
assign detect_max[551][12] = (mid_1[4423:4416] > mid_1[4415:4408]) ? 1 : 0;
assign detect_max[551][13] = (mid_1[4423:4416] > mid_1[4431:4424]) ? 1 : 0;
assign detect_max[551][14] = (mid_1[4423:4416] > mid_2[4415:4408]) ? 1 : 0;
assign detect_max[551][15] = (mid_1[4423:4416] > mid_2[4423:4416]) ? 1 : 0;
assign detect_max[551][16] = (mid_1[4423:4416] > mid_2[4431:4424]) ? 1 : 0;
assign detect_max[551][17] = (mid_1[4423:4416] > btm_0[4415:4408]) ? 1 : 0;
assign detect_max[551][18] = (mid_1[4423:4416] > btm_0[4423:4416]) ? 1 : 0;
assign detect_max[551][19] = (mid_1[4423:4416] > btm_0[4431:4424]) ? 1 : 0;
assign detect_max[551][20] = (mid_1[4423:4416] > btm_1[4415:4408]) ? 1 : 0;
assign detect_max[551][21] = (mid_1[4423:4416] > btm_1[4423:4416]) ? 1 : 0;
assign detect_max[551][22] = (mid_1[4423:4416] > btm_1[4431:4424]) ? 1 : 0;
assign detect_max[551][23] = (mid_1[4423:4416] > btm_2[4415:4408]) ? 1 : 0;
assign detect_max[551][24] = (mid_1[4423:4416] > btm_2[4423:4416]) ? 1 : 0;
assign detect_max[551][25] = (mid_1[4423:4416] > btm_2[4431:4424]) ? 1 : 0;

assign detect_max[552][0] = (mid_1[4431:4424] > top_0[4423:4416]) ? 1 : 0;
assign detect_max[552][1] = (mid_1[4431:4424] > top_0[4431:4424]) ? 1 : 0;
assign detect_max[552][2] = (mid_1[4431:4424] > top_0[4439:4432]) ? 1 : 0;
assign detect_max[552][3] = (mid_1[4431:4424] > top_1[4423:4416]) ? 1 : 0;
assign detect_max[552][4] = (mid_1[4431:4424] > top_1[4431:4424]) ? 1 : 0;
assign detect_max[552][5] = (mid_1[4431:4424] > top_1[4439:4432]) ? 1 : 0;
assign detect_max[552][6] = (mid_1[4431:4424] > top_2[4423:4416]) ? 1 : 0;
assign detect_max[552][7] = (mid_1[4431:4424] > top_2[4431:4424]) ? 1 : 0;
assign detect_max[552][8] = (mid_1[4431:4424] > top_2[4439:4432]) ? 1 : 0;
assign detect_max[552][9] = (mid_1[4431:4424] > mid_0[4423:4416]) ? 1 : 0;
assign detect_max[552][10] = (mid_1[4431:4424] > mid_0[4431:4424]) ? 1 : 0;
assign detect_max[552][11] = (mid_1[4431:4424] > mid_0[4439:4432]) ? 1 : 0;
assign detect_max[552][12] = (mid_1[4431:4424] > mid_1[4423:4416]) ? 1 : 0;
assign detect_max[552][13] = (mid_1[4431:4424] > mid_1[4439:4432]) ? 1 : 0;
assign detect_max[552][14] = (mid_1[4431:4424] > mid_2[4423:4416]) ? 1 : 0;
assign detect_max[552][15] = (mid_1[4431:4424] > mid_2[4431:4424]) ? 1 : 0;
assign detect_max[552][16] = (mid_1[4431:4424] > mid_2[4439:4432]) ? 1 : 0;
assign detect_max[552][17] = (mid_1[4431:4424] > btm_0[4423:4416]) ? 1 : 0;
assign detect_max[552][18] = (mid_1[4431:4424] > btm_0[4431:4424]) ? 1 : 0;
assign detect_max[552][19] = (mid_1[4431:4424] > btm_0[4439:4432]) ? 1 : 0;
assign detect_max[552][20] = (mid_1[4431:4424] > btm_1[4423:4416]) ? 1 : 0;
assign detect_max[552][21] = (mid_1[4431:4424] > btm_1[4431:4424]) ? 1 : 0;
assign detect_max[552][22] = (mid_1[4431:4424] > btm_1[4439:4432]) ? 1 : 0;
assign detect_max[552][23] = (mid_1[4431:4424] > btm_2[4423:4416]) ? 1 : 0;
assign detect_max[552][24] = (mid_1[4431:4424] > btm_2[4431:4424]) ? 1 : 0;
assign detect_max[552][25] = (mid_1[4431:4424] > btm_2[4439:4432]) ? 1 : 0;

assign detect_max[553][0] = (mid_1[4439:4432] > top_0[4431:4424]) ? 1 : 0;
assign detect_max[553][1] = (mid_1[4439:4432] > top_0[4439:4432]) ? 1 : 0;
assign detect_max[553][2] = (mid_1[4439:4432] > top_0[4447:4440]) ? 1 : 0;
assign detect_max[553][3] = (mid_1[4439:4432] > top_1[4431:4424]) ? 1 : 0;
assign detect_max[553][4] = (mid_1[4439:4432] > top_1[4439:4432]) ? 1 : 0;
assign detect_max[553][5] = (mid_1[4439:4432] > top_1[4447:4440]) ? 1 : 0;
assign detect_max[553][6] = (mid_1[4439:4432] > top_2[4431:4424]) ? 1 : 0;
assign detect_max[553][7] = (mid_1[4439:4432] > top_2[4439:4432]) ? 1 : 0;
assign detect_max[553][8] = (mid_1[4439:4432] > top_2[4447:4440]) ? 1 : 0;
assign detect_max[553][9] = (mid_1[4439:4432] > mid_0[4431:4424]) ? 1 : 0;
assign detect_max[553][10] = (mid_1[4439:4432] > mid_0[4439:4432]) ? 1 : 0;
assign detect_max[553][11] = (mid_1[4439:4432] > mid_0[4447:4440]) ? 1 : 0;
assign detect_max[553][12] = (mid_1[4439:4432] > mid_1[4431:4424]) ? 1 : 0;
assign detect_max[553][13] = (mid_1[4439:4432] > mid_1[4447:4440]) ? 1 : 0;
assign detect_max[553][14] = (mid_1[4439:4432] > mid_2[4431:4424]) ? 1 : 0;
assign detect_max[553][15] = (mid_1[4439:4432] > mid_2[4439:4432]) ? 1 : 0;
assign detect_max[553][16] = (mid_1[4439:4432] > mid_2[4447:4440]) ? 1 : 0;
assign detect_max[553][17] = (mid_1[4439:4432] > btm_0[4431:4424]) ? 1 : 0;
assign detect_max[553][18] = (mid_1[4439:4432] > btm_0[4439:4432]) ? 1 : 0;
assign detect_max[553][19] = (mid_1[4439:4432] > btm_0[4447:4440]) ? 1 : 0;
assign detect_max[553][20] = (mid_1[4439:4432] > btm_1[4431:4424]) ? 1 : 0;
assign detect_max[553][21] = (mid_1[4439:4432] > btm_1[4439:4432]) ? 1 : 0;
assign detect_max[553][22] = (mid_1[4439:4432] > btm_1[4447:4440]) ? 1 : 0;
assign detect_max[553][23] = (mid_1[4439:4432] > btm_2[4431:4424]) ? 1 : 0;
assign detect_max[553][24] = (mid_1[4439:4432] > btm_2[4439:4432]) ? 1 : 0;
assign detect_max[553][25] = (mid_1[4439:4432] > btm_2[4447:4440]) ? 1 : 0;

assign detect_max[554][0] = (mid_1[4447:4440] > top_0[4439:4432]) ? 1 : 0;
assign detect_max[554][1] = (mid_1[4447:4440] > top_0[4447:4440]) ? 1 : 0;
assign detect_max[554][2] = (mid_1[4447:4440] > top_0[4455:4448]) ? 1 : 0;
assign detect_max[554][3] = (mid_1[4447:4440] > top_1[4439:4432]) ? 1 : 0;
assign detect_max[554][4] = (mid_1[4447:4440] > top_1[4447:4440]) ? 1 : 0;
assign detect_max[554][5] = (mid_1[4447:4440] > top_1[4455:4448]) ? 1 : 0;
assign detect_max[554][6] = (mid_1[4447:4440] > top_2[4439:4432]) ? 1 : 0;
assign detect_max[554][7] = (mid_1[4447:4440] > top_2[4447:4440]) ? 1 : 0;
assign detect_max[554][8] = (mid_1[4447:4440] > top_2[4455:4448]) ? 1 : 0;
assign detect_max[554][9] = (mid_1[4447:4440] > mid_0[4439:4432]) ? 1 : 0;
assign detect_max[554][10] = (mid_1[4447:4440] > mid_0[4447:4440]) ? 1 : 0;
assign detect_max[554][11] = (mid_1[4447:4440] > mid_0[4455:4448]) ? 1 : 0;
assign detect_max[554][12] = (mid_1[4447:4440] > mid_1[4439:4432]) ? 1 : 0;
assign detect_max[554][13] = (mid_1[4447:4440] > mid_1[4455:4448]) ? 1 : 0;
assign detect_max[554][14] = (mid_1[4447:4440] > mid_2[4439:4432]) ? 1 : 0;
assign detect_max[554][15] = (mid_1[4447:4440] > mid_2[4447:4440]) ? 1 : 0;
assign detect_max[554][16] = (mid_1[4447:4440] > mid_2[4455:4448]) ? 1 : 0;
assign detect_max[554][17] = (mid_1[4447:4440] > btm_0[4439:4432]) ? 1 : 0;
assign detect_max[554][18] = (mid_1[4447:4440] > btm_0[4447:4440]) ? 1 : 0;
assign detect_max[554][19] = (mid_1[4447:4440] > btm_0[4455:4448]) ? 1 : 0;
assign detect_max[554][20] = (mid_1[4447:4440] > btm_1[4439:4432]) ? 1 : 0;
assign detect_max[554][21] = (mid_1[4447:4440] > btm_1[4447:4440]) ? 1 : 0;
assign detect_max[554][22] = (mid_1[4447:4440] > btm_1[4455:4448]) ? 1 : 0;
assign detect_max[554][23] = (mid_1[4447:4440] > btm_2[4439:4432]) ? 1 : 0;
assign detect_max[554][24] = (mid_1[4447:4440] > btm_2[4447:4440]) ? 1 : 0;
assign detect_max[554][25] = (mid_1[4447:4440] > btm_2[4455:4448]) ? 1 : 0;

assign detect_max[555][0] = (mid_1[4455:4448] > top_0[4447:4440]) ? 1 : 0;
assign detect_max[555][1] = (mid_1[4455:4448] > top_0[4455:4448]) ? 1 : 0;
assign detect_max[555][2] = (mid_1[4455:4448] > top_0[4463:4456]) ? 1 : 0;
assign detect_max[555][3] = (mid_1[4455:4448] > top_1[4447:4440]) ? 1 : 0;
assign detect_max[555][4] = (mid_1[4455:4448] > top_1[4455:4448]) ? 1 : 0;
assign detect_max[555][5] = (mid_1[4455:4448] > top_1[4463:4456]) ? 1 : 0;
assign detect_max[555][6] = (mid_1[4455:4448] > top_2[4447:4440]) ? 1 : 0;
assign detect_max[555][7] = (mid_1[4455:4448] > top_2[4455:4448]) ? 1 : 0;
assign detect_max[555][8] = (mid_1[4455:4448] > top_2[4463:4456]) ? 1 : 0;
assign detect_max[555][9] = (mid_1[4455:4448] > mid_0[4447:4440]) ? 1 : 0;
assign detect_max[555][10] = (mid_1[4455:4448] > mid_0[4455:4448]) ? 1 : 0;
assign detect_max[555][11] = (mid_1[4455:4448] > mid_0[4463:4456]) ? 1 : 0;
assign detect_max[555][12] = (mid_1[4455:4448] > mid_1[4447:4440]) ? 1 : 0;
assign detect_max[555][13] = (mid_1[4455:4448] > mid_1[4463:4456]) ? 1 : 0;
assign detect_max[555][14] = (mid_1[4455:4448] > mid_2[4447:4440]) ? 1 : 0;
assign detect_max[555][15] = (mid_1[4455:4448] > mid_2[4455:4448]) ? 1 : 0;
assign detect_max[555][16] = (mid_1[4455:4448] > mid_2[4463:4456]) ? 1 : 0;
assign detect_max[555][17] = (mid_1[4455:4448] > btm_0[4447:4440]) ? 1 : 0;
assign detect_max[555][18] = (mid_1[4455:4448] > btm_0[4455:4448]) ? 1 : 0;
assign detect_max[555][19] = (mid_1[4455:4448] > btm_0[4463:4456]) ? 1 : 0;
assign detect_max[555][20] = (mid_1[4455:4448] > btm_1[4447:4440]) ? 1 : 0;
assign detect_max[555][21] = (mid_1[4455:4448] > btm_1[4455:4448]) ? 1 : 0;
assign detect_max[555][22] = (mid_1[4455:4448] > btm_1[4463:4456]) ? 1 : 0;
assign detect_max[555][23] = (mid_1[4455:4448] > btm_2[4447:4440]) ? 1 : 0;
assign detect_max[555][24] = (mid_1[4455:4448] > btm_2[4455:4448]) ? 1 : 0;
assign detect_max[555][25] = (mid_1[4455:4448] > btm_2[4463:4456]) ? 1 : 0;

assign detect_max[556][0] = (mid_1[4463:4456] > top_0[4455:4448]) ? 1 : 0;
assign detect_max[556][1] = (mid_1[4463:4456] > top_0[4463:4456]) ? 1 : 0;
assign detect_max[556][2] = (mid_1[4463:4456] > top_0[4471:4464]) ? 1 : 0;
assign detect_max[556][3] = (mid_1[4463:4456] > top_1[4455:4448]) ? 1 : 0;
assign detect_max[556][4] = (mid_1[4463:4456] > top_1[4463:4456]) ? 1 : 0;
assign detect_max[556][5] = (mid_1[4463:4456] > top_1[4471:4464]) ? 1 : 0;
assign detect_max[556][6] = (mid_1[4463:4456] > top_2[4455:4448]) ? 1 : 0;
assign detect_max[556][7] = (mid_1[4463:4456] > top_2[4463:4456]) ? 1 : 0;
assign detect_max[556][8] = (mid_1[4463:4456] > top_2[4471:4464]) ? 1 : 0;
assign detect_max[556][9] = (mid_1[4463:4456] > mid_0[4455:4448]) ? 1 : 0;
assign detect_max[556][10] = (mid_1[4463:4456] > mid_0[4463:4456]) ? 1 : 0;
assign detect_max[556][11] = (mid_1[4463:4456] > mid_0[4471:4464]) ? 1 : 0;
assign detect_max[556][12] = (mid_1[4463:4456] > mid_1[4455:4448]) ? 1 : 0;
assign detect_max[556][13] = (mid_1[4463:4456] > mid_1[4471:4464]) ? 1 : 0;
assign detect_max[556][14] = (mid_1[4463:4456] > mid_2[4455:4448]) ? 1 : 0;
assign detect_max[556][15] = (mid_1[4463:4456] > mid_2[4463:4456]) ? 1 : 0;
assign detect_max[556][16] = (mid_1[4463:4456] > mid_2[4471:4464]) ? 1 : 0;
assign detect_max[556][17] = (mid_1[4463:4456] > btm_0[4455:4448]) ? 1 : 0;
assign detect_max[556][18] = (mid_1[4463:4456] > btm_0[4463:4456]) ? 1 : 0;
assign detect_max[556][19] = (mid_1[4463:4456] > btm_0[4471:4464]) ? 1 : 0;
assign detect_max[556][20] = (mid_1[4463:4456] > btm_1[4455:4448]) ? 1 : 0;
assign detect_max[556][21] = (mid_1[4463:4456] > btm_1[4463:4456]) ? 1 : 0;
assign detect_max[556][22] = (mid_1[4463:4456] > btm_1[4471:4464]) ? 1 : 0;
assign detect_max[556][23] = (mid_1[4463:4456] > btm_2[4455:4448]) ? 1 : 0;
assign detect_max[556][24] = (mid_1[4463:4456] > btm_2[4463:4456]) ? 1 : 0;
assign detect_max[556][25] = (mid_1[4463:4456] > btm_2[4471:4464]) ? 1 : 0;

assign detect_max[557][0] = (mid_1[4471:4464] > top_0[4463:4456]) ? 1 : 0;
assign detect_max[557][1] = (mid_1[4471:4464] > top_0[4471:4464]) ? 1 : 0;
assign detect_max[557][2] = (mid_1[4471:4464] > top_0[4479:4472]) ? 1 : 0;
assign detect_max[557][3] = (mid_1[4471:4464] > top_1[4463:4456]) ? 1 : 0;
assign detect_max[557][4] = (mid_1[4471:4464] > top_1[4471:4464]) ? 1 : 0;
assign detect_max[557][5] = (mid_1[4471:4464] > top_1[4479:4472]) ? 1 : 0;
assign detect_max[557][6] = (mid_1[4471:4464] > top_2[4463:4456]) ? 1 : 0;
assign detect_max[557][7] = (mid_1[4471:4464] > top_2[4471:4464]) ? 1 : 0;
assign detect_max[557][8] = (mid_1[4471:4464] > top_2[4479:4472]) ? 1 : 0;
assign detect_max[557][9] = (mid_1[4471:4464] > mid_0[4463:4456]) ? 1 : 0;
assign detect_max[557][10] = (mid_1[4471:4464] > mid_0[4471:4464]) ? 1 : 0;
assign detect_max[557][11] = (mid_1[4471:4464] > mid_0[4479:4472]) ? 1 : 0;
assign detect_max[557][12] = (mid_1[4471:4464] > mid_1[4463:4456]) ? 1 : 0;
assign detect_max[557][13] = (mid_1[4471:4464] > mid_1[4479:4472]) ? 1 : 0;
assign detect_max[557][14] = (mid_1[4471:4464] > mid_2[4463:4456]) ? 1 : 0;
assign detect_max[557][15] = (mid_1[4471:4464] > mid_2[4471:4464]) ? 1 : 0;
assign detect_max[557][16] = (mid_1[4471:4464] > mid_2[4479:4472]) ? 1 : 0;
assign detect_max[557][17] = (mid_1[4471:4464] > btm_0[4463:4456]) ? 1 : 0;
assign detect_max[557][18] = (mid_1[4471:4464] > btm_0[4471:4464]) ? 1 : 0;
assign detect_max[557][19] = (mid_1[4471:4464] > btm_0[4479:4472]) ? 1 : 0;
assign detect_max[557][20] = (mid_1[4471:4464] > btm_1[4463:4456]) ? 1 : 0;
assign detect_max[557][21] = (mid_1[4471:4464] > btm_1[4471:4464]) ? 1 : 0;
assign detect_max[557][22] = (mid_1[4471:4464] > btm_1[4479:4472]) ? 1 : 0;
assign detect_max[557][23] = (mid_1[4471:4464] > btm_2[4463:4456]) ? 1 : 0;
assign detect_max[557][24] = (mid_1[4471:4464] > btm_2[4471:4464]) ? 1 : 0;
assign detect_max[557][25] = (mid_1[4471:4464] > btm_2[4479:4472]) ? 1 : 0;

assign detect_max[558][0] = (mid_1[4479:4472] > top_0[4471:4464]) ? 1 : 0;
assign detect_max[558][1] = (mid_1[4479:4472] > top_0[4479:4472]) ? 1 : 0;
assign detect_max[558][2] = (mid_1[4479:4472] > top_0[4487:4480]) ? 1 : 0;
assign detect_max[558][3] = (mid_1[4479:4472] > top_1[4471:4464]) ? 1 : 0;
assign detect_max[558][4] = (mid_1[4479:4472] > top_1[4479:4472]) ? 1 : 0;
assign detect_max[558][5] = (mid_1[4479:4472] > top_1[4487:4480]) ? 1 : 0;
assign detect_max[558][6] = (mid_1[4479:4472] > top_2[4471:4464]) ? 1 : 0;
assign detect_max[558][7] = (mid_1[4479:4472] > top_2[4479:4472]) ? 1 : 0;
assign detect_max[558][8] = (mid_1[4479:4472] > top_2[4487:4480]) ? 1 : 0;
assign detect_max[558][9] = (mid_1[4479:4472] > mid_0[4471:4464]) ? 1 : 0;
assign detect_max[558][10] = (mid_1[4479:4472] > mid_0[4479:4472]) ? 1 : 0;
assign detect_max[558][11] = (mid_1[4479:4472] > mid_0[4487:4480]) ? 1 : 0;
assign detect_max[558][12] = (mid_1[4479:4472] > mid_1[4471:4464]) ? 1 : 0;
assign detect_max[558][13] = (mid_1[4479:4472] > mid_1[4487:4480]) ? 1 : 0;
assign detect_max[558][14] = (mid_1[4479:4472] > mid_2[4471:4464]) ? 1 : 0;
assign detect_max[558][15] = (mid_1[4479:4472] > mid_2[4479:4472]) ? 1 : 0;
assign detect_max[558][16] = (mid_1[4479:4472] > mid_2[4487:4480]) ? 1 : 0;
assign detect_max[558][17] = (mid_1[4479:4472] > btm_0[4471:4464]) ? 1 : 0;
assign detect_max[558][18] = (mid_1[4479:4472] > btm_0[4479:4472]) ? 1 : 0;
assign detect_max[558][19] = (mid_1[4479:4472] > btm_0[4487:4480]) ? 1 : 0;
assign detect_max[558][20] = (mid_1[4479:4472] > btm_1[4471:4464]) ? 1 : 0;
assign detect_max[558][21] = (mid_1[4479:4472] > btm_1[4479:4472]) ? 1 : 0;
assign detect_max[558][22] = (mid_1[4479:4472] > btm_1[4487:4480]) ? 1 : 0;
assign detect_max[558][23] = (mid_1[4479:4472] > btm_2[4471:4464]) ? 1 : 0;
assign detect_max[558][24] = (mid_1[4479:4472] > btm_2[4479:4472]) ? 1 : 0;
assign detect_max[558][25] = (mid_1[4479:4472] > btm_2[4487:4480]) ? 1 : 0;

assign detect_max[559][0] = (mid_1[4487:4480] > top_0[4479:4472]) ? 1 : 0;
assign detect_max[559][1] = (mid_1[4487:4480] > top_0[4487:4480]) ? 1 : 0;
assign detect_max[559][2] = (mid_1[4487:4480] > top_0[4495:4488]) ? 1 : 0;
assign detect_max[559][3] = (mid_1[4487:4480] > top_1[4479:4472]) ? 1 : 0;
assign detect_max[559][4] = (mid_1[4487:4480] > top_1[4487:4480]) ? 1 : 0;
assign detect_max[559][5] = (mid_1[4487:4480] > top_1[4495:4488]) ? 1 : 0;
assign detect_max[559][6] = (mid_1[4487:4480] > top_2[4479:4472]) ? 1 : 0;
assign detect_max[559][7] = (mid_1[4487:4480] > top_2[4487:4480]) ? 1 : 0;
assign detect_max[559][8] = (mid_1[4487:4480] > top_2[4495:4488]) ? 1 : 0;
assign detect_max[559][9] = (mid_1[4487:4480] > mid_0[4479:4472]) ? 1 : 0;
assign detect_max[559][10] = (mid_1[4487:4480] > mid_0[4487:4480]) ? 1 : 0;
assign detect_max[559][11] = (mid_1[4487:4480] > mid_0[4495:4488]) ? 1 : 0;
assign detect_max[559][12] = (mid_1[4487:4480] > mid_1[4479:4472]) ? 1 : 0;
assign detect_max[559][13] = (mid_1[4487:4480] > mid_1[4495:4488]) ? 1 : 0;
assign detect_max[559][14] = (mid_1[4487:4480] > mid_2[4479:4472]) ? 1 : 0;
assign detect_max[559][15] = (mid_1[4487:4480] > mid_2[4487:4480]) ? 1 : 0;
assign detect_max[559][16] = (mid_1[4487:4480] > mid_2[4495:4488]) ? 1 : 0;
assign detect_max[559][17] = (mid_1[4487:4480] > btm_0[4479:4472]) ? 1 : 0;
assign detect_max[559][18] = (mid_1[4487:4480] > btm_0[4487:4480]) ? 1 : 0;
assign detect_max[559][19] = (mid_1[4487:4480] > btm_0[4495:4488]) ? 1 : 0;
assign detect_max[559][20] = (mid_1[4487:4480] > btm_1[4479:4472]) ? 1 : 0;
assign detect_max[559][21] = (mid_1[4487:4480] > btm_1[4487:4480]) ? 1 : 0;
assign detect_max[559][22] = (mid_1[4487:4480] > btm_1[4495:4488]) ? 1 : 0;
assign detect_max[559][23] = (mid_1[4487:4480] > btm_2[4479:4472]) ? 1 : 0;
assign detect_max[559][24] = (mid_1[4487:4480] > btm_2[4487:4480]) ? 1 : 0;
assign detect_max[559][25] = (mid_1[4487:4480] > btm_2[4495:4488]) ? 1 : 0;

assign detect_max[560][0] = (mid_1[4495:4488] > top_0[4487:4480]) ? 1 : 0;
assign detect_max[560][1] = (mid_1[4495:4488] > top_0[4495:4488]) ? 1 : 0;
assign detect_max[560][2] = (mid_1[4495:4488] > top_0[4503:4496]) ? 1 : 0;
assign detect_max[560][3] = (mid_1[4495:4488] > top_1[4487:4480]) ? 1 : 0;
assign detect_max[560][4] = (mid_1[4495:4488] > top_1[4495:4488]) ? 1 : 0;
assign detect_max[560][5] = (mid_1[4495:4488] > top_1[4503:4496]) ? 1 : 0;
assign detect_max[560][6] = (mid_1[4495:4488] > top_2[4487:4480]) ? 1 : 0;
assign detect_max[560][7] = (mid_1[4495:4488] > top_2[4495:4488]) ? 1 : 0;
assign detect_max[560][8] = (mid_1[4495:4488] > top_2[4503:4496]) ? 1 : 0;
assign detect_max[560][9] = (mid_1[4495:4488] > mid_0[4487:4480]) ? 1 : 0;
assign detect_max[560][10] = (mid_1[4495:4488] > mid_0[4495:4488]) ? 1 : 0;
assign detect_max[560][11] = (mid_1[4495:4488] > mid_0[4503:4496]) ? 1 : 0;
assign detect_max[560][12] = (mid_1[4495:4488] > mid_1[4487:4480]) ? 1 : 0;
assign detect_max[560][13] = (mid_1[4495:4488] > mid_1[4503:4496]) ? 1 : 0;
assign detect_max[560][14] = (mid_1[4495:4488] > mid_2[4487:4480]) ? 1 : 0;
assign detect_max[560][15] = (mid_1[4495:4488] > mid_2[4495:4488]) ? 1 : 0;
assign detect_max[560][16] = (mid_1[4495:4488] > mid_2[4503:4496]) ? 1 : 0;
assign detect_max[560][17] = (mid_1[4495:4488] > btm_0[4487:4480]) ? 1 : 0;
assign detect_max[560][18] = (mid_1[4495:4488] > btm_0[4495:4488]) ? 1 : 0;
assign detect_max[560][19] = (mid_1[4495:4488] > btm_0[4503:4496]) ? 1 : 0;
assign detect_max[560][20] = (mid_1[4495:4488] > btm_1[4487:4480]) ? 1 : 0;
assign detect_max[560][21] = (mid_1[4495:4488] > btm_1[4495:4488]) ? 1 : 0;
assign detect_max[560][22] = (mid_1[4495:4488] > btm_1[4503:4496]) ? 1 : 0;
assign detect_max[560][23] = (mid_1[4495:4488] > btm_2[4487:4480]) ? 1 : 0;
assign detect_max[560][24] = (mid_1[4495:4488] > btm_2[4495:4488]) ? 1 : 0;
assign detect_max[560][25] = (mid_1[4495:4488] > btm_2[4503:4496]) ? 1 : 0;

assign detect_max[561][0] = (mid_1[4503:4496] > top_0[4495:4488]) ? 1 : 0;
assign detect_max[561][1] = (mid_1[4503:4496] > top_0[4503:4496]) ? 1 : 0;
assign detect_max[561][2] = (mid_1[4503:4496] > top_0[4511:4504]) ? 1 : 0;
assign detect_max[561][3] = (mid_1[4503:4496] > top_1[4495:4488]) ? 1 : 0;
assign detect_max[561][4] = (mid_1[4503:4496] > top_1[4503:4496]) ? 1 : 0;
assign detect_max[561][5] = (mid_1[4503:4496] > top_1[4511:4504]) ? 1 : 0;
assign detect_max[561][6] = (mid_1[4503:4496] > top_2[4495:4488]) ? 1 : 0;
assign detect_max[561][7] = (mid_1[4503:4496] > top_2[4503:4496]) ? 1 : 0;
assign detect_max[561][8] = (mid_1[4503:4496] > top_2[4511:4504]) ? 1 : 0;
assign detect_max[561][9] = (mid_1[4503:4496] > mid_0[4495:4488]) ? 1 : 0;
assign detect_max[561][10] = (mid_1[4503:4496] > mid_0[4503:4496]) ? 1 : 0;
assign detect_max[561][11] = (mid_1[4503:4496] > mid_0[4511:4504]) ? 1 : 0;
assign detect_max[561][12] = (mid_1[4503:4496] > mid_1[4495:4488]) ? 1 : 0;
assign detect_max[561][13] = (mid_1[4503:4496] > mid_1[4511:4504]) ? 1 : 0;
assign detect_max[561][14] = (mid_1[4503:4496] > mid_2[4495:4488]) ? 1 : 0;
assign detect_max[561][15] = (mid_1[4503:4496] > mid_2[4503:4496]) ? 1 : 0;
assign detect_max[561][16] = (mid_1[4503:4496] > mid_2[4511:4504]) ? 1 : 0;
assign detect_max[561][17] = (mid_1[4503:4496] > btm_0[4495:4488]) ? 1 : 0;
assign detect_max[561][18] = (mid_1[4503:4496] > btm_0[4503:4496]) ? 1 : 0;
assign detect_max[561][19] = (mid_1[4503:4496] > btm_0[4511:4504]) ? 1 : 0;
assign detect_max[561][20] = (mid_1[4503:4496] > btm_1[4495:4488]) ? 1 : 0;
assign detect_max[561][21] = (mid_1[4503:4496] > btm_1[4503:4496]) ? 1 : 0;
assign detect_max[561][22] = (mid_1[4503:4496] > btm_1[4511:4504]) ? 1 : 0;
assign detect_max[561][23] = (mid_1[4503:4496] > btm_2[4495:4488]) ? 1 : 0;
assign detect_max[561][24] = (mid_1[4503:4496] > btm_2[4503:4496]) ? 1 : 0;
assign detect_max[561][25] = (mid_1[4503:4496] > btm_2[4511:4504]) ? 1 : 0;

assign detect_max[562][0] = (mid_1[4511:4504] > top_0[4503:4496]) ? 1 : 0;
assign detect_max[562][1] = (mid_1[4511:4504] > top_0[4511:4504]) ? 1 : 0;
assign detect_max[562][2] = (mid_1[4511:4504] > top_0[4519:4512]) ? 1 : 0;
assign detect_max[562][3] = (mid_1[4511:4504] > top_1[4503:4496]) ? 1 : 0;
assign detect_max[562][4] = (mid_1[4511:4504] > top_1[4511:4504]) ? 1 : 0;
assign detect_max[562][5] = (mid_1[4511:4504] > top_1[4519:4512]) ? 1 : 0;
assign detect_max[562][6] = (mid_1[4511:4504] > top_2[4503:4496]) ? 1 : 0;
assign detect_max[562][7] = (mid_1[4511:4504] > top_2[4511:4504]) ? 1 : 0;
assign detect_max[562][8] = (mid_1[4511:4504] > top_2[4519:4512]) ? 1 : 0;
assign detect_max[562][9] = (mid_1[4511:4504] > mid_0[4503:4496]) ? 1 : 0;
assign detect_max[562][10] = (mid_1[4511:4504] > mid_0[4511:4504]) ? 1 : 0;
assign detect_max[562][11] = (mid_1[4511:4504] > mid_0[4519:4512]) ? 1 : 0;
assign detect_max[562][12] = (mid_1[4511:4504] > mid_1[4503:4496]) ? 1 : 0;
assign detect_max[562][13] = (mid_1[4511:4504] > mid_1[4519:4512]) ? 1 : 0;
assign detect_max[562][14] = (mid_1[4511:4504] > mid_2[4503:4496]) ? 1 : 0;
assign detect_max[562][15] = (mid_1[4511:4504] > mid_2[4511:4504]) ? 1 : 0;
assign detect_max[562][16] = (mid_1[4511:4504] > mid_2[4519:4512]) ? 1 : 0;
assign detect_max[562][17] = (mid_1[4511:4504] > btm_0[4503:4496]) ? 1 : 0;
assign detect_max[562][18] = (mid_1[4511:4504] > btm_0[4511:4504]) ? 1 : 0;
assign detect_max[562][19] = (mid_1[4511:4504] > btm_0[4519:4512]) ? 1 : 0;
assign detect_max[562][20] = (mid_1[4511:4504] > btm_1[4503:4496]) ? 1 : 0;
assign detect_max[562][21] = (mid_1[4511:4504] > btm_1[4511:4504]) ? 1 : 0;
assign detect_max[562][22] = (mid_1[4511:4504] > btm_1[4519:4512]) ? 1 : 0;
assign detect_max[562][23] = (mid_1[4511:4504] > btm_2[4503:4496]) ? 1 : 0;
assign detect_max[562][24] = (mid_1[4511:4504] > btm_2[4511:4504]) ? 1 : 0;
assign detect_max[562][25] = (mid_1[4511:4504] > btm_2[4519:4512]) ? 1 : 0;

assign detect_max[563][0] = (mid_1[4519:4512] > top_0[4511:4504]) ? 1 : 0;
assign detect_max[563][1] = (mid_1[4519:4512] > top_0[4519:4512]) ? 1 : 0;
assign detect_max[563][2] = (mid_1[4519:4512] > top_0[4527:4520]) ? 1 : 0;
assign detect_max[563][3] = (mid_1[4519:4512] > top_1[4511:4504]) ? 1 : 0;
assign detect_max[563][4] = (mid_1[4519:4512] > top_1[4519:4512]) ? 1 : 0;
assign detect_max[563][5] = (mid_1[4519:4512] > top_1[4527:4520]) ? 1 : 0;
assign detect_max[563][6] = (mid_1[4519:4512] > top_2[4511:4504]) ? 1 : 0;
assign detect_max[563][7] = (mid_1[4519:4512] > top_2[4519:4512]) ? 1 : 0;
assign detect_max[563][8] = (mid_1[4519:4512] > top_2[4527:4520]) ? 1 : 0;
assign detect_max[563][9] = (mid_1[4519:4512] > mid_0[4511:4504]) ? 1 : 0;
assign detect_max[563][10] = (mid_1[4519:4512] > mid_0[4519:4512]) ? 1 : 0;
assign detect_max[563][11] = (mid_1[4519:4512] > mid_0[4527:4520]) ? 1 : 0;
assign detect_max[563][12] = (mid_1[4519:4512] > mid_1[4511:4504]) ? 1 : 0;
assign detect_max[563][13] = (mid_1[4519:4512] > mid_1[4527:4520]) ? 1 : 0;
assign detect_max[563][14] = (mid_1[4519:4512] > mid_2[4511:4504]) ? 1 : 0;
assign detect_max[563][15] = (mid_1[4519:4512] > mid_2[4519:4512]) ? 1 : 0;
assign detect_max[563][16] = (mid_1[4519:4512] > mid_2[4527:4520]) ? 1 : 0;
assign detect_max[563][17] = (mid_1[4519:4512] > btm_0[4511:4504]) ? 1 : 0;
assign detect_max[563][18] = (mid_1[4519:4512] > btm_0[4519:4512]) ? 1 : 0;
assign detect_max[563][19] = (mid_1[4519:4512] > btm_0[4527:4520]) ? 1 : 0;
assign detect_max[563][20] = (mid_1[4519:4512] > btm_1[4511:4504]) ? 1 : 0;
assign detect_max[563][21] = (mid_1[4519:4512] > btm_1[4519:4512]) ? 1 : 0;
assign detect_max[563][22] = (mid_1[4519:4512] > btm_1[4527:4520]) ? 1 : 0;
assign detect_max[563][23] = (mid_1[4519:4512] > btm_2[4511:4504]) ? 1 : 0;
assign detect_max[563][24] = (mid_1[4519:4512] > btm_2[4519:4512]) ? 1 : 0;
assign detect_max[563][25] = (mid_1[4519:4512] > btm_2[4527:4520]) ? 1 : 0;

assign detect_max[564][0] = (mid_1[4527:4520] > top_0[4519:4512]) ? 1 : 0;
assign detect_max[564][1] = (mid_1[4527:4520] > top_0[4527:4520]) ? 1 : 0;
assign detect_max[564][2] = (mid_1[4527:4520] > top_0[4535:4528]) ? 1 : 0;
assign detect_max[564][3] = (mid_1[4527:4520] > top_1[4519:4512]) ? 1 : 0;
assign detect_max[564][4] = (mid_1[4527:4520] > top_1[4527:4520]) ? 1 : 0;
assign detect_max[564][5] = (mid_1[4527:4520] > top_1[4535:4528]) ? 1 : 0;
assign detect_max[564][6] = (mid_1[4527:4520] > top_2[4519:4512]) ? 1 : 0;
assign detect_max[564][7] = (mid_1[4527:4520] > top_2[4527:4520]) ? 1 : 0;
assign detect_max[564][8] = (mid_1[4527:4520] > top_2[4535:4528]) ? 1 : 0;
assign detect_max[564][9] = (mid_1[4527:4520] > mid_0[4519:4512]) ? 1 : 0;
assign detect_max[564][10] = (mid_1[4527:4520] > mid_0[4527:4520]) ? 1 : 0;
assign detect_max[564][11] = (mid_1[4527:4520] > mid_0[4535:4528]) ? 1 : 0;
assign detect_max[564][12] = (mid_1[4527:4520] > mid_1[4519:4512]) ? 1 : 0;
assign detect_max[564][13] = (mid_1[4527:4520] > mid_1[4535:4528]) ? 1 : 0;
assign detect_max[564][14] = (mid_1[4527:4520] > mid_2[4519:4512]) ? 1 : 0;
assign detect_max[564][15] = (mid_1[4527:4520] > mid_2[4527:4520]) ? 1 : 0;
assign detect_max[564][16] = (mid_1[4527:4520] > mid_2[4535:4528]) ? 1 : 0;
assign detect_max[564][17] = (mid_1[4527:4520] > btm_0[4519:4512]) ? 1 : 0;
assign detect_max[564][18] = (mid_1[4527:4520] > btm_0[4527:4520]) ? 1 : 0;
assign detect_max[564][19] = (mid_1[4527:4520] > btm_0[4535:4528]) ? 1 : 0;
assign detect_max[564][20] = (mid_1[4527:4520] > btm_1[4519:4512]) ? 1 : 0;
assign detect_max[564][21] = (mid_1[4527:4520] > btm_1[4527:4520]) ? 1 : 0;
assign detect_max[564][22] = (mid_1[4527:4520] > btm_1[4535:4528]) ? 1 : 0;
assign detect_max[564][23] = (mid_1[4527:4520] > btm_2[4519:4512]) ? 1 : 0;
assign detect_max[564][24] = (mid_1[4527:4520] > btm_2[4527:4520]) ? 1 : 0;
assign detect_max[564][25] = (mid_1[4527:4520] > btm_2[4535:4528]) ? 1 : 0;

assign detect_max[565][0] = (mid_1[4535:4528] > top_0[4527:4520]) ? 1 : 0;
assign detect_max[565][1] = (mid_1[4535:4528] > top_0[4535:4528]) ? 1 : 0;
assign detect_max[565][2] = (mid_1[4535:4528] > top_0[4543:4536]) ? 1 : 0;
assign detect_max[565][3] = (mid_1[4535:4528] > top_1[4527:4520]) ? 1 : 0;
assign detect_max[565][4] = (mid_1[4535:4528] > top_1[4535:4528]) ? 1 : 0;
assign detect_max[565][5] = (mid_1[4535:4528] > top_1[4543:4536]) ? 1 : 0;
assign detect_max[565][6] = (mid_1[4535:4528] > top_2[4527:4520]) ? 1 : 0;
assign detect_max[565][7] = (mid_1[4535:4528] > top_2[4535:4528]) ? 1 : 0;
assign detect_max[565][8] = (mid_1[4535:4528] > top_2[4543:4536]) ? 1 : 0;
assign detect_max[565][9] = (mid_1[4535:4528] > mid_0[4527:4520]) ? 1 : 0;
assign detect_max[565][10] = (mid_1[4535:4528] > mid_0[4535:4528]) ? 1 : 0;
assign detect_max[565][11] = (mid_1[4535:4528] > mid_0[4543:4536]) ? 1 : 0;
assign detect_max[565][12] = (mid_1[4535:4528] > mid_1[4527:4520]) ? 1 : 0;
assign detect_max[565][13] = (mid_1[4535:4528] > mid_1[4543:4536]) ? 1 : 0;
assign detect_max[565][14] = (mid_1[4535:4528] > mid_2[4527:4520]) ? 1 : 0;
assign detect_max[565][15] = (mid_1[4535:4528] > mid_2[4535:4528]) ? 1 : 0;
assign detect_max[565][16] = (mid_1[4535:4528] > mid_2[4543:4536]) ? 1 : 0;
assign detect_max[565][17] = (mid_1[4535:4528] > btm_0[4527:4520]) ? 1 : 0;
assign detect_max[565][18] = (mid_1[4535:4528] > btm_0[4535:4528]) ? 1 : 0;
assign detect_max[565][19] = (mid_1[4535:4528] > btm_0[4543:4536]) ? 1 : 0;
assign detect_max[565][20] = (mid_1[4535:4528] > btm_1[4527:4520]) ? 1 : 0;
assign detect_max[565][21] = (mid_1[4535:4528] > btm_1[4535:4528]) ? 1 : 0;
assign detect_max[565][22] = (mid_1[4535:4528] > btm_1[4543:4536]) ? 1 : 0;
assign detect_max[565][23] = (mid_1[4535:4528] > btm_2[4527:4520]) ? 1 : 0;
assign detect_max[565][24] = (mid_1[4535:4528] > btm_2[4535:4528]) ? 1 : 0;
assign detect_max[565][25] = (mid_1[4535:4528] > btm_2[4543:4536]) ? 1 : 0;

assign detect_max[566][0] = (mid_1[4543:4536] > top_0[4535:4528]) ? 1 : 0;
assign detect_max[566][1] = (mid_1[4543:4536] > top_0[4543:4536]) ? 1 : 0;
assign detect_max[566][2] = (mid_1[4543:4536] > top_0[4551:4544]) ? 1 : 0;
assign detect_max[566][3] = (mid_1[4543:4536] > top_1[4535:4528]) ? 1 : 0;
assign detect_max[566][4] = (mid_1[4543:4536] > top_1[4543:4536]) ? 1 : 0;
assign detect_max[566][5] = (mid_1[4543:4536] > top_1[4551:4544]) ? 1 : 0;
assign detect_max[566][6] = (mid_1[4543:4536] > top_2[4535:4528]) ? 1 : 0;
assign detect_max[566][7] = (mid_1[4543:4536] > top_2[4543:4536]) ? 1 : 0;
assign detect_max[566][8] = (mid_1[4543:4536] > top_2[4551:4544]) ? 1 : 0;
assign detect_max[566][9] = (mid_1[4543:4536] > mid_0[4535:4528]) ? 1 : 0;
assign detect_max[566][10] = (mid_1[4543:4536] > mid_0[4543:4536]) ? 1 : 0;
assign detect_max[566][11] = (mid_1[4543:4536] > mid_0[4551:4544]) ? 1 : 0;
assign detect_max[566][12] = (mid_1[4543:4536] > mid_1[4535:4528]) ? 1 : 0;
assign detect_max[566][13] = (mid_1[4543:4536] > mid_1[4551:4544]) ? 1 : 0;
assign detect_max[566][14] = (mid_1[4543:4536] > mid_2[4535:4528]) ? 1 : 0;
assign detect_max[566][15] = (mid_1[4543:4536] > mid_2[4543:4536]) ? 1 : 0;
assign detect_max[566][16] = (mid_1[4543:4536] > mid_2[4551:4544]) ? 1 : 0;
assign detect_max[566][17] = (mid_1[4543:4536] > btm_0[4535:4528]) ? 1 : 0;
assign detect_max[566][18] = (mid_1[4543:4536] > btm_0[4543:4536]) ? 1 : 0;
assign detect_max[566][19] = (mid_1[4543:4536] > btm_0[4551:4544]) ? 1 : 0;
assign detect_max[566][20] = (mid_1[4543:4536] > btm_1[4535:4528]) ? 1 : 0;
assign detect_max[566][21] = (mid_1[4543:4536] > btm_1[4543:4536]) ? 1 : 0;
assign detect_max[566][22] = (mid_1[4543:4536] > btm_1[4551:4544]) ? 1 : 0;
assign detect_max[566][23] = (mid_1[4543:4536] > btm_2[4535:4528]) ? 1 : 0;
assign detect_max[566][24] = (mid_1[4543:4536] > btm_2[4543:4536]) ? 1 : 0;
assign detect_max[566][25] = (mid_1[4543:4536] > btm_2[4551:4544]) ? 1 : 0;

assign detect_max[567][0] = (mid_1[4551:4544] > top_0[4543:4536]) ? 1 : 0;
assign detect_max[567][1] = (mid_1[4551:4544] > top_0[4551:4544]) ? 1 : 0;
assign detect_max[567][2] = (mid_1[4551:4544] > top_0[4559:4552]) ? 1 : 0;
assign detect_max[567][3] = (mid_1[4551:4544] > top_1[4543:4536]) ? 1 : 0;
assign detect_max[567][4] = (mid_1[4551:4544] > top_1[4551:4544]) ? 1 : 0;
assign detect_max[567][5] = (mid_1[4551:4544] > top_1[4559:4552]) ? 1 : 0;
assign detect_max[567][6] = (mid_1[4551:4544] > top_2[4543:4536]) ? 1 : 0;
assign detect_max[567][7] = (mid_1[4551:4544] > top_2[4551:4544]) ? 1 : 0;
assign detect_max[567][8] = (mid_1[4551:4544] > top_2[4559:4552]) ? 1 : 0;
assign detect_max[567][9] = (mid_1[4551:4544] > mid_0[4543:4536]) ? 1 : 0;
assign detect_max[567][10] = (mid_1[4551:4544] > mid_0[4551:4544]) ? 1 : 0;
assign detect_max[567][11] = (mid_1[4551:4544] > mid_0[4559:4552]) ? 1 : 0;
assign detect_max[567][12] = (mid_1[4551:4544] > mid_1[4543:4536]) ? 1 : 0;
assign detect_max[567][13] = (mid_1[4551:4544] > mid_1[4559:4552]) ? 1 : 0;
assign detect_max[567][14] = (mid_1[4551:4544] > mid_2[4543:4536]) ? 1 : 0;
assign detect_max[567][15] = (mid_1[4551:4544] > mid_2[4551:4544]) ? 1 : 0;
assign detect_max[567][16] = (mid_1[4551:4544] > mid_2[4559:4552]) ? 1 : 0;
assign detect_max[567][17] = (mid_1[4551:4544] > btm_0[4543:4536]) ? 1 : 0;
assign detect_max[567][18] = (mid_1[4551:4544] > btm_0[4551:4544]) ? 1 : 0;
assign detect_max[567][19] = (mid_1[4551:4544] > btm_0[4559:4552]) ? 1 : 0;
assign detect_max[567][20] = (mid_1[4551:4544] > btm_1[4543:4536]) ? 1 : 0;
assign detect_max[567][21] = (mid_1[4551:4544] > btm_1[4551:4544]) ? 1 : 0;
assign detect_max[567][22] = (mid_1[4551:4544] > btm_1[4559:4552]) ? 1 : 0;
assign detect_max[567][23] = (mid_1[4551:4544] > btm_2[4543:4536]) ? 1 : 0;
assign detect_max[567][24] = (mid_1[4551:4544] > btm_2[4551:4544]) ? 1 : 0;
assign detect_max[567][25] = (mid_1[4551:4544] > btm_2[4559:4552]) ? 1 : 0;

assign detect_max[568][0] = (mid_1[4559:4552] > top_0[4551:4544]) ? 1 : 0;
assign detect_max[568][1] = (mid_1[4559:4552] > top_0[4559:4552]) ? 1 : 0;
assign detect_max[568][2] = (mid_1[4559:4552] > top_0[4567:4560]) ? 1 : 0;
assign detect_max[568][3] = (mid_1[4559:4552] > top_1[4551:4544]) ? 1 : 0;
assign detect_max[568][4] = (mid_1[4559:4552] > top_1[4559:4552]) ? 1 : 0;
assign detect_max[568][5] = (mid_1[4559:4552] > top_1[4567:4560]) ? 1 : 0;
assign detect_max[568][6] = (mid_1[4559:4552] > top_2[4551:4544]) ? 1 : 0;
assign detect_max[568][7] = (mid_1[4559:4552] > top_2[4559:4552]) ? 1 : 0;
assign detect_max[568][8] = (mid_1[4559:4552] > top_2[4567:4560]) ? 1 : 0;
assign detect_max[568][9] = (mid_1[4559:4552] > mid_0[4551:4544]) ? 1 : 0;
assign detect_max[568][10] = (mid_1[4559:4552] > mid_0[4559:4552]) ? 1 : 0;
assign detect_max[568][11] = (mid_1[4559:4552] > mid_0[4567:4560]) ? 1 : 0;
assign detect_max[568][12] = (mid_1[4559:4552] > mid_1[4551:4544]) ? 1 : 0;
assign detect_max[568][13] = (mid_1[4559:4552] > mid_1[4567:4560]) ? 1 : 0;
assign detect_max[568][14] = (mid_1[4559:4552] > mid_2[4551:4544]) ? 1 : 0;
assign detect_max[568][15] = (mid_1[4559:4552] > mid_2[4559:4552]) ? 1 : 0;
assign detect_max[568][16] = (mid_1[4559:4552] > mid_2[4567:4560]) ? 1 : 0;
assign detect_max[568][17] = (mid_1[4559:4552] > btm_0[4551:4544]) ? 1 : 0;
assign detect_max[568][18] = (mid_1[4559:4552] > btm_0[4559:4552]) ? 1 : 0;
assign detect_max[568][19] = (mid_1[4559:4552] > btm_0[4567:4560]) ? 1 : 0;
assign detect_max[568][20] = (mid_1[4559:4552] > btm_1[4551:4544]) ? 1 : 0;
assign detect_max[568][21] = (mid_1[4559:4552] > btm_1[4559:4552]) ? 1 : 0;
assign detect_max[568][22] = (mid_1[4559:4552] > btm_1[4567:4560]) ? 1 : 0;
assign detect_max[568][23] = (mid_1[4559:4552] > btm_2[4551:4544]) ? 1 : 0;
assign detect_max[568][24] = (mid_1[4559:4552] > btm_2[4559:4552]) ? 1 : 0;
assign detect_max[568][25] = (mid_1[4559:4552] > btm_2[4567:4560]) ? 1 : 0;

assign detect_max[569][0] = (mid_1[4567:4560] > top_0[4559:4552]) ? 1 : 0;
assign detect_max[569][1] = (mid_1[4567:4560] > top_0[4567:4560]) ? 1 : 0;
assign detect_max[569][2] = (mid_1[4567:4560] > top_0[4575:4568]) ? 1 : 0;
assign detect_max[569][3] = (mid_1[4567:4560] > top_1[4559:4552]) ? 1 : 0;
assign detect_max[569][4] = (mid_1[4567:4560] > top_1[4567:4560]) ? 1 : 0;
assign detect_max[569][5] = (mid_1[4567:4560] > top_1[4575:4568]) ? 1 : 0;
assign detect_max[569][6] = (mid_1[4567:4560] > top_2[4559:4552]) ? 1 : 0;
assign detect_max[569][7] = (mid_1[4567:4560] > top_2[4567:4560]) ? 1 : 0;
assign detect_max[569][8] = (mid_1[4567:4560] > top_2[4575:4568]) ? 1 : 0;
assign detect_max[569][9] = (mid_1[4567:4560] > mid_0[4559:4552]) ? 1 : 0;
assign detect_max[569][10] = (mid_1[4567:4560] > mid_0[4567:4560]) ? 1 : 0;
assign detect_max[569][11] = (mid_1[4567:4560] > mid_0[4575:4568]) ? 1 : 0;
assign detect_max[569][12] = (mid_1[4567:4560] > mid_1[4559:4552]) ? 1 : 0;
assign detect_max[569][13] = (mid_1[4567:4560] > mid_1[4575:4568]) ? 1 : 0;
assign detect_max[569][14] = (mid_1[4567:4560] > mid_2[4559:4552]) ? 1 : 0;
assign detect_max[569][15] = (mid_1[4567:4560] > mid_2[4567:4560]) ? 1 : 0;
assign detect_max[569][16] = (mid_1[4567:4560] > mid_2[4575:4568]) ? 1 : 0;
assign detect_max[569][17] = (mid_1[4567:4560] > btm_0[4559:4552]) ? 1 : 0;
assign detect_max[569][18] = (mid_1[4567:4560] > btm_0[4567:4560]) ? 1 : 0;
assign detect_max[569][19] = (mid_1[4567:4560] > btm_0[4575:4568]) ? 1 : 0;
assign detect_max[569][20] = (mid_1[4567:4560] > btm_1[4559:4552]) ? 1 : 0;
assign detect_max[569][21] = (mid_1[4567:4560] > btm_1[4567:4560]) ? 1 : 0;
assign detect_max[569][22] = (mid_1[4567:4560] > btm_1[4575:4568]) ? 1 : 0;
assign detect_max[569][23] = (mid_1[4567:4560] > btm_2[4559:4552]) ? 1 : 0;
assign detect_max[569][24] = (mid_1[4567:4560] > btm_2[4567:4560]) ? 1 : 0;
assign detect_max[569][25] = (mid_1[4567:4560] > btm_2[4575:4568]) ? 1 : 0;

assign detect_max[570][0] = (mid_1[4575:4568] > top_0[4567:4560]) ? 1 : 0;
assign detect_max[570][1] = (mid_1[4575:4568] > top_0[4575:4568]) ? 1 : 0;
assign detect_max[570][2] = (mid_1[4575:4568] > top_0[4583:4576]) ? 1 : 0;
assign detect_max[570][3] = (mid_1[4575:4568] > top_1[4567:4560]) ? 1 : 0;
assign detect_max[570][4] = (mid_1[4575:4568] > top_1[4575:4568]) ? 1 : 0;
assign detect_max[570][5] = (mid_1[4575:4568] > top_1[4583:4576]) ? 1 : 0;
assign detect_max[570][6] = (mid_1[4575:4568] > top_2[4567:4560]) ? 1 : 0;
assign detect_max[570][7] = (mid_1[4575:4568] > top_2[4575:4568]) ? 1 : 0;
assign detect_max[570][8] = (mid_1[4575:4568] > top_2[4583:4576]) ? 1 : 0;
assign detect_max[570][9] = (mid_1[4575:4568] > mid_0[4567:4560]) ? 1 : 0;
assign detect_max[570][10] = (mid_1[4575:4568] > mid_0[4575:4568]) ? 1 : 0;
assign detect_max[570][11] = (mid_1[4575:4568] > mid_0[4583:4576]) ? 1 : 0;
assign detect_max[570][12] = (mid_1[4575:4568] > mid_1[4567:4560]) ? 1 : 0;
assign detect_max[570][13] = (mid_1[4575:4568] > mid_1[4583:4576]) ? 1 : 0;
assign detect_max[570][14] = (mid_1[4575:4568] > mid_2[4567:4560]) ? 1 : 0;
assign detect_max[570][15] = (mid_1[4575:4568] > mid_2[4575:4568]) ? 1 : 0;
assign detect_max[570][16] = (mid_1[4575:4568] > mid_2[4583:4576]) ? 1 : 0;
assign detect_max[570][17] = (mid_1[4575:4568] > btm_0[4567:4560]) ? 1 : 0;
assign detect_max[570][18] = (mid_1[4575:4568] > btm_0[4575:4568]) ? 1 : 0;
assign detect_max[570][19] = (mid_1[4575:4568] > btm_0[4583:4576]) ? 1 : 0;
assign detect_max[570][20] = (mid_1[4575:4568] > btm_1[4567:4560]) ? 1 : 0;
assign detect_max[570][21] = (mid_1[4575:4568] > btm_1[4575:4568]) ? 1 : 0;
assign detect_max[570][22] = (mid_1[4575:4568] > btm_1[4583:4576]) ? 1 : 0;
assign detect_max[570][23] = (mid_1[4575:4568] > btm_2[4567:4560]) ? 1 : 0;
assign detect_max[570][24] = (mid_1[4575:4568] > btm_2[4575:4568]) ? 1 : 0;
assign detect_max[570][25] = (mid_1[4575:4568] > btm_2[4583:4576]) ? 1 : 0;

assign detect_max[571][0] = (mid_1[4583:4576] > top_0[4575:4568]) ? 1 : 0;
assign detect_max[571][1] = (mid_1[4583:4576] > top_0[4583:4576]) ? 1 : 0;
assign detect_max[571][2] = (mid_1[4583:4576] > top_0[4591:4584]) ? 1 : 0;
assign detect_max[571][3] = (mid_1[4583:4576] > top_1[4575:4568]) ? 1 : 0;
assign detect_max[571][4] = (mid_1[4583:4576] > top_1[4583:4576]) ? 1 : 0;
assign detect_max[571][5] = (mid_1[4583:4576] > top_1[4591:4584]) ? 1 : 0;
assign detect_max[571][6] = (mid_1[4583:4576] > top_2[4575:4568]) ? 1 : 0;
assign detect_max[571][7] = (mid_1[4583:4576] > top_2[4583:4576]) ? 1 : 0;
assign detect_max[571][8] = (mid_1[4583:4576] > top_2[4591:4584]) ? 1 : 0;
assign detect_max[571][9] = (mid_1[4583:4576] > mid_0[4575:4568]) ? 1 : 0;
assign detect_max[571][10] = (mid_1[4583:4576] > mid_0[4583:4576]) ? 1 : 0;
assign detect_max[571][11] = (mid_1[4583:4576] > mid_0[4591:4584]) ? 1 : 0;
assign detect_max[571][12] = (mid_1[4583:4576] > mid_1[4575:4568]) ? 1 : 0;
assign detect_max[571][13] = (mid_1[4583:4576] > mid_1[4591:4584]) ? 1 : 0;
assign detect_max[571][14] = (mid_1[4583:4576] > mid_2[4575:4568]) ? 1 : 0;
assign detect_max[571][15] = (mid_1[4583:4576] > mid_2[4583:4576]) ? 1 : 0;
assign detect_max[571][16] = (mid_1[4583:4576] > mid_2[4591:4584]) ? 1 : 0;
assign detect_max[571][17] = (mid_1[4583:4576] > btm_0[4575:4568]) ? 1 : 0;
assign detect_max[571][18] = (mid_1[4583:4576] > btm_0[4583:4576]) ? 1 : 0;
assign detect_max[571][19] = (mid_1[4583:4576] > btm_0[4591:4584]) ? 1 : 0;
assign detect_max[571][20] = (mid_1[4583:4576] > btm_1[4575:4568]) ? 1 : 0;
assign detect_max[571][21] = (mid_1[4583:4576] > btm_1[4583:4576]) ? 1 : 0;
assign detect_max[571][22] = (mid_1[4583:4576] > btm_1[4591:4584]) ? 1 : 0;
assign detect_max[571][23] = (mid_1[4583:4576] > btm_2[4575:4568]) ? 1 : 0;
assign detect_max[571][24] = (mid_1[4583:4576] > btm_2[4583:4576]) ? 1 : 0;
assign detect_max[571][25] = (mid_1[4583:4576] > btm_2[4591:4584]) ? 1 : 0;

assign detect_max[572][0] = (mid_1[4591:4584] > top_0[4583:4576]) ? 1 : 0;
assign detect_max[572][1] = (mid_1[4591:4584] > top_0[4591:4584]) ? 1 : 0;
assign detect_max[572][2] = (mid_1[4591:4584] > top_0[4599:4592]) ? 1 : 0;
assign detect_max[572][3] = (mid_1[4591:4584] > top_1[4583:4576]) ? 1 : 0;
assign detect_max[572][4] = (mid_1[4591:4584] > top_1[4591:4584]) ? 1 : 0;
assign detect_max[572][5] = (mid_1[4591:4584] > top_1[4599:4592]) ? 1 : 0;
assign detect_max[572][6] = (mid_1[4591:4584] > top_2[4583:4576]) ? 1 : 0;
assign detect_max[572][7] = (mid_1[4591:4584] > top_2[4591:4584]) ? 1 : 0;
assign detect_max[572][8] = (mid_1[4591:4584] > top_2[4599:4592]) ? 1 : 0;
assign detect_max[572][9] = (mid_1[4591:4584] > mid_0[4583:4576]) ? 1 : 0;
assign detect_max[572][10] = (mid_1[4591:4584] > mid_0[4591:4584]) ? 1 : 0;
assign detect_max[572][11] = (mid_1[4591:4584] > mid_0[4599:4592]) ? 1 : 0;
assign detect_max[572][12] = (mid_1[4591:4584] > mid_1[4583:4576]) ? 1 : 0;
assign detect_max[572][13] = (mid_1[4591:4584] > mid_1[4599:4592]) ? 1 : 0;
assign detect_max[572][14] = (mid_1[4591:4584] > mid_2[4583:4576]) ? 1 : 0;
assign detect_max[572][15] = (mid_1[4591:4584] > mid_2[4591:4584]) ? 1 : 0;
assign detect_max[572][16] = (mid_1[4591:4584] > mid_2[4599:4592]) ? 1 : 0;
assign detect_max[572][17] = (mid_1[4591:4584] > btm_0[4583:4576]) ? 1 : 0;
assign detect_max[572][18] = (mid_1[4591:4584] > btm_0[4591:4584]) ? 1 : 0;
assign detect_max[572][19] = (mid_1[4591:4584] > btm_0[4599:4592]) ? 1 : 0;
assign detect_max[572][20] = (mid_1[4591:4584] > btm_1[4583:4576]) ? 1 : 0;
assign detect_max[572][21] = (mid_1[4591:4584] > btm_1[4591:4584]) ? 1 : 0;
assign detect_max[572][22] = (mid_1[4591:4584] > btm_1[4599:4592]) ? 1 : 0;
assign detect_max[572][23] = (mid_1[4591:4584] > btm_2[4583:4576]) ? 1 : 0;
assign detect_max[572][24] = (mid_1[4591:4584] > btm_2[4591:4584]) ? 1 : 0;
assign detect_max[572][25] = (mid_1[4591:4584] > btm_2[4599:4592]) ? 1 : 0;

assign detect_max[573][0] = (mid_1[4599:4592] > top_0[4591:4584]) ? 1 : 0;
assign detect_max[573][1] = (mid_1[4599:4592] > top_0[4599:4592]) ? 1 : 0;
assign detect_max[573][2] = (mid_1[4599:4592] > top_0[4607:4600]) ? 1 : 0;
assign detect_max[573][3] = (mid_1[4599:4592] > top_1[4591:4584]) ? 1 : 0;
assign detect_max[573][4] = (mid_1[4599:4592] > top_1[4599:4592]) ? 1 : 0;
assign detect_max[573][5] = (mid_1[4599:4592] > top_1[4607:4600]) ? 1 : 0;
assign detect_max[573][6] = (mid_1[4599:4592] > top_2[4591:4584]) ? 1 : 0;
assign detect_max[573][7] = (mid_1[4599:4592] > top_2[4599:4592]) ? 1 : 0;
assign detect_max[573][8] = (mid_1[4599:4592] > top_2[4607:4600]) ? 1 : 0;
assign detect_max[573][9] = (mid_1[4599:4592] > mid_0[4591:4584]) ? 1 : 0;
assign detect_max[573][10] = (mid_1[4599:4592] > mid_0[4599:4592]) ? 1 : 0;
assign detect_max[573][11] = (mid_1[4599:4592] > mid_0[4607:4600]) ? 1 : 0;
assign detect_max[573][12] = (mid_1[4599:4592] > mid_1[4591:4584]) ? 1 : 0;
assign detect_max[573][13] = (mid_1[4599:4592] > mid_1[4607:4600]) ? 1 : 0;
assign detect_max[573][14] = (mid_1[4599:4592] > mid_2[4591:4584]) ? 1 : 0;
assign detect_max[573][15] = (mid_1[4599:4592] > mid_2[4599:4592]) ? 1 : 0;
assign detect_max[573][16] = (mid_1[4599:4592] > mid_2[4607:4600]) ? 1 : 0;
assign detect_max[573][17] = (mid_1[4599:4592] > btm_0[4591:4584]) ? 1 : 0;
assign detect_max[573][18] = (mid_1[4599:4592] > btm_0[4599:4592]) ? 1 : 0;
assign detect_max[573][19] = (mid_1[4599:4592] > btm_0[4607:4600]) ? 1 : 0;
assign detect_max[573][20] = (mid_1[4599:4592] > btm_1[4591:4584]) ? 1 : 0;
assign detect_max[573][21] = (mid_1[4599:4592] > btm_1[4599:4592]) ? 1 : 0;
assign detect_max[573][22] = (mid_1[4599:4592] > btm_1[4607:4600]) ? 1 : 0;
assign detect_max[573][23] = (mid_1[4599:4592] > btm_2[4591:4584]) ? 1 : 0;
assign detect_max[573][24] = (mid_1[4599:4592] > btm_2[4599:4592]) ? 1 : 0;
assign detect_max[573][25] = (mid_1[4599:4592] > btm_2[4607:4600]) ? 1 : 0;

assign detect_max[574][0] = (mid_1[4607:4600] > top_0[4599:4592]) ? 1 : 0;
assign detect_max[574][1] = (mid_1[4607:4600] > top_0[4607:4600]) ? 1 : 0;
assign detect_max[574][2] = (mid_1[4607:4600] > top_0[4615:4608]) ? 1 : 0;
assign detect_max[574][3] = (mid_1[4607:4600] > top_1[4599:4592]) ? 1 : 0;
assign detect_max[574][4] = (mid_1[4607:4600] > top_1[4607:4600]) ? 1 : 0;
assign detect_max[574][5] = (mid_1[4607:4600] > top_1[4615:4608]) ? 1 : 0;
assign detect_max[574][6] = (mid_1[4607:4600] > top_2[4599:4592]) ? 1 : 0;
assign detect_max[574][7] = (mid_1[4607:4600] > top_2[4607:4600]) ? 1 : 0;
assign detect_max[574][8] = (mid_1[4607:4600] > top_2[4615:4608]) ? 1 : 0;
assign detect_max[574][9] = (mid_1[4607:4600] > mid_0[4599:4592]) ? 1 : 0;
assign detect_max[574][10] = (mid_1[4607:4600] > mid_0[4607:4600]) ? 1 : 0;
assign detect_max[574][11] = (mid_1[4607:4600] > mid_0[4615:4608]) ? 1 : 0;
assign detect_max[574][12] = (mid_1[4607:4600] > mid_1[4599:4592]) ? 1 : 0;
assign detect_max[574][13] = (mid_1[4607:4600] > mid_1[4615:4608]) ? 1 : 0;
assign detect_max[574][14] = (mid_1[4607:4600] > mid_2[4599:4592]) ? 1 : 0;
assign detect_max[574][15] = (mid_1[4607:4600] > mid_2[4607:4600]) ? 1 : 0;
assign detect_max[574][16] = (mid_1[4607:4600] > mid_2[4615:4608]) ? 1 : 0;
assign detect_max[574][17] = (mid_1[4607:4600] > btm_0[4599:4592]) ? 1 : 0;
assign detect_max[574][18] = (mid_1[4607:4600] > btm_0[4607:4600]) ? 1 : 0;
assign detect_max[574][19] = (mid_1[4607:4600] > btm_0[4615:4608]) ? 1 : 0;
assign detect_max[574][20] = (mid_1[4607:4600] > btm_1[4599:4592]) ? 1 : 0;
assign detect_max[574][21] = (mid_1[4607:4600] > btm_1[4607:4600]) ? 1 : 0;
assign detect_max[574][22] = (mid_1[4607:4600] > btm_1[4615:4608]) ? 1 : 0;
assign detect_max[574][23] = (mid_1[4607:4600] > btm_2[4599:4592]) ? 1 : 0;
assign detect_max[574][24] = (mid_1[4607:4600] > btm_2[4607:4600]) ? 1 : 0;
assign detect_max[574][25] = (mid_1[4607:4600] > btm_2[4615:4608]) ? 1 : 0;

assign detect_max[575][0] = (mid_1[4615:4608] > top_0[4607:4600]) ? 1 : 0;
assign detect_max[575][1] = (mid_1[4615:4608] > top_0[4615:4608]) ? 1 : 0;
assign detect_max[575][2] = (mid_1[4615:4608] > top_0[4623:4616]) ? 1 : 0;
assign detect_max[575][3] = (mid_1[4615:4608] > top_1[4607:4600]) ? 1 : 0;
assign detect_max[575][4] = (mid_1[4615:4608] > top_1[4615:4608]) ? 1 : 0;
assign detect_max[575][5] = (mid_1[4615:4608] > top_1[4623:4616]) ? 1 : 0;
assign detect_max[575][6] = (mid_1[4615:4608] > top_2[4607:4600]) ? 1 : 0;
assign detect_max[575][7] = (mid_1[4615:4608] > top_2[4615:4608]) ? 1 : 0;
assign detect_max[575][8] = (mid_1[4615:4608] > top_2[4623:4616]) ? 1 : 0;
assign detect_max[575][9] = (mid_1[4615:4608] > mid_0[4607:4600]) ? 1 : 0;
assign detect_max[575][10] = (mid_1[4615:4608] > mid_0[4615:4608]) ? 1 : 0;
assign detect_max[575][11] = (mid_1[4615:4608] > mid_0[4623:4616]) ? 1 : 0;
assign detect_max[575][12] = (mid_1[4615:4608] > mid_1[4607:4600]) ? 1 : 0;
assign detect_max[575][13] = (mid_1[4615:4608] > mid_1[4623:4616]) ? 1 : 0;
assign detect_max[575][14] = (mid_1[4615:4608] > mid_2[4607:4600]) ? 1 : 0;
assign detect_max[575][15] = (mid_1[4615:4608] > mid_2[4615:4608]) ? 1 : 0;
assign detect_max[575][16] = (mid_1[4615:4608] > mid_2[4623:4616]) ? 1 : 0;
assign detect_max[575][17] = (mid_1[4615:4608] > btm_0[4607:4600]) ? 1 : 0;
assign detect_max[575][18] = (mid_1[4615:4608] > btm_0[4615:4608]) ? 1 : 0;
assign detect_max[575][19] = (mid_1[4615:4608] > btm_0[4623:4616]) ? 1 : 0;
assign detect_max[575][20] = (mid_1[4615:4608] > btm_1[4607:4600]) ? 1 : 0;
assign detect_max[575][21] = (mid_1[4615:4608] > btm_1[4615:4608]) ? 1 : 0;
assign detect_max[575][22] = (mid_1[4615:4608] > btm_1[4623:4616]) ? 1 : 0;
assign detect_max[575][23] = (mid_1[4615:4608] > btm_2[4607:4600]) ? 1 : 0;
assign detect_max[575][24] = (mid_1[4615:4608] > btm_2[4615:4608]) ? 1 : 0;
assign detect_max[575][25] = (mid_1[4615:4608] > btm_2[4623:4616]) ? 1 : 0;

assign detect_max[576][0] = (mid_1[4623:4616] > top_0[4615:4608]) ? 1 : 0;
assign detect_max[576][1] = (mid_1[4623:4616] > top_0[4623:4616]) ? 1 : 0;
assign detect_max[576][2] = (mid_1[4623:4616] > top_0[4631:4624]) ? 1 : 0;
assign detect_max[576][3] = (mid_1[4623:4616] > top_1[4615:4608]) ? 1 : 0;
assign detect_max[576][4] = (mid_1[4623:4616] > top_1[4623:4616]) ? 1 : 0;
assign detect_max[576][5] = (mid_1[4623:4616] > top_1[4631:4624]) ? 1 : 0;
assign detect_max[576][6] = (mid_1[4623:4616] > top_2[4615:4608]) ? 1 : 0;
assign detect_max[576][7] = (mid_1[4623:4616] > top_2[4623:4616]) ? 1 : 0;
assign detect_max[576][8] = (mid_1[4623:4616] > top_2[4631:4624]) ? 1 : 0;
assign detect_max[576][9] = (mid_1[4623:4616] > mid_0[4615:4608]) ? 1 : 0;
assign detect_max[576][10] = (mid_1[4623:4616] > mid_0[4623:4616]) ? 1 : 0;
assign detect_max[576][11] = (mid_1[4623:4616] > mid_0[4631:4624]) ? 1 : 0;
assign detect_max[576][12] = (mid_1[4623:4616] > mid_1[4615:4608]) ? 1 : 0;
assign detect_max[576][13] = (mid_1[4623:4616] > mid_1[4631:4624]) ? 1 : 0;
assign detect_max[576][14] = (mid_1[4623:4616] > mid_2[4615:4608]) ? 1 : 0;
assign detect_max[576][15] = (mid_1[4623:4616] > mid_2[4623:4616]) ? 1 : 0;
assign detect_max[576][16] = (mid_1[4623:4616] > mid_2[4631:4624]) ? 1 : 0;
assign detect_max[576][17] = (mid_1[4623:4616] > btm_0[4615:4608]) ? 1 : 0;
assign detect_max[576][18] = (mid_1[4623:4616] > btm_0[4623:4616]) ? 1 : 0;
assign detect_max[576][19] = (mid_1[4623:4616] > btm_0[4631:4624]) ? 1 : 0;
assign detect_max[576][20] = (mid_1[4623:4616] > btm_1[4615:4608]) ? 1 : 0;
assign detect_max[576][21] = (mid_1[4623:4616] > btm_1[4623:4616]) ? 1 : 0;
assign detect_max[576][22] = (mid_1[4623:4616] > btm_1[4631:4624]) ? 1 : 0;
assign detect_max[576][23] = (mid_1[4623:4616] > btm_2[4615:4608]) ? 1 : 0;
assign detect_max[576][24] = (mid_1[4623:4616] > btm_2[4623:4616]) ? 1 : 0;
assign detect_max[576][25] = (mid_1[4623:4616] > btm_2[4631:4624]) ? 1 : 0;

assign detect_max[577][0] = (mid_1[4631:4624] > top_0[4623:4616]) ? 1 : 0;
assign detect_max[577][1] = (mid_1[4631:4624] > top_0[4631:4624]) ? 1 : 0;
assign detect_max[577][2] = (mid_1[4631:4624] > top_0[4639:4632]) ? 1 : 0;
assign detect_max[577][3] = (mid_1[4631:4624] > top_1[4623:4616]) ? 1 : 0;
assign detect_max[577][4] = (mid_1[4631:4624] > top_1[4631:4624]) ? 1 : 0;
assign detect_max[577][5] = (mid_1[4631:4624] > top_1[4639:4632]) ? 1 : 0;
assign detect_max[577][6] = (mid_1[4631:4624] > top_2[4623:4616]) ? 1 : 0;
assign detect_max[577][7] = (mid_1[4631:4624] > top_2[4631:4624]) ? 1 : 0;
assign detect_max[577][8] = (mid_1[4631:4624] > top_2[4639:4632]) ? 1 : 0;
assign detect_max[577][9] = (mid_1[4631:4624] > mid_0[4623:4616]) ? 1 : 0;
assign detect_max[577][10] = (mid_1[4631:4624] > mid_0[4631:4624]) ? 1 : 0;
assign detect_max[577][11] = (mid_1[4631:4624] > mid_0[4639:4632]) ? 1 : 0;
assign detect_max[577][12] = (mid_1[4631:4624] > mid_1[4623:4616]) ? 1 : 0;
assign detect_max[577][13] = (mid_1[4631:4624] > mid_1[4639:4632]) ? 1 : 0;
assign detect_max[577][14] = (mid_1[4631:4624] > mid_2[4623:4616]) ? 1 : 0;
assign detect_max[577][15] = (mid_1[4631:4624] > mid_2[4631:4624]) ? 1 : 0;
assign detect_max[577][16] = (mid_1[4631:4624] > mid_2[4639:4632]) ? 1 : 0;
assign detect_max[577][17] = (mid_1[4631:4624] > btm_0[4623:4616]) ? 1 : 0;
assign detect_max[577][18] = (mid_1[4631:4624] > btm_0[4631:4624]) ? 1 : 0;
assign detect_max[577][19] = (mid_1[4631:4624] > btm_0[4639:4632]) ? 1 : 0;
assign detect_max[577][20] = (mid_1[4631:4624] > btm_1[4623:4616]) ? 1 : 0;
assign detect_max[577][21] = (mid_1[4631:4624] > btm_1[4631:4624]) ? 1 : 0;
assign detect_max[577][22] = (mid_1[4631:4624] > btm_1[4639:4632]) ? 1 : 0;
assign detect_max[577][23] = (mid_1[4631:4624] > btm_2[4623:4616]) ? 1 : 0;
assign detect_max[577][24] = (mid_1[4631:4624] > btm_2[4631:4624]) ? 1 : 0;
assign detect_max[577][25] = (mid_1[4631:4624] > btm_2[4639:4632]) ? 1 : 0;

assign detect_max[578][0] = (mid_1[4639:4632] > top_0[4631:4624]) ? 1 : 0;
assign detect_max[578][1] = (mid_1[4639:4632] > top_0[4639:4632]) ? 1 : 0;
assign detect_max[578][2] = (mid_1[4639:4632] > top_0[4647:4640]) ? 1 : 0;
assign detect_max[578][3] = (mid_1[4639:4632] > top_1[4631:4624]) ? 1 : 0;
assign detect_max[578][4] = (mid_1[4639:4632] > top_1[4639:4632]) ? 1 : 0;
assign detect_max[578][5] = (mid_1[4639:4632] > top_1[4647:4640]) ? 1 : 0;
assign detect_max[578][6] = (mid_1[4639:4632] > top_2[4631:4624]) ? 1 : 0;
assign detect_max[578][7] = (mid_1[4639:4632] > top_2[4639:4632]) ? 1 : 0;
assign detect_max[578][8] = (mid_1[4639:4632] > top_2[4647:4640]) ? 1 : 0;
assign detect_max[578][9] = (mid_1[4639:4632] > mid_0[4631:4624]) ? 1 : 0;
assign detect_max[578][10] = (mid_1[4639:4632] > mid_0[4639:4632]) ? 1 : 0;
assign detect_max[578][11] = (mid_1[4639:4632] > mid_0[4647:4640]) ? 1 : 0;
assign detect_max[578][12] = (mid_1[4639:4632] > mid_1[4631:4624]) ? 1 : 0;
assign detect_max[578][13] = (mid_1[4639:4632] > mid_1[4647:4640]) ? 1 : 0;
assign detect_max[578][14] = (mid_1[4639:4632] > mid_2[4631:4624]) ? 1 : 0;
assign detect_max[578][15] = (mid_1[4639:4632] > mid_2[4639:4632]) ? 1 : 0;
assign detect_max[578][16] = (mid_1[4639:4632] > mid_2[4647:4640]) ? 1 : 0;
assign detect_max[578][17] = (mid_1[4639:4632] > btm_0[4631:4624]) ? 1 : 0;
assign detect_max[578][18] = (mid_1[4639:4632] > btm_0[4639:4632]) ? 1 : 0;
assign detect_max[578][19] = (mid_1[4639:4632] > btm_0[4647:4640]) ? 1 : 0;
assign detect_max[578][20] = (mid_1[4639:4632] > btm_1[4631:4624]) ? 1 : 0;
assign detect_max[578][21] = (mid_1[4639:4632] > btm_1[4639:4632]) ? 1 : 0;
assign detect_max[578][22] = (mid_1[4639:4632] > btm_1[4647:4640]) ? 1 : 0;
assign detect_max[578][23] = (mid_1[4639:4632] > btm_2[4631:4624]) ? 1 : 0;
assign detect_max[578][24] = (mid_1[4639:4632] > btm_2[4639:4632]) ? 1 : 0;
assign detect_max[578][25] = (mid_1[4639:4632] > btm_2[4647:4640]) ? 1 : 0;

assign detect_max[579][0] = (mid_1[4647:4640] > top_0[4639:4632]) ? 1 : 0;
assign detect_max[579][1] = (mid_1[4647:4640] > top_0[4647:4640]) ? 1 : 0;
assign detect_max[579][2] = (mid_1[4647:4640] > top_0[4655:4648]) ? 1 : 0;
assign detect_max[579][3] = (mid_1[4647:4640] > top_1[4639:4632]) ? 1 : 0;
assign detect_max[579][4] = (mid_1[4647:4640] > top_1[4647:4640]) ? 1 : 0;
assign detect_max[579][5] = (mid_1[4647:4640] > top_1[4655:4648]) ? 1 : 0;
assign detect_max[579][6] = (mid_1[4647:4640] > top_2[4639:4632]) ? 1 : 0;
assign detect_max[579][7] = (mid_1[4647:4640] > top_2[4647:4640]) ? 1 : 0;
assign detect_max[579][8] = (mid_1[4647:4640] > top_2[4655:4648]) ? 1 : 0;
assign detect_max[579][9] = (mid_1[4647:4640] > mid_0[4639:4632]) ? 1 : 0;
assign detect_max[579][10] = (mid_1[4647:4640] > mid_0[4647:4640]) ? 1 : 0;
assign detect_max[579][11] = (mid_1[4647:4640] > mid_0[4655:4648]) ? 1 : 0;
assign detect_max[579][12] = (mid_1[4647:4640] > mid_1[4639:4632]) ? 1 : 0;
assign detect_max[579][13] = (mid_1[4647:4640] > mid_1[4655:4648]) ? 1 : 0;
assign detect_max[579][14] = (mid_1[4647:4640] > mid_2[4639:4632]) ? 1 : 0;
assign detect_max[579][15] = (mid_1[4647:4640] > mid_2[4647:4640]) ? 1 : 0;
assign detect_max[579][16] = (mid_1[4647:4640] > mid_2[4655:4648]) ? 1 : 0;
assign detect_max[579][17] = (mid_1[4647:4640] > btm_0[4639:4632]) ? 1 : 0;
assign detect_max[579][18] = (mid_1[4647:4640] > btm_0[4647:4640]) ? 1 : 0;
assign detect_max[579][19] = (mid_1[4647:4640] > btm_0[4655:4648]) ? 1 : 0;
assign detect_max[579][20] = (mid_1[4647:4640] > btm_1[4639:4632]) ? 1 : 0;
assign detect_max[579][21] = (mid_1[4647:4640] > btm_1[4647:4640]) ? 1 : 0;
assign detect_max[579][22] = (mid_1[4647:4640] > btm_1[4655:4648]) ? 1 : 0;
assign detect_max[579][23] = (mid_1[4647:4640] > btm_2[4639:4632]) ? 1 : 0;
assign detect_max[579][24] = (mid_1[4647:4640] > btm_2[4647:4640]) ? 1 : 0;
assign detect_max[579][25] = (mid_1[4647:4640] > btm_2[4655:4648]) ? 1 : 0;

assign detect_max[580][0] = (mid_1[4655:4648] > top_0[4647:4640]) ? 1 : 0;
assign detect_max[580][1] = (mid_1[4655:4648] > top_0[4655:4648]) ? 1 : 0;
assign detect_max[580][2] = (mid_1[4655:4648] > top_0[4663:4656]) ? 1 : 0;
assign detect_max[580][3] = (mid_1[4655:4648] > top_1[4647:4640]) ? 1 : 0;
assign detect_max[580][4] = (mid_1[4655:4648] > top_1[4655:4648]) ? 1 : 0;
assign detect_max[580][5] = (mid_1[4655:4648] > top_1[4663:4656]) ? 1 : 0;
assign detect_max[580][6] = (mid_1[4655:4648] > top_2[4647:4640]) ? 1 : 0;
assign detect_max[580][7] = (mid_1[4655:4648] > top_2[4655:4648]) ? 1 : 0;
assign detect_max[580][8] = (mid_1[4655:4648] > top_2[4663:4656]) ? 1 : 0;
assign detect_max[580][9] = (mid_1[4655:4648] > mid_0[4647:4640]) ? 1 : 0;
assign detect_max[580][10] = (mid_1[4655:4648] > mid_0[4655:4648]) ? 1 : 0;
assign detect_max[580][11] = (mid_1[4655:4648] > mid_0[4663:4656]) ? 1 : 0;
assign detect_max[580][12] = (mid_1[4655:4648] > mid_1[4647:4640]) ? 1 : 0;
assign detect_max[580][13] = (mid_1[4655:4648] > mid_1[4663:4656]) ? 1 : 0;
assign detect_max[580][14] = (mid_1[4655:4648] > mid_2[4647:4640]) ? 1 : 0;
assign detect_max[580][15] = (mid_1[4655:4648] > mid_2[4655:4648]) ? 1 : 0;
assign detect_max[580][16] = (mid_1[4655:4648] > mid_2[4663:4656]) ? 1 : 0;
assign detect_max[580][17] = (mid_1[4655:4648] > btm_0[4647:4640]) ? 1 : 0;
assign detect_max[580][18] = (mid_1[4655:4648] > btm_0[4655:4648]) ? 1 : 0;
assign detect_max[580][19] = (mid_1[4655:4648] > btm_0[4663:4656]) ? 1 : 0;
assign detect_max[580][20] = (mid_1[4655:4648] > btm_1[4647:4640]) ? 1 : 0;
assign detect_max[580][21] = (mid_1[4655:4648] > btm_1[4655:4648]) ? 1 : 0;
assign detect_max[580][22] = (mid_1[4655:4648] > btm_1[4663:4656]) ? 1 : 0;
assign detect_max[580][23] = (mid_1[4655:4648] > btm_2[4647:4640]) ? 1 : 0;
assign detect_max[580][24] = (mid_1[4655:4648] > btm_2[4655:4648]) ? 1 : 0;
assign detect_max[580][25] = (mid_1[4655:4648] > btm_2[4663:4656]) ? 1 : 0;

assign detect_max[581][0] = (mid_1[4663:4656] > top_0[4655:4648]) ? 1 : 0;
assign detect_max[581][1] = (mid_1[4663:4656] > top_0[4663:4656]) ? 1 : 0;
assign detect_max[581][2] = (mid_1[4663:4656] > top_0[4671:4664]) ? 1 : 0;
assign detect_max[581][3] = (mid_1[4663:4656] > top_1[4655:4648]) ? 1 : 0;
assign detect_max[581][4] = (mid_1[4663:4656] > top_1[4663:4656]) ? 1 : 0;
assign detect_max[581][5] = (mid_1[4663:4656] > top_1[4671:4664]) ? 1 : 0;
assign detect_max[581][6] = (mid_1[4663:4656] > top_2[4655:4648]) ? 1 : 0;
assign detect_max[581][7] = (mid_1[4663:4656] > top_2[4663:4656]) ? 1 : 0;
assign detect_max[581][8] = (mid_1[4663:4656] > top_2[4671:4664]) ? 1 : 0;
assign detect_max[581][9] = (mid_1[4663:4656] > mid_0[4655:4648]) ? 1 : 0;
assign detect_max[581][10] = (mid_1[4663:4656] > mid_0[4663:4656]) ? 1 : 0;
assign detect_max[581][11] = (mid_1[4663:4656] > mid_0[4671:4664]) ? 1 : 0;
assign detect_max[581][12] = (mid_1[4663:4656] > mid_1[4655:4648]) ? 1 : 0;
assign detect_max[581][13] = (mid_1[4663:4656] > mid_1[4671:4664]) ? 1 : 0;
assign detect_max[581][14] = (mid_1[4663:4656] > mid_2[4655:4648]) ? 1 : 0;
assign detect_max[581][15] = (mid_1[4663:4656] > mid_2[4663:4656]) ? 1 : 0;
assign detect_max[581][16] = (mid_1[4663:4656] > mid_2[4671:4664]) ? 1 : 0;
assign detect_max[581][17] = (mid_1[4663:4656] > btm_0[4655:4648]) ? 1 : 0;
assign detect_max[581][18] = (mid_1[4663:4656] > btm_0[4663:4656]) ? 1 : 0;
assign detect_max[581][19] = (mid_1[4663:4656] > btm_0[4671:4664]) ? 1 : 0;
assign detect_max[581][20] = (mid_1[4663:4656] > btm_1[4655:4648]) ? 1 : 0;
assign detect_max[581][21] = (mid_1[4663:4656] > btm_1[4663:4656]) ? 1 : 0;
assign detect_max[581][22] = (mid_1[4663:4656] > btm_1[4671:4664]) ? 1 : 0;
assign detect_max[581][23] = (mid_1[4663:4656] > btm_2[4655:4648]) ? 1 : 0;
assign detect_max[581][24] = (mid_1[4663:4656] > btm_2[4663:4656]) ? 1 : 0;
assign detect_max[581][25] = (mid_1[4663:4656] > btm_2[4671:4664]) ? 1 : 0;

assign detect_max[582][0] = (mid_1[4671:4664] > top_0[4663:4656]) ? 1 : 0;
assign detect_max[582][1] = (mid_1[4671:4664] > top_0[4671:4664]) ? 1 : 0;
assign detect_max[582][2] = (mid_1[4671:4664] > top_0[4679:4672]) ? 1 : 0;
assign detect_max[582][3] = (mid_1[4671:4664] > top_1[4663:4656]) ? 1 : 0;
assign detect_max[582][4] = (mid_1[4671:4664] > top_1[4671:4664]) ? 1 : 0;
assign detect_max[582][5] = (mid_1[4671:4664] > top_1[4679:4672]) ? 1 : 0;
assign detect_max[582][6] = (mid_1[4671:4664] > top_2[4663:4656]) ? 1 : 0;
assign detect_max[582][7] = (mid_1[4671:4664] > top_2[4671:4664]) ? 1 : 0;
assign detect_max[582][8] = (mid_1[4671:4664] > top_2[4679:4672]) ? 1 : 0;
assign detect_max[582][9] = (mid_1[4671:4664] > mid_0[4663:4656]) ? 1 : 0;
assign detect_max[582][10] = (mid_1[4671:4664] > mid_0[4671:4664]) ? 1 : 0;
assign detect_max[582][11] = (mid_1[4671:4664] > mid_0[4679:4672]) ? 1 : 0;
assign detect_max[582][12] = (mid_1[4671:4664] > mid_1[4663:4656]) ? 1 : 0;
assign detect_max[582][13] = (mid_1[4671:4664] > mid_1[4679:4672]) ? 1 : 0;
assign detect_max[582][14] = (mid_1[4671:4664] > mid_2[4663:4656]) ? 1 : 0;
assign detect_max[582][15] = (mid_1[4671:4664] > mid_2[4671:4664]) ? 1 : 0;
assign detect_max[582][16] = (mid_1[4671:4664] > mid_2[4679:4672]) ? 1 : 0;
assign detect_max[582][17] = (mid_1[4671:4664] > btm_0[4663:4656]) ? 1 : 0;
assign detect_max[582][18] = (mid_1[4671:4664] > btm_0[4671:4664]) ? 1 : 0;
assign detect_max[582][19] = (mid_1[4671:4664] > btm_0[4679:4672]) ? 1 : 0;
assign detect_max[582][20] = (mid_1[4671:4664] > btm_1[4663:4656]) ? 1 : 0;
assign detect_max[582][21] = (mid_1[4671:4664] > btm_1[4671:4664]) ? 1 : 0;
assign detect_max[582][22] = (mid_1[4671:4664] > btm_1[4679:4672]) ? 1 : 0;
assign detect_max[582][23] = (mid_1[4671:4664] > btm_2[4663:4656]) ? 1 : 0;
assign detect_max[582][24] = (mid_1[4671:4664] > btm_2[4671:4664]) ? 1 : 0;
assign detect_max[582][25] = (mid_1[4671:4664] > btm_2[4679:4672]) ? 1 : 0;

assign detect_max[583][0] = (mid_1[4679:4672] > top_0[4671:4664]) ? 1 : 0;
assign detect_max[583][1] = (mid_1[4679:4672] > top_0[4679:4672]) ? 1 : 0;
assign detect_max[583][2] = (mid_1[4679:4672] > top_0[4687:4680]) ? 1 : 0;
assign detect_max[583][3] = (mid_1[4679:4672] > top_1[4671:4664]) ? 1 : 0;
assign detect_max[583][4] = (mid_1[4679:4672] > top_1[4679:4672]) ? 1 : 0;
assign detect_max[583][5] = (mid_1[4679:4672] > top_1[4687:4680]) ? 1 : 0;
assign detect_max[583][6] = (mid_1[4679:4672] > top_2[4671:4664]) ? 1 : 0;
assign detect_max[583][7] = (mid_1[4679:4672] > top_2[4679:4672]) ? 1 : 0;
assign detect_max[583][8] = (mid_1[4679:4672] > top_2[4687:4680]) ? 1 : 0;
assign detect_max[583][9] = (mid_1[4679:4672] > mid_0[4671:4664]) ? 1 : 0;
assign detect_max[583][10] = (mid_1[4679:4672] > mid_0[4679:4672]) ? 1 : 0;
assign detect_max[583][11] = (mid_1[4679:4672] > mid_0[4687:4680]) ? 1 : 0;
assign detect_max[583][12] = (mid_1[4679:4672] > mid_1[4671:4664]) ? 1 : 0;
assign detect_max[583][13] = (mid_1[4679:4672] > mid_1[4687:4680]) ? 1 : 0;
assign detect_max[583][14] = (mid_1[4679:4672] > mid_2[4671:4664]) ? 1 : 0;
assign detect_max[583][15] = (mid_1[4679:4672] > mid_2[4679:4672]) ? 1 : 0;
assign detect_max[583][16] = (mid_1[4679:4672] > mid_2[4687:4680]) ? 1 : 0;
assign detect_max[583][17] = (mid_1[4679:4672] > btm_0[4671:4664]) ? 1 : 0;
assign detect_max[583][18] = (mid_1[4679:4672] > btm_0[4679:4672]) ? 1 : 0;
assign detect_max[583][19] = (mid_1[4679:4672] > btm_0[4687:4680]) ? 1 : 0;
assign detect_max[583][20] = (mid_1[4679:4672] > btm_1[4671:4664]) ? 1 : 0;
assign detect_max[583][21] = (mid_1[4679:4672] > btm_1[4679:4672]) ? 1 : 0;
assign detect_max[583][22] = (mid_1[4679:4672] > btm_1[4687:4680]) ? 1 : 0;
assign detect_max[583][23] = (mid_1[4679:4672] > btm_2[4671:4664]) ? 1 : 0;
assign detect_max[583][24] = (mid_1[4679:4672] > btm_2[4679:4672]) ? 1 : 0;
assign detect_max[583][25] = (mid_1[4679:4672] > btm_2[4687:4680]) ? 1 : 0;

assign detect_max[584][0] = (mid_1[4687:4680] > top_0[4679:4672]) ? 1 : 0;
assign detect_max[584][1] = (mid_1[4687:4680] > top_0[4687:4680]) ? 1 : 0;
assign detect_max[584][2] = (mid_1[4687:4680] > top_0[4695:4688]) ? 1 : 0;
assign detect_max[584][3] = (mid_1[4687:4680] > top_1[4679:4672]) ? 1 : 0;
assign detect_max[584][4] = (mid_1[4687:4680] > top_1[4687:4680]) ? 1 : 0;
assign detect_max[584][5] = (mid_1[4687:4680] > top_1[4695:4688]) ? 1 : 0;
assign detect_max[584][6] = (mid_1[4687:4680] > top_2[4679:4672]) ? 1 : 0;
assign detect_max[584][7] = (mid_1[4687:4680] > top_2[4687:4680]) ? 1 : 0;
assign detect_max[584][8] = (mid_1[4687:4680] > top_2[4695:4688]) ? 1 : 0;
assign detect_max[584][9] = (mid_1[4687:4680] > mid_0[4679:4672]) ? 1 : 0;
assign detect_max[584][10] = (mid_1[4687:4680] > mid_0[4687:4680]) ? 1 : 0;
assign detect_max[584][11] = (mid_1[4687:4680] > mid_0[4695:4688]) ? 1 : 0;
assign detect_max[584][12] = (mid_1[4687:4680] > mid_1[4679:4672]) ? 1 : 0;
assign detect_max[584][13] = (mid_1[4687:4680] > mid_1[4695:4688]) ? 1 : 0;
assign detect_max[584][14] = (mid_1[4687:4680] > mid_2[4679:4672]) ? 1 : 0;
assign detect_max[584][15] = (mid_1[4687:4680] > mid_2[4687:4680]) ? 1 : 0;
assign detect_max[584][16] = (mid_1[4687:4680] > mid_2[4695:4688]) ? 1 : 0;
assign detect_max[584][17] = (mid_1[4687:4680] > btm_0[4679:4672]) ? 1 : 0;
assign detect_max[584][18] = (mid_1[4687:4680] > btm_0[4687:4680]) ? 1 : 0;
assign detect_max[584][19] = (mid_1[4687:4680] > btm_0[4695:4688]) ? 1 : 0;
assign detect_max[584][20] = (mid_1[4687:4680] > btm_1[4679:4672]) ? 1 : 0;
assign detect_max[584][21] = (mid_1[4687:4680] > btm_1[4687:4680]) ? 1 : 0;
assign detect_max[584][22] = (mid_1[4687:4680] > btm_1[4695:4688]) ? 1 : 0;
assign detect_max[584][23] = (mid_1[4687:4680] > btm_2[4679:4672]) ? 1 : 0;
assign detect_max[584][24] = (mid_1[4687:4680] > btm_2[4687:4680]) ? 1 : 0;
assign detect_max[584][25] = (mid_1[4687:4680] > btm_2[4695:4688]) ? 1 : 0;

assign detect_max[585][0] = (mid_1[4695:4688] > top_0[4687:4680]) ? 1 : 0;
assign detect_max[585][1] = (mid_1[4695:4688] > top_0[4695:4688]) ? 1 : 0;
assign detect_max[585][2] = (mid_1[4695:4688] > top_0[4703:4696]) ? 1 : 0;
assign detect_max[585][3] = (mid_1[4695:4688] > top_1[4687:4680]) ? 1 : 0;
assign detect_max[585][4] = (mid_1[4695:4688] > top_1[4695:4688]) ? 1 : 0;
assign detect_max[585][5] = (mid_1[4695:4688] > top_1[4703:4696]) ? 1 : 0;
assign detect_max[585][6] = (mid_1[4695:4688] > top_2[4687:4680]) ? 1 : 0;
assign detect_max[585][7] = (mid_1[4695:4688] > top_2[4695:4688]) ? 1 : 0;
assign detect_max[585][8] = (mid_1[4695:4688] > top_2[4703:4696]) ? 1 : 0;
assign detect_max[585][9] = (mid_1[4695:4688] > mid_0[4687:4680]) ? 1 : 0;
assign detect_max[585][10] = (mid_1[4695:4688] > mid_0[4695:4688]) ? 1 : 0;
assign detect_max[585][11] = (mid_1[4695:4688] > mid_0[4703:4696]) ? 1 : 0;
assign detect_max[585][12] = (mid_1[4695:4688] > mid_1[4687:4680]) ? 1 : 0;
assign detect_max[585][13] = (mid_1[4695:4688] > mid_1[4703:4696]) ? 1 : 0;
assign detect_max[585][14] = (mid_1[4695:4688] > mid_2[4687:4680]) ? 1 : 0;
assign detect_max[585][15] = (mid_1[4695:4688] > mid_2[4695:4688]) ? 1 : 0;
assign detect_max[585][16] = (mid_1[4695:4688] > mid_2[4703:4696]) ? 1 : 0;
assign detect_max[585][17] = (mid_1[4695:4688] > btm_0[4687:4680]) ? 1 : 0;
assign detect_max[585][18] = (mid_1[4695:4688] > btm_0[4695:4688]) ? 1 : 0;
assign detect_max[585][19] = (mid_1[4695:4688] > btm_0[4703:4696]) ? 1 : 0;
assign detect_max[585][20] = (mid_1[4695:4688] > btm_1[4687:4680]) ? 1 : 0;
assign detect_max[585][21] = (mid_1[4695:4688] > btm_1[4695:4688]) ? 1 : 0;
assign detect_max[585][22] = (mid_1[4695:4688] > btm_1[4703:4696]) ? 1 : 0;
assign detect_max[585][23] = (mid_1[4695:4688] > btm_2[4687:4680]) ? 1 : 0;
assign detect_max[585][24] = (mid_1[4695:4688] > btm_2[4695:4688]) ? 1 : 0;
assign detect_max[585][25] = (mid_1[4695:4688] > btm_2[4703:4696]) ? 1 : 0;

assign detect_max[586][0] = (mid_1[4703:4696] > top_0[4695:4688]) ? 1 : 0;
assign detect_max[586][1] = (mid_1[4703:4696] > top_0[4703:4696]) ? 1 : 0;
assign detect_max[586][2] = (mid_1[4703:4696] > top_0[4711:4704]) ? 1 : 0;
assign detect_max[586][3] = (mid_1[4703:4696] > top_1[4695:4688]) ? 1 : 0;
assign detect_max[586][4] = (mid_1[4703:4696] > top_1[4703:4696]) ? 1 : 0;
assign detect_max[586][5] = (mid_1[4703:4696] > top_1[4711:4704]) ? 1 : 0;
assign detect_max[586][6] = (mid_1[4703:4696] > top_2[4695:4688]) ? 1 : 0;
assign detect_max[586][7] = (mid_1[4703:4696] > top_2[4703:4696]) ? 1 : 0;
assign detect_max[586][8] = (mid_1[4703:4696] > top_2[4711:4704]) ? 1 : 0;
assign detect_max[586][9] = (mid_1[4703:4696] > mid_0[4695:4688]) ? 1 : 0;
assign detect_max[586][10] = (mid_1[4703:4696] > mid_0[4703:4696]) ? 1 : 0;
assign detect_max[586][11] = (mid_1[4703:4696] > mid_0[4711:4704]) ? 1 : 0;
assign detect_max[586][12] = (mid_1[4703:4696] > mid_1[4695:4688]) ? 1 : 0;
assign detect_max[586][13] = (mid_1[4703:4696] > mid_1[4711:4704]) ? 1 : 0;
assign detect_max[586][14] = (mid_1[4703:4696] > mid_2[4695:4688]) ? 1 : 0;
assign detect_max[586][15] = (mid_1[4703:4696] > mid_2[4703:4696]) ? 1 : 0;
assign detect_max[586][16] = (mid_1[4703:4696] > mid_2[4711:4704]) ? 1 : 0;
assign detect_max[586][17] = (mid_1[4703:4696] > btm_0[4695:4688]) ? 1 : 0;
assign detect_max[586][18] = (mid_1[4703:4696] > btm_0[4703:4696]) ? 1 : 0;
assign detect_max[586][19] = (mid_1[4703:4696] > btm_0[4711:4704]) ? 1 : 0;
assign detect_max[586][20] = (mid_1[4703:4696] > btm_1[4695:4688]) ? 1 : 0;
assign detect_max[586][21] = (mid_1[4703:4696] > btm_1[4703:4696]) ? 1 : 0;
assign detect_max[586][22] = (mid_1[4703:4696] > btm_1[4711:4704]) ? 1 : 0;
assign detect_max[586][23] = (mid_1[4703:4696] > btm_2[4695:4688]) ? 1 : 0;
assign detect_max[586][24] = (mid_1[4703:4696] > btm_2[4703:4696]) ? 1 : 0;
assign detect_max[586][25] = (mid_1[4703:4696] > btm_2[4711:4704]) ? 1 : 0;

assign detect_max[587][0] = (mid_1[4711:4704] > top_0[4703:4696]) ? 1 : 0;
assign detect_max[587][1] = (mid_1[4711:4704] > top_0[4711:4704]) ? 1 : 0;
assign detect_max[587][2] = (mid_1[4711:4704] > top_0[4719:4712]) ? 1 : 0;
assign detect_max[587][3] = (mid_1[4711:4704] > top_1[4703:4696]) ? 1 : 0;
assign detect_max[587][4] = (mid_1[4711:4704] > top_1[4711:4704]) ? 1 : 0;
assign detect_max[587][5] = (mid_1[4711:4704] > top_1[4719:4712]) ? 1 : 0;
assign detect_max[587][6] = (mid_1[4711:4704] > top_2[4703:4696]) ? 1 : 0;
assign detect_max[587][7] = (mid_1[4711:4704] > top_2[4711:4704]) ? 1 : 0;
assign detect_max[587][8] = (mid_1[4711:4704] > top_2[4719:4712]) ? 1 : 0;
assign detect_max[587][9] = (mid_1[4711:4704] > mid_0[4703:4696]) ? 1 : 0;
assign detect_max[587][10] = (mid_1[4711:4704] > mid_0[4711:4704]) ? 1 : 0;
assign detect_max[587][11] = (mid_1[4711:4704] > mid_0[4719:4712]) ? 1 : 0;
assign detect_max[587][12] = (mid_1[4711:4704] > mid_1[4703:4696]) ? 1 : 0;
assign detect_max[587][13] = (mid_1[4711:4704] > mid_1[4719:4712]) ? 1 : 0;
assign detect_max[587][14] = (mid_1[4711:4704] > mid_2[4703:4696]) ? 1 : 0;
assign detect_max[587][15] = (mid_1[4711:4704] > mid_2[4711:4704]) ? 1 : 0;
assign detect_max[587][16] = (mid_1[4711:4704] > mid_2[4719:4712]) ? 1 : 0;
assign detect_max[587][17] = (mid_1[4711:4704] > btm_0[4703:4696]) ? 1 : 0;
assign detect_max[587][18] = (mid_1[4711:4704] > btm_0[4711:4704]) ? 1 : 0;
assign detect_max[587][19] = (mid_1[4711:4704] > btm_0[4719:4712]) ? 1 : 0;
assign detect_max[587][20] = (mid_1[4711:4704] > btm_1[4703:4696]) ? 1 : 0;
assign detect_max[587][21] = (mid_1[4711:4704] > btm_1[4711:4704]) ? 1 : 0;
assign detect_max[587][22] = (mid_1[4711:4704] > btm_1[4719:4712]) ? 1 : 0;
assign detect_max[587][23] = (mid_1[4711:4704] > btm_2[4703:4696]) ? 1 : 0;
assign detect_max[587][24] = (mid_1[4711:4704] > btm_2[4711:4704]) ? 1 : 0;
assign detect_max[587][25] = (mid_1[4711:4704] > btm_2[4719:4712]) ? 1 : 0;

assign detect_max[588][0] = (mid_1[4719:4712] > top_0[4711:4704]) ? 1 : 0;
assign detect_max[588][1] = (mid_1[4719:4712] > top_0[4719:4712]) ? 1 : 0;
assign detect_max[588][2] = (mid_1[4719:4712] > top_0[4727:4720]) ? 1 : 0;
assign detect_max[588][3] = (mid_1[4719:4712] > top_1[4711:4704]) ? 1 : 0;
assign detect_max[588][4] = (mid_1[4719:4712] > top_1[4719:4712]) ? 1 : 0;
assign detect_max[588][5] = (mid_1[4719:4712] > top_1[4727:4720]) ? 1 : 0;
assign detect_max[588][6] = (mid_1[4719:4712] > top_2[4711:4704]) ? 1 : 0;
assign detect_max[588][7] = (mid_1[4719:4712] > top_2[4719:4712]) ? 1 : 0;
assign detect_max[588][8] = (mid_1[4719:4712] > top_2[4727:4720]) ? 1 : 0;
assign detect_max[588][9] = (mid_1[4719:4712] > mid_0[4711:4704]) ? 1 : 0;
assign detect_max[588][10] = (mid_1[4719:4712] > mid_0[4719:4712]) ? 1 : 0;
assign detect_max[588][11] = (mid_1[4719:4712] > mid_0[4727:4720]) ? 1 : 0;
assign detect_max[588][12] = (mid_1[4719:4712] > mid_1[4711:4704]) ? 1 : 0;
assign detect_max[588][13] = (mid_1[4719:4712] > mid_1[4727:4720]) ? 1 : 0;
assign detect_max[588][14] = (mid_1[4719:4712] > mid_2[4711:4704]) ? 1 : 0;
assign detect_max[588][15] = (mid_1[4719:4712] > mid_2[4719:4712]) ? 1 : 0;
assign detect_max[588][16] = (mid_1[4719:4712] > mid_2[4727:4720]) ? 1 : 0;
assign detect_max[588][17] = (mid_1[4719:4712] > btm_0[4711:4704]) ? 1 : 0;
assign detect_max[588][18] = (mid_1[4719:4712] > btm_0[4719:4712]) ? 1 : 0;
assign detect_max[588][19] = (mid_1[4719:4712] > btm_0[4727:4720]) ? 1 : 0;
assign detect_max[588][20] = (mid_1[4719:4712] > btm_1[4711:4704]) ? 1 : 0;
assign detect_max[588][21] = (mid_1[4719:4712] > btm_1[4719:4712]) ? 1 : 0;
assign detect_max[588][22] = (mid_1[4719:4712] > btm_1[4727:4720]) ? 1 : 0;
assign detect_max[588][23] = (mid_1[4719:4712] > btm_2[4711:4704]) ? 1 : 0;
assign detect_max[588][24] = (mid_1[4719:4712] > btm_2[4719:4712]) ? 1 : 0;
assign detect_max[588][25] = (mid_1[4719:4712] > btm_2[4727:4720]) ? 1 : 0;

assign detect_max[589][0] = (mid_1[4727:4720] > top_0[4719:4712]) ? 1 : 0;
assign detect_max[589][1] = (mid_1[4727:4720] > top_0[4727:4720]) ? 1 : 0;
assign detect_max[589][2] = (mid_1[4727:4720] > top_0[4735:4728]) ? 1 : 0;
assign detect_max[589][3] = (mid_1[4727:4720] > top_1[4719:4712]) ? 1 : 0;
assign detect_max[589][4] = (mid_1[4727:4720] > top_1[4727:4720]) ? 1 : 0;
assign detect_max[589][5] = (mid_1[4727:4720] > top_1[4735:4728]) ? 1 : 0;
assign detect_max[589][6] = (mid_1[4727:4720] > top_2[4719:4712]) ? 1 : 0;
assign detect_max[589][7] = (mid_1[4727:4720] > top_2[4727:4720]) ? 1 : 0;
assign detect_max[589][8] = (mid_1[4727:4720] > top_2[4735:4728]) ? 1 : 0;
assign detect_max[589][9] = (mid_1[4727:4720] > mid_0[4719:4712]) ? 1 : 0;
assign detect_max[589][10] = (mid_1[4727:4720] > mid_0[4727:4720]) ? 1 : 0;
assign detect_max[589][11] = (mid_1[4727:4720] > mid_0[4735:4728]) ? 1 : 0;
assign detect_max[589][12] = (mid_1[4727:4720] > mid_1[4719:4712]) ? 1 : 0;
assign detect_max[589][13] = (mid_1[4727:4720] > mid_1[4735:4728]) ? 1 : 0;
assign detect_max[589][14] = (mid_1[4727:4720] > mid_2[4719:4712]) ? 1 : 0;
assign detect_max[589][15] = (mid_1[4727:4720] > mid_2[4727:4720]) ? 1 : 0;
assign detect_max[589][16] = (mid_1[4727:4720] > mid_2[4735:4728]) ? 1 : 0;
assign detect_max[589][17] = (mid_1[4727:4720] > btm_0[4719:4712]) ? 1 : 0;
assign detect_max[589][18] = (mid_1[4727:4720] > btm_0[4727:4720]) ? 1 : 0;
assign detect_max[589][19] = (mid_1[4727:4720] > btm_0[4735:4728]) ? 1 : 0;
assign detect_max[589][20] = (mid_1[4727:4720] > btm_1[4719:4712]) ? 1 : 0;
assign detect_max[589][21] = (mid_1[4727:4720] > btm_1[4727:4720]) ? 1 : 0;
assign detect_max[589][22] = (mid_1[4727:4720] > btm_1[4735:4728]) ? 1 : 0;
assign detect_max[589][23] = (mid_1[4727:4720] > btm_2[4719:4712]) ? 1 : 0;
assign detect_max[589][24] = (mid_1[4727:4720] > btm_2[4727:4720]) ? 1 : 0;
assign detect_max[589][25] = (mid_1[4727:4720] > btm_2[4735:4728]) ? 1 : 0;

assign detect_max[590][0] = (mid_1[4735:4728] > top_0[4727:4720]) ? 1 : 0;
assign detect_max[590][1] = (mid_1[4735:4728] > top_0[4735:4728]) ? 1 : 0;
assign detect_max[590][2] = (mid_1[4735:4728] > top_0[4743:4736]) ? 1 : 0;
assign detect_max[590][3] = (mid_1[4735:4728] > top_1[4727:4720]) ? 1 : 0;
assign detect_max[590][4] = (mid_1[4735:4728] > top_1[4735:4728]) ? 1 : 0;
assign detect_max[590][5] = (mid_1[4735:4728] > top_1[4743:4736]) ? 1 : 0;
assign detect_max[590][6] = (mid_1[4735:4728] > top_2[4727:4720]) ? 1 : 0;
assign detect_max[590][7] = (mid_1[4735:4728] > top_2[4735:4728]) ? 1 : 0;
assign detect_max[590][8] = (mid_1[4735:4728] > top_2[4743:4736]) ? 1 : 0;
assign detect_max[590][9] = (mid_1[4735:4728] > mid_0[4727:4720]) ? 1 : 0;
assign detect_max[590][10] = (mid_1[4735:4728] > mid_0[4735:4728]) ? 1 : 0;
assign detect_max[590][11] = (mid_1[4735:4728] > mid_0[4743:4736]) ? 1 : 0;
assign detect_max[590][12] = (mid_1[4735:4728] > mid_1[4727:4720]) ? 1 : 0;
assign detect_max[590][13] = (mid_1[4735:4728] > mid_1[4743:4736]) ? 1 : 0;
assign detect_max[590][14] = (mid_1[4735:4728] > mid_2[4727:4720]) ? 1 : 0;
assign detect_max[590][15] = (mid_1[4735:4728] > mid_2[4735:4728]) ? 1 : 0;
assign detect_max[590][16] = (mid_1[4735:4728] > mid_2[4743:4736]) ? 1 : 0;
assign detect_max[590][17] = (mid_1[4735:4728] > btm_0[4727:4720]) ? 1 : 0;
assign detect_max[590][18] = (mid_1[4735:4728] > btm_0[4735:4728]) ? 1 : 0;
assign detect_max[590][19] = (mid_1[4735:4728] > btm_0[4743:4736]) ? 1 : 0;
assign detect_max[590][20] = (mid_1[4735:4728] > btm_1[4727:4720]) ? 1 : 0;
assign detect_max[590][21] = (mid_1[4735:4728] > btm_1[4735:4728]) ? 1 : 0;
assign detect_max[590][22] = (mid_1[4735:4728] > btm_1[4743:4736]) ? 1 : 0;
assign detect_max[590][23] = (mid_1[4735:4728] > btm_2[4727:4720]) ? 1 : 0;
assign detect_max[590][24] = (mid_1[4735:4728] > btm_2[4735:4728]) ? 1 : 0;
assign detect_max[590][25] = (mid_1[4735:4728] > btm_2[4743:4736]) ? 1 : 0;

assign detect_max[591][0] = (mid_1[4743:4736] > top_0[4735:4728]) ? 1 : 0;
assign detect_max[591][1] = (mid_1[4743:4736] > top_0[4743:4736]) ? 1 : 0;
assign detect_max[591][2] = (mid_1[4743:4736] > top_0[4751:4744]) ? 1 : 0;
assign detect_max[591][3] = (mid_1[4743:4736] > top_1[4735:4728]) ? 1 : 0;
assign detect_max[591][4] = (mid_1[4743:4736] > top_1[4743:4736]) ? 1 : 0;
assign detect_max[591][5] = (mid_1[4743:4736] > top_1[4751:4744]) ? 1 : 0;
assign detect_max[591][6] = (mid_1[4743:4736] > top_2[4735:4728]) ? 1 : 0;
assign detect_max[591][7] = (mid_1[4743:4736] > top_2[4743:4736]) ? 1 : 0;
assign detect_max[591][8] = (mid_1[4743:4736] > top_2[4751:4744]) ? 1 : 0;
assign detect_max[591][9] = (mid_1[4743:4736] > mid_0[4735:4728]) ? 1 : 0;
assign detect_max[591][10] = (mid_1[4743:4736] > mid_0[4743:4736]) ? 1 : 0;
assign detect_max[591][11] = (mid_1[4743:4736] > mid_0[4751:4744]) ? 1 : 0;
assign detect_max[591][12] = (mid_1[4743:4736] > mid_1[4735:4728]) ? 1 : 0;
assign detect_max[591][13] = (mid_1[4743:4736] > mid_1[4751:4744]) ? 1 : 0;
assign detect_max[591][14] = (mid_1[4743:4736] > mid_2[4735:4728]) ? 1 : 0;
assign detect_max[591][15] = (mid_1[4743:4736] > mid_2[4743:4736]) ? 1 : 0;
assign detect_max[591][16] = (mid_1[4743:4736] > mid_2[4751:4744]) ? 1 : 0;
assign detect_max[591][17] = (mid_1[4743:4736] > btm_0[4735:4728]) ? 1 : 0;
assign detect_max[591][18] = (mid_1[4743:4736] > btm_0[4743:4736]) ? 1 : 0;
assign detect_max[591][19] = (mid_1[4743:4736] > btm_0[4751:4744]) ? 1 : 0;
assign detect_max[591][20] = (mid_1[4743:4736] > btm_1[4735:4728]) ? 1 : 0;
assign detect_max[591][21] = (mid_1[4743:4736] > btm_1[4743:4736]) ? 1 : 0;
assign detect_max[591][22] = (mid_1[4743:4736] > btm_1[4751:4744]) ? 1 : 0;
assign detect_max[591][23] = (mid_1[4743:4736] > btm_2[4735:4728]) ? 1 : 0;
assign detect_max[591][24] = (mid_1[4743:4736] > btm_2[4743:4736]) ? 1 : 0;
assign detect_max[591][25] = (mid_1[4743:4736] > btm_2[4751:4744]) ? 1 : 0;

assign detect_max[592][0] = (mid_1[4751:4744] > top_0[4743:4736]) ? 1 : 0;
assign detect_max[592][1] = (mid_1[4751:4744] > top_0[4751:4744]) ? 1 : 0;
assign detect_max[592][2] = (mid_1[4751:4744] > top_0[4759:4752]) ? 1 : 0;
assign detect_max[592][3] = (mid_1[4751:4744] > top_1[4743:4736]) ? 1 : 0;
assign detect_max[592][4] = (mid_1[4751:4744] > top_1[4751:4744]) ? 1 : 0;
assign detect_max[592][5] = (mid_1[4751:4744] > top_1[4759:4752]) ? 1 : 0;
assign detect_max[592][6] = (mid_1[4751:4744] > top_2[4743:4736]) ? 1 : 0;
assign detect_max[592][7] = (mid_1[4751:4744] > top_2[4751:4744]) ? 1 : 0;
assign detect_max[592][8] = (mid_1[4751:4744] > top_2[4759:4752]) ? 1 : 0;
assign detect_max[592][9] = (mid_1[4751:4744] > mid_0[4743:4736]) ? 1 : 0;
assign detect_max[592][10] = (mid_1[4751:4744] > mid_0[4751:4744]) ? 1 : 0;
assign detect_max[592][11] = (mid_1[4751:4744] > mid_0[4759:4752]) ? 1 : 0;
assign detect_max[592][12] = (mid_1[4751:4744] > mid_1[4743:4736]) ? 1 : 0;
assign detect_max[592][13] = (mid_1[4751:4744] > mid_1[4759:4752]) ? 1 : 0;
assign detect_max[592][14] = (mid_1[4751:4744] > mid_2[4743:4736]) ? 1 : 0;
assign detect_max[592][15] = (mid_1[4751:4744] > mid_2[4751:4744]) ? 1 : 0;
assign detect_max[592][16] = (mid_1[4751:4744] > mid_2[4759:4752]) ? 1 : 0;
assign detect_max[592][17] = (mid_1[4751:4744] > btm_0[4743:4736]) ? 1 : 0;
assign detect_max[592][18] = (mid_1[4751:4744] > btm_0[4751:4744]) ? 1 : 0;
assign detect_max[592][19] = (mid_1[4751:4744] > btm_0[4759:4752]) ? 1 : 0;
assign detect_max[592][20] = (mid_1[4751:4744] > btm_1[4743:4736]) ? 1 : 0;
assign detect_max[592][21] = (mid_1[4751:4744] > btm_1[4751:4744]) ? 1 : 0;
assign detect_max[592][22] = (mid_1[4751:4744] > btm_1[4759:4752]) ? 1 : 0;
assign detect_max[592][23] = (mid_1[4751:4744] > btm_2[4743:4736]) ? 1 : 0;
assign detect_max[592][24] = (mid_1[4751:4744] > btm_2[4751:4744]) ? 1 : 0;
assign detect_max[592][25] = (mid_1[4751:4744] > btm_2[4759:4752]) ? 1 : 0;

assign detect_max[593][0] = (mid_1[4759:4752] > top_0[4751:4744]) ? 1 : 0;
assign detect_max[593][1] = (mid_1[4759:4752] > top_0[4759:4752]) ? 1 : 0;
assign detect_max[593][2] = (mid_1[4759:4752] > top_0[4767:4760]) ? 1 : 0;
assign detect_max[593][3] = (mid_1[4759:4752] > top_1[4751:4744]) ? 1 : 0;
assign detect_max[593][4] = (mid_1[4759:4752] > top_1[4759:4752]) ? 1 : 0;
assign detect_max[593][5] = (mid_1[4759:4752] > top_1[4767:4760]) ? 1 : 0;
assign detect_max[593][6] = (mid_1[4759:4752] > top_2[4751:4744]) ? 1 : 0;
assign detect_max[593][7] = (mid_1[4759:4752] > top_2[4759:4752]) ? 1 : 0;
assign detect_max[593][8] = (mid_1[4759:4752] > top_2[4767:4760]) ? 1 : 0;
assign detect_max[593][9] = (mid_1[4759:4752] > mid_0[4751:4744]) ? 1 : 0;
assign detect_max[593][10] = (mid_1[4759:4752] > mid_0[4759:4752]) ? 1 : 0;
assign detect_max[593][11] = (mid_1[4759:4752] > mid_0[4767:4760]) ? 1 : 0;
assign detect_max[593][12] = (mid_1[4759:4752] > mid_1[4751:4744]) ? 1 : 0;
assign detect_max[593][13] = (mid_1[4759:4752] > mid_1[4767:4760]) ? 1 : 0;
assign detect_max[593][14] = (mid_1[4759:4752] > mid_2[4751:4744]) ? 1 : 0;
assign detect_max[593][15] = (mid_1[4759:4752] > mid_2[4759:4752]) ? 1 : 0;
assign detect_max[593][16] = (mid_1[4759:4752] > mid_2[4767:4760]) ? 1 : 0;
assign detect_max[593][17] = (mid_1[4759:4752] > btm_0[4751:4744]) ? 1 : 0;
assign detect_max[593][18] = (mid_1[4759:4752] > btm_0[4759:4752]) ? 1 : 0;
assign detect_max[593][19] = (mid_1[4759:4752] > btm_0[4767:4760]) ? 1 : 0;
assign detect_max[593][20] = (mid_1[4759:4752] > btm_1[4751:4744]) ? 1 : 0;
assign detect_max[593][21] = (mid_1[4759:4752] > btm_1[4759:4752]) ? 1 : 0;
assign detect_max[593][22] = (mid_1[4759:4752] > btm_1[4767:4760]) ? 1 : 0;
assign detect_max[593][23] = (mid_1[4759:4752] > btm_2[4751:4744]) ? 1 : 0;
assign detect_max[593][24] = (mid_1[4759:4752] > btm_2[4759:4752]) ? 1 : 0;
assign detect_max[593][25] = (mid_1[4759:4752] > btm_2[4767:4760]) ? 1 : 0;

assign detect_max[594][0] = (mid_1[4767:4760] > top_0[4759:4752]) ? 1 : 0;
assign detect_max[594][1] = (mid_1[4767:4760] > top_0[4767:4760]) ? 1 : 0;
assign detect_max[594][2] = (mid_1[4767:4760] > top_0[4775:4768]) ? 1 : 0;
assign detect_max[594][3] = (mid_1[4767:4760] > top_1[4759:4752]) ? 1 : 0;
assign detect_max[594][4] = (mid_1[4767:4760] > top_1[4767:4760]) ? 1 : 0;
assign detect_max[594][5] = (mid_1[4767:4760] > top_1[4775:4768]) ? 1 : 0;
assign detect_max[594][6] = (mid_1[4767:4760] > top_2[4759:4752]) ? 1 : 0;
assign detect_max[594][7] = (mid_1[4767:4760] > top_2[4767:4760]) ? 1 : 0;
assign detect_max[594][8] = (mid_1[4767:4760] > top_2[4775:4768]) ? 1 : 0;
assign detect_max[594][9] = (mid_1[4767:4760] > mid_0[4759:4752]) ? 1 : 0;
assign detect_max[594][10] = (mid_1[4767:4760] > mid_0[4767:4760]) ? 1 : 0;
assign detect_max[594][11] = (mid_1[4767:4760] > mid_0[4775:4768]) ? 1 : 0;
assign detect_max[594][12] = (mid_1[4767:4760] > mid_1[4759:4752]) ? 1 : 0;
assign detect_max[594][13] = (mid_1[4767:4760] > mid_1[4775:4768]) ? 1 : 0;
assign detect_max[594][14] = (mid_1[4767:4760] > mid_2[4759:4752]) ? 1 : 0;
assign detect_max[594][15] = (mid_1[4767:4760] > mid_2[4767:4760]) ? 1 : 0;
assign detect_max[594][16] = (mid_1[4767:4760] > mid_2[4775:4768]) ? 1 : 0;
assign detect_max[594][17] = (mid_1[4767:4760] > btm_0[4759:4752]) ? 1 : 0;
assign detect_max[594][18] = (mid_1[4767:4760] > btm_0[4767:4760]) ? 1 : 0;
assign detect_max[594][19] = (mid_1[4767:4760] > btm_0[4775:4768]) ? 1 : 0;
assign detect_max[594][20] = (mid_1[4767:4760] > btm_1[4759:4752]) ? 1 : 0;
assign detect_max[594][21] = (mid_1[4767:4760] > btm_1[4767:4760]) ? 1 : 0;
assign detect_max[594][22] = (mid_1[4767:4760] > btm_1[4775:4768]) ? 1 : 0;
assign detect_max[594][23] = (mid_1[4767:4760] > btm_2[4759:4752]) ? 1 : 0;
assign detect_max[594][24] = (mid_1[4767:4760] > btm_2[4767:4760]) ? 1 : 0;
assign detect_max[594][25] = (mid_1[4767:4760] > btm_2[4775:4768]) ? 1 : 0;

assign detect_max[595][0] = (mid_1[4775:4768] > top_0[4767:4760]) ? 1 : 0;
assign detect_max[595][1] = (mid_1[4775:4768] > top_0[4775:4768]) ? 1 : 0;
assign detect_max[595][2] = (mid_1[4775:4768] > top_0[4783:4776]) ? 1 : 0;
assign detect_max[595][3] = (mid_1[4775:4768] > top_1[4767:4760]) ? 1 : 0;
assign detect_max[595][4] = (mid_1[4775:4768] > top_1[4775:4768]) ? 1 : 0;
assign detect_max[595][5] = (mid_1[4775:4768] > top_1[4783:4776]) ? 1 : 0;
assign detect_max[595][6] = (mid_1[4775:4768] > top_2[4767:4760]) ? 1 : 0;
assign detect_max[595][7] = (mid_1[4775:4768] > top_2[4775:4768]) ? 1 : 0;
assign detect_max[595][8] = (mid_1[4775:4768] > top_2[4783:4776]) ? 1 : 0;
assign detect_max[595][9] = (mid_1[4775:4768] > mid_0[4767:4760]) ? 1 : 0;
assign detect_max[595][10] = (mid_1[4775:4768] > mid_0[4775:4768]) ? 1 : 0;
assign detect_max[595][11] = (mid_1[4775:4768] > mid_0[4783:4776]) ? 1 : 0;
assign detect_max[595][12] = (mid_1[4775:4768] > mid_1[4767:4760]) ? 1 : 0;
assign detect_max[595][13] = (mid_1[4775:4768] > mid_1[4783:4776]) ? 1 : 0;
assign detect_max[595][14] = (mid_1[4775:4768] > mid_2[4767:4760]) ? 1 : 0;
assign detect_max[595][15] = (mid_1[4775:4768] > mid_2[4775:4768]) ? 1 : 0;
assign detect_max[595][16] = (mid_1[4775:4768] > mid_2[4783:4776]) ? 1 : 0;
assign detect_max[595][17] = (mid_1[4775:4768] > btm_0[4767:4760]) ? 1 : 0;
assign detect_max[595][18] = (mid_1[4775:4768] > btm_0[4775:4768]) ? 1 : 0;
assign detect_max[595][19] = (mid_1[4775:4768] > btm_0[4783:4776]) ? 1 : 0;
assign detect_max[595][20] = (mid_1[4775:4768] > btm_1[4767:4760]) ? 1 : 0;
assign detect_max[595][21] = (mid_1[4775:4768] > btm_1[4775:4768]) ? 1 : 0;
assign detect_max[595][22] = (mid_1[4775:4768] > btm_1[4783:4776]) ? 1 : 0;
assign detect_max[595][23] = (mid_1[4775:4768] > btm_2[4767:4760]) ? 1 : 0;
assign detect_max[595][24] = (mid_1[4775:4768] > btm_2[4775:4768]) ? 1 : 0;
assign detect_max[595][25] = (mid_1[4775:4768] > btm_2[4783:4776]) ? 1 : 0;

assign detect_max[596][0] = (mid_1[4783:4776] > top_0[4775:4768]) ? 1 : 0;
assign detect_max[596][1] = (mid_1[4783:4776] > top_0[4783:4776]) ? 1 : 0;
assign detect_max[596][2] = (mid_1[4783:4776] > top_0[4791:4784]) ? 1 : 0;
assign detect_max[596][3] = (mid_1[4783:4776] > top_1[4775:4768]) ? 1 : 0;
assign detect_max[596][4] = (mid_1[4783:4776] > top_1[4783:4776]) ? 1 : 0;
assign detect_max[596][5] = (mid_1[4783:4776] > top_1[4791:4784]) ? 1 : 0;
assign detect_max[596][6] = (mid_1[4783:4776] > top_2[4775:4768]) ? 1 : 0;
assign detect_max[596][7] = (mid_1[4783:4776] > top_2[4783:4776]) ? 1 : 0;
assign detect_max[596][8] = (mid_1[4783:4776] > top_2[4791:4784]) ? 1 : 0;
assign detect_max[596][9] = (mid_1[4783:4776] > mid_0[4775:4768]) ? 1 : 0;
assign detect_max[596][10] = (mid_1[4783:4776] > mid_0[4783:4776]) ? 1 : 0;
assign detect_max[596][11] = (mid_1[4783:4776] > mid_0[4791:4784]) ? 1 : 0;
assign detect_max[596][12] = (mid_1[4783:4776] > mid_1[4775:4768]) ? 1 : 0;
assign detect_max[596][13] = (mid_1[4783:4776] > mid_1[4791:4784]) ? 1 : 0;
assign detect_max[596][14] = (mid_1[4783:4776] > mid_2[4775:4768]) ? 1 : 0;
assign detect_max[596][15] = (mid_1[4783:4776] > mid_2[4783:4776]) ? 1 : 0;
assign detect_max[596][16] = (mid_1[4783:4776] > mid_2[4791:4784]) ? 1 : 0;
assign detect_max[596][17] = (mid_1[4783:4776] > btm_0[4775:4768]) ? 1 : 0;
assign detect_max[596][18] = (mid_1[4783:4776] > btm_0[4783:4776]) ? 1 : 0;
assign detect_max[596][19] = (mid_1[4783:4776] > btm_0[4791:4784]) ? 1 : 0;
assign detect_max[596][20] = (mid_1[4783:4776] > btm_1[4775:4768]) ? 1 : 0;
assign detect_max[596][21] = (mid_1[4783:4776] > btm_1[4783:4776]) ? 1 : 0;
assign detect_max[596][22] = (mid_1[4783:4776] > btm_1[4791:4784]) ? 1 : 0;
assign detect_max[596][23] = (mid_1[4783:4776] > btm_2[4775:4768]) ? 1 : 0;
assign detect_max[596][24] = (mid_1[4783:4776] > btm_2[4783:4776]) ? 1 : 0;
assign detect_max[596][25] = (mid_1[4783:4776] > btm_2[4791:4784]) ? 1 : 0;

assign detect_max[597][0] = (mid_1[4791:4784] > top_0[4783:4776]) ? 1 : 0;
assign detect_max[597][1] = (mid_1[4791:4784] > top_0[4791:4784]) ? 1 : 0;
assign detect_max[597][2] = (mid_1[4791:4784] > top_0[4799:4792]) ? 1 : 0;
assign detect_max[597][3] = (mid_1[4791:4784] > top_1[4783:4776]) ? 1 : 0;
assign detect_max[597][4] = (mid_1[4791:4784] > top_1[4791:4784]) ? 1 : 0;
assign detect_max[597][5] = (mid_1[4791:4784] > top_1[4799:4792]) ? 1 : 0;
assign detect_max[597][6] = (mid_1[4791:4784] > top_2[4783:4776]) ? 1 : 0;
assign detect_max[597][7] = (mid_1[4791:4784] > top_2[4791:4784]) ? 1 : 0;
assign detect_max[597][8] = (mid_1[4791:4784] > top_2[4799:4792]) ? 1 : 0;
assign detect_max[597][9] = (mid_1[4791:4784] > mid_0[4783:4776]) ? 1 : 0;
assign detect_max[597][10] = (mid_1[4791:4784] > mid_0[4791:4784]) ? 1 : 0;
assign detect_max[597][11] = (mid_1[4791:4784] > mid_0[4799:4792]) ? 1 : 0;
assign detect_max[597][12] = (mid_1[4791:4784] > mid_1[4783:4776]) ? 1 : 0;
assign detect_max[597][13] = (mid_1[4791:4784] > mid_1[4799:4792]) ? 1 : 0;
assign detect_max[597][14] = (mid_1[4791:4784] > mid_2[4783:4776]) ? 1 : 0;
assign detect_max[597][15] = (mid_1[4791:4784] > mid_2[4791:4784]) ? 1 : 0;
assign detect_max[597][16] = (mid_1[4791:4784] > mid_2[4799:4792]) ? 1 : 0;
assign detect_max[597][17] = (mid_1[4791:4784] > btm_0[4783:4776]) ? 1 : 0;
assign detect_max[597][18] = (mid_1[4791:4784] > btm_0[4791:4784]) ? 1 : 0;
assign detect_max[597][19] = (mid_1[4791:4784] > btm_0[4799:4792]) ? 1 : 0;
assign detect_max[597][20] = (mid_1[4791:4784] > btm_1[4783:4776]) ? 1 : 0;
assign detect_max[597][21] = (mid_1[4791:4784] > btm_1[4791:4784]) ? 1 : 0;
assign detect_max[597][22] = (mid_1[4791:4784] > btm_1[4799:4792]) ? 1 : 0;
assign detect_max[597][23] = (mid_1[4791:4784] > btm_2[4783:4776]) ? 1 : 0;
assign detect_max[597][24] = (mid_1[4791:4784] > btm_2[4791:4784]) ? 1 : 0;
assign detect_max[597][25] = (mid_1[4791:4784] > btm_2[4799:4792]) ? 1 : 0;

assign detect_max[598][0] = (mid_1[4799:4792] > top_0[4791:4784]) ? 1 : 0;
assign detect_max[598][1] = (mid_1[4799:4792] > top_0[4799:4792]) ? 1 : 0;
assign detect_max[598][2] = (mid_1[4799:4792] > top_0[4807:4800]) ? 1 : 0;
assign detect_max[598][3] = (mid_1[4799:4792] > top_1[4791:4784]) ? 1 : 0;
assign detect_max[598][4] = (mid_1[4799:4792] > top_1[4799:4792]) ? 1 : 0;
assign detect_max[598][5] = (mid_1[4799:4792] > top_1[4807:4800]) ? 1 : 0;
assign detect_max[598][6] = (mid_1[4799:4792] > top_2[4791:4784]) ? 1 : 0;
assign detect_max[598][7] = (mid_1[4799:4792] > top_2[4799:4792]) ? 1 : 0;
assign detect_max[598][8] = (mid_1[4799:4792] > top_2[4807:4800]) ? 1 : 0;
assign detect_max[598][9] = (mid_1[4799:4792] > mid_0[4791:4784]) ? 1 : 0;
assign detect_max[598][10] = (mid_1[4799:4792] > mid_0[4799:4792]) ? 1 : 0;
assign detect_max[598][11] = (mid_1[4799:4792] > mid_0[4807:4800]) ? 1 : 0;
assign detect_max[598][12] = (mid_1[4799:4792] > mid_1[4791:4784]) ? 1 : 0;
assign detect_max[598][13] = (mid_1[4799:4792] > mid_1[4807:4800]) ? 1 : 0;
assign detect_max[598][14] = (mid_1[4799:4792] > mid_2[4791:4784]) ? 1 : 0;
assign detect_max[598][15] = (mid_1[4799:4792] > mid_2[4799:4792]) ? 1 : 0;
assign detect_max[598][16] = (mid_1[4799:4792] > mid_2[4807:4800]) ? 1 : 0;
assign detect_max[598][17] = (mid_1[4799:4792] > btm_0[4791:4784]) ? 1 : 0;
assign detect_max[598][18] = (mid_1[4799:4792] > btm_0[4799:4792]) ? 1 : 0;
assign detect_max[598][19] = (mid_1[4799:4792] > btm_0[4807:4800]) ? 1 : 0;
assign detect_max[598][20] = (mid_1[4799:4792] > btm_1[4791:4784]) ? 1 : 0;
assign detect_max[598][21] = (mid_1[4799:4792] > btm_1[4799:4792]) ? 1 : 0;
assign detect_max[598][22] = (mid_1[4799:4792] > btm_1[4807:4800]) ? 1 : 0;
assign detect_max[598][23] = (mid_1[4799:4792] > btm_2[4791:4784]) ? 1 : 0;
assign detect_max[598][24] = (mid_1[4799:4792] > btm_2[4799:4792]) ? 1 : 0;
assign detect_max[598][25] = (mid_1[4799:4792] > btm_2[4807:4800]) ? 1 : 0;

assign detect_max[599][0] = (mid_1[4807:4800] > top_0[4799:4792]) ? 1 : 0;
assign detect_max[599][1] = (mid_1[4807:4800] > top_0[4807:4800]) ? 1 : 0;
assign detect_max[599][2] = (mid_1[4807:4800] > top_0[4815:4808]) ? 1 : 0;
assign detect_max[599][3] = (mid_1[4807:4800] > top_1[4799:4792]) ? 1 : 0;
assign detect_max[599][4] = (mid_1[4807:4800] > top_1[4807:4800]) ? 1 : 0;
assign detect_max[599][5] = (mid_1[4807:4800] > top_1[4815:4808]) ? 1 : 0;
assign detect_max[599][6] = (mid_1[4807:4800] > top_2[4799:4792]) ? 1 : 0;
assign detect_max[599][7] = (mid_1[4807:4800] > top_2[4807:4800]) ? 1 : 0;
assign detect_max[599][8] = (mid_1[4807:4800] > top_2[4815:4808]) ? 1 : 0;
assign detect_max[599][9] = (mid_1[4807:4800] > mid_0[4799:4792]) ? 1 : 0;
assign detect_max[599][10] = (mid_1[4807:4800] > mid_0[4807:4800]) ? 1 : 0;
assign detect_max[599][11] = (mid_1[4807:4800] > mid_0[4815:4808]) ? 1 : 0;
assign detect_max[599][12] = (mid_1[4807:4800] > mid_1[4799:4792]) ? 1 : 0;
assign detect_max[599][13] = (mid_1[4807:4800] > mid_1[4815:4808]) ? 1 : 0;
assign detect_max[599][14] = (mid_1[4807:4800] > mid_2[4799:4792]) ? 1 : 0;
assign detect_max[599][15] = (mid_1[4807:4800] > mid_2[4807:4800]) ? 1 : 0;
assign detect_max[599][16] = (mid_1[4807:4800] > mid_2[4815:4808]) ? 1 : 0;
assign detect_max[599][17] = (mid_1[4807:4800] > btm_0[4799:4792]) ? 1 : 0;
assign detect_max[599][18] = (mid_1[4807:4800] > btm_0[4807:4800]) ? 1 : 0;
assign detect_max[599][19] = (mid_1[4807:4800] > btm_0[4815:4808]) ? 1 : 0;
assign detect_max[599][20] = (mid_1[4807:4800] > btm_1[4799:4792]) ? 1 : 0;
assign detect_max[599][21] = (mid_1[4807:4800] > btm_1[4807:4800]) ? 1 : 0;
assign detect_max[599][22] = (mid_1[4807:4800] > btm_1[4815:4808]) ? 1 : 0;
assign detect_max[599][23] = (mid_1[4807:4800] > btm_2[4799:4792]) ? 1 : 0;
assign detect_max[599][24] = (mid_1[4807:4800] > btm_2[4807:4800]) ? 1 : 0;
assign detect_max[599][25] = (mid_1[4807:4800] > btm_2[4815:4808]) ? 1 : 0;

assign detect_max[600][0] = (mid_1[4815:4808] > top_0[4807:4800]) ? 1 : 0;
assign detect_max[600][1] = (mid_1[4815:4808] > top_0[4815:4808]) ? 1 : 0;
assign detect_max[600][2] = (mid_1[4815:4808] > top_0[4823:4816]) ? 1 : 0;
assign detect_max[600][3] = (mid_1[4815:4808] > top_1[4807:4800]) ? 1 : 0;
assign detect_max[600][4] = (mid_1[4815:4808] > top_1[4815:4808]) ? 1 : 0;
assign detect_max[600][5] = (mid_1[4815:4808] > top_1[4823:4816]) ? 1 : 0;
assign detect_max[600][6] = (mid_1[4815:4808] > top_2[4807:4800]) ? 1 : 0;
assign detect_max[600][7] = (mid_1[4815:4808] > top_2[4815:4808]) ? 1 : 0;
assign detect_max[600][8] = (mid_1[4815:4808] > top_2[4823:4816]) ? 1 : 0;
assign detect_max[600][9] = (mid_1[4815:4808] > mid_0[4807:4800]) ? 1 : 0;
assign detect_max[600][10] = (mid_1[4815:4808] > mid_0[4815:4808]) ? 1 : 0;
assign detect_max[600][11] = (mid_1[4815:4808] > mid_0[4823:4816]) ? 1 : 0;
assign detect_max[600][12] = (mid_1[4815:4808] > mid_1[4807:4800]) ? 1 : 0;
assign detect_max[600][13] = (mid_1[4815:4808] > mid_1[4823:4816]) ? 1 : 0;
assign detect_max[600][14] = (mid_1[4815:4808] > mid_2[4807:4800]) ? 1 : 0;
assign detect_max[600][15] = (mid_1[4815:4808] > mid_2[4815:4808]) ? 1 : 0;
assign detect_max[600][16] = (mid_1[4815:4808] > mid_2[4823:4816]) ? 1 : 0;
assign detect_max[600][17] = (mid_1[4815:4808] > btm_0[4807:4800]) ? 1 : 0;
assign detect_max[600][18] = (mid_1[4815:4808] > btm_0[4815:4808]) ? 1 : 0;
assign detect_max[600][19] = (mid_1[4815:4808] > btm_0[4823:4816]) ? 1 : 0;
assign detect_max[600][20] = (mid_1[4815:4808] > btm_1[4807:4800]) ? 1 : 0;
assign detect_max[600][21] = (mid_1[4815:4808] > btm_1[4815:4808]) ? 1 : 0;
assign detect_max[600][22] = (mid_1[4815:4808] > btm_1[4823:4816]) ? 1 : 0;
assign detect_max[600][23] = (mid_1[4815:4808] > btm_2[4807:4800]) ? 1 : 0;
assign detect_max[600][24] = (mid_1[4815:4808] > btm_2[4815:4808]) ? 1 : 0;
assign detect_max[600][25] = (mid_1[4815:4808] > btm_2[4823:4816]) ? 1 : 0;

assign detect_max[601][0] = (mid_1[4823:4816] > top_0[4815:4808]) ? 1 : 0;
assign detect_max[601][1] = (mid_1[4823:4816] > top_0[4823:4816]) ? 1 : 0;
assign detect_max[601][2] = (mid_1[4823:4816] > top_0[4831:4824]) ? 1 : 0;
assign detect_max[601][3] = (mid_1[4823:4816] > top_1[4815:4808]) ? 1 : 0;
assign detect_max[601][4] = (mid_1[4823:4816] > top_1[4823:4816]) ? 1 : 0;
assign detect_max[601][5] = (mid_1[4823:4816] > top_1[4831:4824]) ? 1 : 0;
assign detect_max[601][6] = (mid_1[4823:4816] > top_2[4815:4808]) ? 1 : 0;
assign detect_max[601][7] = (mid_1[4823:4816] > top_2[4823:4816]) ? 1 : 0;
assign detect_max[601][8] = (mid_1[4823:4816] > top_2[4831:4824]) ? 1 : 0;
assign detect_max[601][9] = (mid_1[4823:4816] > mid_0[4815:4808]) ? 1 : 0;
assign detect_max[601][10] = (mid_1[4823:4816] > mid_0[4823:4816]) ? 1 : 0;
assign detect_max[601][11] = (mid_1[4823:4816] > mid_0[4831:4824]) ? 1 : 0;
assign detect_max[601][12] = (mid_1[4823:4816] > mid_1[4815:4808]) ? 1 : 0;
assign detect_max[601][13] = (mid_1[4823:4816] > mid_1[4831:4824]) ? 1 : 0;
assign detect_max[601][14] = (mid_1[4823:4816] > mid_2[4815:4808]) ? 1 : 0;
assign detect_max[601][15] = (mid_1[4823:4816] > mid_2[4823:4816]) ? 1 : 0;
assign detect_max[601][16] = (mid_1[4823:4816] > mid_2[4831:4824]) ? 1 : 0;
assign detect_max[601][17] = (mid_1[4823:4816] > btm_0[4815:4808]) ? 1 : 0;
assign detect_max[601][18] = (mid_1[4823:4816] > btm_0[4823:4816]) ? 1 : 0;
assign detect_max[601][19] = (mid_1[4823:4816] > btm_0[4831:4824]) ? 1 : 0;
assign detect_max[601][20] = (mid_1[4823:4816] > btm_1[4815:4808]) ? 1 : 0;
assign detect_max[601][21] = (mid_1[4823:4816] > btm_1[4823:4816]) ? 1 : 0;
assign detect_max[601][22] = (mid_1[4823:4816] > btm_1[4831:4824]) ? 1 : 0;
assign detect_max[601][23] = (mid_1[4823:4816] > btm_2[4815:4808]) ? 1 : 0;
assign detect_max[601][24] = (mid_1[4823:4816] > btm_2[4823:4816]) ? 1 : 0;
assign detect_max[601][25] = (mid_1[4823:4816] > btm_2[4831:4824]) ? 1 : 0;

assign detect_max[602][0] = (mid_1[4831:4824] > top_0[4823:4816]) ? 1 : 0;
assign detect_max[602][1] = (mid_1[4831:4824] > top_0[4831:4824]) ? 1 : 0;
assign detect_max[602][2] = (mid_1[4831:4824] > top_0[4839:4832]) ? 1 : 0;
assign detect_max[602][3] = (mid_1[4831:4824] > top_1[4823:4816]) ? 1 : 0;
assign detect_max[602][4] = (mid_1[4831:4824] > top_1[4831:4824]) ? 1 : 0;
assign detect_max[602][5] = (mid_1[4831:4824] > top_1[4839:4832]) ? 1 : 0;
assign detect_max[602][6] = (mid_1[4831:4824] > top_2[4823:4816]) ? 1 : 0;
assign detect_max[602][7] = (mid_1[4831:4824] > top_2[4831:4824]) ? 1 : 0;
assign detect_max[602][8] = (mid_1[4831:4824] > top_2[4839:4832]) ? 1 : 0;
assign detect_max[602][9] = (mid_1[4831:4824] > mid_0[4823:4816]) ? 1 : 0;
assign detect_max[602][10] = (mid_1[4831:4824] > mid_0[4831:4824]) ? 1 : 0;
assign detect_max[602][11] = (mid_1[4831:4824] > mid_0[4839:4832]) ? 1 : 0;
assign detect_max[602][12] = (mid_1[4831:4824] > mid_1[4823:4816]) ? 1 : 0;
assign detect_max[602][13] = (mid_1[4831:4824] > mid_1[4839:4832]) ? 1 : 0;
assign detect_max[602][14] = (mid_1[4831:4824] > mid_2[4823:4816]) ? 1 : 0;
assign detect_max[602][15] = (mid_1[4831:4824] > mid_2[4831:4824]) ? 1 : 0;
assign detect_max[602][16] = (mid_1[4831:4824] > mid_2[4839:4832]) ? 1 : 0;
assign detect_max[602][17] = (mid_1[4831:4824] > btm_0[4823:4816]) ? 1 : 0;
assign detect_max[602][18] = (mid_1[4831:4824] > btm_0[4831:4824]) ? 1 : 0;
assign detect_max[602][19] = (mid_1[4831:4824] > btm_0[4839:4832]) ? 1 : 0;
assign detect_max[602][20] = (mid_1[4831:4824] > btm_1[4823:4816]) ? 1 : 0;
assign detect_max[602][21] = (mid_1[4831:4824] > btm_1[4831:4824]) ? 1 : 0;
assign detect_max[602][22] = (mid_1[4831:4824] > btm_1[4839:4832]) ? 1 : 0;
assign detect_max[602][23] = (mid_1[4831:4824] > btm_2[4823:4816]) ? 1 : 0;
assign detect_max[602][24] = (mid_1[4831:4824] > btm_2[4831:4824]) ? 1 : 0;
assign detect_max[602][25] = (mid_1[4831:4824] > btm_2[4839:4832]) ? 1 : 0;

assign detect_max[603][0] = (mid_1[4839:4832] > top_0[4831:4824]) ? 1 : 0;
assign detect_max[603][1] = (mid_1[4839:4832] > top_0[4839:4832]) ? 1 : 0;
assign detect_max[603][2] = (mid_1[4839:4832] > top_0[4847:4840]) ? 1 : 0;
assign detect_max[603][3] = (mid_1[4839:4832] > top_1[4831:4824]) ? 1 : 0;
assign detect_max[603][4] = (mid_1[4839:4832] > top_1[4839:4832]) ? 1 : 0;
assign detect_max[603][5] = (mid_1[4839:4832] > top_1[4847:4840]) ? 1 : 0;
assign detect_max[603][6] = (mid_1[4839:4832] > top_2[4831:4824]) ? 1 : 0;
assign detect_max[603][7] = (mid_1[4839:4832] > top_2[4839:4832]) ? 1 : 0;
assign detect_max[603][8] = (mid_1[4839:4832] > top_2[4847:4840]) ? 1 : 0;
assign detect_max[603][9] = (mid_1[4839:4832] > mid_0[4831:4824]) ? 1 : 0;
assign detect_max[603][10] = (mid_1[4839:4832] > mid_0[4839:4832]) ? 1 : 0;
assign detect_max[603][11] = (mid_1[4839:4832] > mid_0[4847:4840]) ? 1 : 0;
assign detect_max[603][12] = (mid_1[4839:4832] > mid_1[4831:4824]) ? 1 : 0;
assign detect_max[603][13] = (mid_1[4839:4832] > mid_1[4847:4840]) ? 1 : 0;
assign detect_max[603][14] = (mid_1[4839:4832] > mid_2[4831:4824]) ? 1 : 0;
assign detect_max[603][15] = (mid_1[4839:4832] > mid_2[4839:4832]) ? 1 : 0;
assign detect_max[603][16] = (mid_1[4839:4832] > mid_2[4847:4840]) ? 1 : 0;
assign detect_max[603][17] = (mid_1[4839:4832] > btm_0[4831:4824]) ? 1 : 0;
assign detect_max[603][18] = (mid_1[4839:4832] > btm_0[4839:4832]) ? 1 : 0;
assign detect_max[603][19] = (mid_1[4839:4832] > btm_0[4847:4840]) ? 1 : 0;
assign detect_max[603][20] = (mid_1[4839:4832] > btm_1[4831:4824]) ? 1 : 0;
assign detect_max[603][21] = (mid_1[4839:4832] > btm_1[4839:4832]) ? 1 : 0;
assign detect_max[603][22] = (mid_1[4839:4832] > btm_1[4847:4840]) ? 1 : 0;
assign detect_max[603][23] = (mid_1[4839:4832] > btm_2[4831:4824]) ? 1 : 0;
assign detect_max[603][24] = (mid_1[4839:4832] > btm_2[4839:4832]) ? 1 : 0;
assign detect_max[603][25] = (mid_1[4839:4832] > btm_2[4847:4840]) ? 1 : 0;

assign detect_max[604][0] = (mid_1[4847:4840] > top_0[4839:4832]) ? 1 : 0;
assign detect_max[604][1] = (mid_1[4847:4840] > top_0[4847:4840]) ? 1 : 0;
assign detect_max[604][2] = (mid_1[4847:4840] > top_0[4855:4848]) ? 1 : 0;
assign detect_max[604][3] = (mid_1[4847:4840] > top_1[4839:4832]) ? 1 : 0;
assign detect_max[604][4] = (mid_1[4847:4840] > top_1[4847:4840]) ? 1 : 0;
assign detect_max[604][5] = (mid_1[4847:4840] > top_1[4855:4848]) ? 1 : 0;
assign detect_max[604][6] = (mid_1[4847:4840] > top_2[4839:4832]) ? 1 : 0;
assign detect_max[604][7] = (mid_1[4847:4840] > top_2[4847:4840]) ? 1 : 0;
assign detect_max[604][8] = (mid_1[4847:4840] > top_2[4855:4848]) ? 1 : 0;
assign detect_max[604][9] = (mid_1[4847:4840] > mid_0[4839:4832]) ? 1 : 0;
assign detect_max[604][10] = (mid_1[4847:4840] > mid_0[4847:4840]) ? 1 : 0;
assign detect_max[604][11] = (mid_1[4847:4840] > mid_0[4855:4848]) ? 1 : 0;
assign detect_max[604][12] = (mid_1[4847:4840] > mid_1[4839:4832]) ? 1 : 0;
assign detect_max[604][13] = (mid_1[4847:4840] > mid_1[4855:4848]) ? 1 : 0;
assign detect_max[604][14] = (mid_1[4847:4840] > mid_2[4839:4832]) ? 1 : 0;
assign detect_max[604][15] = (mid_1[4847:4840] > mid_2[4847:4840]) ? 1 : 0;
assign detect_max[604][16] = (mid_1[4847:4840] > mid_2[4855:4848]) ? 1 : 0;
assign detect_max[604][17] = (mid_1[4847:4840] > btm_0[4839:4832]) ? 1 : 0;
assign detect_max[604][18] = (mid_1[4847:4840] > btm_0[4847:4840]) ? 1 : 0;
assign detect_max[604][19] = (mid_1[4847:4840] > btm_0[4855:4848]) ? 1 : 0;
assign detect_max[604][20] = (mid_1[4847:4840] > btm_1[4839:4832]) ? 1 : 0;
assign detect_max[604][21] = (mid_1[4847:4840] > btm_1[4847:4840]) ? 1 : 0;
assign detect_max[604][22] = (mid_1[4847:4840] > btm_1[4855:4848]) ? 1 : 0;
assign detect_max[604][23] = (mid_1[4847:4840] > btm_2[4839:4832]) ? 1 : 0;
assign detect_max[604][24] = (mid_1[4847:4840] > btm_2[4847:4840]) ? 1 : 0;
assign detect_max[604][25] = (mid_1[4847:4840] > btm_2[4855:4848]) ? 1 : 0;

assign detect_max[605][0] = (mid_1[4855:4848] > top_0[4847:4840]) ? 1 : 0;
assign detect_max[605][1] = (mid_1[4855:4848] > top_0[4855:4848]) ? 1 : 0;
assign detect_max[605][2] = (mid_1[4855:4848] > top_0[4863:4856]) ? 1 : 0;
assign detect_max[605][3] = (mid_1[4855:4848] > top_1[4847:4840]) ? 1 : 0;
assign detect_max[605][4] = (mid_1[4855:4848] > top_1[4855:4848]) ? 1 : 0;
assign detect_max[605][5] = (mid_1[4855:4848] > top_1[4863:4856]) ? 1 : 0;
assign detect_max[605][6] = (mid_1[4855:4848] > top_2[4847:4840]) ? 1 : 0;
assign detect_max[605][7] = (mid_1[4855:4848] > top_2[4855:4848]) ? 1 : 0;
assign detect_max[605][8] = (mid_1[4855:4848] > top_2[4863:4856]) ? 1 : 0;
assign detect_max[605][9] = (mid_1[4855:4848] > mid_0[4847:4840]) ? 1 : 0;
assign detect_max[605][10] = (mid_1[4855:4848] > mid_0[4855:4848]) ? 1 : 0;
assign detect_max[605][11] = (mid_1[4855:4848] > mid_0[4863:4856]) ? 1 : 0;
assign detect_max[605][12] = (mid_1[4855:4848] > mid_1[4847:4840]) ? 1 : 0;
assign detect_max[605][13] = (mid_1[4855:4848] > mid_1[4863:4856]) ? 1 : 0;
assign detect_max[605][14] = (mid_1[4855:4848] > mid_2[4847:4840]) ? 1 : 0;
assign detect_max[605][15] = (mid_1[4855:4848] > mid_2[4855:4848]) ? 1 : 0;
assign detect_max[605][16] = (mid_1[4855:4848] > mid_2[4863:4856]) ? 1 : 0;
assign detect_max[605][17] = (mid_1[4855:4848] > btm_0[4847:4840]) ? 1 : 0;
assign detect_max[605][18] = (mid_1[4855:4848] > btm_0[4855:4848]) ? 1 : 0;
assign detect_max[605][19] = (mid_1[4855:4848] > btm_0[4863:4856]) ? 1 : 0;
assign detect_max[605][20] = (mid_1[4855:4848] > btm_1[4847:4840]) ? 1 : 0;
assign detect_max[605][21] = (mid_1[4855:4848] > btm_1[4855:4848]) ? 1 : 0;
assign detect_max[605][22] = (mid_1[4855:4848] > btm_1[4863:4856]) ? 1 : 0;
assign detect_max[605][23] = (mid_1[4855:4848] > btm_2[4847:4840]) ? 1 : 0;
assign detect_max[605][24] = (mid_1[4855:4848] > btm_2[4855:4848]) ? 1 : 0;
assign detect_max[605][25] = (mid_1[4855:4848] > btm_2[4863:4856]) ? 1 : 0;

assign detect_max[606][0] = (mid_1[4863:4856] > top_0[4855:4848]) ? 1 : 0;
assign detect_max[606][1] = (mid_1[4863:4856] > top_0[4863:4856]) ? 1 : 0;
assign detect_max[606][2] = (mid_1[4863:4856] > top_0[4871:4864]) ? 1 : 0;
assign detect_max[606][3] = (mid_1[4863:4856] > top_1[4855:4848]) ? 1 : 0;
assign detect_max[606][4] = (mid_1[4863:4856] > top_1[4863:4856]) ? 1 : 0;
assign detect_max[606][5] = (mid_1[4863:4856] > top_1[4871:4864]) ? 1 : 0;
assign detect_max[606][6] = (mid_1[4863:4856] > top_2[4855:4848]) ? 1 : 0;
assign detect_max[606][7] = (mid_1[4863:4856] > top_2[4863:4856]) ? 1 : 0;
assign detect_max[606][8] = (mid_1[4863:4856] > top_2[4871:4864]) ? 1 : 0;
assign detect_max[606][9] = (mid_1[4863:4856] > mid_0[4855:4848]) ? 1 : 0;
assign detect_max[606][10] = (mid_1[4863:4856] > mid_0[4863:4856]) ? 1 : 0;
assign detect_max[606][11] = (mid_1[4863:4856] > mid_0[4871:4864]) ? 1 : 0;
assign detect_max[606][12] = (mid_1[4863:4856] > mid_1[4855:4848]) ? 1 : 0;
assign detect_max[606][13] = (mid_1[4863:4856] > mid_1[4871:4864]) ? 1 : 0;
assign detect_max[606][14] = (mid_1[4863:4856] > mid_2[4855:4848]) ? 1 : 0;
assign detect_max[606][15] = (mid_1[4863:4856] > mid_2[4863:4856]) ? 1 : 0;
assign detect_max[606][16] = (mid_1[4863:4856] > mid_2[4871:4864]) ? 1 : 0;
assign detect_max[606][17] = (mid_1[4863:4856] > btm_0[4855:4848]) ? 1 : 0;
assign detect_max[606][18] = (mid_1[4863:4856] > btm_0[4863:4856]) ? 1 : 0;
assign detect_max[606][19] = (mid_1[4863:4856] > btm_0[4871:4864]) ? 1 : 0;
assign detect_max[606][20] = (mid_1[4863:4856] > btm_1[4855:4848]) ? 1 : 0;
assign detect_max[606][21] = (mid_1[4863:4856] > btm_1[4863:4856]) ? 1 : 0;
assign detect_max[606][22] = (mid_1[4863:4856] > btm_1[4871:4864]) ? 1 : 0;
assign detect_max[606][23] = (mid_1[4863:4856] > btm_2[4855:4848]) ? 1 : 0;
assign detect_max[606][24] = (mid_1[4863:4856] > btm_2[4863:4856]) ? 1 : 0;
assign detect_max[606][25] = (mid_1[4863:4856] > btm_2[4871:4864]) ? 1 : 0;

assign detect_max[607][0] = (mid_1[4871:4864] > top_0[4863:4856]) ? 1 : 0;
assign detect_max[607][1] = (mid_1[4871:4864] > top_0[4871:4864]) ? 1 : 0;
assign detect_max[607][2] = (mid_1[4871:4864] > top_0[4879:4872]) ? 1 : 0;
assign detect_max[607][3] = (mid_1[4871:4864] > top_1[4863:4856]) ? 1 : 0;
assign detect_max[607][4] = (mid_1[4871:4864] > top_1[4871:4864]) ? 1 : 0;
assign detect_max[607][5] = (mid_1[4871:4864] > top_1[4879:4872]) ? 1 : 0;
assign detect_max[607][6] = (mid_1[4871:4864] > top_2[4863:4856]) ? 1 : 0;
assign detect_max[607][7] = (mid_1[4871:4864] > top_2[4871:4864]) ? 1 : 0;
assign detect_max[607][8] = (mid_1[4871:4864] > top_2[4879:4872]) ? 1 : 0;
assign detect_max[607][9] = (mid_1[4871:4864] > mid_0[4863:4856]) ? 1 : 0;
assign detect_max[607][10] = (mid_1[4871:4864] > mid_0[4871:4864]) ? 1 : 0;
assign detect_max[607][11] = (mid_1[4871:4864] > mid_0[4879:4872]) ? 1 : 0;
assign detect_max[607][12] = (mid_1[4871:4864] > mid_1[4863:4856]) ? 1 : 0;
assign detect_max[607][13] = (mid_1[4871:4864] > mid_1[4879:4872]) ? 1 : 0;
assign detect_max[607][14] = (mid_1[4871:4864] > mid_2[4863:4856]) ? 1 : 0;
assign detect_max[607][15] = (mid_1[4871:4864] > mid_2[4871:4864]) ? 1 : 0;
assign detect_max[607][16] = (mid_1[4871:4864] > mid_2[4879:4872]) ? 1 : 0;
assign detect_max[607][17] = (mid_1[4871:4864] > btm_0[4863:4856]) ? 1 : 0;
assign detect_max[607][18] = (mid_1[4871:4864] > btm_0[4871:4864]) ? 1 : 0;
assign detect_max[607][19] = (mid_1[4871:4864] > btm_0[4879:4872]) ? 1 : 0;
assign detect_max[607][20] = (mid_1[4871:4864] > btm_1[4863:4856]) ? 1 : 0;
assign detect_max[607][21] = (mid_1[4871:4864] > btm_1[4871:4864]) ? 1 : 0;
assign detect_max[607][22] = (mid_1[4871:4864] > btm_1[4879:4872]) ? 1 : 0;
assign detect_max[607][23] = (mid_1[4871:4864] > btm_2[4863:4856]) ? 1 : 0;
assign detect_max[607][24] = (mid_1[4871:4864] > btm_2[4871:4864]) ? 1 : 0;
assign detect_max[607][25] = (mid_1[4871:4864] > btm_2[4879:4872]) ? 1 : 0;

assign detect_max[608][0] = (mid_1[4879:4872] > top_0[4871:4864]) ? 1 : 0;
assign detect_max[608][1] = (mid_1[4879:4872] > top_0[4879:4872]) ? 1 : 0;
assign detect_max[608][2] = (mid_1[4879:4872] > top_0[4887:4880]) ? 1 : 0;
assign detect_max[608][3] = (mid_1[4879:4872] > top_1[4871:4864]) ? 1 : 0;
assign detect_max[608][4] = (mid_1[4879:4872] > top_1[4879:4872]) ? 1 : 0;
assign detect_max[608][5] = (mid_1[4879:4872] > top_1[4887:4880]) ? 1 : 0;
assign detect_max[608][6] = (mid_1[4879:4872] > top_2[4871:4864]) ? 1 : 0;
assign detect_max[608][7] = (mid_1[4879:4872] > top_2[4879:4872]) ? 1 : 0;
assign detect_max[608][8] = (mid_1[4879:4872] > top_2[4887:4880]) ? 1 : 0;
assign detect_max[608][9] = (mid_1[4879:4872] > mid_0[4871:4864]) ? 1 : 0;
assign detect_max[608][10] = (mid_1[4879:4872] > mid_0[4879:4872]) ? 1 : 0;
assign detect_max[608][11] = (mid_1[4879:4872] > mid_0[4887:4880]) ? 1 : 0;
assign detect_max[608][12] = (mid_1[4879:4872] > mid_1[4871:4864]) ? 1 : 0;
assign detect_max[608][13] = (mid_1[4879:4872] > mid_1[4887:4880]) ? 1 : 0;
assign detect_max[608][14] = (mid_1[4879:4872] > mid_2[4871:4864]) ? 1 : 0;
assign detect_max[608][15] = (mid_1[4879:4872] > mid_2[4879:4872]) ? 1 : 0;
assign detect_max[608][16] = (mid_1[4879:4872] > mid_2[4887:4880]) ? 1 : 0;
assign detect_max[608][17] = (mid_1[4879:4872] > btm_0[4871:4864]) ? 1 : 0;
assign detect_max[608][18] = (mid_1[4879:4872] > btm_0[4879:4872]) ? 1 : 0;
assign detect_max[608][19] = (mid_1[4879:4872] > btm_0[4887:4880]) ? 1 : 0;
assign detect_max[608][20] = (mid_1[4879:4872] > btm_1[4871:4864]) ? 1 : 0;
assign detect_max[608][21] = (mid_1[4879:4872] > btm_1[4879:4872]) ? 1 : 0;
assign detect_max[608][22] = (mid_1[4879:4872] > btm_1[4887:4880]) ? 1 : 0;
assign detect_max[608][23] = (mid_1[4879:4872] > btm_2[4871:4864]) ? 1 : 0;
assign detect_max[608][24] = (mid_1[4879:4872] > btm_2[4879:4872]) ? 1 : 0;
assign detect_max[608][25] = (mid_1[4879:4872] > btm_2[4887:4880]) ? 1 : 0;

assign detect_max[609][0] = (mid_1[4887:4880] > top_0[4879:4872]) ? 1 : 0;
assign detect_max[609][1] = (mid_1[4887:4880] > top_0[4887:4880]) ? 1 : 0;
assign detect_max[609][2] = (mid_1[4887:4880] > top_0[4895:4888]) ? 1 : 0;
assign detect_max[609][3] = (mid_1[4887:4880] > top_1[4879:4872]) ? 1 : 0;
assign detect_max[609][4] = (mid_1[4887:4880] > top_1[4887:4880]) ? 1 : 0;
assign detect_max[609][5] = (mid_1[4887:4880] > top_1[4895:4888]) ? 1 : 0;
assign detect_max[609][6] = (mid_1[4887:4880] > top_2[4879:4872]) ? 1 : 0;
assign detect_max[609][7] = (mid_1[4887:4880] > top_2[4887:4880]) ? 1 : 0;
assign detect_max[609][8] = (mid_1[4887:4880] > top_2[4895:4888]) ? 1 : 0;
assign detect_max[609][9] = (mid_1[4887:4880] > mid_0[4879:4872]) ? 1 : 0;
assign detect_max[609][10] = (mid_1[4887:4880] > mid_0[4887:4880]) ? 1 : 0;
assign detect_max[609][11] = (mid_1[4887:4880] > mid_0[4895:4888]) ? 1 : 0;
assign detect_max[609][12] = (mid_1[4887:4880] > mid_1[4879:4872]) ? 1 : 0;
assign detect_max[609][13] = (mid_1[4887:4880] > mid_1[4895:4888]) ? 1 : 0;
assign detect_max[609][14] = (mid_1[4887:4880] > mid_2[4879:4872]) ? 1 : 0;
assign detect_max[609][15] = (mid_1[4887:4880] > mid_2[4887:4880]) ? 1 : 0;
assign detect_max[609][16] = (mid_1[4887:4880] > mid_2[4895:4888]) ? 1 : 0;
assign detect_max[609][17] = (mid_1[4887:4880] > btm_0[4879:4872]) ? 1 : 0;
assign detect_max[609][18] = (mid_1[4887:4880] > btm_0[4887:4880]) ? 1 : 0;
assign detect_max[609][19] = (mid_1[4887:4880] > btm_0[4895:4888]) ? 1 : 0;
assign detect_max[609][20] = (mid_1[4887:4880] > btm_1[4879:4872]) ? 1 : 0;
assign detect_max[609][21] = (mid_1[4887:4880] > btm_1[4887:4880]) ? 1 : 0;
assign detect_max[609][22] = (mid_1[4887:4880] > btm_1[4895:4888]) ? 1 : 0;
assign detect_max[609][23] = (mid_1[4887:4880] > btm_2[4879:4872]) ? 1 : 0;
assign detect_max[609][24] = (mid_1[4887:4880] > btm_2[4887:4880]) ? 1 : 0;
assign detect_max[609][25] = (mid_1[4887:4880] > btm_2[4895:4888]) ? 1 : 0;

assign detect_max[610][0] = (mid_1[4895:4888] > top_0[4887:4880]) ? 1 : 0;
assign detect_max[610][1] = (mid_1[4895:4888] > top_0[4895:4888]) ? 1 : 0;
assign detect_max[610][2] = (mid_1[4895:4888] > top_0[4903:4896]) ? 1 : 0;
assign detect_max[610][3] = (mid_1[4895:4888] > top_1[4887:4880]) ? 1 : 0;
assign detect_max[610][4] = (mid_1[4895:4888] > top_1[4895:4888]) ? 1 : 0;
assign detect_max[610][5] = (mid_1[4895:4888] > top_1[4903:4896]) ? 1 : 0;
assign detect_max[610][6] = (mid_1[4895:4888] > top_2[4887:4880]) ? 1 : 0;
assign detect_max[610][7] = (mid_1[4895:4888] > top_2[4895:4888]) ? 1 : 0;
assign detect_max[610][8] = (mid_1[4895:4888] > top_2[4903:4896]) ? 1 : 0;
assign detect_max[610][9] = (mid_1[4895:4888] > mid_0[4887:4880]) ? 1 : 0;
assign detect_max[610][10] = (mid_1[4895:4888] > mid_0[4895:4888]) ? 1 : 0;
assign detect_max[610][11] = (mid_1[4895:4888] > mid_0[4903:4896]) ? 1 : 0;
assign detect_max[610][12] = (mid_1[4895:4888] > mid_1[4887:4880]) ? 1 : 0;
assign detect_max[610][13] = (mid_1[4895:4888] > mid_1[4903:4896]) ? 1 : 0;
assign detect_max[610][14] = (mid_1[4895:4888] > mid_2[4887:4880]) ? 1 : 0;
assign detect_max[610][15] = (mid_1[4895:4888] > mid_2[4895:4888]) ? 1 : 0;
assign detect_max[610][16] = (mid_1[4895:4888] > mid_2[4903:4896]) ? 1 : 0;
assign detect_max[610][17] = (mid_1[4895:4888] > btm_0[4887:4880]) ? 1 : 0;
assign detect_max[610][18] = (mid_1[4895:4888] > btm_0[4895:4888]) ? 1 : 0;
assign detect_max[610][19] = (mid_1[4895:4888] > btm_0[4903:4896]) ? 1 : 0;
assign detect_max[610][20] = (mid_1[4895:4888] > btm_1[4887:4880]) ? 1 : 0;
assign detect_max[610][21] = (mid_1[4895:4888] > btm_1[4895:4888]) ? 1 : 0;
assign detect_max[610][22] = (mid_1[4895:4888] > btm_1[4903:4896]) ? 1 : 0;
assign detect_max[610][23] = (mid_1[4895:4888] > btm_2[4887:4880]) ? 1 : 0;
assign detect_max[610][24] = (mid_1[4895:4888] > btm_2[4895:4888]) ? 1 : 0;
assign detect_max[610][25] = (mid_1[4895:4888] > btm_2[4903:4896]) ? 1 : 0;

assign detect_max[611][0] = (mid_1[4903:4896] > top_0[4895:4888]) ? 1 : 0;
assign detect_max[611][1] = (mid_1[4903:4896] > top_0[4903:4896]) ? 1 : 0;
assign detect_max[611][2] = (mid_1[4903:4896] > top_0[4911:4904]) ? 1 : 0;
assign detect_max[611][3] = (mid_1[4903:4896] > top_1[4895:4888]) ? 1 : 0;
assign detect_max[611][4] = (mid_1[4903:4896] > top_1[4903:4896]) ? 1 : 0;
assign detect_max[611][5] = (mid_1[4903:4896] > top_1[4911:4904]) ? 1 : 0;
assign detect_max[611][6] = (mid_1[4903:4896] > top_2[4895:4888]) ? 1 : 0;
assign detect_max[611][7] = (mid_1[4903:4896] > top_2[4903:4896]) ? 1 : 0;
assign detect_max[611][8] = (mid_1[4903:4896] > top_2[4911:4904]) ? 1 : 0;
assign detect_max[611][9] = (mid_1[4903:4896] > mid_0[4895:4888]) ? 1 : 0;
assign detect_max[611][10] = (mid_1[4903:4896] > mid_0[4903:4896]) ? 1 : 0;
assign detect_max[611][11] = (mid_1[4903:4896] > mid_0[4911:4904]) ? 1 : 0;
assign detect_max[611][12] = (mid_1[4903:4896] > mid_1[4895:4888]) ? 1 : 0;
assign detect_max[611][13] = (mid_1[4903:4896] > mid_1[4911:4904]) ? 1 : 0;
assign detect_max[611][14] = (mid_1[4903:4896] > mid_2[4895:4888]) ? 1 : 0;
assign detect_max[611][15] = (mid_1[4903:4896] > mid_2[4903:4896]) ? 1 : 0;
assign detect_max[611][16] = (mid_1[4903:4896] > mid_2[4911:4904]) ? 1 : 0;
assign detect_max[611][17] = (mid_1[4903:4896] > btm_0[4895:4888]) ? 1 : 0;
assign detect_max[611][18] = (mid_1[4903:4896] > btm_0[4903:4896]) ? 1 : 0;
assign detect_max[611][19] = (mid_1[4903:4896] > btm_0[4911:4904]) ? 1 : 0;
assign detect_max[611][20] = (mid_1[4903:4896] > btm_1[4895:4888]) ? 1 : 0;
assign detect_max[611][21] = (mid_1[4903:4896] > btm_1[4903:4896]) ? 1 : 0;
assign detect_max[611][22] = (mid_1[4903:4896] > btm_1[4911:4904]) ? 1 : 0;
assign detect_max[611][23] = (mid_1[4903:4896] > btm_2[4895:4888]) ? 1 : 0;
assign detect_max[611][24] = (mid_1[4903:4896] > btm_2[4903:4896]) ? 1 : 0;
assign detect_max[611][25] = (mid_1[4903:4896] > btm_2[4911:4904]) ? 1 : 0;

assign detect_max[612][0] = (mid_1[4911:4904] > top_0[4903:4896]) ? 1 : 0;
assign detect_max[612][1] = (mid_1[4911:4904] > top_0[4911:4904]) ? 1 : 0;
assign detect_max[612][2] = (mid_1[4911:4904] > top_0[4919:4912]) ? 1 : 0;
assign detect_max[612][3] = (mid_1[4911:4904] > top_1[4903:4896]) ? 1 : 0;
assign detect_max[612][4] = (mid_1[4911:4904] > top_1[4911:4904]) ? 1 : 0;
assign detect_max[612][5] = (mid_1[4911:4904] > top_1[4919:4912]) ? 1 : 0;
assign detect_max[612][6] = (mid_1[4911:4904] > top_2[4903:4896]) ? 1 : 0;
assign detect_max[612][7] = (mid_1[4911:4904] > top_2[4911:4904]) ? 1 : 0;
assign detect_max[612][8] = (mid_1[4911:4904] > top_2[4919:4912]) ? 1 : 0;
assign detect_max[612][9] = (mid_1[4911:4904] > mid_0[4903:4896]) ? 1 : 0;
assign detect_max[612][10] = (mid_1[4911:4904] > mid_0[4911:4904]) ? 1 : 0;
assign detect_max[612][11] = (mid_1[4911:4904] > mid_0[4919:4912]) ? 1 : 0;
assign detect_max[612][12] = (mid_1[4911:4904] > mid_1[4903:4896]) ? 1 : 0;
assign detect_max[612][13] = (mid_1[4911:4904] > mid_1[4919:4912]) ? 1 : 0;
assign detect_max[612][14] = (mid_1[4911:4904] > mid_2[4903:4896]) ? 1 : 0;
assign detect_max[612][15] = (mid_1[4911:4904] > mid_2[4911:4904]) ? 1 : 0;
assign detect_max[612][16] = (mid_1[4911:4904] > mid_2[4919:4912]) ? 1 : 0;
assign detect_max[612][17] = (mid_1[4911:4904] > btm_0[4903:4896]) ? 1 : 0;
assign detect_max[612][18] = (mid_1[4911:4904] > btm_0[4911:4904]) ? 1 : 0;
assign detect_max[612][19] = (mid_1[4911:4904] > btm_0[4919:4912]) ? 1 : 0;
assign detect_max[612][20] = (mid_1[4911:4904] > btm_1[4903:4896]) ? 1 : 0;
assign detect_max[612][21] = (mid_1[4911:4904] > btm_1[4911:4904]) ? 1 : 0;
assign detect_max[612][22] = (mid_1[4911:4904] > btm_1[4919:4912]) ? 1 : 0;
assign detect_max[612][23] = (mid_1[4911:4904] > btm_2[4903:4896]) ? 1 : 0;
assign detect_max[612][24] = (mid_1[4911:4904] > btm_2[4911:4904]) ? 1 : 0;
assign detect_max[612][25] = (mid_1[4911:4904] > btm_2[4919:4912]) ? 1 : 0;

assign detect_max[613][0] = (mid_1[4919:4912] > top_0[4911:4904]) ? 1 : 0;
assign detect_max[613][1] = (mid_1[4919:4912] > top_0[4919:4912]) ? 1 : 0;
assign detect_max[613][2] = (mid_1[4919:4912] > top_0[4927:4920]) ? 1 : 0;
assign detect_max[613][3] = (mid_1[4919:4912] > top_1[4911:4904]) ? 1 : 0;
assign detect_max[613][4] = (mid_1[4919:4912] > top_1[4919:4912]) ? 1 : 0;
assign detect_max[613][5] = (mid_1[4919:4912] > top_1[4927:4920]) ? 1 : 0;
assign detect_max[613][6] = (mid_1[4919:4912] > top_2[4911:4904]) ? 1 : 0;
assign detect_max[613][7] = (mid_1[4919:4912] > top_2[4919:4912]) ? 1 : 0;
assign detect_max[613][8] = (mid_1[4919:4912] > top_2[4927:4920]) ? 1 : 0;
assign detect_max[613][9] = (mid_1[4919:4912] > mid_0[4911:4904]) ? 1 : 0;
assign detect_max[613][10] = (mid_1[4919:4912] > mid_0[4919:4912]) ? 1 : 0;
assign detect_max[613][11] = (mid_1[4919:4912] > mid_0[4927:4920]) ? 1 : 0;
assign detect_max[613][12] = (mid_1[4919:4912] > mid_1[4911:4904]) ? 1 : 0;
assign detect_max[613][13] = (mid_1[4919:4912] > mid_1[4927:4920]) ? 1 : 0;
assign detect_max[613][14] = (mid_1[4919:4912] > mid_2[4911:4904]) ? 1 : 0;
assign detect_max[613][15] = (mid_1[4919:4912] > mid_2[4919:4912]) ? 1 : 0;
assign detect_max[613][16] = (mid_1[4919:4912] > mid_2[4927:4920]) ? 1 : 0;
assign detect_max[613][17] = (mid_1[4919:4912] > btm_0[4911:4904]) ? 1 : 0;
assign detect_max[613][18] = (mid_1[4919:4912] > btm_0[4919:4912]) ? 1 : 0;
assign detect_max[613][19] = (mid_1[4919:4912] > btm_0[4927:4920]) ? 1 : 0;
assign detect_max[613][20] = (mid_1[4919:4912] > btm_1[4911:4904]) ? 1 : 0;
assign detect_max[613][21] = (mid_1[4919:4912] > btm_1[4919:4912]) ? 1 : 0;
assign detect_max[613][22] = (mid_1[4919:4912] > btm_1[4927:4920]) ? 1 : 0;
assign detect_max[613][23] = (mid_1[4919:4912] > btm_2[4911:4904]) ? 1 : 0;
assign detect_max[613][24] = (mid_1[4919:4912] > btm_2[4919:4912]) ? 1 : 0;
assign detect_max[613][25] = (mid_1[4919:4912] > btm_2[4927:4920]) ? 1 : 0;

assign detect_max[614][0] = (mid_1[4927:4920] > top_0[4919:4912]) ? 1 : 0;
assign detect_max[614][1] = (mid_1[4927:4920] > top_0[4927:4920]) ? 1 : 0;
assign detect_max[614][2] = (mid_1[4927:4920] > top_0[4935:4928]) ? 1 : 0;
assign detect_max[614][3] = (mid_1[4927:4920] > top_1[4919:4912]) ? 1 : 0;
assign detect_max[614][4] = (mid_1[4927:4920] > top_1[4927:4920]) ? 1 : 0;
assign detect_max[614][5] = (mid_1[4927:4920] > top_1[4935:4928]) ? 1 : 0;
assign detect_max[614][6] = (mid_1[4927:4920] > top_2[4919:4912]) ? 1 : 0;
assign detect_max[614][7] = (mid_1[4927:4920] > top_2[4927:4920]) ? 1 : 0;
assign detect_max[614][8] = (mid_1[4927:4920] > top_2[4935:4928]) ? 1 : 0;
assign detect_max[614][9] = (mid_1[4927:4920] > mid_0[4919:4912]) ? 1 : 0;
assign detect_max[614][10] = (mid_1[4927:4920] > mid_0[4927:4920]) ? 1 : 0;
assign detect_max[614][11] = (mid_1[4927:4920] > mid_0[4935:4928]) ? 1 : 0;
assign detect_max[614][12] = (mid_1[4927:4920] > mid_1[4919:4912]) ? 1 : 0;
assign detect_max[614][13] = (mid_1[4927:4920] > mid_1[4935:4928]) ? 1 : 0;
assign detect_max[614][14] = (mid_1[4927:4920] > mid_2[4919:4912]) ? 1 : 0;
assign detect_max[614][15] = (mid_1[4927:4920] > mid_2[4927:4920]) ? 1 : 0;
assign detect_max[614][16] = (mid_1[4927:4920] > mid_2[4935:4928]) ? 1 : 0;
assign detect_max[614][17] = (mid_1[4927:4920] > btm_0[4919:4912]) ? 1 : 0;
assign detect_max[614][18] = (mid_1[4927:4920] > btm_0[4927:4920]) ? 1 : 0;
assign detect_max[614][19] = (mid_1[4927:4920] > btm_0[4935:4928]) ? 1 : 0;
assign detect_max[614][20] = (mid_1[4927:4920] > btm_1[4919:4912]) ? 1 : 0;
assign detect_max[614][21] = (mid_1[4927:4920] > btm_1[4927:4920]) ? 1 : 0;
assign detect_max[614][22] = (mid_1[4927:4920] > btm_1[4935:4928]) ? 1 : 0;
assign detect_max[614][23] = (mid_1[4927:4920] > btm_2[4919:4912]) ? 1 : 0;
assign detect_max[614][24] = (mid_1[4927:4920] > btm_2[4927:4920]) ? 1 : 0;
assign detect_max[614][25] = (mid_1[4927:4920] > btm_2[4935:4928]) ? 1 : 0;

assign detect_max[615][0] = (mid_1[4935:4928] > top_0[4927:4920]) ? 1 : 0;
assign detect_max[615][1] = (mid_1[4935:4928] > top_0[4935:4928]) ? 1 : 0;
assign detect_max[615][2] = (mid_1[4935:4928] > top_0[4943:4936]) ? 1 : 0;
assign detect_max[615][3] = (mid_1[4935:4928] > top_1[4927:4920]) ? 1 : 0;
assign detect_max[615][4] = (mid_1[4935:4928] > top_1[4935:4928]) ? 1 : 0;
assign detect_max[615][5] = (mid_1[4935:4928] > top_1[4943:4936]) ? 1 : 0;
assign detect_max[615][6] = (mid_1[4935:4928] > top_2[4927:4920]) ? 1 : 0;
assign detect_max[615][7] = (mid_1[4935:4928] > top_2[4935:4928]) ? 1 : 0;
assign detect_max[615][8] = (mid_1[4935:4928] > top_2[4943:4936]) ? 1 : 0;
assign detect_max[615][9] = (mid_1[4935:4928] > mid_0[4927:4920]) ? 1 : 0;
assign detect_max[615][10] = (mid_1[4935:4928] > mid_0[4935:4928]) ? 1 : 0;
assign detect_max[615][11] = (mid_1[4935:4928] > mid_0[4943:4936]) ? 1 : 0;
assign detect_max[615][12] = (mid_1[4935:4928] > mid_1[4927:4920]) ? 1 : 0;
assign detect_max[615][13] = (mid_1[4935:4928] > mid_1[4943:4936]) ? 1 : 0;
assign detect_max[615][14] = (mid_1[4935:4928] > mid_2[4927:4920]) ? 1 : 0;
assign detect_max[615][15] = (mid_1[4935:4928] > mid_2[4935:4928]) ? 1 : 0;
assign detect_max[615][16] = (mid_1[4935:4928] > mid_2[4943:4936]) ? 1 : 0;
assign detect_max[615][17] = (mid_1[4935:4928] > btm_0[4927:4920]) ? 1 : 0;
assign detect_max[615][18] = (mid_1[4935:4928] > btm_0[4935:4928]) ? 1 : 0;
assign detect_max[615][19] = (mid_1[4935:4928] > btm_0[4943:4936]) ? 1 : 0;
assign detect_max[615][20] = (mid_1[4935:4928] > btm_1[4927:4920]) ? 1 : 0;
assign detect_max[615][21] = (mid_1[4935:4928] > btm_1[4935:4928]) ? 1 : 0;
assign detect_max[615][22] = (mid_1[4935:4928] > btm_1[4943:4936]) ? 1 : 0;
assign detect_max[615][23] = (mid_1[4935:4928] > btm_2[4927:4920]) ? 1 : 0;
assign detect_max[615][24] = (mid_1[4935:4928] > btm_2[4935:4928]) ? 1 : 0;
assign detect_max[615][25] = (mid_1[4935:4928] > btm_2[4943:4936]) ? 1 : 0;

assign detect_max[616][0] = (mid_1[4943:4936] > top_0[4935:4928]) ? 1 : 0;
assign detect_max[616][1] = (mid_1[4943:4936] > top_0[4943:4936]) ? 1 : 0;
assign detect_max[616][2] = (mid_1[4943:4936] > top_0[4951:4944]) ? 1 : 0;
assign detect_max[616][3] = (mid_1[4943:4936] > top_1[4935:4928]) ? 1 : 0;
assign detect_max[616][4] = (mid_1[4943:4936] > top_1[4943:4936]) ? 1 : 0;
assign detect_max[616][5] = (mid_1[4943:4936] > top_1[4951:4944]) ? 1 : 0;
assign detect_max[616][6] = (mid_1[4943:4936] > top_2[4935:4928]) ? 1 : 0;
assign detect_max[616][7] = (mid_1[4943:4936] > top_2[4943:4936]) ? 1 : 0;
assign detect_max[616][8] = (mid_1[4943:4936] > top_2[4951:4944]) ? 1 : 0;
assign detect_max[616][9] = (mid_1[4943:4936] > mid_0[4935:4928]) ? 1 : 0;
assign detect_max[616][10] = (mid_1[4943:4936] > mid_0[4943:4936]) ? 1 : 0;
assign detect_max[616][11] = (mid_1[4943:4936] > mid_0[4951:4944]) ? 1 : 0;
assign detect_max[616][12] = (mid_1[4943:4936] > mid_1[4935:4928]) ? 1 : 0;
assign detect_max[616][13] = (mid_1[4943:4936] > mid_1[4951:4944]) ? 1 : 0;
assign detect_max[616][14] = (mid_1[4943:4936] > mid_2[4935:4928]) ? 1 : 0;
assign detect_max[616][15] = (mid_1[4943:4936] > mid_2[4943:4936]) ? 1 : 0;
assign detect_max[616][16] = (mid_1[4943:4936] > mid_2[4951:4944]) ? 1 : 0;
assign detect_max[616][17] = (mid_1[4943:4936] > btm_0[4935:4928]) ? 1 : 0;
assign detect_max[616][18] = (mid_1[4943:4936] > btm_0[4943:4936]) ? 1 : 0;
assign detect_max[616][19] = (mid_1[4943:4936] > btm_0[4951:4944]) ? 1 : 0;
assign detect_max[616][20] = (mid_1[4943:4936] > btm_1[4935:4928]) ? 1 : 0;
assign detect_max[616][21] = (mid_1[4943:4936] > btm_1[4943:4936]) ? 1 : 0;
assign detect_max[616][22] = (mid_1[4943:4936] > btm_1[4951:4944]) ? 1 : 0;
assign detect_max[616][23] = (mid_1[4943:4936] > btm_2[4935:4928]) ? 1 : 0;
assign detect_max[616][24] = (mid_1[4943:4936] > btm_2[4943:4936]) ? 1 : 0;
assign detect_max[616][25] = (mid_1[4943:4936] > btm_2[4951:4944]) ? 1 : 0;

assign detect_max[617][0] = (mid_1[4951:4944] > top_0[4943:4936]) ? 1 : 0;
assign detect_max[617][1] = (mid_1[4951:4944] > top_0[4951:4944]) ? 1 : 0;
assign detect_max[617][2] = (mid_1[4951:4944] > top_0[4959:4952]) ? 1 : 0;
assign detect_max[617][3] = (mid_1[4951:4944] > top_1[4943:4936]) ? 1 : 0;
assign detect_max[617][4] = (mid_1[4951:4944] > top_1[4951:4944]) ? 1 : 0;
assign detect_max[617][5] = (mid_1[4951:4944] > top_1[4959:4952]) ? 1 : 0;
assign detect_max[617][6] = (mid_1[4951:4944] > top_2[4943:4936]) ? 1 : 0;
assign detect_max[617][7] = (mid_1[4951:4944] > top_2[4951:4944]) ? 1 : 0;
assign detect_max[617][8] = (mid_1[4951:4944] > top_2[4959:4952]) ? 1 : 0;
assign detect_max[617][9] = (mid_1[4951:4944] > mid_0[4943:4936]) ? 1 : 0;
assign detect_max[617][10] = (mid_1[4951:4944] > mid_0[4951:4944]) ? 1 : 0;
assign detect_max[617][11] = (mid_1[4951:4944] > mid_0[4959:4952]) ? 1 : 0;
assign detect_max[617][12] = (mid_1[4951:4944] > mid_1[4943:4936]) ? 1 : 0;
assign detect_max[617][13] = (mid_1[4951:4944] > mid_1[4959:4952]) ? 1 : 0;
assign detect_max[617][14] = (mid_1[4951:4944] > mid_2[4943:4936]) ? 1 : 0;
assign detect_max[617][15] = (mid_1[4951:4944] > mid_2[4951:4944]) ? 1 : 0;
assign detect_max[617][16] = (mid_1[4951:4944] > mid_2[4959:4952]) ? 1 : 0;
assign detect_max[617][17] = (mid_1[4951:4944] > btm_0[4943:4936]) ? 1 : 0;
assign detect_max[617][18] = (mid_1[4951:4944] > btm_0[4951:4944]) ? 1 : 0;
assign detect_max[617][19] = (mid_1[4951:4944] > btm_0[4959:4952]) ? 1 : 0;
assign detect_max[617][20] = (mid_1[4951:4944] > btm_1[4943:4936]) ? 1 : 0;
assign detect_max[617][21] = (mid_1[4951:4944] > btm_1[4951:4944]) ? 1 : 0;
assign detect_max[617][22] = (mid_1[4951:4944] > btm_1[4959:4952]) ? 1 : 0;
assign detect_max[617][23] = (mid_1[4951:4944] > btm_2[4943:4936]) ? 1 : 0;
assign detect_max[617][24] = (mid_1[4951:4944] > btm_2[4951:4944]) ? 1 : 0;
assign detect_max[617][25] = (mid_1[4951:4944] > btm_2[4959:4952]) ? 1 : 0;

assign detect_max[618][0] = (mid_1[4959:4952] > top_0[4951:4944]) ? 1 : 0;
assign detect_max[618][1] = (mid_1[4959:4952] > top_0[4959:4952]) ? 1 : 0;
assign detect_max[618][2] = (mid_1[4959:4952] > top_0[4967:4960]) ? 1 : 0;
assign detect_max[618][3] = (mid_1[4959:4952] > top_1[4951:4944]) ? 1 : 0;
assign detect_max[618][4] = (mid_1[4959:4952] > top_1[4959:4952]) ? 1 : 0;
assign detect_max[618][5] = (mid_1[4959:4952] > top_1[4967:4960]) ? 1 : 0;
assign detect_max[618][6] = (mid_1[4959:4952] > top_2[4951:4944]) ? 1 : 0;
assign detect_max[618][7] = (mid_1[4959:4952] > top_2[4959:4952]) ? 1 : 0;
assign detect_max[618][8] = (mid_1[4959:4952] > top_2[4967:4960]) ? 1 : 0;
assign detect_max[618][9] = (mid_1[4959:4952] > mid_0[4951:4944]) ? 1 : 0;
assign detect_max[618][10] = (mid_1[4959:4952] > mid_0[4959:4952]) ? 1 : 0;
assign detect_max[618][11] = (mid_1[4959:4952] > mid_0[4967:4960]) ? 1 : 0;
assign detect_max[618][12] = (mid_1[4959:4952] > mid_1[4951:4944]) ? 1 : 0;
assign detect_max[618][13] = (mid_1[4959:4952] > mid_1[4967:4960]) ? 1 : 0;
assign detect_max[618][14] = (mid_1[4959:4952] > mid_2[4951:4944]) ? 1 : 0;
assign detect_max[618][15] = (mid_1[4959:4952] > mid_2[4959:4952]) ? 1 : 0;
assign detect_max[618][16] = (mid_1[4959:4952] > mid_2[4967:4960]) ? 1 : 0;
assign detect_max[618][17] = (mid_1[4959:4952] > btm_0[4951:4944]) ? 1 : 0;
assign detect_max[618][18] = (mid_1[4959:4952] > btm_0[4959:4952]) ? 1 : 0;
assign detect_max[618][19] = (mid_1[4959:4952] > btm_0[4967:4960]) ? 1 : 0;
assign detect_max[618][20] = (mid_1[4959:4952] > btm_1[4951:4944]) ? 1 : 0;
assign detect_max[618][21] = (mid_1[4959:4952] > btm_1[4959:4952]) ? 1 : 0;
assign detect_max[618][22] = (mid_1[4959:4952] > btm_1[4967:4960]) ? 1 : 0;
assign detect_max[618][23] = (mid_1[4959:4952] > btm_2[4951:4944]) ? 1 : 0;
assign detect_max[618][24] = (mid_1[4959:4952] > btm_2[4959:4952]) ? 1 : 0;
assign detect_max[618][25] = (mid_1[4959:4952] > btm_2[4967:4960]) ? 1 : 0;

assign detect_max[619][0] = (mid_1[4967:4960] > top_0[4959:4952]) ? 1 : 0;
assign detect_max[619][1] = (mid_1[4967:4960] > top_0[4967:4960]) ? 1 : 0;
assign detect_max[619][2] = (mid_1[4967:4960] > top_0[4975:4968]) ? 1 : 0;
assign detect_max[619][3] = (mid_1[4967:4960] > top_1[4959:4952]) ? 1 : 0;
assign detect_max[619][4] = (mid_1[4967:4960] > top_1[4967:4960]) ? 1 : 0;
assign detect_max[619][5] = (mid_1[4967:4960] > top_1[4975:4968]) ? 1 : 0;
assign detect_max[619][6] = (mid_1[4967:4960] > top_2[4959:4952]) ? 1 : 0;
assign detect_max[619][7] = (mid_1[4967:4960] > top_2[4967:4960]) ? 1 : 0;
assign detect_max[619][8] = (mid_1[4967:4960] > top_2[4975:4968]) ? 1 : 0;
assign detect_max[619][9] = (mid_1[4967:4960] > mid_0[4959:4952]) ? 1 : 0;
assign detect_max[619][10] = (mid_1[4967:4960] > mid_0[4967:4960]) ? 1 : 0;
assign detect_max[619][11] = (mid_1[4967:4960] > mid_0[4975:4968]) ? 1 : 0;
assign detect_max[619][12] = (mid_1[4967:4960] > mid_1[4959:4952]) ? 1 : 0;
assign detect_max[619][13] = (mid_1[4967:4960] > mid_1[4975:4968]) ? 1 : 0;
assign detect_max[619][14] = (mid_1[4967:4960] > mid_2[4959:4952]) ? 1 : 0;
assign detect_max[619][15] = (mid_1[4967:4960] > mid_2[4967:4960]) ? 1 : 0;
assign detect_max[619][16] = (mid_1[4967:4960] > mid_2[4975:4968]) ? 1 : 0;
assign detect_max[619][17] = (mid_1[4967:4960] > btm_0[4959:4952]) ? 1 : 0;
assign detect_max[619][18] = (mid_1[4967:4960] > btm_0[4967:4960]) ? 1 : 0;
assign detect_max[619][19] = (mid_1[4967:4960] > btm_0[4975:4968]) ? 1 : 0;
assign detect_max[619][20] = (mid_1[4967:4960] > btm_1[4959:4952]) ? 1 : 0;
assign detect_max[619][21] = (mid_1[4967:4960] > btm_1[4967:4960]) ? 1 : 0;
assign detect_max[619][22] = (mid_1[4967:4960] > btm_1[4975:4968]) ? 1 : 0;
assign detect_max[619][23] = (mid_1[4967:4960] > btm_2[4959:4952]) ? 1 : 0;
assign detect_max[619][24] = (mid_1[4967:4960] > btm_2[4967:4960]) ? 1 : 0;
assign detect_max[619][25] = (mid_1[4967:4960] > btm_2[4975:4968]) ? 1 : 0;

assign detect_max[620][0] = (mid_1[4975:4968] > top_0[4967:4960]) ? 1 : 0;
assign detect_max[620][1] = (mid_1[4975:4968] > top_0[4975:4968]) ? 1 : 0;
assign detect_max[620][2] = (mid_1[4975:4968] > top_0[4983:4976]) ? 1 : 0;
assign detect_max[620][3] = (mid_1[4975:4968] > top_1[4967:4960]) ? 1 : 0;
assign detect_max[620][4] = (mid_1[4975:4968] > top_1[4975:4968]) ? 1 : 0;
assign detect_max[620][5] = (mid_1[4975:4968] > top_1[4983:4976]) ? 1 : 0;
assign detect_max[620][6] = (mid_1[4975:4968] > top_2[4967:4960]) ? 1 : 0;
assign detect_max[620][7] = (mid_1[4975:4968] > top_2[4975:4968]) ? 1 : 0;
assign detect_max[620][8] = (mid_1[4975:4968] > top_2[4983:4976]) ? 1 : 0;
assign detect_max[620][9] = (mid_1[4975:4968] > mid_0[4967:4960]) ? 1 : 0;
assign detect_max[620][10] = (mid_1[4975:4968] > mid_0[4975:4968]) ? 1 : 0;
assign detect_max[620][11] = (mid_1[4975:4968] > mid_0[4983:4976]) ? 1 : 0;
assign detect_max[620][12] = (mid_1[4975:4968] > mid_1[4967:4960]) ? 1 : 0;
assign detect_max[620][13] = (mid_1[4975:4968] > mid_1[4983:4976]) ? 1 : 0;
assign detect_max[620][14] = (mid_1[4975:4968] > mid_2[4967:4960]) ? 1 : 0;
assign detect_max[620][15] = (mid_1[4975:4968] > mid_2[4975:4968]) ? 1 : 0;
assign detect_max[620][16] = (mid_1[4975:4968] > mid_2[4983:4976]) ? 1 : 0;
assign detect_max[620][17] = (mid_1[4975:4968] > btm_0[4967:4960]) ? 1 : 0;
assign detect_max[620][18] = (mid_1[4975:4968] > btm_0[4975:4968]) ? 1 : 0;
assign detect_max[620][19] = (mid_1[4975:4968] > btm_0[4983:4976]) ? 1 : 0;
assign detect_max[620][20] = (mid_1[4975:4968] > btm_1[4967:4960]) ? 1 : 0;
assign detect_max[620][21] = (mid_1[4975:4968] > btm_1[4975:4968]) ? 1 : 0;
assign detect_max[620][22] = (mid_1[4975:4968] > btm_1[4983:4976]) ? 1 : 0;
assign detect_max[620][23] = (mid_1[4975:4968] > btm_2[4967:4960]) ? 1 : 0;
assign detect_max[620][24] = (mid_1[4975:4968] > btm_2[4975:4968]) ? 1 : 0;
assign detect_max[620][25] = (mid_1[4975:4968] > btm_2[4983:4976]) ? 1 : 0;

assign detect_max[621][0] = (mid_1[4983:4976] > top_0[4975:4968]) ? 1 : 0;
assign detect_max[621][1] = (mid_1[4983:4976] > top_0[4983:4976]) ? 1 : 0;
assign detect_max[621][2] = (mid_1[4983:4976] > top_0[4991:4984]) ? 1 : 0;
assign detect_max[621][3] = (mid_1[4983:4976] > top_1[4975:4968]) ? 1 : 0;
assign detect_max[621][4] = (mid_1[4983:4976] > top_1[4983:4976]) ? 1 : 0;
assign detect_max[621][5] = (mid_1[4983:4976] > top_1[4991:4984]) ? 1 : 0;
assign detect_max[621][6] = (mid_1[4983:4976] > top_2[4975:4968]) ? 1 : 0;
assign detect_max[621][7] = (mid_1[4983:4976] > top_2[4983:4976]) ? 1 : 0;
assign detect_max[621][8] = (mid_1[4983:4976] > top_2[4991:4984]) ? 1 : 0;
assign detect_max[621][9] = (mid_1[4983:4976] > mid_0[4975:4968]) ? 1 : 0;
assign detect_max[621][10] = (mid_1[4983:4976] > mid_0[4983:4976]) ? 1 : 0;
assign detect_max[621][11] = (mid_1[4983:4976] > mid_0[4991:4984]) ? 1 : 0;
assign detect_max[621][12] = (mid_1[4983:4976] > mid_1[4975:4968]) ? 1 : 0;
assign detect_max[621][13] = (mid_1[4983:4976] > mid_1[4991:4984]) ? 1 : 0;
assign detect_max[621][14] = (mid_1[4983:4976] > mid_2[4975:4968]) ? 1 : 0;
assign detect_max[621][15] = (mid_1[4983:4976] > mid_2[4983:4976]) ? 1 : 0;
assign detect_max[621][16] = (mid_1[4983:4976] > mid_2[4991:4984]) ? 1 : 0;
assign detect_max[621][17] = (mid_1[4983:4976] > btm_0[4975:4968]) ? 1 : 0;
assign detect_max[621][18] = (mid_1[4983:4976] > btm_0[4983:4976]) ? 1 : 0;
assign detect_max[621][19] = (mid_1[4983:4976] > btm_0[4991:4984]) ? 1 : 0;
assign detect_max[621][20] = (mid_1[4983:4976] > btm_1[4975:4968]) ? 1 : 0;
assign detect_max[621][21] = (mid_1[4983:4976] > btm_1[4983:4976]) ? 1 : 0;
assign detect_max[621][22] = (mid_1[4983:4976] > btm_1[4991:4984]) ? 1 : 0;
assign detect_max[621][23] = (mid_1[4983:4976] > btm_2[4975:4968]) ? 1 : 0;
assign detect_max[621][24] = (mid_1[4983:4976] > btm_2[4983:4976]) ? 1 : 0;
assign detect_max[621][25] = (mid_1[4983:4976] > btm_2[4991:4984]) ? 1 : 0;

assign detect_max[622][0] = (mid_1[4991:4984] > top_0[4983:4976]) ? 1 : 0;
assign detect_max[622][1] = (mid_1[4991:4984] > top_0[4991:4984]) ? 1 : 0;
assign detect_max[622][2] = (mid_1[4991:4984] > top_0[4999:4992]) ? 1 : 0;
assign detect_max[622][3] = (mid_1[4991:4984] > top_1[4983:4976]) ? 1 : 0;
assign detect_max[622][4] = (mid_1[4991:4984] > top_1[4991:4984]) ? 1 : 0;
assign detect_max[622][5] = (mid_1[4991:4984] > top_1[4999:4992]) ? 1 : 0;
assign detect_max[622][6] = (mid_1[4991:4984] > top_2[4983:4976]) ? 1 : 0;
assign detect_max[622][7] = (mid_1[4991:4984] > top_2[4991:4984]) ? 1 : 0;
assign detect_max[622][8] = (mid_1[4991:4984] > top_2[4999:4992]) ? 1 : 0;
assign detect_max[622][9] = (mid_1[4991:4984] > mid_0[4983:4976]) ? 1 : 0;
assign detect_max[622][10] = (mid_1[4991:4984] > mid_0[4991:4984]) ? 1 : 0;
assign detect_max[622][11] = (mid_1[4991:4984] > mid_0[4999:4992]) ? 1 : 0;
assign detect_max[622][12] = (mid_1[4991:4984] > mid_1[4983:4976]) ? 1 : 0;
assign detect_max[622][13] = (mid_1[4991:4984] > mid_1[4999:4992]) ? 1 : 0;
assign detect_max[622][14] = (mid_1[4991:4984] > mid_2[4983:4976]) ? 1 : 0;
assign detect_max[622][15] = (mid_1[4991:4984] > mid_2[4991:4984]) ? 1 : 0;
assign detect_max[622][16] = (mid_1[4991:4984] > mid_2[4999:4992]) ? 1 : 0;
assign detect_max[622][17] = (mid_1[4991:4984] > btm_0[4983:4976]) ? 1 : 0;
assign detect_max[622][18] = (mid_1[4991:4984] > btm_0[4991:4984]) ? 1 : 0;
assign detect_max[622][19] = (mid_1[4991:4984] > btm_0[4999:4992]) ? 1 : 0;
assign detect_max[622][20] = (mid_1[4991:4984] > btm_1[4983:4976]) ? 1 : 0;
assign detect_max[622][21] = (mid_1[4991:4984] > btm_1[4991:4984]) ? 1 : 0;
assign detect_max[622][22] = (mid_1[4991:4984] > btm_1[4999:4992]) ? 1 : 0;
assign detect_max[622][23] = (mid_1[4991:4984] > btm_2[4983:4976]) ? 1 : 0;
assign detect_max[622][24] = (mid_1[4991:4984] > btm_2[4991:4984]) ? 1 : 0;
assign detect_max[622][25] = (mid_1[4991:4984] > btm_2[4999:4992]) ? 1 : 0;

assign detect_max[623][0] = (mid_1[4999:4992] > top_0[4991:4984]) ? 1 : 0;
assign detect_max[623][1] = (mid_1[4999:4992] > top_0[4999:4992]) ? 1 : 0;
assign detect_max[623][2] = (mid_1[4999:4992] > top_0[5007:5000]) ? 1 : 0;
assign detect_max[623][3] = (mid_1[4999:4992] > top_1[4991:4984]) ? 1 : 0;
assign detect_max[623][4] = (mid_1[4999:4992] > top_1[4999:4992]) ? 1 : 0;
assign detect_max[623][5] = (mid_1[4999:4992] > top_1[5007:5000]) ? 1 : 0;
assign detect_max[623][6] = (mid_1[4999:4992] > top_2[4991:4984]) ? 1 : 0;
assign detect_max[623][7] = (mid_1[4999:4992] > top_2[4999:4992]) ? 1 : 0;
assign detect_max[623][8] = (mid_1[4999:4992] > top_2[5007:5000]) ? 1 : 0;
assign detect_max[623][9] = (mid_1[4999:4992] > mid_0[4991:4984]) ? 1 : 0;
assign detect_max[623][10] = (mid_1[4999:4992] > mid_0[4999:4992]) ? 1 : 0;
assign detect_max[623][11] = (mid_1[4999:4992] > mid_0[5007:5000]) ? 1 : 0;
assign detect_max[623][12] = (mid_1[4999:4992] > mid_1[4991:4984]) ? 1 : 0;
assign detect_max[623][13] = (mid_1[4999:4992] > mid_1[5007:5000]) ? 1 : 0;
assign detect_max[623][14] = (mid_1[4999:4992] > mid_2[4991:4984]) ? 1 : 0;
assign detect_max[623][15] = (mid_1[4999:4992] > mid_2[4999:4992]) ? 1 : 0;
assign detect_max[623][16] = (mid_1[4999:4992] > mid_2[5007:5000]) ? 1 : 0;
assign detect_max[623][17] = (mid_1[4999:4992] > btm_0[4991:4984]) ? 1 : 0;
assign detect_max[623][18] = (mid_1[4999:4992] > btm_0[4999:4992]) ? 1 : 0;
assign detect_max[623][19] = (mid_1[4999:4992] > btm_0[5007:5000]) ? 1 : 0;
assign detect_max[623][20] = (mid_1[4999:4992] > btm_1[4991:4984]) ? 1 : 0;
assign detect_max[623][21] = (mid_1[4999:4992] > btm_1[4999:4992]) ? 1 : 0;
assign detect_max[623][22] = (mid_1[4999:4992] > btm_1[5007:5000]) ? 1 : 0;
assign detect_max[623][23] = (mid_1[4999:4992] > btm_2[4991:4984]) ? 1 : 0;
assign detect_max[623][24] = (mid_1[4999:4992] > btm_2[4999:4992]) ? 1 : 0;
assign detect_max[623][25] = (mid_1[4999:4992] > btm_2[5007:5000]) ? 1 : 0;

assign detect_max[624][0] = (mid_1[5007:5000] > top_0[4999:4992]) ? 1 : 0;
assign detect_max[624][1] = (mid_1[5007:5000] > top_0[5007:5000]) ? 1 : 0;
assign detect_max[624][2] = (mid_1[5007:5000] > top_0[5015:5008]) ? 1 : 0;
assign detect_max[624][3] = (mid_1[5007:5000] > top_1[4999:4992]) ? 1 : 0;
assign detect_max[624][4] = (mid_1[5007:5000] > top_1[5007:5000]) ? 1 : 0;
assign detect_max[624][5] = (mid_1[5007:5000] > top_1[5015:5008]) ? 1 : 0;
assign detect_max[624][6] = (mid_1[5007:5000] > top_2[4999:4992]) ? 1 : 0;
assign detect_max[624][7] = (mid_1[5007:5000] > top_2[5007:5000]) ? 1 : 0;
assign detect_max[624][8] = (mid_1[5007:5000] > top_2[5015:5008]) ? 1 : 0;
assign detect_max[624][9] = (mid_1[5007:5000] > mid_0[4999:4992]) ? 1 : 0;
assign detect_max[624][10] = (mid_1[5007:5000] > mid_0[5007:5000]) ? 1 : 0;
assign detect_max[624][11] = (mid_1[5007:5000] > mid_0[5015:5008]) ? 1 : 0;
assign detect_max[624][12] = (mid_1[5007:5000] > mid_1[4999:4992]) ? 1 : 0;
assign detect_max[624][13] = (mid_1[5007:5000] > mid_1[5015:5008]) ? 1 : 0;
assign detect_max[624][14] = (mid_1[5007:5000] > mid_2[4999:4992]) ? 1 : 0;
assign detect_max[624][15] = (mid_1[5007:5000] > mid_2[5007:5000]) ? 1 : 0;
assign detect_max[624][16] = (mid_1[5007:5000] > mid_2[5015:5008]) ? 1 : 0;
assign detect_max[624][17] = (mid_1[5007:5000] > btm_0[4999:4992]) ? 1 : 0;
assign detect_max[624][18] = (mid_1[5007:5000] > btm_0[5007:5000]) ? 1 : 0;
assign detect_max[624][19] = (mid_1[5007:5000] > btm_0[5015:5008]) ? 1 : 0;
assign detect_max[624][20] = (mid_1[5007:5000] > btm_1[4999:4992]) ? 1 : 0;
assign detect_max[624][21] = (mid_1[5007:5000] > btm_1[5007:5000]) ? 1 : 0;
assign detect_max[624][22] = (mid_1[5007:5000] > btm_1[5015:5008]) ? 1 : 0;
assign detect_max[624][23] = (mid_1[5007:5000] > btm_2[4999:4992]) ? 1 : 0;
assign detect_max[624][24] = (mid_1[5007:5000] > btm_2[5007:5000]) ? 1 : 0;
assign detect_max[624][25] = (mid_1[5007:5000] > btm_2[5015:5008]) ? 1 : 0;

assign detect_max[625][0] = (mid_1[5015:5008] > top_0[5007:5000]) ? 1 : 0;
assign detect_max[625][1] = (mid_1[5015:5008] > top_0[5015:5008]) ? 1 : 0;
assign detect_max[625][2] = (mid_1[5015:5008] > top_0[5023:5016]) ? 1 : 0;
assign detect_max[625][3] = (mid_1[5015:5008] > top_1[5007:5000]) ? 1 : 0;
assign detect_max[625][4] = (mid_1[5015:5008] > top_1[5015:5008]) ? 1 : 0;
assign detect_max[625][5] = (mid_1[5015:5008] > top_1[5023:5016]) ? 1 : 0;
assign detect_max[625][6] = (mid_1[5015:5008] > top_2[5007:5000]) ? 1 : 0;
assign detect_max[625][7] = (mid_1[5015:5008] > top_2[5015:5008]) ? 1 : 0;
assign detect_max[625][8] = (mid_1[5015:5008] > top_2[5023:5016]) ? 1 : 0;
assign detect_max[625][9] = (mid_1[5015:5008] > mid_0[5007:5000]) ? 1 : 0;
assign detect_max[625][10] = (mid_1[5015:5008] > mid_0[5015:5008]) ? 1 : 0;
assign detect_max[625][11] = (mid_1[5015:5008] > mid_0[5023:5016]) ? 1 : 0;
assign detect_max[625][12] = (mid_1[5015:5008] > mid_1[5007:5000]) ? 1 : 0;
assign detect_max[625][13] = (mid_1[5015:5008] > mid_1[5023:5016]) ? 1 : 0;
assign detect_max[625][14] = (mid_1[5015:5008] > mid_2[5007:5000]) ? 1 : 0;
assign detect_max[625][15] = (mid_1[5015:5008] > mid_2[5015:5008]) ? 1 : 0;
assign detect_max[625][16] = (mid_1[5015:5008] > mid_2[5023:5016]) ? 1 : 0;
assign detect_max[625][17] = (mid_1[5015:5008] > btm_0[5007:5000]) ? 1 : 0;
assign detect_max[625][18] = (mid_1[5015:5008] > btm_0[5015:5008]) ? 1 : 0;
assign detect_max[625][19] = (mid_1[5015:5008] > btm_0[5023:5016]) ? 1 : 0;
assign detect_max[625][20] = (mid_1[5015:5008] > btm_1[5007:5000]) ? 1 : 0;
assign detect_max[625][21] = (mid_1[5015:5008] > btm_1[5015:5008]) ? 1 : 0;
assign detect_max[625][22] = (mid_1[5015:5008] > btm_1[5023:5016]) ? 1 : 0;
assign detect_max[625][23] = (mid_1[5015:5008] > btm_2[5007:5000]) ? 1 : 0;
assign detect_max[625][24] = (mid_1[5015:5008] > btm_2[5015:5008]) ? 1 : 0;
assign detect_max[625][25] = (mid_1[5015:5008] > btm_2[5023:5016]) ? 1 : 0;

assign detect_max[626][0] = (mid_1[5023:5016] > top_0[5015:5008]) ? 1 : 0;
assign detect_max[626][1] = (mid_1[5023:5016] > top_0[5023:5016]) ? 1 : 0;
assign detect_max[626][2] = (mid_1[5023:5016] > top_0[5031:5024]) ? 1 : 0;
assign detect_max[626][3] = (mid_1[5023:5016] > top_1[5015:5008]) ? 1 : 0;
assign detect_max[626][4] = (mid_1[5023:5016] > top_1[5023:5016]) ? 1 : 0;
assign detect_max[626][5] = (mid_1[5023:5016] > top_1[5031:5024]) ? 1 : 0;
assign detect_max[626][6] = (mid_1[5023:5016] > top_2[5015:5008]) ? 1 : 0;
assign detect_max[626][7] = (mid_1[5023:5016] > top_2[5023:5016]) ? 1 : 0;
assign detect_max[626][8] = (mid_1[5023:5016] > top_2[5031:5024]) ? 1 : 0;
assign detect_max[626][9] = (mid_1[5023:5016] > mid_0[5015:5008]) ? 1 : 0;
assign detect_max[626][10] = (mid_1[5023:5016] > mid_0[5023:5016]) ? 1 : 0;
assign detect_max[626][11] = (mid_1[5023:5016] > mid_0[5031:5024]) ? 1 : 0;
assign detect_max[626][12] = (mid_1[5023:5016] > mid_1[5015:5008]) ? 1 : 0;
assign detect_max[626][13] = (mid_1[5023:5016] > mid_1[5031:5024]) ? 1 : 0;
assign detect_max[626][14] = (mid_1[5023:5016] > mid_2[5015:5008]) ? 1 : 0;
assign detect_max[626][15] = (mid_1[5023:5016] > mid_2[5023:5016]) ? 1 : 0;
assign detect_max[626][16] = (mid_1[5023:5016] > mid_2[5031:5024]) ? 1 : 0;
assign detect_max[626][17] = (mid_1[5023:5016] > btm_0[5015:5008]) ? 1 : 0;
assign detect_max[626][18] = (mid_1[5023:5016] > btm_0[5023:5016]) ? 1 : 0;
assign detect_max[626][19] = (mid_1[5023:5016] > btm_0[5031:5024]) ? 1 : 0;
assign detect_max[626][20] = (mid_1[5023:5016] > btm_1[5015:5008]) ? 1 : 0;
assign detect_max[626][21] = (mid_1[5023:5016] > btm_1[5023:5016]) ? 1 : 0;
assign detect_max[626][22] = (mid_1[5023:5016] > btm_1[5031:5024]) ? 1 : 0;
assign detect_max[626][23] = (mid_1[5023:5016] > btm_2[5015:5008]) ? 1 : 0;
assign detect_max[626][24] = (mid_1[5023:5016] > btm_2[5023:5016]) ? 1 : 0;
assign detect_max[626][25] = (mid_1[5023:5016] > btm_2[5031:5024]) ? 1 : 0;

assign detect_max[627][0] = (mid_1[5031:5024] > top_0[5023:5016]) ? 1 : 0;
assign detect_max[627][1] = (mid_1[5031:5024] > top_0[5031:5024]) ? 1 : 0;
assign detect_max[627][2] = (mid_1[5031:5024] > top_0[5039:5032]) ? 1 : 0;
assign detect_max[627][3] = (mid_1[5031:5024] > top_1[5023:5016]) ? 1 : 0;
assign detect_max[627][4] = (mid_1[5031:5024] > top_1[5031:5024]) ? 1 : 0;
assign detect_max[627][5] = (mid_1[5031:5024] > top_1[5039:5032]) ? 1 : 0;
assign detect_max[627][6] = (mid_1[5031:5024] > top_2[5023:5016]) ? 1 : 0;
assign detect_max[627][7] = (mid_1[5031:5024] > top_2[5031:5024]) ? 1 : 0;
assign detect_max[627][8] = (mid_1[5031:5024] > top_2[5039:5032]) ? 1 : 0;
assign detect_max[627][9] = (mid_1[5031:5024] > mid_0[5023:5016]) ? 1 : 0;
assign detect_max[627][10] = (mid_1[5031:5024] > mid_0[5031:5024]) ? 1 : 0;
assign detect_max[627][11] = (mid_1[5031:5024] > mid_0[5039:5032]) ? 1 : 0;
assign detect_max[627][12] = (mid_1[5031:5024] > mid_1[5023:5016]) ? 1 : 0;
assign detect_max[627][13] = (mid_1[5031:5024] > mid_1[5039:5032]) ? 1 : 0;
assign detect_max[627][14] = (mid_1[5031:5024] > mid_2[5023:5016]) ? 1 : 0;
assign detect_max[627][15] = (mid_1[5031:5024] > mid_2[5031:5024]) ? 1 : 0;
assign detect_max[627][16] = (mid_1[5031:5024] > mid_2[5039:5032]) ? 1 : 0;
assign detect_max[627][17] = (mid_1[5031:5024] > btm_0[5023:5016]) ? 1 : 0;
assign detect_max[627][18] = (mid_1[5031:5024] > btm_0[5031:5024]) ? 1 : 0;
assign detect_max[627][19] = (mid_1[5031:5024] > btm_0[5039:5032]) ? 1 : 0;
assign detect_max[627][20] = (mid_1[5031:5024] > btm_1[5023:5016]) ? 1 : 0;
assign detect_max[627][21] = (mid_1[5031:5024] > btm_1[5031:5024]) ? 1 : 0;
assign detect_max[627][22] = (mid_1[5031:5024] > btm_1[5039:5032]) ? 1 : 0;
assign detect_max[627][23] = (mid_1[5031:5024] > btm_2[5023:5016]) ? 1 : 0;
assign detect_max[627][24] = (mid_1[5031:5024] > btm_2[5031:5024]) ? 1 : 0;
assign detect_max[627][25] = (mid_1[5031:5024] > btm_2[5039:5032]) ? 1 : 0;

assign detect_max[628][0] = (mid_1[5039:5032] > top_0[5031:5024]) ? 1 : 0;
assign detect_max[628][1] = (mid_1[5039:5032] > top_0[5039:5032]) ? 1 : 0;
assign detect_max[628][2] = (mid_1[5039:5032] > top_0[5047:5040]) ? 1 : 0;
assign detect_max[628][3] = (mid_1[5039:5032] > top_1[5031:5024]) ? 1 : 0;
assign detect_max[628][4] = (mid_1[5039:5032] > top_1[5039:5032]) ? 1 : 0;
assign detect_max[628][5] = (mid_1[5039:5032] > top_1[5047:5040]) ? 1 : 0;
assign detect_max[628][6] = (mid_1[5039:5032] > top_2[5031:5024]) ? 1 : 0;
assign detect_max[628][7] = (mid_1[5039:5032] > top_2[5039:5032]) ? 1 : 0;
assign detect_max[628][8] = (mid_1[5039:5032] > top_2[5047:5040]) ? 1 : 0;
assign detect_max[628][9] = (mid_1[5039:5032] > mid_0[5031:5024]) ? 1 : 0;
assign detect_max[628][10] = (mid_1[5039:5032] > mid_0[5039:5032]) ? 1 : 0;
assign detect_max[628][11] = (mid_1[5039:5032] > mid_0[5047:5040]) ? 1 : 0;
assign detect_max[628][12] = (mid_1[5039:5032] > mid_1[5031:5024]) ? 1 : 0;
assign detect_max[628][13] = (mid_1[5039:5032] > mid_1[5047:5040]) ? 1 : 0;
assign detect_max[628][14] = (mid_1[5039:5032] > mid_2[5031:5024]) ? 1 : 0;
assign detect_max[628][15] = (mid_1[5039:5032] > mid_2[5039:5032]) ? 1 : 0;
assign detect_max[628][16] = (mid_1[5039:5032] > mid_2[5047:5040]) ? 1 : 0;
assign detect_max[628][17] = (mid_1[5039:5032] > btm_0[5031:5024]) ? 1 : 0;
assign detect_max[628][18] = (mid_1[5039:5032] > btm_0[5039:5032]) ? 1 : 0;
assign detect_max[628][19] = (mid_1[5039:5032] > btm_0[5047:5040]) ? 1 : 0;
assign detect_max[628][20] = (mid_1[5039:5032] > btm_1[5031:5024]) ? 1 : 0;
assign detect_max[628][21] = (mid_1[5039:5032] > btm_1[5039:5032]) ? 1 : 0;
assign detect_max[628][22] = (mid_1[5039:5032] > btm_1[5047:5040]) ? 1 : 0;
assign detect_max[628][23] = (mid_1[5039:5032] > btm_2[5031:5024]) ? 1 : 0;
assign detect_max[628][24] = (mid_1[5039:5032] > btm_2[5039:5032]) ? 1 : 0;
assign detect_max[628][25] = (mid_1[5039:5032] > btm_2[5047:5040]) ? 1 : 0;

assign detect_max[629][0] = (mid_1[5047:5040] > top_0[5039:5032]) ? 1 : 0;
assign detect_max[629][1] = (mid_1[5047:5040] > top_0[5047:5040]) ? 1 : 0;
assign detect_max[629][2] = (mid_1[5047:5040] > top_0[5055:5048]) ? 1 : 0;
assign detect_max[629][3] = (mid_1[5047:5040] > top_1[5039:5032]) ? 1 : 0;
assign detect_max[629][4] = (mid_1[5047:5040] > top_1[5047:5040]) ? 1 : 0;
assign detect_max[629][5] = (mid_1[5047:5040] > top_1[5055:5048]) ? 1 : 0;
assign detect_max[629][6] = (mid_1[5047:5040] > top_2[5039:5032]) ? 1 : 0;
assign detect_max[629][7] = (mid_1[5047:5040] > top_2[5047:5040]) ? 1 : 0;
assign detect_max[629][8] = (mid_1[5047:5040] > top_2[5055:5048]) ? 1 : 0;
assign detect_max[629][9] = (mid_1[5047:5040] > mid_0[5039:5032]) ? 1 : 0;
assign detect_max[629][10] = (mid_1[5047:5040] > mid_0[5047:5040]) ? 1 : 0;
assign detect_max[629][11] = (mid_1[5047:5040] > mid_0[5055:5048]) ? 1 : 0;
assign detect_max[629][12] = (mid_1[5047:5040] > mid_1[5039:5032]) ? 1 : 0;
assign detect_max[629][13] = (mid_1[5047:5040] > mid_1[5055:5048]) ? 1 : 0;
assign detect_max[629][14] = (mid_1[5047:5040] > mid_2[5039:5032]) ? 1 : 0;
assign detect_max[629][15] = (mid_1[5047:5040] > mid_2[5047:5040]) ? 1 : 0;
assign detect_max[629][16] = (mid_1[5047:5040] > mid_2[5055:5048]) ? 1 : 0;
assign detect_max[629][17] = (mid_1[5047:5040] > btm_0[5039:5032]) ? 1 : 0;
assign detect_max[629][18] = (mid_1[5047:5040] > btm_0[5047:5040]) ? 1 : 0;
assign detect_max[629][19] = (mid_1[5047:5040] > btm_0[5055:5048]) ? 1 : 0;
assign detect_max[629][20] = (mid_1[5047:5040] > btm_1[5039:5032]) ? 1 : 0;
assign detect_max[629][21] = (mid_1[5047:5040] > btm_1[5047:5040]) ? 1 : 0;
assign detect_max[629][22] = (mid_1[5047:5040] > btm_1[5055:5048]) ? 1 : 0;
assign detect_max[629][23] = (mid_1[5047:5040] > btm_2[5039:5032]) ? 1 : 0;
assign detect_max[629][24] = (mid_1[5047:5040] > btm_2[5047:5040]) ? 1 : 0;
assign detect_max[629][25] = (mid_1[5047:5040] > btm_2[5055:5048]) ? 1 : 0;

assign detect_max[630][0] = (mid_1[5055:5048] > top_0[5047:5040]) ? 1 : 0;
assign detect_max[630][1] = (mid_1[5055:5048] > top_0[5055:5048]) ? 1 : 0;
assign detect_max[630][2] = (mid_1[5055:5048] > top_0[5063:5056]) ? 1 : 0;
assign detect_max[630][3] = (mid_1[5055:5048] > top_1[5047:5040]) ? 1 : 0;
assign detect_max[630][4] = (mid_1[5055:5048] > top_1[5055:5048]) ? 1 : 0;
assign detect_max[630][5] = (mid_1[5055:5048] > top_1[5063:5056]) ? 1 : 0;
assign detect_max[630][6] = (mid_1[5055:5048] > top_2[5047:5040]) ? 1 : 0;
assign detect_max[630][7] = (mid_1[5055:5048] > top_2[5055:5048]) ? 1 : 0;
assign detect_max[630][8] = (mid_1[5055:5048] > top_2[5063:5056]) ? 1 : 0;
assign detect_max[630][9] = (mid_1[5055:5048] > mid_0[5047:5040]) ? 1 : 0;
assign detect_max[630][10] = (mid_1[5055:5048] > mid_0[5055:5048]) ? 1 : 0;
assign detect_max[630][11] = (mid_1[5055:5048] > mid_0[5063:5056]) ? 1 : 0;
assign detect_max[630][12] = (mid_1[5055:5048] > mid_1[5047:5040]) ? 1 : 0;
assign detect_max[630][13] = (mid_1[5055:5048] > mid_1[5063:5056]) ? 1 : 0;
assign detect_max[630][14] = (mid_1[5055:5048] > mid_2[5047:5040]) ? 1 : 0;
assign detect_max[630][15] = (mid_1[5055:5048] > mid_2[5055:5048]) ? 1 : 0;
assign detect_max[630][16] = (mid_1[5055:5048] > mid_2[5063:5056]) ? 1 : 0;
assign detect_max[630][17] = (mid_1[5055:5048] > btm_0[5047:5040]) ? 1 : 0;
assign detect_max[630][18] = (mid_1[5055:5048] > btm_0[5055:5048]) ? 1 : 0;
assign detect_max[630][19] = (mid_1[5055:5048] > btm_0[5063:5056]) ? 1 : 0;
assign detect_max[630][20] = (mid_1[5055:5048] > btm_1[5047:5040]) ? 1 : 0;
assign detect_max[630][21] = (mid_1[5055:5048] > btm_1[5055:5048]) ? 1 : 0;
assign detect_max[630][22] = (mid_1[5055:5048] > btm_1[5063:5056]) ? 1 : 0;
assign detect_max[630][23] = (mid_1[5055:5048] > btm_2[5047:5040]) ? 1 : 0;
assign detect_max[630][24] = (mid_1[5055:5048] > btm_2[5055:5048]) ? 1 : 0;
assign detect_max[630][25] = (mid_1[5055:5048] > btm_2[5063:5056]) ? 1 : 0;

assign detect_max[631][0] = (mid_1[5063:5056] > top_0[5055:5048]) ? 1 : 0;
assign detect_max[631][1] = (mid_1[5063:5056] > top_0[5063:5056]) ? 1 : 0;
assign detect_max[631][2] = (mid_1[5063:5056] > top_0[5071:5064]) ? 1 : 0;
assign detect_max[631][3] = (mid_1[5063:5056] > top_1[5055:5048]) ? 1 : 0;
assign detect_max[631][4] = (mid_1[5063:5056] > top_1[5063:5056]) ? 1 : 0;
assign detect_max[631][5] = (mid_1[5063:5056] > top_1[5071:5064]) ? 1 : 0;
assign detect_max[631][6] = (mid_1[5063:5056] > top_2[5055:5048]) ? 1 : 0;
assign detect_max[631][7] = (mid_1[5063:5056] > top_2[5063:5056]) ? 1 : 0;
assign detect_max[631][8] = (mid_1[5063:5056] > top_2[5071:5064]) ? 1 : 0;
assign detect_max[631][9] = (mid_1[5063:5056] > mid_0[5055:5048]) ? 1 : 0;
assign detect_max[631][10] = (mid_1[5063:5056] > mid_0[5063:5056]) ? 1 : 0;
assign detect_max[631][11] = (mid_1[5063:5056] > mid_0[5071:5064]) ? 1 : 0;
assign detect_max[631][12] = (mid_1[5063:5056] > mid_1[5055:5048]) ? 1 : 0;
assign detect_max[631][13] = (mid_1[5063:5056] > mid_1[5071:5064]) ? 1 : 0;
assign detect_max[631][14] = (mid_1[5063:5056] > mid_2[5055:5048]) ? 1 : 0;
assign detect_max[631][15] = (mid_1[5063:5056] > mid_2[5063:5056]) ? 1 : 0;
assign detect_max[631][16] = (mid_1[5063:5056] > mid_2[5071:5064]) ? 1 : 0;
assign detect_max[631][17] = (mid_1[5063:5056] > btm_0[5055:5048]) ? 1 : 0;
assign detect_max[631][18] = (mid_1[5063:5056] > btm_0[5063:5056]) ? 1 : 0;
assign detect_max[631][19] = (mid_1[5063:5056] > btm_0[5071:5064]) ? 1 : 0;
assign detect_max[631][20] = (mid_1[5063:5056] > btm_1[5055:5048]) ? 1 : 0;
assign detect_max[631][21] = (mid_1[5063:5056] > btm_1[5063:5056]) ? 1 : 0;
assign detect_max[631][22] = (mid_1[5063:5056] > btm_1[5071:5064]) ? 1 : 0;
assign detect_max[631][23] = (mid_1[5063:5056] > btm_2[5055:5048]) ? 1 : 0;
assign detect_max[631][24] = (mid_1[5063:5056] > btm_2[5063:5056]) ? 1 : 0;
assign detect_max[631][25] = (mid_1[5063:5056] > btm_2[5071:5064]) ? 1 : 0;

assign detect_max[632][0] = (mid_1[5071:5064] > top_0[5063:5056]) ? 1 : 0;
assign detect_max[632][1] = (mid_1[5071:5064] > top_0[5071:5064]) ? 1 : 0;
assign detect_max[632][2] = (mid_1[5071:5064] > top_0[5079:5072]) ? 1 : 0;
assign detect_max[632][3] = (mid_1[5071:5064] > top_1[5063:5056]) ? 1 : 0;
assign detect_max[632][4] = (mid_1[5071:5064] > top_1[5071:5064]) ? 1 : 0;
assign detect_max[632][5] = (mid_1[5071:5064] > top_1[5079:5072]) ? 1 : 0;
assign detect_max[632][6] = (mid_1[5071:5064] > top_2[5063:5056]) ? 1 : 0;
assign detect_max[632][7] = (mid_1[5071:5064] > top_2[5071:5064]) ? 1 : 0;
assign detect_max[632][8] = (mid_1[5071:5064] > top_2[5079:5072]) ? 1 : 0;
assign detect_max[632][9] = (mid_1[5071:5064] > mid_0[5063:5056]) ? 1 : 0;
assign detect_max[632][10] = (mid_1[5071:5064] > mid_0[5071:5064]) ? 1 : 0;
assign detect_max[632][11] = (mid_1[5071:5064] > mid_0[5079:5072]) ? 1 : 0;
assign detect_max[632][12] = (mid_1[5071:5064] > mid_1[5063:5056]) ? 1 : 0;
assign detect_max[632][13] = (mid_1[5071:5064] > mid_1[5079:5072]) ? 1 : 0;
assign detect_max[632][14] = (mid_1[5071:5064] > mid_2[5063:5056]) ? 1 : 0;
assign detect_max[632][15] = (mid_1[5071:5064] > mid_2[5071:5064]) ? 1 : 0;
assign detect_max[632][16] = (mid_1[5071:5064] > mid_2[5079:5072]) ? 1 : 0;
assign detect_max[632][17] = (mid_1[5071:5064] > btm_0[5063:5056]) ? 1 : 0;
assign detect_max[632][18] = (mid_1[5071:5064] > btm_0[5071:5064]) ? 1 : 0;
assign detect_max[632][19] = (mid_1[5071:5064] > btm_0[5079:5072]) ? 1 : 0;
assign detect_max[632][20] = (mid_1[5071:5064] > btm_1[5063:5056]) ? 1 : 0;
assign detect_max[632][21] = (mid_1[5071:5064] > btm_1[5071:5064]) ? 1 : 0;
assign detect_max[632][22] = (mid_1[5071:5064] > btm_1[5079:5072]) ? 1 : 0;
assign detect_max[632][23] = (mid_1[5071:5064] > btm_2[5063:5056]) ? 1 : 0;
assign detect_max[632][24] = (mid_1[5071:5064] > btm_2[5071:5064]) ? 1 : 0;
assign detect_max[632][25] = (mid_1[5071:5064] > btm_2[5079:5072]) ? 1 : 0;

assign detect_max[633][0] = (mid_1[5079:5072] > top_0[5071:5064]) ? 1 : 0;
assign detect_max[633][1] = (mid_1[5079:5072] > top_0[5079:5072]) ? 1 : 0;
assign detect_max[633][2] = (mid_1[5079:5072] > top_0[5087:5080]) ? 1 : 0;
assign detect_max[633][3] = (mid_1[5079:5072] > top_1[5071:5064]) ? 1 : 0;
assign detect_max[633][4] = (mid_1[5079:5072] > top_1[5079:5072]) ? 1 : 0;
assign detect_max[633][5] = (mid_1[5079:5072] > top_1[5087:5080]) ? 1 : 0;
assign detect_max[633][6] = (mid_1[5079:5072] > top_2[5071:5064]) ? 1 : 0;
assign detect_max[633][7] = (mid_1[5079:5072] > top_2[5079:5072]) ? 1 : 0;
assign detect_max[633][8] = (mid_1[5079:5072] > top_2[5087:5080]) ? 1 : 0;
assign detect_max[633][9] = (mid_1[5079:5072] > mid_0[5071:5064]) ? 1 : 0;
assign detect_max[633][10] = (mid_1[5079:5072] > mid_0[5079:5072]) ? 1 : 0;
assign detect_max[633][11] = (mid_1[5079:5072] > mid_0[5087:5080]) ? 1 : 0;
assign detect_max[633][12] = (mid_1[5079:5072] > mid_1[5071:5064]) ? 1 : 0;
assign detect_max[633][13] = (mid_1[5079:5072] > mid_1[5087:5080]) ? 1 : 0;
assign detect_max[633][14] = (mid_1[5079:5072] > mid_2[5071:5064]) ? 1 : 0;
assign detect_max[633][15] = (mid_1[5079:5072] > mid_2[5079:5072]) ? 1 : 0;
assign detect_max[633][16] = (mid_1[5079:5072] > mid_2[5087:5080]) ? 1 : 0;
assign detect_max[633][17] = (mid_1[5079:5072] > btm_0[5071:5064]) ? 1 : 0;
assign detect_max[633][18] = (mid_1[5079:5072] > btm_0[5079:5072]) ? 1 : 0;
assign detect_max[633][19] = (mid_1[5079:5072] > btm_0[5087:5080]) ? 1 : 0;
assign detect_max[633][20] = (mid_1[5079:5072] > btm_1[5071:5064]) ? 1 : 0;
assign detect_max[633][21] = (mid_1[5079:5072] > btm_1[5079:5072]) ? 1 : 0;
assign detect_max[633][22] = (mid_1[5079:5072] > btm_1[5087:5080]) ? 1 : 0;
assign detect_max[633][23] = (mid_1[5079:5072] > btm_2[5071:5064]) ? 1 : 0;
assign detect_max[633][24] = (mid_1[5079:5072] > btm_2[5079:5072]) ? 1 : 0;
assign detect_max[633][25] = (mid_1[5079:5072] > btm_2[5087:5080]) ? 1 : 0;

assign detect_max[634][0] = (mid_1[5087:5080] > top_0[5079:5072]) ? 1 : 0;
assign detect_max[634][1] = (mid_1[5087:5080] > top_0[5087:5080]) ? 1 : 0;
assign detect_max[634][2] = (mid_1[5087:5080] > top_0[5095:5088]) ? 1 : 0;
assign detect_max[634][3] = (mid_1[5087:5080] > top_1[5079:5072]) ? 1 : 0;
assign detect_max[634][4] = (mid_1[5087:5080] > top_1[5087:5080]) ? 1 : 0;
assign detect_max[634][5] = (mid_1[5087:5080] > top_1[5095:5088]) ? 1 : 0;
assign detect_max[634][6] = (mid_1[5087:5080] > top_2[5079:5072]) ? 1 : 0;
assign detect_max[634][7] = (mid_1[5087:5080] > top_2[5087:5080]) ? 1 : 0;
assign detect_max[634][8] = (mid_1[5087:5080] > top_2[5095:5088]) ? 1 : 0;
assign detect_max[634][9] = (mid_1[5087:5080] > mid_0[5079:5072]) ? 1 : 0;
assign detect_max[634][10] = (mid_1[5087:5080] > mid_0[5087:5080]) ? 1 : 0;
assign detect_max[634][11] = (mid_1[5087:5080] > mid_0[5095:5088]) ? 1 : 0;
assign detect_max[634][12] = (mid_1[5087:5080] > mid_1[5079:5072]) ? 1 : 0;
assign detect_max[634][13] = (mid_1[5087:5080] > mid_1[5095:5088]) ? 1 : 0;
assign detect_max[634][14] = (mid_1[5087:5080] > mid_2[5079:5072]) ? 1 : 0;
assign detect_max[634][15] = (mid_1[5087:5080] > mid_2[5087:5080]) ? 1 : 0;
assign detect_max[634][16] = (mid_1[5087:5080] > mid_2[5095:5088]) ? 1 : 0;
assign detect_max[634][17] = (mid_1[5087:5080] > btm_0[5079:5072]) ? 1 : 0;
assign detect_max[634][18] = (mid_1[5087:5080] > btm_0[5087:5080]) ? 1 : 0;
assign detect_max[634][19] = (mid_1[5087:5080] > btm_0[5095:5088]) ? 1 : 0;
assign detect_max[634][20] = (mid_1[5087:5080] > btm_1[5079:5072]) ? 1 : 0;
assign detect_max[634][21] = (mid_1[5087:5080] > btm_1[5087:5080]) ? 1 : 0;
assign detect_max[634][22] = (mid_1[5087:5080] > btm_1[5095:5088]) ? 1 : 0;
assign detect_max[634][23] = (mid_1[5087:5080] > btm_2[5079:5072]) ? 1 : 0;
assign detect_max[634][24] = (mid_1[5087:5080] > btm_2[5087:5080]) ? 1 : 0;
assign detect_max[634][25] = (mid_1[5087:5080] > btm_2[5095:5088]) ? 1 : 0;

assign detect_max[635][0] = (mid_1[5095:5088] > top_0[5087:5080]) ? 1 : 0;
assign detect_max[635][1] = (mid_1[5095:5088] > top_0[5095:5088]) ? 1 : 0;
assign detect_max[635][2] = (mid_1[5095:5088] > top_0[5103:5096]) ? 1 : 0;
assign detect_max[635][3] = (mid_1[5095:5088] > top_1[5087:5080]) ? 1 : 0;
assign detect_max[635][4] = (mid_1[5095:5088] > top_1[5095:5088]) ? 1 : 0;
assign detect_max[635][5] = (mid_1[5095:5088] > top_1[5103:5096]) ? 1 : 0;
assign detect_max[635][6] = (mid_1[5095:5088] > top_2[5087:5080]) ? 1 : 0;
assign detect_max[635][7] = (mid_1[5095:5088] > top_2[5095:5088]) ? 1 : 0;
assign detect_max[635][8] = (mid_1[5095:5088] > top_2[5103:5096]) ? 1 : 0;
assign detect_max[635][9] = (mid_1[5095:5088] > mid_0[5087:5080]) ? 1 : 0;
assign detect_max[635][10] = (mid_1[5095:5088] > mid_0[5095:5088]) ? 1 : 0;
assign detect_max[635][11] = (mid_1[5095:5088] > mid_0[5103:5096]) ? 1 : 0;
assign detect_max[635][12] = (mid_1[5095:5088] > mid_1[5087:5080]) ? 1 : 0;
assign detect_max[635][13] = (mid_1[5095:5088] > mid_1[5103:5096]) ? 1 : 0;
assign detect_max[635][14] = (mid_1[5095:5088] > mid_2[5087:5080]) ? 1 : 0;
assign detect_max[635][15] = (mid_1[5095:5088] > mid_2[5095:5088]) ? 1 : 0;
assign detect_max[635][16] = (mid_1[5095:5088] > mid_2[5103:5096]) ? 1 : 0;
assign detect_max[635][17] = (mid_1[5095:5088] > btm_0[5087:5080]) ? 1 : 0;
assign detect_max[635][18] = (mid_1[5095:5088] > btm_0[5095:5088]) ? 1 : 0;
assign detect_max[635][19] = (mid_1[5095:5088] > btm_0[5103:5096]) ? 1 : 0;
assign detect_max[635][20] = (mid_1[5095:5088] > btm_1[5087:5080]) ? 1 : 0;
assign detect_max[635][21] = (mid_1[5095:5088] > btm_1[5095:5088]) ? 1 : 0;
assign detect_max[635][22] = (mid_1[5095:5088] > btm_1[5103:5096]) ? 1 : 0;
assign detect_max[635][23] = (mid_1[5095:5088] > btm_2[5087:5080]) ? 1 : 0;
assign detect_max[635][24] = (mid_1[5095:5088] > btm_2[5095:5088]) ? 1 : 0;
assign detect_max[635][25] = (mid_1[5095:5088] > btm_2[5103:5096]) ? 1 : 0;

assign detect_max[636][0] = (mid_1[5103:5096] > top_0[5095:5088]) ? 1 : 0;
assign detect_max[636][1] = (mid_1[5103:5096] > top_0[5103:5096]) ? 1 : 0;
assign detect_max[636][2] = (mid_1[5103:5096] > top_0[5111:5104]) ? 1 : 0;
assign detect_max[636][3] = (mid_1[5103:5096] > top_1[5095:5088]) ? 1 : 0;
assign detect_max[636][4] = (mid_1[5103:5096] > top_1[5103:5096]) ? 1 : 0;
assign detect_max[636][5] = (mid_1[5103:5096] > top_1[5111:5104]) ? 1 : 0;
assign detect_max[636][6] = (mid_1[5103:5096] > top_2[5095:5088]) ? 1 : 0;
assign detect_max[636][7] = (mid_1[5103:5096] > top_2[5103:5096]) ? 1 : 0;
assign detect_max[636][8] = (mid_1[5103:5096] > top_2[5111:5104]) ? 1 : 0;
assign detect_max[636][9] = (mid_1[5103:5096] > mid_0[5095:5088]) ? 1 : 0;
assign detect_max[636][10] = (mid_1[5103:5096] > mid_0[5103:5096]) ? 1 : 0;
assign detect_max[636][11] = (mid_1[5103:5096] > mid_0[5111:5104]) ? 1 : 0;
assign detect_max[636][12] = (mid_1[5103:5096] > mid_1[5095:5088]) ? 1 : 0;
assign detect_max[636][13] = (mid_1[5103:5096] > mid_1[5111:5104]) ? 1 : 0;
assign detect_max[636][14] = (mid_1[5103:5096] > mid_2[5095:5088]) ? 1 : 0;
assign detect_max[636][15] = (mid_1[5103:5096] > mid_2[5103:5096]) ? 1 : 0;
assign detect_max[636][16] = (mid_1[5103:5096] > mid_2[5111:5104]) ? 1 : 0;
assign detect_max[636][17] = (mid_1[5103:5096] > btm_0[5095:5088]) ? 1 : 0;
assign detect_max[636][18] = (mid_1[5103:5096] > btm_0[5103:5096]) ? 1 : 0;
assign detect_max[636][19] = (mid_1[5103:5096] > btm_0[5111:5104]) ? 1 : 0;
assign detect_max[636][20] = (mid_1[5103:5096] > btm_1[5095:5088]) ? 1 : 0;
assign detect_max[636][21] = (mid_1[5103:5096] > btm_1[5103:5096]) ? 1 : 0;
assign detect_max[636][22] = (mid_1[5103:5096] > btm_1[5111:5104]) ? 1 : 0;
assign detect_max[636][23] = (mid_1[5103:5096] > btm_2[5095:5088]) ? 1 : 0;
assign detect_max[636][24] = (mid_1[5103:5096] > btm_2[5103:5096]) ? 1 : 0;
assign detect_max[636][25] = (mid_1[5103:5096] > btm_2[5111:5104]) ? 1 : 0;

assign detect_max[637][0] = (mid_1[5111:5104] > top_0[5103:5096]) ? 1 : 0;
assign detect_max[637][1] = (mid_1[5111:5104] > top_0[5111:5104]) ? 1 : 0;
assign detect_max[637][2] = (mid_1[5111:5104] > top_0[5119:5112]) ? 1 : 0;
assign detect_max[637][3] = (mid_1[5111:5104] > top_1[5103:5096]) ? 1 : 0;
assign detect_max[637][4] = (mid_1[5111:5104] > top_1[5111:5104]) ? 1 : 0;
assign detect_max[637][5] = (mid_1[5111:5104] > top_1[5119:5112]) ? 1 : 0;
assign detect_max[637][6] = (mid_1[5111:5104] > top_2[5103:5096]) ? 1 : 0;
assign detect_max[637][7] = (mid_1[5111:5104] > top_2[5111:5104]) ? 1 : 0;
assign detect_max[637][8] = (mid_1[5111:5104] > top_2[5119:5112]) ? 1 : 0;
assign detect_max[637][9] = (mid_1[5111:5104] > mid_0[5103:5096]) ? 1 : 0;
assign detect_max[637][10] = (mid_1[5111:5104] > mid_0[5111:5104]) ? 1 : 0;
assign detect_max[637][11] = (mid_1[5111:5104] > mid_0[5119:5112]) ? 1 : 0;
assign detect_max[637][12] = (mid_1[5111:5104] > mid_1[5103:5096]) ? 1 : 0;
assign detect_max[637][13] = (mid_1[5111:5104] > mid_1[5119:5112]) ? 1 : 0;
assign detect_max[637][14] = (mid_1[5111:5104] > mid_2[5103:5096]) ? 1 : 0;
assign detect_max[637][15] = (mid_1[5111:5104] > mid_2[5111:5104]) ? 1 : 0;
assign detect_max[637][16] = (mid_1[5111:5104] > mid_2[5119:5112]) ? 1 : 0;
assign detect_max[637][17] = (mid_1[5111:5104] > btm_0[5103:5096]) ? 1 : 0;
assign detect_max[637][18] = (mid_1[5111:5104] > btm_0[5111:5104]) ? 1 : 0;
assign detect_max[637][19] = (mid_1[5111:5104] > btm_0[5119:5112]) ? 1 : 0;
assign detect_max[637][20] = (mid_1[5111:5104] > btm_1[5103:5096]) ? 1 : 0;
assign detect_max[637][21] = (mid_1[5111:5104] > btm_1[5111:5104]) ? 1 : 0;
assign detect_max[637][22] = (mid_1[5111:5104] > btm_1[5119:5112]) ? 1 : 0;
assign detect_max[637][23] = (mid_1[5111:5104] > btm_2[5103:5096]) ? 1 : 0;
assign detect_max[637][24] = (mid_1[5111:5104] > btm_2[5111:5104]) ? 1 : 0;
assign detect_max[637][25] = (mid_1[5111:5104] > btm_2[5119:5112]) ? 1 : 0;

wire [637:0] is_max;
assign is_max[0] = (&detect_max[0]) ? 1:0;
assign is_max[1] = (&detect_max[1]) ? 1:0;
assign is_max[2] = (&detect_max[2]) ? 1:0;
assign is_max[3] = (&detect_max[3]) ? 1:0;
assign is_max[4] = (&detect_max[4]) ? 1:0;
assign is_max[5] = (&detect_max[5]) ? 1:0;
assign is_max[6] = (&detect_max[6]) ? 1:0;
assign is_max[7] = (&detect_max[7]) ? 1:0;
assign is_max[8] = (&detect_max[8]) ? 1:0;
assign is_max[9] = (&detect_max[9]) ? 1:0;
assign is_max[10] = (&detect_max[10]) ? 1:0;
assign is_max[11] = (&detect_max[11]) ? 1:0;
assign is_max[12] = (&detect_max[12]) ? 1:0;
assign is_max[13] = (&detect_max[13]) ? 1:0;
assign is_max[14] = (&detect_max[14]) ? 1:0;
assign is_max[15] = (&detect_max[15]) ? 1:0;
assign is_max[16] = (&detect_max[16]) ? 1:0;
assign is_max[17] = (&detect_max[17]) ? 1:0;
assign is_max[18] = (&detect_max[18]) ? 1:0;
assign is_max[19] = (&detect_max[19]) ? 1:0;
assign is_max[20] = (&detect_max[20]) ? 1:0;
assign is_max[21] = (&detect_max[21]) ? 1:0;
assign is_max[22] = (&detect_max[22]) ? 1:0;
assign is_max[23] = (&detect_max[23]) ? 1:0;
assign is_max[24] = (&detect_max[24]) ? 1:0;
assign is_max[25] = (&detect_max[25]) ? 1:0;
assign is_max[26] = (&detect_max[26]) ? 1:0;
assign is_max[27] = (&detect_max[27]) ? 1:0;
assign is_max[28] = (&detect_max[28]) ? 1:0;
assign is_max[29] = (&detect_max[29]) ? 1:0;
assign is_max[30] = (&detect_max[30]) ? 1:0;
assign is_max[31] = (&detect_max[31]) ? 1:0;
assign is_max[32] = (&detect_max[32]) ? 1:0;
assign is_max[33] = (&detect_max[33]) ? 1:0;
assign is_max[34] = (&detect_max[34]) ? 1:0;
assign is_max[35] = (&detect_max[35]) ? 1:0;
assign is_max[36] = (&detect_max[36]) ? 1:0;
assign is_max[37] = (&detect_max[37]) ? 1:0;
assign is_max[38] = (&detect_max[38]) ? 1:0;
assign is_max[39] = (&detect_max[39]) ? 1:0;
assign is_max[40] = (&detect_max[40]) ? 1:0;
assign is_max[41] = (&detect_max[41]) ? 1:0;
assign is_max[42] = (&detect_max[42]) ? 1:0;
assign is_max[43] = (&detect_max[43]) ? 1:0;
assign is_max[44] = (&detect_max[44]) ? 1:0;
assign is_max[45] = (&detect_max[45]) ? 1:0;
assign is_max[46] = (&detect_max[46]) ? 1:0;
assign is_max[47] = (&detect_max[47]) ? 1:0;
assign is_max[48] = (&detect_max[48]) ? 1:0;
assign is_max[49] = (&detect_max[49]) ? 1:0;
assign is_max[50] = (&detect_max[50]) ? 1:0;
assign is_max[51] = (&detect_max[51]) ? 1:0;
assign is_max[52] = (&detect_max[52]) ? 1:0;
assign is_max[53] = (&detect_max[53]) ? 1:0;
assign is_max[54] = (&detect_max[54]) ? 1:0;
assign is_max[55] = (&detect_max[55]) ? 1:0;
assign is_max[56] = (&detect_max[56]) ? 1:0;
assign is_max[57] = (&detect_max[57]) ? 1:0;
assign is_max[58] = (&detect_max[58]) ? 1:0;
assign is_max[59] = (&detect_max[59]) ? 1:0;
assign is_max[60] = (&detect_max[60]) ? 1:0;
assign is_max[61] = (&detect_max[61]) ? 1:0;
assign is_max[62] = (&detect_max[62]) ? 1:0;
assign is_max[63] = (&detect_max[63]) ? 1:0;
assign is_max[64] = (&detect_max[64]) ? 1:0;
assign is_max[65] = (&detect_max[65]) ? 1:0;
assign is_max[66] = (&detect_max[66]) ? 1:0;
assign is_max[67] = (&detect_max[67]) ? 1:0;
assign is_max[68] = (&detect_max[68]) ? 1:0;
assign is_max[69] = (&detect_max[69]) ? 1:0;
assign is_max[70] = (&detect_max[70]) ? 1:0;
assign is_max[71] = (&detect_max[71]) ? 1:0;
assign is_max[72] = (&detect_max[72]) ? 1:0;
assign is_max[73] = (&detect_max[73]) ? 1:0;
assign is_max[74] = (&detect_max[74]) ? 1:0;
assign is_max[75] = (&detect_max[75]) ? 1:0;
assign is_max[76] = (&detect_max[76]) ? 1:0;
assign is_max[77] = (&detect_max[77]) ? 1:0;
assign is_max[78] = (&detect_max[78]) ? 1:0;
assign is_max[79] = (&detect_max[79]) ? 1:0;
assign is_max[80] = (&detect_max[80]) ? 1:0;
assign is_max[81] = (&detect_max[81]) ? 1:0;
assign is_max[82] = (&detect_max[82]) ? 1:0;
assign is_max[83] = (&detect_max[83]) ? 1:0;
assign is_max[84] = (&detect_max[84]) ? 1:0;
assign is_max[85] = (&detect_max[85]) ? 1:0;
assign is_max[86] = (&detect_max[86]) ? 1:0;
assign is_max[87] = (&detect_max[87]) ? 1:0;
assign is_max[88] = (&detect_max[88]) ? 1:0;
assign is_max[89] = (&detect_max[89]) ? 1:0;
assign is_max[90] = (&detect_max[90]) ? 1:0;
assign is_max[91] = (&detect_max[91]) ? 1:0;
assign is_max[92] = (&detect_max[92]) ? 1:0;
assign is_max[93] = (&detect_max[93]) ? 1:0;
assign is_max[94] = (&detect_max[94]) ? 1:0;
assign is_max[95] = (&detect_max[95]) ? 1:0;
assign is_max[96] = (&detect_max[96]) ? 1:0;
assign is_max[97] = (&detect_max[97]) ? 1:0;
assign is_max[98] = (&detect_max[98]) ? 1:0;
assign is_max[99] = (&detect_max[99]) ? 1:0;
assign is_max[100] = (&detect_max[100]) ? 1:0;
assign is_max[101] = (&detect_max[101]) ? 1:0;
assign is_max[102] = (&detect_max[102]) ? 1:0;
assign is_max[103] = (&detect_max[103]) ? 1:0;
assign is_max[104] = (&detect_max[104]) ? 1:0;
assign is_max[105] = (&detect_max[105]) ? 1:0;
assign is_max[106] = (&detect_max[106]) ? 1:0;
assign is_max[107] = (&detect_max[107]) ? 1:0;
assign is_max[108] = (&detect_max[108]) ? 1:0;
assign is_max[109] = (&detect_max[109]) ? 1:0;
assign is_max[110] = (&detect_max[110]) ? 1:0;
assign is_max[111] = (&detect_max[111]) ? 1:0;
assign is_max[112] = (&detect_max[112]) ? 1:0;
assign is_max[113] = (&detect_max[113]) ? 1:0;
assign is_max[114] = (&detect_max[114]) ? 1:0;
assign is_max[115] = (&detect_max[115]) ? 1:0;
assign is_max[116] = (&detect_max[116]) ? 1:0;
assign is_max[117] = (&detect_max[117]) ? 1:0;
assign is_max[118] = (&detect_max[118]) ? 1:0;
assign is_max[119] = (&detect_max[119]) ? 1:0;
assign is_max[120] = (&detect_max[120]) ? 1:0;
assign is_max[121] = (&detect_max[121]) ? 1:0;
assign is_max[122] = (&detect_max[122]) ? 1:0;
assign is_max[123] = (&detect_max[123]) ? 1:0;
assign is_max[124] = (&detect_max[124]) ? 1:0;
assign is_max[125] = (&detect_max[125]) ? 1:0;
assign is_max[126] = (&detect_max[126]) ? 1:0;
assign is_max[127] = (&detect_max[127]) ? 1:0;
assign is_max[128] = (&detect_max[128]) ? 1:0;
assign is_max[129] = (&detect_max[129]) ? 1:0;
assign is_max[130] = (&detect_max[130]) ? 1:0;
assign is_max[131] = (&detect_max[131]) ? 1:0;
assign is_max[132] = (&detect_max[132]) ? 1:0;
assign is_max[133] = (&detect_max[133]) ? 1:0;
assign is_max[134] = (&detect_max[134]) ? 1:0;
assign is_max[135] = (&detect_max[135]) ? 1:0;
assign is_max[136] = (&detect_max[136]) ? 1:0;
assign is_max[137] = (&detect_max[137]) ? 1:0;
assign is_max[138] = (&detect_max[138]) ? 1:0;
assign is_max[139] = (&detect_max[139]) ? 1:0;
assign is_max[140] = (&detect_max[140]) ? 1:0;
assign is_max[141] = (&detect_max[141]) ? 1:0;
assign is_max[142] = (&detect_max[142]) ? 1:0;
assign is_max[143] = (&detect_max[143]) ? 1:0;
assign is_max[144] = (&detect_max[144]) ? 1:0;
assign is_max[145] = (&detect_max[145]) ? 1:0;
assign is_max[146] = (&detect_max[146]) ? 1:0;
assign is_max[147] = (&detect_max[147]) ? 1:0;
assign is_max[148] = (&detect_max[148]) ? 1:0;
assign is_max[149] = (&detect_max[149]) ? 1:0;
assign is_max[150] = (&detect_max[150]) ? 1:0;
assign is_max[151] = (&detect_max[151]) ? 1:0;
assign is_max[152] = (&detect_max[152]) ? 1:0;
assign is_max[153] = (&detect_max[153]) ? 1:0;
assign is_max[154] = (&detect_max[154]) ? 1:0;
assign is_max[155] = (&detect_max[155]) ? 1:0;
assign is_max[156] = (&detect_max[156]) ? 1:0;
assign is_max[157] = (&detect_max[157]) ? 1:0;
assign is_max[158] = (&detect_max[158]) ? 1:0;
assign is_max[159] = (&detect_max[159]) ? 1:0;
assign is_max[160] = (&detect_max[160]) ? 1:0;
assign is_max[161] = (&detect_max[161]) ? 1:0;
assign is_max[162] = (&detect_max[162]) ? 1:0;
assign is_max[163] = (&detect_max[163]) ? 1:0;
assign is_max[164] = (&detect_max[164]) ? 1:0;
assign is_max[165] = (&detect_max[165]) ? 1:0;
assign is_max[166] = (&detect_max[166]) ? 1:0;
assign is_max[167] = (&detect_max[167]) ? 1:0;
assign is_max[168] = (&detect_max[168]) ? 1:0;
assign is_max[169] = (&detect_max[169]) ? 1:0;
assign is_max[170] = (&detect_max[170]) ? 1:0;
assign is_max[171] = (&detect_max[171]) ? 1:0;
assign is_max[172] = (&detect_max[172]) ? 1:0;
assign is_max[173] = (&detect_max[173]) ? 1:0;
assign is_max[174] = (&detect_max[174]) ? 1:0;
assign is_max[175] = (&detect_max[175]) ? 1:0;
assign is_max[176] = (&detect_max[176]) ? 1:0;
assign is_max[177] = (&detect_max[177]) ? 1:0;
assign is_max[178] = (&detect_max[178]) ? 1:0;
assign is_max[179] = (&detect_max[179]) ? 1:0;
assign is_max[180] = (&detect_max[180]) ? 1:0;
assign is_max[181] = (&detect_max[181]) ? 1:0;
assign is_max[182] = (&detect_max[182]) ? 1:0;
assign is_max[183] = (&detect_max[183]) ? 1:0;
assign is_max[184] = (&detect_max[184]) ? 1:0;
assign is_max[185] = (&detect_max[185]) ? 1:0;
assign is_max[186] = (&detect_max[186]) ? 1:0;
assign is_max[187] = (&detect_max[187]) ? 1:0;
assign is_max[188] = (&detect_max[188]) ? 1:0;
assign is_max[189] = (&detect_max[189]) ? 1:0;
assign is_max[190] = (&detect_max[190]) ? 1:0;
assign is_max[191] = (&detect_max[191]) ? 1:0;
assign is_max[192] = (&detect_max[192]) ? 1:0;
assign is_max[193] = (&detect_max[193]) ? 1:0;
assign is_max[194] = (&detect_max[194]) ? 1:0;
assign is_max[195] = (&detect_max[195]) ? 1:0;
assign is_max[196] = (&detect_max[196]) ? 1:0;
assign is_max[197] = (&detect_max[197]) ? 1:0;
assign is_max[198] = (&detect_max[198]) ? 1:0;
assign is_max[199] = (&detect_max[199]) ? 1:0;
assign is_max[200] = (&detect_max[200]) ? 1:0;
assign is_max[201] = (&detect_max[201]) ? 1:0;
assign is_max[202] = (&detect_max[202]) ? 1:0;
assign is_max[203] = (&detect_max[203]) ? 1:0;
assign is_max[204] = (&detect_max[204]) ? 1:0;
assign is_max[205] = (&detect_max[205]) ? 1:0;
assign is_max[206] = (&detect_max[206]) ? 1:0;
assign is_max[207] = (&detect_max[207]) ? 1:0;
assign is_max[208] = (&detect_max[208]) ? 1:0;
assign is_max[209] = (&detect_max[209]) ? 1:0;
assign is_max[210] = (&detect_max[210]) ? 1:0;
assign is_max[211] = (&detect_max[211]) ? 1:0;
assign is_max[212] = (&detect_max[212]) ? 1:0;
assign is_max[213] = (&detect_max[213]) ? 1:0;
assign is_max[214] = (&detect_max[214]) ? 1:0;
assign is_max[215] = (&detect_max[215]) ? 1:0;
assign is_max[216] = (&detect_max[216]) ? 1:0;
assign is_max[217] = (&detect_max[217]) ? 1:0;
assign is_max[218] = (&detect_max[218]) ? 1:0;
assign is_max[219] = (&detect_max[219]) ? 1:0;
assign is_max[220] = (&detect_max[220]) ? 1:0;
assign is_max[221] = (&detect_max[221]) ? 1:0;
assign is_max[222] = (&detect_max[222]) ? 1:0;
assign is_max[223] = (&detect_max[223]) ? 1:0;
assign is_max[224] = (&detect_max[224]) ? 1:0;
assign is_max[225] = (&detect_max[225]) ? 1:0;
assign is_max[226] = (&detect_max[226]) ? 1:0;
assign is_max[227] = (&detect_max[227]) ? 1:0;
assign is_max[228] = (&detect_max[228]) ? 1:0;
assign is_max[229] = (&detect_max[229]) ? 1:0;
assign is_max[230] = (&detect_max[230]) ? 1:0;
assign is_max[231] = (&detect_max[231]) ? 1:0;
assign is_max[232] = (&detect_max[232]) ? 1:0;
assign is_max[233] = (&detect_max[233]) ? 1:0;
assign is_max[234] = (&detect_max[234]) ? 1:0;
assign is_max[235] = (&detect_max[235]) ? 1:0;
assign is_max[236] = (&detect_max[236]) ? 1:0;
assign is_max[237] = (&detect_max[237]) ? 1:0;
assign is_max[238] = (&detect_max[238]) ? 1:0;
assign is_max[239] = (&detect_max[239]) ? 1:0;
assign is_max[240] = (&detect_max[240]) ? 1:0;
assign is_max[241] = (&detect_max[241]) ? 1:0;
assign is_max[242] = (&detect_max[242]) ? 1:0;
assign is_max[243] = (&detect_max[243]) ? 1:0;
assign is_max[244] = (&detect_max[244]) ? 1:0;
assign is_max[245] = (&detect_max[245]) ? 1:0;
assign is_max[246] = (&detect_max[246]) ? 1:0;
assign is_max[247] = (&detect_max[247]) ? 1:0;
assign is_max[248] = (&detect_max[248]) ? 1:0;
assign is_max[249] = (&detect_max[249]) ? 1:0;
assign is_max[250] = (&detect_max[250]) ? 1:0;
assign is_max[251] = (&detect_max[251]) ? 1:0;
assign is_max[252] = (&detect_max[252]) ? 1:0;
assign is_max[253] = (&detect_max[253]) ? 1:0;
assign is_max[254] = (&detect_max[254]) ? 1:0;
assign is_max[255] = (&detect_max[255]) ? 1:0;
assign is_max[256] = (&detect_max[256]) ? 1:0;
assign is_max[257] = (&detect_max[257]) ? 1:0;
assign is_max[258] = (&detect_max[258]) ? 1:0;
assign is_max[259] = (&detect_max[259]) ? 1:0;
assign is_max[260] = (&detect_max[260]) ? 1:0;
assign is_max[261] = (&detect_max[261]) ? 1:0;
assign is_max[262] = (&detect_max[262]) ? 1:0;
assign is_max[263] = (&detect_max[263]) ? 1:0;
assign is_max[264] = (&detect_max[264]) ? 1:0;
assign is_max[265] = (&detect_max[265]) ? 1:0;
assign is_max[266] = (&detect_max[266]) ? 1:0;
assign is_max[267] = (&detect_max[267]) ? 1:0;
assign is_max[268] = (&detect_max[268]) ? 1:0;
assign is_max[269] = (&detect_max[269]) ? 1:0;
assign is_max[270] = (&detect_max[270]) ? 1:0;
assign is_max[271] = (&detect_max[271]) ? 1:0;
assign is_max[272] = (&detect_max[272]) ? 1:0;
assign is_max[273] = (&detect_max[273]) ? 1:0;
assign is_max[274] = (&detect_max[274]) ? 1:0;
assign is_max[275] = (&detect_max[275]) ? 1:0;
assign is_max[276] = (&detect_max[276]) ? 1:0;
assign is_max[277] = (&detect_max[277]) ? 1:0;
assign is_max[278] = (&detect_max[278]) ? 1:0;
assign is_max[279] = (&detect_max[279]) ? 1:0;
assign is_max[280] = (&detect_max[280]) ? 1:0;
assign is_max[281] = (&detect_max[281]) ? 1:0;
assign is_max[282] = (&detect_max[282]) ? 1:0;
assign is_max[283] = (&detect_max[283]) ? 1:0;
assign is_max[284] = (&detect_max[284]) ? 1:0;
assign is_max[285] = (&detect_max[285]) ? 1:0;
assign is_max[286] = (&detect_max[286]) ? 1:0;
assign is_max[287] = (&detect_max[287]) ? 1:0;
assign is_max[288] = (&detect_max[288]) ? 1:0;
assign is_max[289] = (&detect_max[289]) ? 1:0;
assign is_max[290] = (&detect_max[290]) ? 1:0;
assign is_max[291] = (&detect_max[291]) ? 1:0;
assign is_max[292] = (&detect_max[292]) ? 1:0;
assign is_max[293] = (&detect_max[293]) ? 1:0;
assign is_max[294] = (&detect_max[294]) ? 1:0;
assign is_max[295] = (&detect_max[295]) ? 1:0;
assign is_max[296] = (&detect_max[296]) ? 1:0;
assign is_max[297] = (&detect_max[297]) ? 1:0;
assign is_max[298] = (&detect_max[298]) ? 1:0;
assign is_max[299] = (&detect_max[299]) ? 1:0;
assign is_max[300] = (&detect_max[300]) ? 1:0;
assign is_max[301] = (&detect_max[301]) ? 1:0;
assign is_max[302] = (&detect_max[302]) ? 1:0;
assign is_max[303] = (&detect_max[303]) ? 1:0;
assign is_max[304] = (&detect_max[304]) ? 1:0;
assign is_max[305] = (&detect_max[305]) ? 1:0;
assign is_max[306] = (&detect_max[306]) ? 1:0;
assign is_max[307] = (&detect_max[307]) ? 1:0;
assign is_max[308] = (&detect_max[308]) ? 1:0;
assign is_max[309] = (&detect_max[309]) ? 1:0;
assign is_max[310] = (&detect_max[310]) ? 1:0;
assign is_max[311] = (&detect_max[311]) ? 1:0;
assign is_max[312] = (&detect_max[312]) ? 1:0;
assign is_max[313] = (&detect_max[313]) ? 1:0;
assign is_max[314] = (&detect_max[314]) ? 1:0;
assign is_max[315] = (&detect_max[315]) ? 1:0;
assign is_max[316] = (&detect_max[316]) ? 1:0;
assign is_max[317] = (&detect_max[317]) ? 1:0;
assign is_max[318] = (&detect_max[318]) ? 1:0;
assign is_max[319] = (&detect_max[319]) ? 1:0;
assign is_max[320] = (&detect_max[320]) ? 1:0;
assign is_max[321] = (&detect_max[321]) ? 1:0;
assign is_max[322] = (&detect_max[322]) ? 1:0;
assign is_max[323] = (&detect_max[323]) ? 1:0;
assign is_max[324] = (&detect_max[324]) ? 1:0;
assign is_max[325] = (&detect_max[325]) ? 1:0;
assign is_max[326] = (&detect_max[326]) ? 1:0;
assign is_max[327] = (&detect_max[327]) ? 1:0;
assign is_max[328] = (&detect_max[328]) ? 1:0;
assign is_max[329] = (&detect_max[329]) ? 1:0;
assign is_max[330] = (&detect_max[330]) ? 1:0;
assign is_max[331] = (&detect_max[331]) ? 1:0;
assign is_max[332] = (&detect_max[332]) ? 1:0;
assign is_max[333] = (&detect_max[333]) ? 1:0;
assign is_max[334] = (&detect_max[334]) ? 1:0;
assign is_max[335] = (&detect_max[335]) ? 1:0;
assign is_max[336] = (&detect_max[336]) ? 1:0;
assign is_max[337] = (&detect_max[337]) ? 1:0;
assign is_max[338] = (&detect_max[338]) ? 1:0;
assign is_max[339] = (&detect_max[339]) ? 1:0;
assign is_max[340] = (&detect_max[340]) ? 1:0;
assign is_max[341] = (&detect_max[341]) ? 1:0;
assign is_max[342] = (&detect_max[342]) ? 1:0;
assign is_max[343] = (&detect_max[343]) ? 1:0;
assign is_max[344] = (&detect_max[344]) ? 1:0;
assign is_max[345] = (&detect_max[345]) ? 1:0;
assign is_max[346] = (&detect_max[346]) ? 1:0;
assign is_max[347] = (&detect_max[347]) ? 1:0;
assign is_max[348] = (&detect_max[348]) ? 1:0;
assign is_max[349] = (&detect_max[349]) ? 1:0;
assign is_max[350] = (&detect_max[350]) ? 1:0;
assign is_max[351] = (&detect_max[351]) ? 1:0;
assign is_max[352] = (&detect_max[352]) ? 1:0;
assign is_max[353] = (&detect_max[353]) ? 1:0;
assign is_max[354] = (&detect_max[354]) ? 1:0;
assign is_max[355] = (&detect_max[355]) ? 1:0;
assign is_max[356] = (&detect_max[356]) ? 1:0;
assign is_max[357] = (&detect_max[357]) ? 1:0;
assign is_max[358] = (&detect_max[358]) ? 1:0;
assign is_max[359] = (&detect_max[359]) ? 1:0;
assign is_max[360] = (&detect_max[360]) ? 1:0;
assign is_max[361] = (&detect_max[361]) ? 1:0;
assign is_max[362] = (&detect_max[362]) ? 1:0;
assign is_max[363] = (&detect_max[363]) ? 1:0;
assign is_max[364] = (&detect_max[364]) ? 1:0;
assign is_max[365] = (&detect_max[365]) ? 1:0;
assign is_max[366] = (&detect_max[366]) ? 1:0;
assign is_max[367] = (&detect_max[367]) ? 1:0;
assign is_max[368] = (&detect_max[368]) ? 1:0;
assign is_max[369] = (&detect_max[369]) ? 1:0;
assign is_max[370] = (&detect_max[370]) ? 1:0;
assign is_max[371] = (&detect_max[371]) ? 1:0;
assign is_max[372] = (&detect_max[372]) ? 1:0;
assign is_max[373] = (&detect_max[373]) ? 1:0;
assign is_max[374] = (&detect_max[374]) ? 1:0;
assign is_max[375] = (&detect_max[375]) ? 1:0;
assign is_max[376] = (&detect_max[376]) ? 1:0;
assign is_max[377] = (&detect_max[377]) ? 1:0;
assign is_max[378] = (&detect_max[378]) ? 1:0;
assign is_max[379] = (&detect_max[379]) ? 1:0;
assign is_max[380] = (&detect_max[380]) ? 1:0;
assign is_max[381] = (&detect_max[381]) ? 1:0;
assign is_max[382] = (&detect_max[382]) ? 1:0;
assign is_max[383] = (&detect_max[383]) ? 1:0;
assign is_max[384] = (&detect_max[384]) ? 1:0;
assign is_max[385] = (&detect_max[385]) ? 1:0;
assign is_max[386] = (&detect_max[386]) ? 1:0;
assign is_max[387] = (&detect_max[387]) ? 1:0;
assign is_max[388] = (&detect_max[388]) ? 1:0;
assign is_max[389] = (&detect_max[389]) ? 1:0;
assign is_max[390] = (&detect_max[390]) ? 1:0;
assign is_max[391] = (&detect_max[391]) ? 1:0;
assign is_max[392] = (&detect_max[392]) ? 1:0;
assign is_max[393] = (&detect_max[393]) ? 1:0;
assign is_max[394] = (&detect_max[394]) ? 1:0;
assign is_max[395] = (&detect_max[395]) ? 1:0;
assign is_max[396] = (&detect_max[396]) ? 1:0;
assign is_max[397] = (&detect_max[397]) ? 1:0;
assign is_max[398] = (&detect_max[398]) ? 1:0;
assign is_max[399] = (&detect_max[399]) ? 1:0;
assign is_max[400] = (&detect_max[400]) ? 1:0;
assign is_max[401] = (&detect_max[401]) ? 1:0;
assign is_max[402] = (&detect_max[402]) ? 1:0;
assign is_max[403] = (&detect_max[403]) ? 1:0;
assign is_max[404] = (&detect_max[404]) ? 1:0;
assign is_max[405] = (&detect_max[405]) ? 1:0;
assign is_max[406] = (&detect_max[406]) ? 1:0;
assign is_max[407] = (&detect_max[407]) ? 1:0;
assign is_max[408] = (&detect_max[408]) ? 1:0;
assign is_max[409] = (&detect_max[409]) ? 1:0;
assign is_max[410] = (&detect_max[410]) ? 1:0;
assign is_max[411] = (&detect_max[411]) ? 1:0;
assign is_max[412] = (&detect_max[412]) ? 1:0;
assign is_max[413] = (&detect_max[413]) ? 1:0;
assign is_max[414] = (&detect_max[414]) ? 1:0;
assign is_max[415] = (&detect_max[415]) ? 1:0;
assign is_max[416] = (&detect_max[416]) ? 1:0;
assign is_max[417] = (&detect_max[417]) ? 1:0;
assign is_max[418] = (&detect_max[418]) ? 1:0;
assign is_max[419] = (&detect_max[419]) ? 1:0;
assign is_max[420] = (&detect_max[420]) ? 1:0;
assign is_max[421] = (&detect_max[421]) ? 1:0;
assign is_max[422] = (&detect_max[422]) ? 1:0;
assign is_max[423] = (&detect_max[423]) ? 1:0;
assign is_max[424] = (&detect_max[424]) ? 1:0;
assign is_max[425] = (&detect_max[425]) ? 1:0;
assign is_max[426] = (&detect_max[426]) ? 1:0;
assign is_max[427] = (&detect_max[427]) ? 1:0;
assign is_max[428] = (&detect_max[428]) ? 1:0;
assign is_max[429] = (&detect_max[429]) ? 1:0;
assign is_max[430] = (&detect_max[430]) ? 1:0;
assign is_max[431] = (&detect_max[431]) ? 1:0;
assign is_max[432] = (&detect_max[432]) ? 1:0;
assign is_max[433] = (&detect_max[433]) ? 1:0;
assign is_max[434] = (&detect_max[434]) ? 1:0;
assign is_max[435] = (&detect_max[435]) ? 1:0;
assign is_max[436] = (&detect_max[436]) ? 1:0;
assign is_max[437] = (&detect_max[437]) ? 1:0;
assign is_max[438] = (&detect_max[438]) ? 1:0;
assign is_max[439] = (&detect_max[439]) ? 1:0;
assign is_max[440] = (&detect_max[440]) ? 1:0;
assign is_max[441] = (&detect_max[441]) ? 1:0;
assign is_max[442] = (&detect_max[442]) ? 1:0;
assign is_max[443] = (&detect_max[443]) ? 1:0;
assign is_max[444] = (&detect_max[444]) ? 1:0;
assign is_max[445] = (&detect_max[445]) ? 1:0;
assign is_max[446] = (&detect_max[446]) ? 1:0;
assign is_max[447] = (&detect_max[447]) ? 1:0;
assign is_max[448] = (&detect_max[448]) ? 1:0;
assign is_max[449] = (&detect_max[449]) ? 1:0;
assign is_max[450] = (&detect_max[450]) ? 1:0;
assign is_max[451] = (&detect_max[451]) ? 1:0;
assign is_max[452] = (&detect_max[452]) ? 1:0;
assign is_max[453] = (&detect_max[453]) ? 1:0;
assign is_max[454] = (&detect_max[454]) ? 1:0;
assign is_max[455] = (&detect_max[455]) ? 1:0;
assign is_max[456] = (&detect_max[456]) ? 1:0;
assign is_max[457] = (&detect_max[457]) ? 1:0;
assign is_max[458] = (&detect_max[458]) ? 1:0;
assign is_max[459] = (&detect_max[459]) ? 1:0;
assign is_max[460] = (&detect_max[460]) ? 1:0;
assign is_max[461] = (&detect_max[461]) ? 1:0;
assign is_max[462] = (&detect_max[462]) ? 1:0;
assign is_max[463] = (&detect_max[463]) ? 1:0;
assign is_max[464] = (&detect_max[464]) ? 1:0;
assign is_max[465] = (&detect_max[465]) ? 1:0;
assign is_max[466] = (&detect_max[466]) ? 1:0;
assign is_max[467] = (&detect_max[467]) ? 1:0;
assign is_max[468] = (&detect_max[468]) ? 1:0;
assign is_max[469] = (&detect_max[469]) ? 1:0;
assign is_max[470] = (&detect_max[470]) ? 1:0;
assign is_max[471] = (&detect_max[471]) ? 1:0;
assign is_max[472] = (&detect_max[472]) ? 1:0;
assign is_max[473] = (&detect_max[473]) ? 1:0;
assign is_max[474] = (&detect_max[474]) ? 1:0;
assign is_max[475] = (&detect_max[475]) ? 1:0;
assign is_max[476] = (&detect_max[476]) ? 1:0;
assign is_max[477] = (&detect_max[477]) ? 1:0;
assign is_max[478] = (&detect_max[478]) ? 1:0;
assign is_max[479] = (&detect_max[479]) ? 1:0;
assign is_max[480] = (&detect_max[480]) ? 1:0;
assign is_max[481] = (&detect_max[481]) ? 1:0;
assign is_max[482] = (&detect_max[482]) ? 1:0;
assign is_max[483] = (&detect_max[483]) ? 1:0;
assign is_max[484] = (&detect_max[484]) ? 1:0;
assign is_max[485] = (&detect_max[485]) ? 1:0;
assign is_max[486] = (&detect_max[486]) ? 1:0;
assign is_max[487] = (&detect_max[487]) ? 1:0;
assign is_max[488] = (&detect_max[488]) ? 1:0;
assign is_max[489] = (&detect_max[489]) ? 1:0;
assign is_max[490] = (&detect_max[490]) ? 1:0;
assign is_max[491] = (&detect_max[491]) ? 1:0;
assign is_max[492] = (&detect_max[492]) ? 1:0;
assign is_max[493] = (&detect_max[493]) ? 1:0;
assign is_max[494] = (&detect_max[494]) ? 1:0;
assign is_max[495] = (&detect_max[495]) ? 1:0;
assign is_max[496] = (&detect_max[496]) ? 1:0;
assign is_max[497] = (&detect_max[497]) ? 1:0;
assign is_max[498] = (&detect_max[498]) ? 1:0;
assign is_max[499] = (&detect_max[499]) ? 1:0;
assign is_max[500] = (&detect_max[500]) ? 1:0;
assign is_max[501] = (&detect_max[501]) ? 1:0;
assign is_max[502] = (&detect_max[502]) ? 1:0;
assign is_max[503] = (&detect_max[503]) ? 1:0;
assign is_max[504] = (&detect_max[504]) ? 1:0;
assign is_max[505] = (&detect_max[505]) ? 1:0;
assign is_max[506] = (&detect_max[506]) ? 1:0;
assign is_max[507] = (&detect_max[507]) ? 1:0;
assign is_max[508] = (&detect_max[508]) ? 1:0;
assign is_max[509] = (&detect_max[509]) ? 1:0;
assign is_max[510] = (&detect_max[510]) ? 1:0;
assign is_max[511] = (&detect_max[511]) ? 1:0;
assign is_max[512] = (&detect_max[512]) ? 1:0;
assign is_max[513] = (&detect_max[513]) ? 1:0;
assign is_max[514] = (&detect_max[514]) ? 1:0;
assign is_max[515] = (&detect_max[515]) ? 1:0;
assign is_max[516] = (&detect_max[516]) ? 1:0;
assign is_max[517] = (&detect_max[517]) ? 1:0;
assign is_max[518] = (&detect_max[518]) ? 1:0;
assign is_max[519] = (&detect_max[519]) ? 1:0;
assign is_max[520] = (&detect_max[520]) ? 1:0;
assign is_max[521] = (&detect_max[521]) ? 1:0;
assign is_max[522] = (&detect_max[522]) ? 1:0;
assign is_max[523] = (&detect_max[523]) ? 1:0;
assign is_max[524] = (&detect_max[524]) ? 1:0;
assign is_max[525] = (&detect_max[525]) ? 1:0;
assign is_max[526] = (&detect_max[526]) ? 1:0;
assign is_max[527] = (&detect_max[527]) ? 1:0;
assign is_max[528] = (&detect_max[528]) ? 1:0;
assign is_max[529] = (&detect_max[529]) ? 1:0;
assign is_max[530] = (&detect_max[530]) ? 1:0;
assign is_max[531] = (&detect_max[531]) ? 1:0;
assign is_max[532] = (&detect_max[532]) ? 1:0;
assign is_max[533] = (&detect_max[533]) ? 1:0;
assign is_max[534] = (&detect_max[534]) ? 1:0;
assign is_max[535] = (&detect_max[535]) ? 1:0;
assign is_max[536] = (&detect_max[536]) ? 1:0;
assign is_max[537] = (&detect_max[537]) ? 1:0;
assign is_max[538] = (&detect_max[538]) ? 1:0;
assign is_max[539] = (&detect_max[539]) ? 1:0;
assign is_max[540] = (&detect_max[540]) ? 1:0;
assign is_max[541] = (&detect_max[541]) ? 1:0;
assign is_max[542] = (&detect_max[542]) ? 1:0;
assign is_max[543] = (&detect_max[543]) ? 1:0;
assign is_max[544] = (&detect_max[544]) ? 1:0;
assign is_max[545] = (&detect_max[545]) ? 1:0;
assign is_max[546] = (&detect_max[546]) ? 1:0;
assign is_max[547] = (&detect_max[547]) ? 1:0;
assign is_max[548] = (&detect_max[548]) ? 1:0;
assign is_max[549] = (&detect_max[549]) ? 1:0;
assign is_max[550] = (&detect_max[550]) ? 1:0;
assign is_max[551] = (&detect_max[551]) ? 1:0;
assign is_max[552] = (&detect_max[552]) ? 1:0;
assign is_max[553] = (&detect_max[553]) ? 1:0;
assign is_max[554] = (&detect_max[554]) ? 1:0;
assign is_max[555] = (&detect_max[555]) ? 1:0;
assign is_max[556] = (&detect_max[556]) ? 1:0;
assign is_max[557] = (&detect_max[557]) ? 1:0;
assign is_max[558] = (&detect_max[558]) ? 1:0;
assign is_max[559] = (&detect_max[559]) ? 1:0;
assign is_max[560] = (&detect_max[560]) ? 1:0;
assign is_max[561] = (&detect_max[561]) ? 1:0;
assign is_max[562] = (&detect_max[562]) ? 1:0;
assign is_max[563] = (&detect_max[563]) ? 1:0;
assign is_max[564] = (&detect_max[564]) ? 1:0;
assign is_max[565] = (&detect_max[565]) ? 1:0;
assign is_max[566] = (&detect_max[566]) ? 1:0;
assign is_max[567] = (&detect_max[567]) ? 1:0;
assign is_max[568] = (&detect_max[568]) ? 1:0;
assign is_max[569] = (&detect_max[569]) ? 1:0;
assign is_max[570] = (&detect_max[570]) ? 1:0;
assign is_max[571] = (&detect_max[571]) ? 1:0;
assign is_max[572] = (&detect_max[572]) ? 1:0;
assign is_max[573] = (&detect_max[573]) ? 1:0;
assign is_max[574] = (&detect_max[574]) ? 1:0;
assign is_max[575] = (&detect_max[575]) ? 1:0;
assign is_max[576] = (&detect_max[576]) ? 1:0;
assign is_max[577] = (&detect_max[577]) ? 1:0;
assign is_max[578] = (&detect_max[578]) ? 1:0;
assign is_max[579] = (&detect_max[579]) ? 1:0;
assign is_max[580] = (&detect_max[580]) ? 1:0;
assign is_max[581] = (&detect_max[581]) ? 1:0;
assign is_max[582] = (&detect_max[582]) ? 1:0;
assign is_max[583] = (&detect_max[583]) ? 1:0;
assign is_max[584] = (&detect_max[584]) ? 1:0;
assign is_max[585] = (&detect_max[585]) ? 1:0;
assign is_max[586] = (&detect_max[586]) ? 1:0;
assign is_max[587] = (&detect_max[587]) ? 1:0;
assign is_max[588] = (&detect_max[588]) ? 1:0;
assign is_max[589] = (&detect_max[589]) ? 1:0;
assign is_max[590] = (&detect_max[590]) ? 1:0;
assign is_max[591] = (&detect_max[591]) ? 1:0;
assign is_max[592] = (&detect_max[592]) ? 1:0;
assign is_max[593] = (&detect_max[593]) ? 1:0;
assign is_max[594] = (&detect_max[594]) ? 1:0;
assign is_max[595] = (&detect_max[595]) ? 1:0;
assign is_max[596] = (&detect_max[596]) ? 1:0;
assign is_max[597] = (&detect_max[597]) ? 1:0;
assign is_max[598] = (&detect_max[598]) ? 1:0;
assign is_max[599] = (&detect_max[599]) ? 1:0;
assign is_max[600] = (&detect_max[600]) ? 1:0;
assign is_max[601] = (&detect_max[601]) ? 1:0;
assign is_max[602] = (&detect_max[602]) ? 1:0;
assign is_max[603] = (&detect_max[603]) ? 1:0;
assign is_max[604] = (&detect_max[604]) ? 1:0;
assign is_max[605] = (&detect_max[605]) ? 1:0;
assign is_max[606] = (&detect_max[606]) ? 1:0;
assign is_max[607] = (&detect_max[607]) ? 1:0;
assign is_max[608] = (&detect_max[608]) ? 1:0;
assign is_max[609] = (&detect_max[609]) ? 1:0;
assign is_max[610] = (&detect_max[610]) ? 1:0;
assign is_max[611] = (&detect_max[611]) ? 1:0;
assign is_max[612] = (&detect_max[612]) ? 1:0;
assign is_max[613] = (&detect_max[613]) ? 1:0;
assign is_max[614] = (&detect_max[614]) ? 1:0;
assign is_max[615] = (&detect_max[615]) ? 1:0;
assign is_max[616] = (&detect_max[616]) ? 1:0;
assign is_max[617] = (&detect_max[617]) ? 1:0;
assign is_max[618] = (&detect_max[618]) ? 1:0;
assign is_max[619] = (&detect_max[619]) ? 1:0;
assign is_max[620] = (&detect_max[620]) ? 1:0;
assign is_max[621] = (&detect_max[621]) ? 1:0;
assign is_max[622] = (&detect_max[622]) ? 1:0;
assign is_max[623] = (&detect_max[623]) ? 1:0;
assign is_max[624] = (&detect_max[624]) ? 1:0;
assign is_max[625] = (&detect_max[625]) ? 1:0;
assign is_max[626] = (&detect_max[626]) ? 1:0;
assign is_max[627] = (&detect_max[627]) ? 1:0;
assign is_max[628] = (&detect_max[628]) ? 1:0;
assign is_max[629] = (&detect_max[629]) ? 1:0;
assign is_max[630] = (&detect_max[630]) ? 1:0;
assign is_max[631] = (&detect_max[631]) ? 1:0;
assign is_max[632] = (&detect_max[632]) ? 1:0;
assign is_max[633] = (&detect_max[633]) ? 1:0;
assign is_max[634] = (&detect_max[634]) ? 1:0;
assign is_max[635] = (&detect_max[635]) ? 1:0;
assign is_max[636] = (&detect_max[636]) ? 1:0;
assign is_max[637] = (&detect_max[637]) ? 1:0;

wire	[25:0]		detect_min[0:637];
assign detect_min[0][0] = (mid_1[15:8] < top_0[7:0]) ? 1 : 0;
assign detect_min[0][1] = (mid_1[15:8] < top_0[15:8]) ? 1 : 0;
assign detect_min[0][2] = (mid_1[15:8] < top_0[23:16]) ? 1 : 0;
assign detect_min[0][3] = (mid_1[15:8] < top_1[7:0]) ? 1 : 0;
assign detect_min[0][4] = (mid_1[15:8] < top_1[15:8]) ? 1 : 0;
assign detect_min[0][5] = (mid_1[15:8] < top_1[23:16]) ? 1 : 0;
assign detect_min[0][6] = (mid_1[15:8] < top_2[7:0]) ? 1 : 0;
assign detect_min[0][7] = (mid_1[15:8] < top_2[15:8]) ? 1 : 0;
assign detect_min[0][8] = (mid_1[15:8] < top_2[23:16]) ? 1 : 0;
assign detect_min[0][9] = (mid_1[15:8] < mid_0[7:0]) ? 1 : 0;
assign detect_min[0][10] = (mid_1[15:8] < mid_0[15:8]) ? 1 : 0;
assign detect_min[0][11] = (mid_1[15:8] < mid_0[23:16]) ? 1 : 0;
assign detect_min[0][12] = (mid_1[15:8] < mid_1[7:0]) ? 1 : 0;
assign detect_min[0][13] = (mid_1[15:8] < mid_1[23:16]) ? 1 : 0;
assign detect_min[0][14] = (mid_1[15:8] < mid_2[7:0]) ? 1 : 0;
assign detect_min[0][15] = (mid_1[15:8] < mid_2[15:8]) ? 1 : 0;
assign detect_min[0][16] = (mid_1[15:8] < mid_2[23:16]) ? 1 : 0;
assign detect_min[0][17] = (mid_1[15:8] < btm_0[7:0]) ? 1 : 0;
assign detect_min[0][18] = (mid_1[15:8] < btm_0[15:8]) ? 1 : 0;
assign detect_min[0][19] = (mid_1[15:8] < btm_0[23:16]) ? 1 : 0;
assign detect_min[0][20] = (mid_1[15:8] < btm_1[7:0]) ? 1 : 0;
assign detect_min[0][21] = (mid_1[15:8] < btm_1[15:8]) ? 1 : 0;
assign detect_min[0][22] = (mid_1[15:8] < btm_1[23:16]) ? 1 : 0;
assign detect_min[0][23] = (mid_1[15:8] < btm_2[7:0]) ? 1 : 0;
assign detect_min[0][24] = (mid_1[15:8] < btm_2[15:8]) ? 1 : 0;
assign detect_min[0][25] = (mid_1[15:8] < btm_2[23:16]) ? 1 : 0;

assign detect_min[1][0] = (mid_1[23:16] < top_0[15:8]) ? 1 : 0;
assign detect_min[1][1] = (mid_1[23:16] < top_0[23:16]) ? 1 : 0;
assign detect_min[1][2] = (mid_1[23:16] < top_0[31:24]) ? 1 : 0;
assign detect_min[1][3] = (mid_1[23:16] < top_1[15:8]) ? 1 : 0;
assign detect_min[1][4] = (mid_1[23:16] < top_1[23:16]) ? 1 : 0;
assign detect_min[1][5] = (mid_1[23:16] < top_1[31:24]) ? 1 : 0;
assign detect_min[1][6] = (mid_1[23:16] < top_2[15:8]) ? 1 : 0;
assign detect_min[1][7] = (mid_1[23:16] < top_2[23:16]) ? 1 : 0;
assign detect_min[1][8] = (mid_1[23:16] < top_2[31:24]) ? 1 : 0;
assign detect_min[1][9] = (mid_1[23:16] < mid_0[15:8]) ? 1 : 0;
assign detect_min[1][10] = (mid_1[23:16] < mid_0[23:16]) ? 1 : 0;
assign detect_min[1][11] = (mid_1[23:16] < mid_0[31:24]) ? 1 : 0;
assign detect_min[1][12] = (mid_1[23:16] < mid_1[15:8]) ? 1 : 0;
assign detect_min[1][13] = (mid_1[23:16] < mid_1[31:24]) ? 1 : 0;
assign detect_min[1][14] = (mid_1[23:16] < mid_2[15:8]) ? 1 : 0;
assign detect_min[1][15] = (mid_1[23:16] < mid_2[23:16]) ? 1 : 0;
assign detect_min[1][16] = (mid_1[23:16] < mid_2[31:24]) ? 1 : 0;
assign detect_min[1][17] = (mid_1[23:16] < btm_0[15:8]) ? 1 : 0;
assign detect_min[1][18] = (mid_1[23:16] < btm_0[23:16]) ? 1 : 0;
assign detect_min[1][19] = (mid_1[23:16] < btm_0[31:24]) ? 1 : 0;
assign detect_min[1][20] = (mid_1[23:16] < btm_1[15:8]) ? 1 : 0;
assign detect_min[1][21] = (mid_1[23:16] < btm_1[23:16]) ? 1 : 0;
assign detect_min[1][22] = (mid_1[23:16] < btm_1[31:24]) ? 1 : 0;
assign detect_min[1][23] = (mid_1[23:16] < btm_2[15:8]) ? 1 : 0;
assign detect_min[1][24] = (mid_1[23:16] < btm_2[23:16]) ? 1 : 0;
assign detect_min[1][25] = (mid_1[23:16] < btm_2[31:24]) ? 1 : 0;

assign detect_min[2][0] = (mid_1[31:24] < top_0[23:16]) ? 1 : 0;
assign detect_min[2][1] = (mid_1[31:24] < top_0[31:24]) ? 1 : 0;
assign detect_min[2][2] = (mid_1[31:24] < top_0[39:32]) ? 1 : 0;
assign detect_min[2][3] = (mid_1[31:24] < top_1[23:16]) ? 1 : 0;
assign detect_min[2][4] = (mid_1[31:24] < top_1[31:24]) ? 1 : 0;
assign detect_min[2][5] = (mid_1[31:24] < top_1[39:32]) ? 1 : 0;
assign detect_min[2][6] = (mid_1[31:24] < top_2[23:16]) ? 1 : 0;
assign detect_min[2][7] = (mid_1[31:24] < top_2[31:24]) ? 1 : 0;
assign detect_min[2][8] = (mid_1[31:24] < top_2[39:32]) ? 1 : 0;
assign detect_min[2][9] = (mid_1[31:24] < mid_0[23:16]) ? 1 : 0;
assign detect_min[2][10] = (mid_1[31:24] < mid_0[31:24]) ? 1 : 0;
assign detect_min[2][11] = (mid_1[31:24] < mid_0[39:32]) ? 1 : 0;
assign detect_min[2][12] = (mid_1[31:24] < mid_1[23:16]) ? 1 : 0;
assign detect_min[2][13] = (mid_1[31:24] < mid_1[39:32]) ? 1 : 0;
assign detect_min[2][14] = (mid_1[31:24] < mid_2[23:16]) ? 1 : 0;
assign detect_min[2][15] = (mid_1[31:24] < mid_2[31:24]) ? 1 : 0;
assign detect_min[2][16] = (mid_1[31:24] < mid_2[39:32]) ? 1 : 0;
assign detect_min[2][17] = (mid_1[31:24] < btm_0[23:16]) ? 1 : 0;
assign detect_min[2][18] = (mid_1[31:24] < btm_0[31:24]) ? 1 : 0;
assign detect_min[2][19] = (mid_1[31:24] < btm_0[39:32]) ? 1 : 0;
assign detect_min[2][20] = (mid_1[31:24] < btm_1[23:16]) ? 1 : 0;
assign detect_min[2][21] = (mid_1[31:24] < btm_1[31:24]) ? 1 : 0;
assign detect_min[2][22] = (mid_1[31:24] < btm_1[39:32]) ? 1 : 0;
assign detect_min[2][23] = (mid_1[31:24] < btm_2[23:16]) ? 1 : 0;
assign detect_min[2][24] = (mid_1[31:24] < btm_2[31:24]) ? 1 : 0;
assign detect_min[2][25] = (mid_1[31:24] < btm_2[39:32]) ? 1 : 0;

assign detect_min[3][0] = (mid_1[39:32] < top_0[31:24]) ? 1 : 0;
assign detect_min[3][1] = (mid_1[39:32] < top_0[39:32]) ? 1 : 0;
assign detect_min[3][2] = (mid_1[39:32] < top_0[47:40]) ? 1 : 0;
assign detect_min[3][3] = (mid_1[39:32] < top_1[31:24]) ? 1 : 0;
assign detect_min[3][4] = (mid_1[39:32] < top_1[39:32]) ? 1 : 0;
assign detect_min[3][5] = (mid_1[39:32] < top_1[47:40]) ? 1 : 0;
assign detect_min[3][6] = (mid_1[39:32] < top_2[31:24]) ? 1 : 0;
assign detect_min[3][7] = (mid_1[39:32] < top_2[39:32]) ? 1 : 0;
assign detect_min[3][8] = (mid_1[39:32] < top_2[47:40]) ? 1 : 0;
assign detect_min[3][9] = (mid_1[39:32] < mid_0[31:24]) ? 1 : 0;
assign detect_min[3][10] = (mid_1[39:32] < mid_0[39:32]) ? 1 : 0;
assign detect_min[3][11] = (mid_1[39:32] < mid_0[47:40]) ? 1 : 0;
assign detect_min[3][12] = (mid_1[39:32] < mid_1[31:24]) ? 1 : 0;
assign detect_min[3][13] = (mid_1[39:32] < mid_1[47:40]) ? 1 : 0;
assign detect_min[3][14] = (mid_1[39:32] < mid_2[31:24]) ? 1 : 0;
assign detect_min[3][15] = (mid_1[39:32] < mid_2[39:32]) ? 1 : 0;
assign detect_min[3][16] = (mid_1[39:32] < mid_2[47:40]) ? 1 : 0;
assign detect_min[3][17] = (mid_1[39:32] < btm_0[31:24]) ? 1 : 0;
assign detect_min[3][18] = (mid_1[39:32] < btm_0[39:32]) ? 1 : 0;
assign detect_min[3][19] = (mid_1[39:32] < btm_0[47:40]) ? 1 : 0;
assign detect_min[3][20] = (mid_1[39:32] < btm_1[31:24]) ? 1 : 0;
assign detect_min[3][21] = (mid_1[39:32] < btm_1[39:32]) ? 1 : 0;
assign detect_min[3][22] = (mid_1[39:32] < btm_1[47:40]) ? 1 : 0;
assign detect_min[3][23] = (mid_1[39:32] < btm_2[31:24]) ? 1 : 0;
assign detect_min[3][24] = (mid_1[39:32] < btm_2[39:32]) ? 1 : 0;
assign detect_min[3][25] = (mid_1[39:32] < btm_2[47:40]) ? 1 : 0;

assign detect_min[4][0] = (mid_1[47:40] < top_0[39:32]) ? 1 : 0;
assign detect_min[4][1] = (mid_1[47:40] < top_0[47:40]) ? 1 : 0;
assign detect_min[4][2] = (mid_1[47:40] < top_0[55:48]) ? 1 : 0;
assign detect_min[4][3] = (mid_1[47:40] < top_1[39:32]) ? 1 : 0;
assign detect_min[4][4] = (mid_1[47:40] < top_1[47:40]) ? 1 : 0;
assign detect_min[4][5] = (mid_1[47:40] < top_1[55:48]) ? 1 : 0;
assign detect_min[4][6] = (mid_1[47:40] < top_2[39:32]) ? 1 : 0;
assign detect_min[4][7] = (mid_1[47:40] < top_2[47:40]) ? 1 : 0;
assign detect_min[4][8] = (mid_1[47:40] < top_2[55:48]) ? 1 : 0;
assign detect_min[4][9] = (mid_1[47:40] < mid_0[39:32]) ? 1 : 0;
assign detect_min[4][10] = (mid_1[47:40] < mid_0[47:40]) ? 1 : 0;
assign detect_min[4][11] = (mid_1[47:40] < mid_0[55:48]) ? 1 : 0;
assign detect_min[4][12] = (mid_1[47:40] < mid_1[39:32]) ? 1 : 0;
assign detect_min[4][13] = (mid_1[47:40] < mid_1[55:48]) ? 1 : 0;
assign detect_min[4][14] = (mid_1[47:40] < mid_2[39:32]) ? 1 : 0;
assign detect_min[4][15] = (mid_1[47:40] < mid_2[47:40]) ? 1 : 0;
assign detect_min[4][16] = (mid_1[47:40] < mid_2[55:48]) ? 1 : 0;
assign detect_min[4][17] = (mid_1[47:40] < btm_0[39:32]) ? 1 : 0;
assign detect_min[4][18] = (mid_1[47:40] < btm_0[47:40]) ? 1 : 0;
assign detect_min[4][19] = (mid_1[47:40] < btm_0[55:48]) ? 1 : 0;
assign detect_min[4][20] = (mid_1[47:40] < btm_1[39:32]) ? 1 : 0;
assign detect_min[4][21] = (mid_1[47:40] < btm_1[47:40]) ? 1 : 0;
assign detect_min[4][22] = (mid_1[47:40] < btm_1[55:48]) ? 1 : 0;
assign detect_min[4][23] = (mid_1[47:40] < btm_2[39:32]) ? 1 : 0;
assign detect_min[4][24] = (mid_1[47:40] < btm_2[47:40]) ? 1 : 0;
assign detect_min[4][25] = (mid_1[47:40] < btm_2[55:48]) ? 1 : 0;

assign detect_min[5][0] = (mid_1[55:48] < top_0[47:40]) ? 1 : 0;
assign detect_min[5][1] = (mid_1[55:48] < top_0[55:48]) ? 1 : 0;
assign detect_min[5][2] = (mid_1[55:48] < top_0[63:56]) ? 1 : 0;
assign detect_min[5][3] = (mid_1[55:48] < top_1[47:40]) ? 1 : 0;
assign detect_min[5][4] = (mid_1[55:48] < top_1[55:48]) ? 1 : 0;
assign detect_min[5][5] = (mid_1[55:48] < top_1[63:56]) ? 1 : 0;
assign detect_min[5][6] = (mid_1[55:48] < top_2[47:40]) ? 1 : 0;
assign detect_min[5][7] = (mid_1[55:48] < top_2[55:48]) ? 1 : 0;
assign detect_min[5][8] = (mid_1[55:48] < top_2[63:56]) ? 1 : 0;
assign detect_min[5][9] = (mid_1[55:48] < mid_0[47:40]) ? 1 : 0;
assign detect_min[5][10] = (mid_1[55:48] < mid_0[55:48]) ? 1 : 0;
assign detect_min[5][11] = (mid_1[55:48] < mid_0[63:56]) ? 1 : 0;
assign detect_min[5][12] = (mid_1[55:48] < mid_1[47:40]) ? 1 : 0;
assign detect_min[5][13] = (mid_1[55:48] < mid_1[63:56]) ? 1 : 0;
assign detect_min[5][14] = (mid_1[55:48] < mid_2[47:40]) ? 1 : 0;
assign detect_min[5][15] = (mid_1[55:48] < mid_2[55:48]) ? 1 : 0;
assign detect_min[5][16] = (mid_1[55:48] < mid_2[63:56]) ? 1 : 0;
assign detect_min[5][17] = (mid_1[55:48] < btm_0[47:40]) ? 1 : 0;
assign detect_min[5][18] = (mid_1[55:48] < btm_0[55:48]) ? 1 : 0;
assign detect_min[5][19] = (mid_1[55:48] < btm_0[63:56]) ? 1 : 0;
assign detect_min[5][20] = (mid_1[55:48] < btm_1[47:40]) ? 1 : 0;
assign detect_min[5][21] = (mid_1[55:48] < btm_1[55:48]) ? 1 : 0;
assign detect_min[5][22] = (mid_1[55:48] < btm_1[63:56]) ? 1 : 0;
assign detect_min[5][23] = (mid_1[55:48] < btm_2[47:40]) ? 1 : 0;
assign detect_min[5][24] = (mid_1[55:48] < btm_2[55:48]) ? 1 : 0;
assign detect_min[5][25] = (mid_1[55:48] < btm_2[63:56]) ? 1 : 0;

assign detect_min[6][0] = (mid_1[63:56] < top_0[55:48]) ? 1 : 0;
assign detect_min[6][1] = (mid_1[63:56] < top_0[63:56]) ? 1 : 0;
assign detect_min[6][2] = (mid_1[63:56] < top_0[71:64]) ? 1 : 0;
assign detect_min[6][3] = (mid_1[63:56] < top_1[55:48]) ? 1 : 0;
assign detect_min[6][4] = (mid_1[63:56] < top_1[63:56]) ? 1 : 0;
assign detect_min[6][5] = (mid_1[63:56] < top_1[71:64]) ? 1 : 0;
assign detect_min[6][6] = (mid_1[63:56] < top_2[55:48]) ? 1 : 0;
assign detect_min[6][7] = (mid_1[63:56] < top_2[63:56]) ? 1 : 0;
assign detect_min[6][8] = (mid_1[63:56] < top_2[71:64]) ? 1 : 0;
assign detect_min[6][9] = (mid_1[63:56] < mid_0[55:48]) ? 1 : 0;
assign detect_min[6][10] = (mid_1[63:56] < mid_0[63:56]) ? 1 : 0;
assign detect_min[6][11] = (mid_1[63:56] < mid_0[71:64]) ? 1 : 0;
assign detect_min[6][12] = (mid_1[63:56] < mid_1[55:48]) ? 1 : 0;
assign detect_min[6][13] = (mid_1[63:56] < mid_1[71:64]) ? 1 : 0;
assign detect_min[6][14] = (mid_1[63:56] < mid_2[55:48]) ? 1 : 0;
assign detect_min[6][15] = (mid_1[63:56] < mid_2[63:56]) ? 1 : 0;
assign detect_min[6][16] = (mid_1[63:56] < mid_2[71:64]) ? 1 : 0;
assign detect_min[6][17] = (mid_1[63:56] < btm_0[55:48]) ? 1 : 0;
assign detect_min[6][18] = (mid_1[63:56] < btm_0[63:56]) ? 1 : 0;
assign detect_min[6][19] = (mid_1[63:56] < btm_0[71:64]) ? 1 : 0;
assign detect_min[6][20] = (mid_1[63:56] < btm_1[55:48]) ? 1 : 0;
assign detect_min[6][21] = (mid_1[63:56] < btm_1[63:56]) ? 1 : 0;
assign detect_min[6][22] = (mid_1[63:56] < btm_1[71:64]) ? 1 : 0;
assign detect_min[6][23] = (mid_1[63:56] < btm_2[55:48]) ? 1 : 0;
assign detect_min[6][24] = (mid_1[63:56] < btm_2[63:56]) ? 1 : 0;
assign detect_min[6][25] = (mid_1[63:56] < btm_2[71:64]) ? 1 : 0;

assign detect_min[7][0] = (mid_1[71:64] < top_0[63:56]) ? 1 : 0;
assign detect_min[7][1] = (mid_1[71:64] < top_0[71:64]) ? 1 : 0;
assign detect_min[7][2] = (mid_1[71:64] < top_0[79:72]) ? 1 : 0;
assign detect_min[7][3] = (mid_1[71:64] < top_1[63:56]) ? 1 : 0;
assign detect_min[7][4] = (mid_1[71:64] < top_1[71:64]) ? 1 : 0;
assign detect_min[7][5] = (mid_1[71:64] < top_1[79:72]) ? 1 : 0;
assign detect_min[7][6] = (mid_1[71:64] < top_2[63:56]) ? 1 : 0;
assign detect_min[7][7] = (mid_1[71:64] < top_2[71:64]) ? 1 : 0;
assign detect_min[7][8] = (mid_1[71:64] < top_2[79:72]) ? 1 : 0;
assign detect_min[7][9] = (mid_1[71:64] < mid_0[63:56]) ? 1 : 0;
assign detect_min[7][10] = (mid_1[71:64] < mid_0[71:64]) ? 1 : 0;
assign detect_min[7][11] = (mid_1[71:64] < mid_0[79:72]) ? 1 : 0;
assign detect_min[7][12] = (mid_1[71:64] < mid_1[63:56]) ? 1 : 0;
assign detect_min[7][13] = (mid_1[71:64] < mid_1[79:72]) ? 1 : 0;
assign detect_min[7][14] = (mid_1[71:64] < mid_2[63:56]) ? 1 : 0;
assign detect_min[7][15] = (mid_1[71:64] < mid_2[71:64]) ? 1 : 0;
assign detect_min[7][16] = (mid_1[71:64] < mid_2[79:72]) ? 1 : 0;
assign detect_min[7][17] = (mid_1[71:64] < btm_0[63:56]) ? 1 : 0;
assign detect_min[7][18] = (mid_1[71:64] < btm_0[71:64]) ? 1 : 0;
assign detect_min[7][19] = (mid_1[71:64] < btm_0[79:72]) ? 1 : 0;
assign detect_min[7][20] = (mid_1[71:64] < btm_1[63:56]) ? 1 : 0;
assign detect_min[7][21] = (mid_1[71:64] < btm_1[71:64]) ? 1 : 0;
assign detect_min[7][22] = (mid_1[71:64] < btm_1[79:72]) ? 1 : 0;
assign detect_min[7][23] = (mid_1[71:64] < btm_2[63:56]) ? 1 : 0;
assign detect_min[7][24] = (mid_1[71:64] < btm_2[71:64]) ? 1 : 0;
assign detect_min[7][25] = (mid_1[71:64] < btm_2[79:72]) ? 1 : 0;

assign detect_min[8][0] = (mid_1[79:72] < top_0[71:64]) ? 1 : 0;
assign detect_min[8][1] = (mid_1[79:72] < top_0[79:72]) ? 1 : 0;
assign detect_min[8][2] = (mid_1[79:72] < top_0[87:80]) ? 1 : 0;
assign detect_min[8][3] = (mid_1[79:72] < top_1[71:64]) ? 1 : 0;
assign detect_min[8][4] = (mid_1[79:72] < top_1[79:72]) ? 1 : 0;
assign detect_min[8][5] = (mid_1[79:72] < top_1[87:80]) ? 1 : 0;
assign detect_min[8][6] = (mid_1[79:72] < top_2[71:64]) ? 1 : 0;
assign detect_min[8][7] = (mid_1[79:72] < top_2[79:72]) ? 1 : 0;
assign detect_min[8][8] = (mid_1[79:72] < top_2[87:80]) ? 1 : 0;
assign detect_min[8][9] = (mid_1[79:72] < mid_0[71:64]) ? 1 : 0;
assign detect_min[8][10] = (mid_1[79:72] < mid_0[79:72]) ? 1 : 0;
assign detect_min[8][11] = (mid_1[79:72] < mid_0[87:80]) ? 1 : 0;
assign detect_min[8][12] = (mid_1[79:72] < mid_1[71:64]) ? 1 : 0;
assign detect_min[8][13] = (mid_1[79:72] < mid_1[87:80]) ? 1 : 0;
assign detect_min[8][14] = (mid_1[79:72] < mid_2[71:64]) ? 1 : 0;
assign detect_min[8][15] = (mid_1[79:72] < mid_2[79:72]) ? 1 : 0;
assign detect_min[8][16] = (mid_1[79:72] < mid_2[87:80]) ? 1 : 0;
assign detect_min[8][17] = (mid_1[79:72] < btm_0[71:64]) ? 1 : 0;
assign detect_min[8][18] = (mid_1[79:72] < btm_0[79:72]) ? 1 : 0;
assign detect_min[8][19] = (mid_1[79:72] < btm_0[87:80]) ? 1 : 0;
assign detect_min[8][20] = (mid_1[79:72] < btm_1[71:64]) ? 1 : 0;
assign detect_min[8][21] = (mid_1[79:72] < btm_1[79:72]) ? 1 : 0;
assign detect_min[8][22] = (mid_1[79:72] < btm_1[87:80]) ? 1 : 0;
assign detect_min[8][23] = (mid_1[79:72] < btm_2[71:64]) ? 1 : 0;
assign detect_min[8][24] = (mid_1[79:72] < btm_2[79:72]) ? 1 : 0;
assign detect_min[8][25] = (mid_1[79:72] < btm_2[87:80]) ? 1 : 0;

assign detect_min[9][0] = (mid_1[87:80] < top_0[79:72]) ? 1 : 0;
assign detect_min[9][1] = (mid_1[87:80] < top_0[87:80]) ? 1 : 0;
assign detect_min[9][2] = (mid_1[87:80] < top_0[95:88]) ? 1 : 0;
assign detect_min[9][3] = (mid_1[87:80] < top_1[79:72]) ? 1 : 0;
assign detect_min[9][4] = (mid_1[87:80] < top_1[87:80]) ? 1 : 0;
assign detect_min[9][5] = (mid_1[87:80] < top_1[95:88]) ? 1 : 0;
assign detect_min[9][6] = (mid_1[87:80] < top_2[79:72]) ? 1 : 0;
assign detect_min[9][7] = (mid_1[87:80] < top_2[87:80]) ? 1 : 0;
assign detect_min[9][8] = (mid_1[87:80] < top_2[95:88]) ? 1 : 0;
assign detect_min[9][9] = (mid_1[87:80] < mid_0[79:72]) ? 1 : 0;
assign detect_min[9][10] = (mid_1[87:80] < mid_0[87:80]) ? 1 : 0;
assign detect_min[9][11] = (mid_1[87:80] < mid_0[95:88]) ? 1 : 0;
assign detect_min[9][12] = (mid_1[87:80] < mid_1[79:72]) ? 1 : 0;
assign detect_min[9][13] = (mid_1[87:80] < mid_1[95:88]) ? 1 : 0;
assign detect_min[9][14] = (mid_1[87:80] < mid_2[79:72]) ? 1 : 0;
assign detect_min[9][15] = (mid_1[87:80] < mid_2[87:80]) ? 1 : 0;
assign detect_min[9][16] = (mid_1[87:80] < mid_2[95:88]) ? 1 : 0;
assign detect_min[9][17] = (mid_1[87:80] < btm_0[79:72]) ? 1 : 0;
assign detect_min[9][18] = (mid_1[87:80] < btm_0[87:80]) ? 1 : 0;
assign detect_min[9][19] = (mid_1[87:80] < btm_0[95:88]) ? 1 : 0;
assign detect_min[9][20] = (mid_1[87:80] < btm_1[79:72]) ? 1 : 0;
assign detect_min[9][21] = (mid_1[87:80] < btm_1[87:80]) ? 1 : 0;
assign detect_min[9][22] = (mid_1[87:80] < btm_1[95:88]) ? 1 : 0;
assign detect_min[9][23] = (mid_1[87:80] < btm_2[79:72]) ? 1 : 0;
assign detect_min[9][24] = (mid_1[87:80] < btm_2[87:80]) ? 1 : 0;
assign detect_min[9][25] = (mid_1[87:80] < btm_2[95:88]) ? 1 : 0;

assign detect_min[10][0] = (mid_1[95:88] < top_0[87:80]) ? 1 : 0;
assign detect_min[10][1] = (mid_1[95:88] < top_0[95:88]) ? 1 : 0;
assign detect_min[10][2] = (mid_1[95:88] < top_0[103:96]) ? 1 : 0;
assign detect_min[10][3] = (mid_1[95:88] < top_1[87:80]) ? 1 : 0;
assign detect_min[10][4] = (mid_1[95:88] < top_1[95:88]) ? 1 : 0;
assign detect_min[10][5] = (mid_1[95:88] < top_1[103:96]) ? 1 : 0;
assign detect_min[10][6] = (mid_1[95:88] < top_2[87:80]) ? 1 : 0;
assign detect_min[10][7] = (mid_1[95:88] < top_2[95:88]) ? 1 : 0;
assign detect_min[10][8] = (mid_1[95:88] < top_2[103:96]) ? 1 : 0;
assign detect_min[10][9] = (mid_1[95:88] < mid_0[87:80]) ? 1 : 0;
assign detect_min[10][10] = (mid_1[95:88] < mid_0[95:88]) ? 1 : 0;
assign detect_min[10][11] = (mid_1[95:88] < mid_0[103:96]) ? 1 : 0;
assign detect_min[10][12] = (mid_1[95:88] < mid_1[87:80]) ? 1 : 0;
assign detect_min[10][13] = (mid_1[95:88] < mid_1[103:96]) ? 1 : 0;
assign detect_min[10][14] = (mid_1[95:88] < mid_2[87:80]) ? 1 : 0;
assign detect_min[10][15] = (mid_1[95:88] < mid_2[95:88]) ? 1 : 0;
assign detect_min[10][16] = (mid_1[95:88] < mid_2[103:96]) ? 1 : 0;
assign detect_min[10][17] = (mid_1[95:88] < btm_0[87:80]) ? 1 : 0;
assign detect_min[10][18] = (mid_1[95:88] < btm_0[95:88]) ? 1 : 0;
assign detect_min[10][19] = (mid_1[95:88] < btm_0[103:96]) ? 1 : 0;
assign detect_min[10][20] = (mid_1[95:88] < btm_1[87:80]) ? 1 : 0;
assign detect_min[10][21] = (mid_1[95:88] < btm_1[95:88]) ? 1 : 0;
assign detect_min[10][22] = (mid_1[95:88] < btm_1[103:96]) ? 1 : 0;
assign detect_min[10][23] = (mid_1[95:88] < btm_2[87:80]) ? 1 : 0;
assign detect_min[10][24] = (mid_1[95:88] < btm_2[95:88]) ? 1 : 0;
assign detect_min[10][25] = (mid_1[95:88] < btm_2[103:96]) ? 1 : 0;

assign detect_min[11][0] = (mid_1[103:96] < top_0[95:88]) ? 1 : 0;
assign detect_min[11][1] = (mid_1[103:96] < top_0[103:96]) ? 1 : 0;
assign detect_min[11][2] = (mid_1[103:96] < top_0[111:104]) ? 1 : 0;
assign detect_min[11][3] = (mid_1[103:96] < top_1[95:88]) ? 1 : 0;
assign detect_min[11][4] = (mid_1[103:96] < top_1[103:96]) ? 1 : 0;
assign detect_min[11][5] = (mid_1[103:96] < top_1[111:104]) ? 1 : 0;
assign detect_min[11][6] = (mid_1[103:96] < top_2[95:88]) ? 1 : 0;
assign detect_min[11][7] = (mid_1[103:96] < top_2[103:96]) ? 1 : 0;
assign detect_min[11][8] = (mid_1[103:96] < top_2[111:104]) ? 1 : 0;
assign detect_min[11][9] = (mid_1[103:96] < mid_0[95:88]) ? 1 : 0;
assign detect_min[11][10] = (mid_1[103:96] < mid_0[103:96]) ? 1 : 0;
assign detect_min[11][11] = (mid_1[103:96] < mid_0[111:104]) ? 1 : 0;
assign detect_min[11][12] = (mid_1[103:96] < mid_1[95:88]) ? 1 : 0;
assign detect_min[11][13] = (mid_1[103:96] < mid_1[111:104]) ? 1 : 0;
assign detect_min[11][14] = (mid_1[103:96] < mid_2[95:88]) ? 1 : 0;
assign detect_min[11][15] = (mid_1[103:96] < mid_2[103:96]) ? 1 : 0;
assign detect_min[11][16] = (mid_1[103:96] < mid_2[111:104]) ? 1 : 0;
assign detect_min[11][17] = (mid_1[103:96] < btm_0[95:88]) ? 1 : 0;
assign detect_min[11][18] = (mid_1[103:96] < btm_0[103:96]) ? 1 : 0;
assign detect_min[11][19] = (mid_1[103:96] < btm_0[111:104]) ? 1 : 0;
assign detect_min[11][20] = (mid_1[103:96] < btm_1[95:88]) ? 1 : 0;
assign detect_min[11][21] = (mid_1[103:96] < btm_1[103:96]) ? 1 : 0;
assign detect_min[11][22] = (mid_1[103:96] < btm_1[111:104]) ? 1 : 0;
assign detect_min[11][23] = (mid_1[103:96] < btm_2[95:88]) ? 1 : 0;
assign detect_min[11][24] = (mid_1[103:96] < btm_2[103:96]) ? 1 : 0;
assign detect_min[11][25] = (mid_1[103:96] < btm_2[111:104]) ? 1 : 0;

assign detect_min[12][0] = (mid_1[111:104] < top_0[103:96]) ? 1 : 0;
assign detect_min[12][1] = (mid_1[111:104] < top_0[111:104]) ? 1 : 0;
assign detect_min[12][2] = (mid_1[111:104] < top_0[119:112]) ? 1 : 0;
assign detect_min[12][3] = (mid_1[111:104] < top_1[103:96]) ? 1 : 0;
assign detect_min[12][4] = (mid_1[111:104] < top_1[111:104]) ? 1 : 0;
assign detect_min[12][5] = (mid_1[111:104] < top_1[119:112]) ? 1 : 0;
assign detect_min[12][6] = (mid_1[111:104] < top_2[103:96]) ? 1 : 0;
assign detect_min[12][7] = (mid_1[111:104] < top_2[111:104]) ? 1 : 0;
assign detect_min[12][8] = (mid_1[111:104] < top_2[119:112]) ? 1 : 0;
assign detect_min[12][9] = (mid_1[111:104] < mid_0[103:96]) ? 1 : 0;
assign detect_min[12][10] = (mid_1[111:104] < mid_0[111:104]) ? 1 : 0;
assign detect_min[12][11] = (mid_1[111:104] < mid_0[119:112]) ? 1 : 0;
assign detect_min[12][12] = (mid_1[111:104] < mid_1[103:96]) ? 1 : 0;
assign detect_min[12][13] = (mid_1[111:104] < mid_1[119:112]) ? 1 : 0;
assign detect_min[12][14] = (mid_1[111:104] < mid_2[103:96]) ? 1 : 0;
assign detect_min[12][15] = (mid_1[111:104] < mid_2[111:104]) ? 1 : 0;
assign detect_min[12][16] = (mid_1[111:104] < mid_2[119:112]) ? 1 : 0;
assign detect_min[12][17] = (mid_1[111:104] < btm_0[103:96]) ? 1 : 0;
assign detect_min[12][18] = (mid_1[111:104] < btm_0[111:104]) ? 1 : 0;
assign detect_min[12][19] = (mid_1[111:104] < btm_0[119:112]) ? 1 : 0;
assign detect_min[12][20] = (mid_1[111:104] < btm_1[103:96]) ? 1 : 0;
assign detect_min[12][21] = (mid_1[111:104] < btm_1[111:104]) ? 1 : 0;
assign detect_min[12][22] = (mid_1[111:104] < btm_1[119:112]) ? 1 : 0;
assign detect_min[12][23] = (mid_1[111:104] < btm_2[103:96]) ? 1 : 0;
assign detect_min[12][24] = (mid_1[111:104] < btm_2[111:104]) ? 1 : 0;
assign detect_min[12][25] = (mid_1[111:104] < btm_2[119:112]) ? 1 : 0;

assign detect_min[13][0] = (mid_1[119:112] < top_0[111:104]) ? 1 : 0;
assign detect_min[13][1] = (mid_1[119:112] < top_0[119:112]) ? 1 : 0;
assign detect_min[13][2] = (mid_1[119:112] < top_0[127:120]) ? 1 : 0;
assign detect_min[13][3] = (mid_1[119:112] < top_1[111:104]) ? 1 : 0;
assign detect_min[13][4] = (mid_1[119:112] < top_1[119:112]) ? 1 : 0;
assign detect_min[13][5] = (mid_1[119:112] < top_1[127:120]) ? 1 : 0;
assign detect_min[13][6] = (mid_1[119:112] < top_2[111:104]) ? 1 : 0;
assign detect_min[13][7] = (mid_1[119:112] < top_2[119:112]) ? 1 : 0;
assign detect_min[13][8] = (mid_1[119:112] < top_2[127:120]) ? 1 : 0;
assign detect_min[13][9] = (mid_1[119:112] < mid_0[111:104]) ? 1 : 0;
assign detect_min[13][10] = (mid_1[119:112] < mid_0[119:112]) ? 1 : 0;
assign detect_min[13][11] = (mid_1[119:112] < mid_0[127:120]) ? 1 : 0;
assign detect_min[13][12] = (mid_1[119:112] < mid_1[111:104]) ? 1 : 0;
assign detect_min[13][13] = (mid_1[119:112] < mid_1[127:120]) ? 1 : 0;
assign detect_min[13][14] = (mid_1[119:112] < mid_2[111:104]) ? 1 : 0;
assign detect_min[13][15] = (mid_1[119:112] < mid_2[119:112]) ? 1 : 0;
assign detect_min[13][16] = (mid_1[119:112] < mid_2[127:120]) ? 1 : 0;
assign detect_min[13][17] = (mid_1[119:112] < btm_0[111:104]) ? 1 : 0;
assign detect_min[13][18] = (mid_1[119:112] < btm_0[119:112]) ? 1 : 0;
assign detect_min[13][19] = (mid_1[119:112] < btm_0[127:120]) ? 1 : 0;
assign detect_min[13][20] = (mid_1[119:112] < btm_1[111:104]) ? 1 : 0;
assign detect_min[13][21] = (mid_1[119:112] < btm_1[119:112]) ? 1 : 0;
assign detect_min[13][22] = (mid_1[119:112] < btm_1[127:120]) ? 1 : 0;
assign detect_min[13][23] = (mid_1[119:112] < btm_2[111:104]) ? 1 : 0;
assign detect_min[13][24] = (mid_1[119:112] < btm_2[119:112]) ? 1 : 0;
assign detect_min[13][25] = (mid_1[119:112] < btm_2[127:120]) ? 1 : 0;

assign detect_min[14][0] = (mid_1[127:120] < top_0[119:112]) ? 1 : 0;
assign detect_min[14][1] = (mid_1[127:120] < top_0[127:120]) ? 1 : 0;
assign detect_min[14][2] = (mid_1[127:120] < top_0[135:128]) ? 1 : 0;
assign detect_min[14][3] = (mid_1[127:120] < top_1[119:112]) ? 1 : 0;
assign detect_min[14][4] = (mid_1[127:120] < top_1[127:120]) ? 1 : 0;
assign detect_min[14][5] = (mid_1[127:120] < top_1[135:128]) ? 1 : 0;
assign detect_min[14][6] = (mid_1[127:120] < top_2[119:112]) ? 1 : 0;
assign detect_min[14][7] = (mid_1[127:120] < top_2[127:120]) ? 1 : 0;
assign detect_min[14][8] = (mid_1[127:120] < top_2[135:128]) ? 1 : 0;
assign detect_min[14][9] = (mid_1[127:120] < mid_0[119:112]) ? 1 : 0;
assign detect_min[14][10] = (mid_1[127:120] < mid_0[127:120]) ? 1 : 0;
assign detect_min[14][11] = (mid_1[127:120] < mid_0[135:128]) ? 1 : 0;
assign detect_min[14][12] = (mid_1[127:120] < mid_1[119:112]) ? 1 : 0;
assign detect_min[14][13] = (mid_1[127:120] < mid_1[135:128]) ? 1 : 0;
assign detect_min[14][14] = (mid_1[127:120] < mid_2[119:112]) ? 1 : 0;
assign detect_min[14][15] = (mid_1[127:120] < mid_2[127:120]) ? 1 : 0;
assign detect_min[14][16] = (mid_1[127:120] < mid_2[135:128]) ? 1 : 0;
assign detect_min[14][17] = (mid_1[127:120] < btm_0[119:112]) ? 1 : 0;
assign detect_min[14][18] = (mid_1[127:120] < btm_0[127:120]) ? 1 : 0;
assign detect_min[14][19] = (mid_1[127:120] < btm_0[135:128]) ? 1 : 0;
assign detect_min[14][20] = (mid_1[127:120] < btm_1[119:112]) ? 1 : 0;
assign detect_min[14][21] = (mid_1[127:120] < btm_1[127:120]) ? 1 : 0;
assign detect_min[14][22] = (mid_1[127:120] < btm_1[135:128]) ? 1 : 0;
assign detect_min[14][23] = (mid_1[127:120] < btm_2[119:112]) ? 1 : 0;
assign detect_min[14][24] = (mid_1[127:120] < btm_2[127:120]) ? 1 : 0;
assign detect_min[14][25] = (mid_1[127:120] < btm_2[135:128]) ? 1 : 0;

assign detect_min[15][0] = (mid_1[135:128] < top_0[127:120]) ? 1 : 0;
assign detect_min[15][1] = (mid_1[135:128] < top_0[135:128]) ? 1 : 0;
assign detect_min[15][2] = (mid_1[135:128] < top_0[143:136]) ? 1 : 0;
assign detect_min[15][3] = (mid_1[135:128] < top_1[127:120]) ? 1 : 0;
assign detect_min[15][4] = (mid_1[135:128] < top_1[135:128]) ? 1 : 0;
assign detect_min[15][5] = (mid_1[135:128] < top_1[143:136]) ? 1 : 0;
assign detect_min[15][6] = (mid_1[135:128] < top_2[127:120]) ? 1 : 0;
assign detect_min[15][7] = (mid_1[135:128] < top_2[135:128]) ? 1 : 0;
assign detect_min[15][8] = (mid_1[135:128] < top_2[143:136]) ? 1 : 0;
assign detect_min[15][9] = (mid_1[135:128] < mid_0[127:120]) ? 1 : 0;
assign detect_min[15][10] = (mid_1[135:128] < mid_0[135:128]) ? 1 : 0;
assign detect_min[15][11] = (mid_1[135:128] < mid_0[143:136]) ? 1 : 0;
assign detect_min[15][12] = (mid_1[135:128] < mid_1[127:120]) ? 1 : 0;
assign detect_min[15][13] = (mid_1[135:128] < mid_1[143:136]) ? 1 : 0;
assign detect_min[15][14] = (mid_1[135:128] < mid_2[127:120]) ? 1 : 0;
assign detect_min[15][15] = (mid_1[135:128] < mid_2[135:128]) ? 1 : 0;
assign detect_min[15][16] = (mid_1[135:128] < mid_2[143:136]) ? 1 : 0;
assign detect_min[15][17] = (mid_1[135:128] < btm_0[127:120]) ? 1 : 0;
assign detect_min[15][18] = (mid_1[135:128] < btm_0[135:128]) ? 1 : 0;
assign detect_min[15][19] = (mid_1[135:128] < btm_0[143:136]) ? 1 : 0;
assign detect_min[15][20] = (mid_1[135:128] < btm_1[127:120]) ? 1 : 0;
assign detect_min[15][21] = (mid_1[135:128] < btm_1[135:128]) ? 1 : 0;
assign detect_min[15][22] = (mid_1[135:128] < btm_1[143:136]) ? 1 : 0;
assign detect_min[15][23] = (mid_1[135:128] < btm_2[127:120]) ? 1 : 0;
assign detect_min[15][24] = (mid_1[135:128] < btm_2[135:128]) ? 1 : 0;
assign detect_min[15][25] = (mid_1[135:128] < btm_2[143:136]) ? 1 : 0;

assign detect_min[16][0] = (mid_1[143:136] < top_0[135:128]) ? 1 : 0;
assign detect_min[16][1] = (mid_1[143:136] < top_0[143:136]) ? 1 : 0;
assign detect_min[16][2] = (mid_1[143:136] < top_0[151:144]) ? 1 : 0;
assign detect_min[16][3] = (mid_1[143:136] < top_1[135:128]) ? 1 : 0;
assign detect_min[16][4] = (mid_1[143:136] < top_1[143:136]) ? 1 : 0;
assign detect_min[16][5] = (mid_1[143:136] < top_1[151:144]) ? 1 : 0;
assign detect_min[16][6] = (mid_1[143:136] < top_2[135:128]) ? 1 : 0;
assign detect_min[16][7] = (mid_1[143:136] < top_2[143:136]) ? 1 : 0;
assign detect_min[16][8] = (mid_1[143:136] < top_2[151:144]) ? 1 : 0;
assign detect_min[16][9] = (mid_1[143:136] < mid_0[135:128]) ? 1 : 0;
assign detect_min[16][10] = (mid_1[143:136] < mid_0[143:136]) ? 1 : 0;
assign detect_min[16][11] = (mid_1[143:136] < mid_0[151:144]) ? 1 : 0;
assign detect_min[16][12] = (mid_1[143:136] < mid_1[135:128]) ? 1 : 0;
assign detect_min[16][13] = (mid_1[143:136] < mid_1[151:144]) ? 1 : 0;
assign detect_min[16][14] = (mid_1[143:136] < mid_2[135:128]) ? 1 : 0;
assign detect_min[16][15] = (mid_1[143:136] < mid_2[143:136]) ? 1 : 0;
assign detect_min[16][16] = (mid_1[143:136] < mid_2[151:144]) ? 1 : 0;
assign detect_min[16][17] = (mid_1[143:136] < btm_0[135:128]) ? 1 : 0;
assign detect_min[16][18] = (mid_1[143:136] < btm_0[143:136]) ? 1 : 0;
assign detect_min[16][19] = (mid_1[143:136] < btm_0[151:144]) ? 1 : 0;
assign detect_min[16][20] = (mid_1[143:136] < btm_1[135:128]) ? 1 : 0;
assign detect_min[16][21] = (mid_1[143:136] < btm_1[143:136]) ? 1 : 0;
assign detect_min[16][22] = (mid_1[143:136] < btm_1[151:144]) ? 1 : 0;
assign detect_min[16][23] = (mid_1[143:136] < btm_2[135:128]) ? 1 : 0;
assign detect_min[16][24] = (mid_1[143:136] < btm_2[143:136]) ? 1 : 0;
assign detect_min[16][25] = (mid_1[143:136] < btm_2[151:144]) ? 1 : 0;

assign detect_min[17][0] = (mid_1[151:144] < top_0[143:136]) ? 1 : 0;
assign detect_min[17][1] = (mid_1[151:144] < top_0[151:144]) ? 1 : 0;
assign detect_min[17][2] = (mid_1[151:144] < top_0[159:152]) ? 1 : 0;
assign detect_min[17][3] = (mid_1[151:144] < top_1[143:136]) ? 1 : 0;
assign detect_min[17][4] = (mid_1[151:144] < top_1[151:144]) ? 1 : 0;
assign detect_min[17][5] = (mid_1[151:144] < top_1[159:152]) ? 1 : 0;
assign detect_min[17][6] = (mid_1[151:144] < top_2[143:136]) ? 1 : 0;
assign detect_min[17][7] = (mid_1[151:144] < top_2[151:144]) ? 1 : 0;
assign detect_min[17][8] = (mid_1[151:144] < top_2[159:152]) ? 1 : 0;
assign detect_min[17][9] = (mid_1[151:144] < mid_0[143:136]) ? 1 : 0;
assign detect_min[17][10] = (mid_1[151:144] < mid_0[151:144]) ? 1 : 0;
assign detect_min[17][11] = (mid_1[151:144] < mid_0[159:152]) ? 1 : 0;
assign detect_min[17][12] = (mid_1[151:144] < mid_1[143:136]) ? 1 : 0;
assign detect_min[17][13] = (mid_1[151:144] < mid_1[159:152]) ? 1 : 0;
assign detect_min[17][14] = (mid_1[151:144] < mid_2[143:136]) ? 1 : 0;
assign detect_min[17][15] = (mid_1[151:144] < mid_2[151:144]) ? 1 : 0;
assign detect_min[17][16] = (mid_1[151:144] < mid_2[159:152]) ? 1 : 0;
assign detect_min[17][17] = (mid_1[151:144] < btm_0[143:136]) ? 1 : 0;
assign detect_min[17][18] = (mid_1[151:144] < btm_0[151:144]) ? 1 : 0;
assign detect_min[17][19] = (mid_1[151:144] < btm_0[159:152]) ? 1 : 0;
assign detect_min[17][20] = (mid_1[151:144] < btm_1[143:136]) ? 1 : 0;
assign detect_min[17][21] = (mid_1[151:144] < btm_1[151:144]) ? 1 : 0;
assign detect_min[17][22] = (mid_1[151:144] < btm_1[159:152]) ? 1 : 0;
assign detect_min[17][23] = (mid_1[151:144] < btm_2[143:136]) ? 1 : 0;
assign detect_min[17][24] = (mid_1[151:144] < btm_2[151:144]) ? 1 : 0;
assign detect_min[17][25] = (mid_1[151:144] < btm_2[159:152]) ? 1 : 0;

assign detect_min[18][0] = (mid_1[159:152] < top_0[151:144]) ? 1 : 0;
assign detect_min[18][1] = (mid_1[159:152] < top_0[159:152]) ? 1 : 0;
assign detect_min[18][2] = (mid_1[159:152] < top_0[167:160]) ? 1 : 0;
assign detect_min[18][3] = (mid_1[159:152] < top_1[151:144]) ? 1 : 0;
assign detect_min[18][4] = (mid_1[159:152] < top_1[159:152]) ? 1 : 0;
assign detect_min[18][5] = (mid_1[159:152] < top_1[167:160]) ? 1 : 0;
assign detect_min[18][6] = (mid_1[159:152] < top_2[151:144]) ? 1 : 0;
assign detect_min[18][7] = (mid_1[159:152] < top_2[159:152]) ? 1 : 0;
assign detect_min[18][8] = (mid_1[159:152] < top_2[167:160]) ? 1 : 0;
assign detect_min[18][9] = (mid_1[159:152] < mid_0[151:144]) ? 1 : 0;
assign detect_min[18][10] = (mid_1[159:152] < mid_0[159:152]) ? 1 : 0;
assign detect_min[18][11] = (mid_1[159:152] < mid_0[167:160]) ? 1 : 0;
assign detect_min[18][12] = (mid_1[159:152] < mid_1[151:144]) ? 1 : 0;
assign detect_min[18][13] = (mid_1[159:152] < mid_1[167:160]) ? 1 : 0;
assign detect_min[18][14] = (mid_1[159:152] < mid_2[151:144]) ? 1 : 0;
assign detect_min[18][15] = (mid_1[159:152] < mid_2[159:152]) ? 1 : 0;
assign detect_min[18][16] = (mid_1[159:152] < mid_2[167:160]) ? 1 : 0;
assign detect_min[18][17] = (mid_1[159:152] < btm_0[151:144]) ? 1 : 0;
assign detect_min[18][18] = (mid_1[159:152] < btm_0[159:152]) ? 1 : 0;
assign detect_min[18][19] = (mid_1[159:152] < btm_0[167:160]) ? 1 : 0;
assign detect_min[18][20] = (mid_1[159:152] < btm_1[151:144]) ? 1 : 0;
assign detect_min[18][21] = (mid_1[159:152] < btm_1[159:152]) ? 1 : 0;
assign detect_min[18][22] = (mid_1[159:152] < btm_1[167:160]) ? 1 : 0;
assign detect_min[18][23] = (mid_1[159:152] < btm_2[151:144]) ? 1 : 0;
assign detect_min[18][24] = (mid_1[159:152] < btm_2[159:152]) ? 1 : 0;
assign detect_min[18][25] = (mid_1[159:152] < btm_2[167:160]) ? 1 : 0;

assign detect_min[19][0] = (mid_1[167:160] < top_0[159:152]) ? 1 : 0;
assign detect_min[19][1] = (mid_1[167:160] < top_0[167:160]) ? 1 : 0;
assign detect_min[19][2] = (mid_1[167:160] < top_0[175:168]) ? 1 : 0;
assign detect_min[19][3] = (mid_1[167:160] < top_1[159:152]) ? 1 : 0;
assign detect_min[19][4] = (mid_1[167:160] < top_1[167:160]) ? 1 : 0;
assign detect_min[19][5] = (mid_1[167:160] < top_1[175:168]) ? 1 : 0;
assign detect_min[19][6] = (mid_1[167:160] < top_2[159:152]) ? 1 : 0;
assign detect_min[19][7] = (mid_1[167:160] < top_2[167:160]) ? 1 : 0;
assign detect_min[19][8] = (mid_1[167:160] < top_2[175:168]) ? 1 : 0;
assign detect_min[19][9] = (mid_1[167:160] < mid_0[159:152]) ? 1 : 0;
assign detect_min[19][10] = (mid_1[167:160] < mid_0[167:160]) ? 1 : 0;
assign detect_min[19][11] = (mid_1[167:160] < mid_0[175:168]) ? 1 : 0;
assign detect_min[19][12] = (mid_1[167:160] < mid_1[159:152]) ? 1 : 0;
assign detect_min[19][13] = (mid_1[167:160] < mid_1[175:168]) ? 1 : 0;
assign detect_min[19][14] = (mid_1[167:160] < mid_2[159:152]) ? 1 : 0;
assign detect_min[19][15] = (mid_1[167:160] < mid_2[167:160]) ? 1 : 0;
assign detect_min[19][16] = (mid_1[167:160] < mid_2[175:168]) ? 1 : 0;
assign detect_min[19][17] = (mid_1[167:160] < btm_0[159:152]) ? 1 : 0;
assign detect_min[19][18] = (mid_1[167:160] < btm_0[167:160]) ? 1 : 0;
assign detect_min[19][19] = (mid_1[167:160] < btm_0[175:168]) ? 1 : 0;
assign detect_min[19][20] = (mid_1[167:160] < btm_1[159:152]) ? 1 : 0;
assign detect_min[19][21] = (mid_1[167:160] < btm_1[167:160]) ? 1 : 0;
assign detect_min[19][22] = (mid_1[167:160] < btm_1[175:168]) ? 1 : 0;
assign detect_min[19][23] = (mid_1[167:160] < btm_2[159:152]) ? 1 : 0;
assign detect_min[19][24] = (mid_1[167:160] < btm_2[167:160]) ? 1 : 0;
assign detect_min[19][25] = (mid_1[167:160] < btm_2[175:168]) ? 1 : 0;

assign detect_min[20][0] = (mid_1[175:168] < top_0[167:160]) ? 1 : 0;
assign detect_min[20][1] = (mid_1[175:168] < top_0[175:168]) ? 1 : 0;
assign detect_min[20][2] = (mid_1[175:168] < top_0[183:176]) ? 1 : 0;
assign detect_min[20][3] = (mid_1[175:168] < top_1[167:160]) ? 1 : 0;
assign detect_min[20][4] = (mid_1[175:168] < top_1[175:168]) ? 1 : 0;
assign detect_min[20][5] = (mid_1[175:168] < top_1[183:176]) ? 1 : 0;
assign detect_min[20][6] = (mid_1[175:168] < top_2[167:160]) ? 1 : 0;
assign detect_min[20][7] = (mid_1[175:168] < top_2[175:168]) ? 1 : 0;
assign detect_min[20][8] = (mid_1[175:168] < top_2[183:176]) ? 1 : 0;
assign detect_min[20][9] = (mid_1[175:168] < mid_0[167:160]) ? 1 : 0;
assign detect_min[20][10] = (mid_1[175:168] < mid_0[175:168]) ? 1 : 0;
assign detect_min[20][11] = (mid_1[175:168] < mid_0[183:176]) ? 1 : 0;
assign detect_min[20][12] = (mid_1[175:168] < mid_1[167:160]) ? 1 : 0;
assign detect_min[20][13] = (mid_1[175:168] < mid_1[183:176]) ? 1 : 0;
assign detect_min[20][14] = (mid_1[175:168] < mid_2[167:160]) ? 1 : 0;
assign detect_min[20][15] = (mid_1[175:168] < mid_2[175:168]) ? 1 : 0;
assign detect_min[20][16] = (mid_1[175:168] < mid_2[183:176]) ? 1 : 0;
assign detect_min[20][17] = (mid_1[175:168] < btm_0[167:160]) ? 1 : 0;
assign detect_min[20][18] = (mid_1[175:168] < btm_0[175:168]) ? 1 : 0;
assign detect_min[20][19] = (mid_1[175:168] < btm_0[183:176]) ? 1 : 0;
assign detect_min[20][20] = (mid_1[175:168] < btm_1[167:160]) ? 1 : 0;
assign detect_min[20][21] = (mid_1[175:168] < btm_1[175:168]) ? 1 : 0;
assign detect_min[20][22] = (mid_1[175:168] < btm_1[183:176]) ? 1 : 0;
assign detect_min[20][23] = (mid_1[175:168] < btm_2[167:160]) ? 1 : 0;
assign detect_min[20][24] = (mid_1[175:168] < btm_2[175:168]) ? 1 : 0;
assign detect_min[20][25] = (mid_1[175:168] < btm_2[183:176]) ? 1 : 0;

assign detect_min[21][0] = (mid_1[183:176] < top_0[175:168]) ? 1 : 0;
assign detect_min[21][1] = (mid_1[183:176] < top_0[183:176]) ? 1 : 0;
assign detect_min[21][2] = (mid_1[183:176] < top_0[191:184]) ? 1 : 0;
assign detect_min[21][3] = (mid_1[183:176] < top_1[175:168]) ? 1 : 0;
assign detect_min[21][4] = (mid_1[183:176] < top_1[183:176]) ? 1 : 0;
assign detect_min[21][5] = (mid_1[183:176] < top_1[191:184]) ? 1 : 0;
assign detect_min[21][6] = (mid_1[183:176] < top_2[175:168]) ? 1 : 0;
assign detect_min[21][7] = (mid_1[183:176] < top_2[183:176]) ? 1 : 0;
assign detect_min[21][8] = (mid_1[183:176] < top_2[191:184]) ? 1 : 0;
assign detect_min[21][9] = (mid_1[183:176] < mid_0[175:168]) ? 1 : 0;
assign detect_min[21][10] = (mid_1[183:176] < mid_0[183:176]) ? 1 : 0;
assign detect_min[21][11] = (mid_1[183:176] < mid_0[191:184]) ? 1 : 0;
assign detect_min[21][12] = (mid_1[183:176] < mid_1[175:168]) ? 1 : 0;
assign detect_min[21][13] = (mid_1[183:176] < mid_1[191:184]) ? 1 : 0;
assign detect_min[21][14] = (mid_1[183:176] < mid_2[175:168]) ? 1 : 0;
assign detect_min[21][15] = (mid_1[183:176] < mid_2[183:176]) ? 1 : 0;
assign detect_min[21][16] = (mid_1[183:176] < mid_2[191:184]) ? 1 : 0;
assign detect_min[21][17] = (mid_1[183:176] < btm_0[175:168]) ? 1 : 0;
assign detect_min[21][18] = (mid_1[183:176] < btm_0[183:176]) ? 1 : 0;
assign detect_min[21][19] = (mid_1[183:176] < btm_0[191:184]) ? 1 : 0;
assign detect_min[21][20] = (mid_1[183:176] < btm_1[175:168]) ? 1 : 0;
assign detect_min[21][21] = (mid_1[183:176] < btm_1[183:176]) ? 1 : 0;
assign detect_min[21][22] = (mid_1[183:176] < btm_1[191:184]) ? 1 : 0;
assign detect_min[21][23] = (mid_1[183:176] < btm_2[175:168]) ? 1 : 0;
assign detect_min[21][24] = (mid_1[183:176] < btm_2[183:176]) ? 1 : 0;
assign detect_min[21][25] = (mid_1[183:176] < btm_2[191:184]) ? 1 : 0;

assign detect_min[22][0] = (mid_1[191:184] < top_0[183:176]) ? 1 : 0;
assign detect_min[22][1] = (mid_1[191:184] < top_0[191:184]) ? 1 : 0;
assign detect_min[22][2] = (mid_1[191:184] < top_0[199:192]) ? 1 : 0;
assign detect_min[22][3] = (mid_1[191:184] < top_1[183:176]) ? 1 : 0;
assign detect_min[22][4] = (mid_1[191:184] < top_1[191:184]) ? 1 : 0;
assign detect_min[22][5] = (mid_1[191:184] < top_1[199:192]) ? 1 : 0;
assign detect_min[22][6] = (mid_1[191:184] < top_2[183:176]) ? 1 : 0;
assign detect_min[22][7] = (mid_1[191:184] < top_2[191:184]) ? 1 : 0;
assign detect_min[22][8] = (mid_1[191:184] < top_2[199:192]) ? 1 : 0;
assign detect_min[22][9] = (mid_1[191:184] < mid_0[183:176]) ? 1 : 0;
assign detect_min[22][10] = (mid_1[191:184] < mid_0[191:184]) ? 1 : 0;
assign detect_min[22][11] = (mid_1[191:184] < mid_0[199:192]) ? 1 : 0;
assign detect_min[22][12] = (mid_1[191:184] < mid_1[183:176]) ? 1 : 0;
assign detect_min[22][13] = (mid_1[191:184] < mid_1[199:192]) ? 1 : 0;
assign detect_min[22][14] = (mid_1[191:184] < mid_2[183:176]) ? 1 : 0;
assign detect_min[22][15] = (mid_1[191:184] < mid_2[191:184]) ? 1 : 0;
assign detect_min[22][16] = (mid_1[191:184] < mid_2[199:192]) ? 1 : 0;
assign detect_min[22][17] = (mid_1[191:184] < btm_0[183:176]) ? 1 : 0;
assign detect_min[22][18] = (mid_1[191:184] < btm_0[191:184]) ? 1 : 0;
assign detect_min[22][19] = (mid_1[191:184] < btm_0[199:192]) ? 1 : 0;
assign detect_min[22][20] = (mid_1[191:184] < btm_1[183:176]) ? 1 : 0;
assign detect_min[22][21] = (mid_1[191:184] < btm_1[191:184]) ? 1 : 0;
assign detect_min[22][22] = (mid_1[191:184] < btm_1[199:192]) ? 1 : 0;
assign detect_min[22][23] = (mid_1[191:184] < btm_2[183:176]) ? 1 : 0;
assign detect_min[22][24] = (mid_1[191:184] < btm_2[191:184]) ? 1 : 0;
assign detect_min[22][25] = (mid_1[191:184] < btm_2[199:192]) ? 1 : 0;

assign detect_min[23][0] = (mid_1[199:192] < top_0[191:184]) ? 1 : 0;
assign detect_min[23][1] = (mid_1[199:192] < top_0[199:192]) ? 1 : 0;
assign detect_min[23][2] = (mid_1[199:192] < top_0[207:200]) ? 1 : 0;
assign detect_min[23][3] = (mid_1[199:192] < top_1[191:184]) ? 1 : 0;
assign detect_min[23][4] = (mid_1[199:192] < top_1[199:192]) ? 1 : 0;
assign detect_min[23][5] = (mid_1[199:192] < top_1[207:200]) ? 1 : 0;
assign detect_min[23][6] = (mid_1[199:192] < top_2[191:184]) ? 1 : 0;
assign detect_min[23][7] = (mid_1[199:192] < top_2[199:192]) ? 1 : 0;
assign detect_min[23][8] = (mid_1[199:192] < top_2[207:200]) ? 1 : 0;
assign detect_min[23][9] = (mid_1[199:192] < mid_0[191:184]) ? 1 : 0;
assign detect_min[23][10] = (mid_1[199:192] < mid_0[199:192]) ? 1 : 0;
assign detect_min[23][11] = (mid_1[199:192] < mid_0[207:200]) ? 1 : 0;
assign detect_min[23][12] = (mid_1[199:192] < mid_1[191:184]) ? 1 : 0;
assign detect_min[23][13] = (mid_1[199:192] < mid_1[207:200]) ? 1 : 0;
assign detect_min[23][14] = (mid_1[199:192] < mid_2[191:184]) ? 1 : 0;
assign detect_min[23][15] = (mid_1[199:192] < mid_2[199:192]) ? 1 : 0;
assign detect_min[23][16] = (mid_1[199:192] < mid_2[207:200]) ? 1 : 0;
assign detect_min[23][17] = (mid_1[199:192] < btm_0[191:184]) ? 1 : 0;
assign detect_min[23][18] = (mid_1[199:192] < btm_0[199:192]) ? 1 : 0;
assign detect_min[23][19] = (mid_1[199:192] < btm_0[207:200]) ? 1 : 0;
assign detect_min[23][20] = (mid_1[199:192] < btm_1[191:184]) ? 1 : 0;
assign detect_min[23][21] = (mid_1[199:192] < btm_1[199:192]) ? 1 : 0;
assign detect_min[23][22] = (mid_1[199:192] < btm_1[207:200]) ? 1 : 0;
assign detect_min[23][23] = (mid_1[199:192] < btm_2[191:184]) ? 1 : 0;
assign detect_min[23][24] = (mid_1[199:192] < btm_2[199:192]) ? 1 : 0;
assign detect_min[23][25] = (mid_1[199:192] < btm_2[207:200]) ? 1 : 0;

assign detect_min[24][0] = (mid_1[207:200] < top_0[199:192]) ? 1 : 0;
assign detect_min[24][1] = (mid_1[207:200] < top_0[207:200]) ? 1 : 0;
assign detect_min[24][2] = (mid_1[207:200] < top_0[215:208]) ? 1 : 0;
assign detect_min[24][3] = (mid_1[207:200] < top_1[199:192]) ? 1 : 0;
assign detect_min[24][4] = (mid_1[207:200] < top_1[207:200]) ? 1 : 0;
assign detect_min[24][5] = (mid_1[207:200] < top_1[215:208]) ? 1 : 0;
assign detect_min[24][6] = (mid_1[207:200] < top_2[199:192]) ? 1 : 0;
assign detect_min[24][7] = (mid_1[207:200] < top_2[207:200]) ? 1 : 0;
assign detect_min[24][8] = (mid_1[207:200] < top_2[215:208]) ? 1 : 0;
assign detect_min[24][9] = (mid_1[207:200] < mid_0[199:192]) ? 1 : 0;
assign detect_min[24][10] = (mid_1[207:200] < mid_0[207:200]) ? 1 : 0;
assign detect_min[24][11] = (mid_1[207:200] < mid_0[215:208]) ? 1 : 0;
assign detect_min[24][12] = (mid_1[207:200] < mid_1[199:192]) ? 1 : 0;
assign detect_min[24][13] = (mid_1[207:200] < mid_1[215:208]) ? 1 : 0;
assign detect_min[24][14] = (mid_1[207:200] < mid_2[199:192]) ? 1 : 0;
assign detect_min[24][15] = (mid_1[207:200] < mid_2[207:200]) ? 1 : 0;
assign detect_min[24][16] = (mid_1[207:200] < mid_2[215:208]) ? 1 : 0;
assign detect_min[24][17] = (mid_1[207:200] < btm_0[199:192]) ? 1 : 0;
assign detect_min[24][18] = (mid_1[207:200] < btm_0[207:200]) ? 1 : 0;
assign detect_min[24][19] = (mid_1[207:200] < btm_0[215:208]) ? 1 : 0;
assign detect_min[24][20] = (mid_1[207:200] < btm_1[199:192]) ? 1 : 0;
assign detect_min[24][21] = (mid_1[207:200] < btm_1[207:200]) ? 1 : 0;
assign detect_min[24][22] = (mid_1[207:200] < btm_1[215:208]) ? 1 : 0;
assign detect_min[24][23] = (mid_1[207:200] < btm_2[199:192]) ? 1 : 0;
assign detect_min[24][24] = (mid_1[207:200] < btm_2[207:200]) ? 1 : 0;
assign detect_min[24][25] = (mid_1[207:200] < btm_2[215:208]) ? 1 : 0;

assign detect_min[25][0] = (mid_1[215:208] < top_0[207:200]) ? 1 : 0;
assign detect_min[25][1] = (mid_1[215:208] < top_0[215:208]) ? 1 : 0;
assign detect_min[25][2] = (mid_1[215:208] < top_0[223:216]) ? 1 : 0;
assign detect_min[25][3] = (mid_1[215:208] < top_1[207:200]) ? 1 : 0;
assign detect_min[25][4] = (mid_1[215:208] < top_1[215:208]) ? 1 : 0;
assign detect_min[25][5] = (mid_1[215:208] < top_1[223:216]) ? 1 : 0;
assign detect_min[25][6] = (mid_1[215:208] < top_2[207:200]) ? 1 : 0;
assign detect_min[25][7] = (mid_1[215:208] < top_2[215:208]) ? 1 : 0;
assign detect_min[25][8] = (mid_1[215:208] < top_2[223:216]) ? 1 : 0;
assign detect_min[25][9] = (mid_1[215:208] < mid_0[207:200]) ? 1 : 0;
assign detect_min[25][10] = (mid_1[215:208] < mid_0[215:208]) ? 1 : 0;
assign detect_min[25][11] = (mid_1[215:208] < mid_0[223:216]) ? 1 : 0;
assign detect_min[25][12] = (mid_1[215:208] < mid_1[207:200]) ? 1 : 0;
assign detect_min[25][13] = (mid_1[215:208] < mid_1[223:216]) ? 1 : 0;
assign detect_min[25][14] = (mid_1[215:208] < mid_2[207:200]) ? 1 : 0;
assign detect_min[25][15] = (mid_1[215:208] < mid_2[215:208]) ? 1 : 0;
assign detect_min[25][16] = (mid_1[215:208] < mid_2[223:216]) ? 1 : 0;
assign detect_min[25][17] = (mid_1[215:208] < btm_0[207:200]) ? 1 : 0;
assign detect_min[25][18] = (mid_1[215:208] < btm_0[215:208]) ? 1 : 0;
assign detect_min[25][19] = (mid_1[215:208] < btm_0[223:216]) ? 1 : 0;
assign detect_min[25][20] = (mid_1[215:208] < btm_1[207:200]) ? 1 : 0;
assign detect_min[25][21] = (mid_1[215:208] < btm_1[215:208]) ? 1 : 0;
assign detect_min[25][22] = (mid_1[215:208] < btm_1[223:216]) ? 1 : 0;
assign detect_min[25][23] = (mid_1[215:208] < btm_2[207:200]) ? 1 : 0;
assign detect_min[25][24] = (mid_1[215:208] < btm_2[215:208]) ? 1 : 0;
assign detect_min[25][25] = (mid_1[215:208] < btm_2[223:216]) ? 1 : 0;

assign detect_min[26][0] = (mid_1[223:216] < top_0[215:208]) ? 1 : 0;
assign detect_min[26][1] = (mid_1[223:216] < top_0[223:216]) ? 1 : 0;
assign detect_min[26][2] = (mid_1[223:216] < top_0[231:224]) ? 1 : 0;
assign detect_min[26][3] = (mid_1[223:216] < top_1[215:208]) ? 1 : 0;
assign detect_min[26][4] = (mid_1[223:216] < top_1[223:216]) ? 1 : 0;
assign detect_min[26][5] = (mid_1[223:216] < top_1[231:224]) ? 1 : 0;
assign detect_min[26][6] = (mid_1[223:216] < top_2[215:208]) ? 1 : 0;
assign detect_min[26][7] = (mid_1[223:216] < top_2[223:216]) ? 1 : 0;
assign detect_min[26][8] = (mid_1[223:216] < top_2[231:224]) ? 1 : 0;
assign detect_min[26][9] = (mid_1[223:216] < mid_0[215:208]) ? 1 : 0;
assign detect_min[26][10] = (mid_1[223:216] < mid_0[223:216]) ? 1 : 0;
assign detect_min[26][11] = (mid_1[223:216] < mid_0[231:224]) ? 1 : 0;
assign detect_min[26][12] = (mid_1[223:216] < mid_1[215:208]) ? 1 : 0;
assign detect_min[26][13] = (mid_1[223:216] < mid_1[231:224]) ? 1 : 0;
assign detect_min[26][14] = (mid_1[223:216] < mid_2[215:208]) ? 1 : 0;
assign detect_min[26][15] = (mid_1[223:216] < mid_2[223:216]) ? 1 : 0;
assign detect_min[26][16] = (mid_1[223:216] < mid_2[231:224]) ? 1 : 0;
assign detect_min[26][17] = (mid_1[223:216] < btm_0[215:208]) ? 1 : 0;
assign detect_min[26][18] = (mid_1[223:216] < btm_0[223:216]) ? 1 : 0;
assign detect_min[26][19] = (mid_1[223:216] < btm_0[231:224]) ? 1 : 0;
assign detect_min[26][20] = (mid_1[223:216] < btm_1[215:208]) ? 1 : 0;
assign detect_min[26][21] = (mid_1[223:216] < btm_1[223:216]) ? 1 : 0;
assign detect_min[26][22] = (mid_1[223:216] < btm_1[231:224]) ? 1 : 0;
assign detect_min[26][23] = (mid_1[223:216] < btm_2[215:208]) ? 1 : 0;
assign detect_min[26][24] = (mid_1[223:216] < btm_2[223:216]) ? 1 : 0;
assign detect_min[26][25] = (mid_1[223:216] < btm_2[231:224]) ? 1 : 0;

assign detect_min[27][0] = (mid_1[231:224] < top_0[223:216]) ? 1 : 0;
assign detect_min[27][1] = (mid_1[231:224] < top_0[231:224]) ? 1 : 0;
assign detect_min[27][2] = (mid_1[231:224] < top_0[239:232]) ? 1 : 0;
assign detect_min[27][3] = (mid_1[231:224] < top_1[223:216]) ? 1 : 0;
assign detect_min[27][4] = (mid_1[231:224] < top_1[231:224]) ? 1 : 0;
assign detect_min[27][5] = (mid_1[231:224] < top_1[239:232]) ? 1 : 0;
assign detect_min[27][6] = (mid_1[231:224] < top_2[223:216]) ? 1 : 0;
assign detect_min[27][7] = (mid_1[231:224] < top_2[231:224]) ? 1 : 0;
assign detect_min[27][8] = (mid_1[231:224] < top_2[239:232]) ? 1 : 0;
assign detect_min[27][9] = (mid_1[231:224] < mid_0[223:216]) ? 1 : 0;
assign detect_min[27][10] = (mid_1[231:224] < mid_0[231:224]) ? 1 : 0;
assign detect_min[27][11] = (mid_1[231:224] < mid_0[239:232]) ? 1 : 0;
assign detect_min[27][12] = (mid_1[231:224] < mid_1[223:216]) ? 1 : 0;
assign detect_min[27][13] = (mid_1[231:224] < mid_1[239:232]) ? 1 : 0;
assign detect_min[27][14] = (mid_1[231:224] < mid_2[223:216]) ? 1 : 0;
assign detect_min[27][15] = (mid_1[231:224] < mid_2[231:224]) ? 1 : 0;
assign detect_min[27][16] = (mid_1[231:224] < mid_2[239:232]) ? 1 : 0;
assign detect_min[27][17] = (mid_1[231:224] < btm_0[223:216]) ? 1 : 0;
assign detect_min[27][18] = (mid_1[231:224] < btm_0[231:224]) ? 1 : 0;
assign detect_min[27][19] = (mid_1[231:224] < btm_0[239:232]) ? 1 : 0;
assign detect_min[27][20] = (mid_1[231:224] < btm_1[223:216]) ? 1 : 0;
assign detect_min[27][21] = (mid_1[231:224] < btm_1[231:224]) ? 1 : 0;
assign detect_min[27][22] = (mid_1[231:224] < btm_1[239:232]) ? 1 : 0;
assign detect_min[27][23] = (mid_1[231:224] < btm_2[223:216]) ? 1 : 0;
assign detect_min[27][24] = (mid_1[231:224] < btm_2[231:224]) ? 1 : 0;
assign detect_min[27][25] = (mid_1[231:224] < btm_2[239:232]) ? 1 : 0;

assign detect_min[28][0] = (mid_1[239:232] < top_0[231:224]) ? 1 : 0;
assign detect_min[28][1] = (mid_1[239:232] < top_0[239:232]) ? 1 : 0;
assign detect_min[28][2] = (mid_1[239:232] < top_0[247:240]) ? 1 : 0;
assign detect_min[28][3] = (mid_1[239:232] < top_1[231:224]) ? 1 : 0;
assign detect_min[28][4] = (mid_1[239:232] < top_1[239:232]) ? 1 : 0;
assign detect_min[28][5] = (mid_1[239:232] < top_1[247:240]) ? 1 : 0;
assign detect_min[28][6] = (mid_1[239:232] < top_2[231:224]) ? 1 : 0;
assign detect_min[28][7] = (mid_1[239:232] < top_2[239:232]) ? 1 : 0;
assign detect_min[28][8] = (mid_1[239:232] < top_2[247:240]) ? 1 : 0;
assign detect_min[28][9] = (mid_1[239:232] < mid_0[231:224]) ? 1 : 0;
assign detect_min[28][10] = (mid_1[239:232] < mid_0[239:232]) ? 1 : 0;
assign detect_min[28][11] = (mid_1[239:232] < mid_0[247:240]) ? 1 : 0;
assign detect_min[28][12] = (mid_1[239:232] < mid_1[231:224]) ? 1 : 0;
assign detect_min[28][13] = (mid_1[239:232] < mid_1[247:240]) ? 1 : 0;
assign detect_min[28][14] = (mid_1[239:232] < mid_2[231:224]) ? 1 : 0;
assign detect_min[28][15] = (mid_1[239:232] < mid_2[239:232]) ? 1 : 0;
assign detect_min[28][16] = (mid_1[239:232] < mid_2[247:240]) ? 1 : 0;
assign detect_min[28][17] = (mid_1[239:232] < btm_0[231:224]) ? 1 : 0;
assign detect_min[28][18] = (mid_1[239:232] < btm_0[239:232]) ? 1 : 0;
assign detect_min[28][19] = (mid_1[239:232] < btm_0[247:240]) ? 1 : 0;
assign detect_min[28][20] = (mid_1[239:232] < btm_1[231:224]) ? 1 : 0;
assign detect_min[28][21] = (mid_1[239:232] < btm_1[239:232]) ? 1 : 0;
assign detect_min[28][22] = (mid_1[239:232] < btm_1[247:240]) ? 1 : 0;
assign detect_min[28][23] = (mid_1[239:232] < btm_2[231:224]) ? 1 : 0;
assign detect_min[28][24] = (mid_1[239:232] < btm_2[239:232]) ? 1 : 0;
assign detect_min[28][25] = (mid_1[239:232] < btm_2[247:240]) ? 1 : 0;

assign detect_min[29][0] = (mid_1[247:240] < top_0[239:232]) ? 1 : 0;
assign detect_min[29][1] = (mid_1[247:240] < top_0[247:240]) ? 1 : 0;
assign detect_min[29][2] = (mid_1[247:240] < top_0[255:248]) ? 1 : 0;
assign detect_min[29][3] = (mid_1[247:240] < top_1[239:232]) ? 1 : 0;
assign detect_min[29][4] = (mid_1[247:240] < top_1[247:240]) ? 1 : 0;
assign detect_min[29][5] = (mid_1[247:240] < top_1[255:248]) ? 1 : 0;
assign detect_min[29][6] = (mid_1[247:240] < top_2[239:232]) ? 1 : 0;
assign detect_min[29][7] = (mid_1[247:240] < top_2[247:240]) ? 1 : 0;
assign detect_min[29][8] = (mid_1[247:240] < top_2[255:248]) ? 1 : 0;
assign detect_min[29][9] = (mid_1[247:240] < mid_0[239:232]) ? 1 : 0;
assign detect_min[29][10] = (mid_1[247:240] < mid_0[247:240]) ? 1 : 0;
assign detect_min[29][11] = (mid_1[247:240] < mid_0[255:248]) ? 1 : 0;
assign detect_min[29][12] = (mid_1[247:240] < mid_1[239:232]) ? 1 : 0;
assign detect_min[29][13] = (mid_1[247:240] < mid_1[255:248]) ? 1 : 0;
assign detect_min[29][14] = (mid_1[247:240] < mid_2[239:232]) ? 1 : 0;
assign detect_min[29][15] = (mid_1[247:240] < mid_2[247:240]) ? 1 : 0;
assign detect_min[29][16] = (mid_1[247:240] < mid_2[255:248]) ? 1 : 0;
assign detect_min[29][17] = (mid_1[247:240] < btm_0[239:232]) ? 1 : 0;
assign detect_min[29][18] = (mid_1[247:240] < btm_0[247:240]) ? 1 : 0;
assign detect_min[29][19] = (mid_1[247:240] < btm_0[255:248]) ? 1 : 0;
assign detect_min[29][20] = (mid_1[247:240] < btm_1[239:232]) ? 1 : 0;
assign detect_min[29][21] = (mid_1[247:240] < btm_1[247:240]) ? 1 : 0;
assign detect_min[29][22] = (mid_1[247:240] < btm_1[255:248]) ? 1 : 0;
assign detect_min[29][23] = (mid_1[247:240] < btm_2[239:232]) ? 1 : 0;
assign detect_min[29][24] = (mid_1[247:240] < btm_2[247:240]) ? 1 : 0;
assign detect_min[29][25] = (mid_1[247:240] < btm_2[255:248]) ? 1 : 0;

assign detect_min[30][0] = (mid_1[255:248] < top_0[247:240]) ? 1 : 0;
assign detect_min[30][1] = (mid_1[255:248] < top_0[255:248]) ? 1 : 0;
assign detect_min[30][2] = (mid_1[255:248] < top_0[263:256]) ? 1 : 0;
assign detect_min[30][3] = (mid_1[255:248] < top_1[247:240]) ? 1 : 0;
assign detect_min[30][4] = (mid_1[255:248] < top_1[255:248]) ? 1 : 0;
assign detect_min[30][5] = (mid_1[255:248] < top_1[263:256]) ? 1 : 0;
assign detect_min[30][6] = (mid_1[255:248] < top_2[247:240]) ? 1 : 0;
assign detect_min[30][7] = (mid_1[255:248] < top_2[255:248]) ? 1 : 0;
assign detect_min[30][8] = (mid_1[255:248] < top_2[263:256]) ? 1 : 0;
assign detect_min[30][9] = (mid_1[255:248] < mid_0[247:240]) ? 1 : 0;
assign detect_min[30][10] = (mid_1[255:248] < mid_0[255:248]) ? 1 : 0;
assign detect_min[30][11] = (mid_1[255:248] < mid_0[263:256]) ? 1 : 0;
assign detect_min[30][12] = (mid_1[255:248] < mid_1[247:240]) ? 1 : 0;
assign detect_min[30][13] = (mid_1[255:248] < mid_1[263:256]) ? 1 : 0;
assign detect_min[30][14] = (mid_1[255:248] < mid_2[247:240]) ? 1 : 0;
assign detect_min[30][15] = (mid_1[255:248] < mid_2[255:248]) ? 1 : 0;
assign detect_min[30][16] = (mid_1[255:248] < mid_2[263:256]) ? 1 : 0;
assign detect_min[30][17] = (mid_1[255:248] < btm_0[247:240]) ? 1 : 0;
assign detect_min[30][18] = (mid_1[255:248] < btm_0[255:248]) ? 1 : 0;
assign detect_min[30][19] = (mid_1[255:248] < btm_0[263:256]) ? 1 : 0;
assign detect_min[30][20] = (mid_1[255:248] < btm_1[247:240]) ? 1 : 0;
assign detect_min[30][21] = (mid_1[255:248] < btm_1[255:248]) ? 1 : 0;
assign detect_min[30][22] = (mid_1[255:248] < btm_1[263:256]) ? 1 : 0;
assign detect_min[30][23] = (mid_1[255:248] < btm_2[247:240]) ? 1 : 0;
assign detect_min[30][24] = (mid_1[255:248] < btm_2[255:248]) ? 1 : 0;
assign detect_min[30][25] = (mid_1[255:248] < btm_2[263:256]) ? 1 : 0;

assign detect_min[31][0] = (mid_1[263:256] < top_0[255:248]) ? 1 : 0;
assign detect_min[31][1] = (mid_1[263:256] < top_0[263:256]) ? 1 : 0;
assign detect_min[31][2] = (mid_1[263:256] < top_0[271:264]) ? 1 : 0;
assign detect_min[31][3] = (mid_1[263:256] < top_1[255:248]) ? 1 : 0;
assign detect_min[31][4] = (mid_1[263:256] < top_1[263:256]) ? 1 : 0;
assign detect_min[31][5] = (mid_1[263:256] < top_1[271:264]) ? 1 : 0;
assign detect_min[31][6] = (mid_1[263:256] < top_2[255:248]) ? 1 : 0;
assign detect_min[31][7] = (mid_1[263:256] < top_2[263:256]) ? 1 : 0;
assign detect_min[31][8] = (mid_1[263:256] < top_2[271:264]) ? 1 : 0;
assign detect_min[31][9] = (mid_1[263:256] < mid_0[255:248]) ? 1 : 0;
assign detect_min[31][10] = (mid_1[263:256] < mid_0[263:256]) ? 1 : 0;
assign detect_min[31][11] = (mid_1[263:256] < mid_0[271:264]) ? 1 : 0;
assign detect_min[31][12] = (mid_1[263:256] < mid_1[255:248]) ? 1 : 0;
assign detect_min[31][13] = (mid_1[263:256] < mid_1[271:264]) ? 1 : 0;
assign detect_min[31][14] = (mid_1[263:256] < mid_2[255:248]) ? 1 : 0;
assign detect_min[31][15] = (mid_1[263:256] < mid_2[263:256]) ? 1 : 0;
assign detect_min[31][16] = (mid_1[263:256] < mid_2[271:264]) ? 1 : 0;
assign detect_min[31][17] = (mid_1[263:256] < btm_0[255:248]) ? 1 : 0;
assign detect_min[31][18] = (mid_1[263:256] < btm_0[263:256]) ? 1 : 0;
assign detect_min[31][19] = (mid_1[263:256] < btm_0[271:264]) ? 1 : 0;
assign detect_min[31][20] = (mid_1[263:256] < btm_1[255:248]) ? 1 : 0;
assign detect_min[31][21] = (mid_1[263:256] < btm_1[263:256]) ? 1 : 0;
assign detect_min[31][22] = (mid_1[263:256] < btm_1[271:264]) ? 1 : 0;
assign detect_min[31][23] = (mid_1[263:256] < btm_2[255:248]) ? 1 : 0;
assign detect_min[31][24] = (mid_1[263:256] < btm_2[263:256]) ? 1 : 0;
assign detect_min[31][25] = (mid_1[263:256] < btm_2[271:264]) ? 1 : 0;

assign detect_min[32][0] = (mid_1[271:264] < top_0[263:256]) ? 1 : 0;
assign detect_min[32][1] = (mid_1[271:264] < top_0[271:264]) ? 1 : 0;
assign detect_min[32][2] = (mid_1[271:264] < top_0[279:272]) ? 1 : 0;
assign detect_min[32][3] = (mid_1[271:264] < top_1[263:256]) ? 1 : 0;
assign detect_min[32][4] = (mid_1[271:264] < top_1[271:264]) ? 1 : 0;
assign detect_min[32][5] = (mid_1[271:264] < top_1[279:272]) ? 1 : 0;
assign detect_min[32][6] = (mid_1[271:264] < top_2[263:256]) ? 1 : 0;
assign detect_min[32][7] = (mid_1[271:264] < top_2[271:264]) ? 1 : 0;
assign detect_min[32][8] = (mid_1[271:264] < top_2[279:272]) ? 1 : 0;
assign detect_min[32][9] = (mid_1[271:264] < mid_0[263:256]) ? 1 : 0;
assign detect_min[32][10] = (mid_1[271:264] < mid_0[271:264]) ? 1 : 0;
assign detect_min[32][11] = (mid_1[271:264] < mid_0[279:272]) ? 1 : 0;
assign detect_min[32][12] = (mid_1[271:264] < mid_1[263:256]) ? 1 : 0;
assign detect_min[32][13] = (mid_1[271:264] < mid_1[279:272]) ? 1 : 0;
assign detect_min[32][14] = (mid_1[271:264] < mid_2[263:256]) ? 1 : 0;
assign detect_min[32][15] = (mid_1[271:264] < mid_2[271:264]) ? 1 : 0;
assign detect_min[32][16] = (mid_1[271:264] < mid_2[279:272]) ? 1 : 0;
assign detect_min[32][17] = (mid_1[271:264] < btm_0[263:256]) ? 1 : 0;
assign detect_min[32][18] = (mid_1[271:264] < btm_0[271:264]) ? 1 : 0;
assign detect_min[32][19] = (mid_1[271:264] < btm_0[279:272]) ? 1 : 0;
assign detect_min[32][20] = (mid_1[271:264] < btm_1[263:256]) ? 1 : 0;
assign detect_min[32][21] = (mid_1[271:264] < btm_1[271:264]) ? 1 : 0;
assign detect_min[32][22] = (mid_1[271:264] < btm_1[279:272]) ? 1 : 0;
assign detect_min[32][23] = (mid_1[271:264] < btm_2[263:256]) ? 1 : 0;
assign detect_min[32][24] = (mid_1[271:264] < btm_2[271:264]) ? 1 : 0;
assign detect_min[32][25] = (mid_1[271:264] < btm_2[279:272]) ? 1 : 0;

assign detect_min[33][0] = (mid_1[279:272] < top_0[271:264]) ? 1 : 0;
assign detect_min[33][1] = (mid_1[279:272] < top_0[279:272]) ? 1 : 0;
assign detect_min[33][2] = (mid_1[279:272] < top_0[287:280]) ? 1 : 0;
assign detect_min[33][3] = (mid_1[279:272] < top_1[271:264]) ? 1 : 0;
assign detect_min[33][4] = (mid_1[279:272] < top_1[279:272]) ? 1 : 0;
assign detect_min[33][5] = (mid_1[279:272] < top_1[287:280]) ? 1 : 0;
assign detect_min[33][6] = (mid_1[279:272] < top_2[271:264]) ? 1 : 0;
assign detect_min[33][7] = (mid_1[279:272] < top_2[279:272]) ? 1 : 0;
assign detect_min[33][8] = (mid_1[279:272] < top_2[287:280]) ? 1 : 0;
assign detect_min[33][9] = (mid_1[279:272] < mid_0[271:264]) ? 1 : 0;
assign detect_min[33][10] = (mid_1[279:272] < mid_0[279:272]) ? 1 : 0;
assign detect_min[33][11] = (mid_1[279:272] < mid_0[287:280]) ? 1 : 0;
assign detect_min[33][12] = (mid_1[279:272] < mid_1[271:264]) ? 1 : 0;
assign detect_min[33][13] = (mid_1[279:272] < mid_1[287:280]) ? 1 : 0;
assign detect_min[33][14] = (mid_1[279:272] < mid_2[271:264]) ? 1 : 0;
assign detect_min[33][15] = (mid_1[279:272] < mid_2[279:272]) ? 1 : 0;
assign detect_min[33][16] = (mid_1[279:272] < mid_2[287:280]) ? 1 : 0;
assign detect_min[33][17] = (mid_1[279:272] < btm_0[271:264]) ? 1 : 0;
assign detect_min[33][18] = (mid_1[279:272] < btm_0[279:272]) ? 1 : 0;
assign detect_min[33][19] = (mid_1[279:272] < btm_0[287:280]) ? 1 : 0;
assign detect_min[33][20] = (mid_1[279:272] < btm_1[271:264]) ? 1 : 0;
assign detect_min[33][21] = (mid_1[279:272] < btm_1[279:272]) ? 1 : 0;
assign detect_min[33][22] = (mid_1[279:272] < btm_1[287:280]) ? 1 : 0;
assign detect_min[33][23] = (mid_1[279:272] < btm_2[271:264]) ? 1 : 0;
assign detect_min[33][24] = (mid_1[279:272] < btm_2[279:272]) ? 1 : 0;
assign detect_min[33][25] = (mid_1[279:272] < btm_2[287:280]) ? 1 : 0;

assign detect_min[34][0] = (mid_1[287:280] < top_0[279:272]) ? 1 : 0;
assign detect_min[34][1] = (mid_1[287:280] < top_0[287:280]) ? 1 : 0;
assign detect_min[34][2] = (mid_1[287:280] < top_0[295:288]) ? 1 : 0;
assign detect_min[34][3] = (mid_1[287:280] < top_1[279:272]) ? 1 : 0;
assign detect_min[34][4] = (mid_1[287:280] < top_1[287:280]) ? 1 : 0;
assign detect_min[34][5] = (mid_1[287:280] < top_1[295:288]) ? 1 : 0;
assign detect_min[34][6] = (mid_1[287:280] < top_2[279:272]) ? 1 : 0;
assign detect_min[34][7] = (mid_1[287:280] < top_2[287:280]) ? 1 : 0;
assign detect_min[34][8] = (mid_1[287:280] < top_2[295:288]) ? 1 : 0;
assign detect_min[34][9] = (mid_1[287:280] < mid_0[279:272]) ? 1 : 0;
assign detect_min[34][10] = (mid_1[287:280] < mid_0[287:280]) ? 1 : 0;
assign detect_min[34][11] = (mid_1[287:280] < mid_0[295:288]) ? 1 : 0;
assign detect_min[34][12] = (mid_1[287:280] < mid_1[279:272]) ? 1 : 0;
assign detect_min[34][13] = (mid_1[287:280] < mid_1[295:288]) ? 1 : 0;
assign detect_min[34][14] = (mid_1[287:280] < mid_2[279:272]) ? 1 : 0;
assign detect_min[34][15] = (mid_1[287:280] < mid_2[287:280]) ? 1 : 0;
assign detect_min[34][16] = (mid_1[287:280] < mid_2[295:288]) ? 1 : 0;
assign detect_min[34][17] = (mid_1[287:280] < btm_0[279:272]) ? 1 : 0;
assign detect_min[34][18] = (mid_1[287:280] < btm_0[287:280]) ? 1 : 0;
assign detect_min[34][19] = (mid_1[287:280] < btm_0[295:288]) ? 1 : 0;
assign detect_min[34][20] = (mid_1[287:280] < btm_1[279:272]) ? 1 : 0;
assign detect_min[34][21] = (mid_1[287:280] < btm_1[287:280]) ? 1 : 0;
assign detect_min[34][22] = (mid_1[287:280] < btm_1[295:288]) ? 1 : 0;
assign detect_min[34][23] = (mid_1[287:280] < btm_2[279:272]) ? 1 : 0;
assign detect_min[34][24] = (mid_1[287:280] < btm_2[287:280]) ? 1 : 0;
assign detect_min[34][25] = (mid_1[287:280] < btm_2[295:288]) ? 1 : 0;

assign detect_min[35][0] = (mid_1[295:288] < top_0[287:280]) ? 1 : 0;
assign detect_min[35][1] = (mid_1[295:288] < top_0[295:288]) ? 1 : 0;
assign detect_min[35][2] = (mid_1[295:288] < top_0[303:296]) ? 1 : 0;
assign detect_min[35][3] = (mid_1[295:288] < top_1[287:280]) ? 1 : 0;
assign detect_min[35][4] = (mid_1[295:288] < top_1[295:288]) ? 1 : 0;
assign detect_min[35][5] = (mid_1[295:288] < top_1[303:296]) ? 1 : 0;
assign detect_min[35][6] = (mid_1[295:288] < top_2[287:280]) ? 1 : 0;
assign detect_min[35][7] = (mid_1[295:288] < top_2[295:288]) ? 1 : 0;
assign detect_min[35][8] = (mid_1[295:288] < top_2[303:296]) ? 1 : 0;
assign detect_min[35][9] = (mid_1[295:288] < mid_0[287:280]) ? 1 : 0;
assign detect_min[35][10] = (mid_1[295:288] < mid_0[295:288]) ? 1 : 0;
assign detect_min[35][11] = (mid_1[295:288] < mid_0[303:296]) ? 1 : 0;
assign detect_min[35][12] = (mid_1[295:288] < mid_1[287:280]) ? 1 : 0;
assign detect_min[35][13] = (mid_1[295:288] < mid_1[303:296]) ? 1 : 0;
assign detect_min[35][14] = (mid_1[295:288] < mid_2[287:280]) ? 1 : 0;
assign detect_min[35][15] = (mid_1[295:288] < mid_2[295:288]) ? 1 : 0;
assign detect_min[35][16] = (mid_1[295:288] < mid_2[303:296]) ? 1 : 0;
assign detect_min[35][17] = (mid_1[295:288] < btm_0[287:280]) ? 1 : 0;
assign detect_min[35][18] = (mid_1[295:288] < btm_0[295:288]) ? 1 : 0;
assign detect_min[35][19] = (mid_1[295:288] < btm_0[303:296]) ? 1 : 0;
assign detect_min[35][20] = (mid_1[295:288] < btm_1[287:280]) ? 1 : 0;
assign detect_min[35][21] = (mid_1[295:288] < btm_1[295:288]) ? 1 : 0;
assign detect_min[35][22] = (mid_1[295:288] < btm_1[303:296]) ? 1 : 0;
assign detect_min[35][23] = (mid_1[295:288] < btm_2[287:280]) ? 1 : 0;
assign detect_min[35][24] = (mid_1[295:288] < btm_2[295:288]) ? 1 : 0;
assign detect_min[35][25] = (mid_1[295:288] < btm_2[303:296]) ? 1 : 0;

assign detect_min[36][0] = (mid_1[303:296] < top_0[295:288]) ? 1 : 0;
assign detect_min[36][1] = (mid_1[303:296] < top_0[303:296]) ? 1 : 0;
assign detect_min[36][2] = (mid_1[303:296] < top_0[311:304]) ? 1 : 0;
assign detect_min[36][3] = (mid_1[303:296] < top_1[295:288]) ? 1 : 0;
assign detect_min[36][4] = (mid_1[303:296] < top_1[303:296]) ? 1 : 0;
assign detect_min[36][5] = (mid_1[303:296] < top_1[311:304]) ? 1 : 0;
assign detect_min[36][6] = (mid_1[303:296] < top_2[295:288]) ? 1 : 0;
assign detect_min[36][7] = (mid_1[303:296] < top_2[303:296]) ? 1 : 0;
assign detect_min[36][8] = (mid_1[303:296] < top_2[311:304]) ? 1 : 0;
assign detect_min[36][9] = (mid_1[303:296] < mid_0[295:288]) ? 1 : 0;
assign detect_min[36][10] = (mid_1[303:296] < mid_0[303:296]) ? 1 : 0;
assign detect_min[36][11] = (mid_1[303:296] < mid_0[311:304]) ? 1 : 0;
assign detect_min[36][12] = (mid_1[303:296] < mid_1[295:288]) ? 1 : 0;
assign detect_min[36][13] = (mid_1[303:296] < mid_1[311:304]) ? 1 : 0;
assign detect_min[36][14] = (mid_1[303:296] < mid_2[295:288]) ? 1 : 0;
assign detect_min[36][15] = (mid_1[303:296] < mid_2[303:296]) ? 1 : 0;
assign detect_min[36][16] = (mid_1[303:296] < mid_2[311:304]) ? 1 : 0;
assign detect_min[36][17] = (mid_1[303:296] < btm_0[295:288]) ? 1 : 0;
assign detect_min[36][18] = (mid_1[303:296] < btm_0[303:296]) ? 1 : 0;
assign detect_min[36][19] = (mid_1[303:296] < btm_0[311:304]) ? 1 : 0;
assign detect_min[36][20] = (mid_1[303:296] < btm_1[295:288]) ? 1 : 0;
assign detect_min[36][21] = (mid_1[303:296] < btm_1[303:296]) ? 1 : 0;
assign detect_min[36][22] = (mid_1[303:296] < btm_1[311:304]) ? 1 : 0;
assign detect_min[36][23] = (mid_1[303:296] < btm_2[295:288]) ? 1 : 0;
assign detect_min[36][24] = (mid_1[303:296] < btm_2[303:296]) ? 1 : 0;
assign detect_min[36][25] = (mid_1[303:296] < btm_2[311:304]) ? 1 : 0;

assign detect_min[37][0] = (mid_1[311:304] < top_0[303:296]) ? 1 : 0;
assign detect_min[37][1] = (mid_1[311:304] < top_0[311:304]) ? 1 : 0;
assign detect_min[37][2] = (mid_1[311:304] < top_0[319:312]) ? 1 : 0;
assign detect_min[37][3] = (mid_1[311:304] < top_1[303:296]) ? 1 : 0;
assign detect_min[37][4] = (mid_1[311:304] < top_1[311:304]) ? 1 : 0;
assign detect_min[37][5] = (mid_1[311:304] < top_1[319:312]) ? 1 : 0;
assign detect_min[37][6] = (mid_1[311:304] < top_2[303:296]) ? 1 : 0;
assign detect_min[37][7] = (mid_1[311:304] < top_2[311:304]) ? 1 : 0;
assign detect_min[37][8] = (mid_1[311:304] < top_2[319:312]) ? 1 : 0;
assign detect_min[37][9] = (mid_1[311:304] < mid_0[303:296]) ? 1 : 0;
assign detect_min[37][10] = (mid_1[311:304] < mid_0[311:304]) ? 1 : 0;
assign detect_min[37][11] = (mid_1[311:304] < mid_0[319:312]) ? 1 : 0;
assign detect_min[37][12] = (mid_1[311:304] < mid_1[303:296]) ? 1 : 0;
assign detect_min[37][13] = (mid_1[311:304] < mid_1[319:312]) ? 1 : 0;
assign detect_min[37][14] = (mid_1[311:304] < mid_2[303:296]) ? 1 : 0;
assign detect_min[37][15] = (mid_1[311:304] < mid_2[311:304]) ? 1 : 0;
assign detect_min[37][16] = (mid_1[311:304] < mid_2[319:312]) ? 1 : 0;
assign detect_min[37][17] = (mid_1[311:304] < btm_0[303:296]) ? 1 : 0;
assign detect_min[37][18] = (mid_1[311:304] < btm_0[311:304]) ? 1 : 0;
assign detect_min[37][19] = (mid_1[311:304] < btm_0[319:312]) ? 1 : 0;
assign detect_min[37][20] = (mid_1[311:304] < btm_1[303:296]) ? 1 : 0;
assign detect_min[37][21] = (mid_1[311:304] < btm_1[311:304]) ? 1 : 0;
assign detect_min[37][22] = (mid_1[311:304] < btm_1[319:312]) ? 1 : 0;
assign detect_min[37][23] = (mid_1[311:304] < btm_2[303:296]) ? 1 : 0;
assign detect_min[37][24] = (mid_1[311:304] < btm_2[311:304]) ? 1 : 0;
assign detect_min[37][25] = (mid_1[311:304] < btm_2[319:312]) ? 1 : 0;

assign detect_min[38][0] = (mid_1[319:312] < top_0[311:304]) ? 1 : 0;
assign detect_min[38][1] = (mid_1[319:312] < top_0[319:312]) ? 1 : 0;
assign detect_min[38][2] = (mid_1[319:312] < top_0[327:320]) ? 1 : 0;
assign detect_min[38][3] = (mid_1[319:312] < top_1[311:304]) ? 1 : 0;
assign detect_min[38][4] = (mid_1[319:312] < top_1[319:312]) ? 1 : 0;
assign detect_min[38][5] = (mid_1[319:312] < top_1[327:320]) ? 1 : 0;
assign detect_min[38][6] = (mid_1[319:312] < top_2[311:304]) ? 1 : 0;
assign detect_min[38][7] = (mid_1[319:312] < top_2[319:312]) ? 1 : 0;
assign detect_min[38][8] = (mid_1[319:312] < top_2[327:320]) ? 1 : 0;
assign detect_min[38][9] = (mid_1[319:312] < mid_0[311:304]) ? 1 : 0;
assign detect_min[38][10] = (mid_1[319:312] < mid_0[319:312]) ? 1 : 0;
assign detect_min[38][11] = (mid_1[319:312] < mid_0[327:320]) ? 1 : 0;
assign detect_min[38][12] = (mid_1[319:312] < mid_1[311:304]) ? 1 : 0;
assign detect_min[38][13] = (mid_1[319:312] < mid_1[327:320]) ? 1 : 0;
assign detect_min[38][14] = (mid_1[319:312] < mid_2[311:304]) ? 1 : 0;
assign detect_min[38][15] = (mid_1[319:312] < mid_2[319:312]) ? 1 : 0;
assign detect_min[38][16] = (mid_1[319:312] < mid_2[327:320]) ? 1 : 0;
assign detect_min[38][17] = (mid_1[319:312] < btm_0[311:304]) ? 1 : 0;
assign detect_min[38][18] = (mid_1[319:312] < btm_0[319:312]) ? 1 : 0;
assign detect_min[38][19] = (mid_1[319:312] < btm_0[327:320]) ? 1 : 0;
assign detect_min[38][20] = (mid_1[319:312] < btm_1[311:304]) ? 1 : 0;
assign detect_min[38][21] = (mid_1[319:312] < btm_1[319:312]) ? 1 : 0;
assign detect_min[38][22] = (mid_1[319:312] < btm_1[327:320]) ? 1 : 0;
assign detect_min[38][23] = (mid_1[319:312] < btm_2[311:304]) ? 1 : 0;
assign detect_min[38][24] = (mid_1[319:312] < btm_2[319:312]) ? 1 : 0;
assign detect_min[38][25] = (mid_1[319:312] < btm_2[327:320]) ? 1 : 0;

assign detect_min[39][0] = (mid_1[327:320] < top_0[319:312]) ? 1 : 0;
assign detect_min[39][1] = (mid_1[327:320] < top_0[327:320]) ? 1 : 0;
assign detect_min[39][2] = (mid_1[327:320] < top_0[335:328]) ? 1 : 0;
assign detect_min[39][3] = (mid_1[327:320] < top_1[319:312]) ? 1 : 0;
assign detect_min[39][4] = (mid_1[327:320] < top_1[327:320]) ? 1 : 0;
assign detect_min[39][5] = (mid_1[327:320] < top_1[335:328]) ? 1 : 0;
assign detect_min[39][6] = (mid_1[327:320] < top_2[319:312]) ? 1 : 0;
assign detect_min[39][7] = (mid_1[327:320] < top_2[327:320]) ? 1 : 0;
assign detect_min[39][8] = (mid_1[327:320] < top_2[335:328]) ? 1 : 0;
assign detect_min[39][9] = (mid_1[327:320] < mid_0[319:312]) ? 1 : 0;
assign detect_min[39][10] = (mid_1[327:320] < mid_0[327:320]) ? 1 : 0;
assign detect_min[39][11] = (mid_1[327:320] < mid_0[335:328]) ? 1 : 0;
assign detect_min[39][12] = (mid_1[327:320] < mid_1[319:312]) ? 1 : 0;
assign detect_min[39][13] = (mid_1[327:320] < mid_1[335:328]) ? 1 : 0;
assign detect_min[39][14] = (mid_1[327:320] < mid_2[319:312]) ? 1 : 0;
assign detect_min[39][15] = (mid_1[327:320] < mid_2[327:320]) ? 1 : 0;
assign detect_min[39][16] = (mid_1[327:320] < mid_2[335:328]) ? 1 : 0;
assign detect_min[39][17] = (mid_1[327:320] < btm_0[319:312]) ? 1 : 0;
assign detect_min[39][18] = (mid_1[327:320] < btm_0[327:320]) ? 1 : 0;
assign detect_min[39][19] = (mid_1[327:320] < btm_0[335:328]) ? 1 : 0;
assign detect_min[39][20] = (mid_1[327:320] < btm_1[319:312]) ? 1 : 0;
assign detect_min[39][21] = (mid_1[327:320] < btm_1[327:320]) ? 1 : 0;
assign detect_min[39][22] = (mid_1[327:320] < btm_1[335:328]) ? 1 : 0;
assign detect_min[39][23] = (mid_1[327:320] < btm_2[319:312]) ? 1 : 0;
assign detect_min[39][24] = (mid_1[327:320] < btm_2[327:320]) ? 1 : 0;
assign detect_min[39][25] = (mid_1[327:320] < btm_2[335:328]) ? 1 : 0;

assign detect_min[40][0] = (mid_1[335:328] < top_0[327:320]) ? 1 : 0;
assign detect_min[40][1] = (mid_1[335:328] < top_0[335:328]) ? 1 : 0;
assign detect_min[40][2] = (mid_1[335:328] < top_0[343:336]) ? 1 : 0;
assign detect_min[40][3] = (mid_1[335:328] < top_1[327:320]) ? 1 : 0;
assign detect_min[40][4] = (mid_1[335:328] < top_1[335:328]) ? 1 : 0;
assign detect_min[40][5] = (mid_1[335:328] < top_1[343:336]) ? 1 : 0;
assign detect_min[40][6] = (mid_1[335:328] < top_2[327:320]) ? 1 : 0;
assign detect_min[40][7] = (mid_1[335:328] < top_2[335:328]) ? 1 : 0;
assign detect_min[40][8] = (mid_1[335:328] < top_2[343:336]) ? 1 : 0;
assign detect_min[40][9] = (mid_1[335:328] < mid_0[327:320]) ? 1 : 0;
assign detect_min[40][10] = (mid_1[335:328] < mid_0[335:328]) ? 1 : 0;
assign detect_min[40][11] = (mid_1[335:328] < mid_0[343:336]) ? 1 : 0;
assign detect_min[40][12] = (mid_1[335:328] < mid_1[327:320]) ? 1 : 0;
assign detect_min[40][13] = (mid_1[335:328] < mid_1[343:336]) ? 1 : 0;
assign detect_min[40][14] = (mid_1[335:328] < mid_2[327:320]) ? 1 : 0;
assign detect_min[40][15] = (mid_1[335:328] < mid_2[335:328]) ? 1 : 0;
assign detect_min[40][16] = (mid_1[335:328] < mid_2[343:336]) ? 1 : 0;
assign detect_min[40][17] = (mid_1[335:328] < btm_0[327:320]) ? 1 : 0;
assign detect_min[40][18] = (mid_1[335:328] < btm_0[335:328]) ? 1 : 0;
assign detect_min[40][19] = (mid_1[335:328] < btm_0[343:336]) ? 1 : 0;
assign detect_min[40][20] = (mid_1[335:328] < btm_1[327:320]) ? 1 : 0;
assign detect_min[40][21] = (mid_1[335:328] < btm_1[335:328]) ? 1 : 0;
assign detect_min[40][22] = (mid_1[335:328] < btm_1[343:336]) ? 1 : 0;
assign detect_min[40][23] = (mid_1[335:328] < btm_2[327:320]) ? 1 : 0;
assign detect_min[40][24] = (mid_1[335:328] < btm_2[335:328]) ? 1 : 0;
assign detect_min[40][25] = (mid_1[335:328] < btm_2[343:336]) ? 1 : 0;

assign detect_min[41][0] = (mid_1[343:336] < top_0[335:328]) ? 1 : 0;
assign detect_min[41][1] = (mid_1[343:336] < top_0[343:336]) ? 1 : 0;
assign detect_min[41][2] = (mid_1[343:336] < top_0[351:344]) ? 1 : 0;
assign detect_min[41][3] = (mid_1[343:336] < top_1[335:328]) ? 1 : 0;
assign detect_min[41][4] = (mid_1[343:336] < top_1[343:336]) ? 1 : 0;
assign detect_min[41][5] = (mid_1[343:336] < top_1[351:344]) ? 1 : 0;
assign detect_min[41][6] = (mid_1[343:336] < top_2[335:328]) ? 1 : 0;
assign detect_min[41][7] = (mid_1[343:336] < top_2[343:336]) ? 1 : 0;
assign detect_min[41][8] = (mid_1[343:336] < top_2[351:344]) ? 1 : 0;
assign detect_min[41][9] = (mid_1[343:336] < mid_0[335:328]) ? 1 : 0;
assign detect_min[41][10] = (mid_1[343:336] < mid_0[343:336]) ? 1 : 0;
assign detect_min[41][11] = (mid_1[343:336] < mid_0[351:344]) ? 1 : 0;
assign detect_min[41][12] = (mid_1[343:336] < mid_1[335:328]) ? 1 : 0;
assign detect_min[41][13] = (mid_1[343:336] < mid_1[351:344]) ? 1 : 0;
assign detect_min[41][14] = (mid_1[343:336] < mid_2[335:328]) ? 1 : 0;
assign detect_min[41][15] = (mid_1[343:336] < mid_2[343:336]) ? 1 : 0;
assign detect_min[41][16] = (mid_1[343:336] < mid_2[351:344]) ? 1 : 0;
assign detect_min[41][17] = (mid_1[343:336] < btm_0[335:328]) ? 1 : 0;
assign detect_min[41][18] = (mid_1[343:336] < btm_0[343:336]) ? 1 : 0;
assign detect_min[41][19] = (mid_1[343:336] < btm_0[351:344]) ? 1 : 0;
assign detect_min[41][20] = (mid_1[343:336] < btm_1[335:328]) ? 1 : 0;
assign detect_min[41][21] = (mid_1[343:336] < btm_1[343:336]) ? 1 : 0;
assign detect_min[41][22] = (mid_1[343:336] < btm_1[351:344]) ? 1 : 0;
assign detect_min[41][23] = (mid_1[343:336] < btm_2[335:328]) ? 1 : 0;
assign detect_min[41][24] = (mid_1[343:336] < btm_2[343:336]) ? 1 : 0;
assign detect_min[41][25] = (mid_1[343:336] < btm_2[351:344]) ? 1 : 0;

assign detect_min[42][0] = (mid_1[351:344] < top_0[343:336]) ? 1 : 0;
assign detect_min[42][1] = (mid_1[351:344] < top_0[351:344]) ? 1 : 0;
assign detect_min[42][2] = (mid_1[351:344] < top_0[359:352]) ? 1 : 0;
assign detect_min[42][3] = (mid_1[351:344] < top_1[343:336]) ? 1 : 0;
assign detect_min[42][4] = (mid_1[351:344] < top_1[351:344]) ? 1 : 0;
assign detect_min[42][5] = (mid_1[351:344] < top_1[359:352]) ? 1 : 0;
assign detect_min[42][6] = (mid_1[351:344] < top_2[343:336]) ? 1 : 0;
assign detect_min[42][7] = (mid_1[351:344] < top_2[351:344]) ? 1 : 0;
assign detect_min[42][8] = (mid_1[351:344] < top_2[359:352]) ? 1 : 0;
assign detect_min[42][9] = (mid_1[351:344] < mid_0[343:336]) ? 1 : 0;
assign detect_min[42][10] = (mid_1[351:344] < mid_0[351:344]) ? 1 : 0;
assign detect_min[42][11] = (mid_1[351:344] < mid_0[359:352]) ? 1 : 0;
assign detect_min[42][12] = (mid_1[351:344] < mid_1[343:336]) ? 1 : 0;
assign detect_min[42][13] = (mid_1[351:344] < mid_1[359:352]) ? 1 : 0;
assign detect_min[42][14] = (mid_1[351:344] < mid_2[343:336]) ? 1 : 0;
assign detect_min[42][15] = (mid_1[351:344] < mid_2[351:344]) ? 1 : 0;
assign detect_min[42][16] = (mid_1[351:344] < mid_2[359:352]) ? 1 : 0;
assign detect_min[42][17] = (mid_1[351:344] < btm_0[343:336]) ? 1 : 0;
assign detect_min[42][18] = (mid_1[351:344] < btm_0[351:344]) ? 1 : 0;
assign detect_min[42][19] = (mid_1[351:344] < btm_0[359:352]) ? 1 : 0;
assign detect_min[42][20] = (mid_1[351:344] < btm_1[343:336]) ? 1 : 0;
assign detect_min[42][21] = (mid_1[351:344] < btm_1[351:344]) ? 1 : 0;
assign detect_min[42][22] = (mid_1[351:344] < btm_1[359:352]) ? 1 : 0;
assign detect_min[42][23] = (mid_1[351:344] < btm_2[343:336]) ? 1 : 0;
assign detect_min[42][24] = (mid_1[351:344] < btm_2[351:344]) ? 1 : 0;
assign detect_min[42][25] = (mid_1[351:344] < btm_2[359:352]) ? 1 : 0;

assign detect_min[43][0] = (mid_1[359:352] < top_0[351:344]) ? 1 : 0;
assign detect_min[43][1] = (mid_1[359:352] < top_0[359:352]) ? 1 : 0;
assign detect_min[43][2] = (mid_1[359:352] < top_0[367:360]) ? 1 : 0;
assign detect_min[43][3] = (mid_1[359:352] < top_1[351:344]) ? 1 : 0;
assign detect_min[43][4] = (mid_1[359:352] < top_1[359:352]) ? 1 : 0;
assign detect_min[43][5] = (mid_1[359:352] < top_1[367:360]) ? 1 : 0;
assign detect_min[43][6] = (mid_1[359:352] < top_2[351:344]) ? 1 : 0;
assign detect_min[43][7] = (mid_1[359:352] < top_2[359:352]) ? 1 : 0;
assign detect_min[43][8] = (mid_1[359:352] < top_2[367:360]) ? 1 : 0;
assign detect_min[43][9] = (mid_1[359:352] < mid_0[351:344]) ? 1 : 0;
assign detect_min[43][10] = (mid_1[359:352] < mid_0[359:352]) ? 1 : 0;
assign detect_min[43][11] = (mid_1[359:352] < mid_0[367:360]) ? 1 : 0;
assign detect_min[43][12] = (mid_1[359:352] < mid_1[351:344]) ? 1 : 0;
assign detect_min[43][13] = (mid_1[359:352] < mid_1[367:360]) ? 1 : 0;
assign detect_min[43][14] = (mid_1[359:352] < mid_2[351:344]) ? 1 : 0;
assign detect_min[43][15] = (mid_1[359:352] < mid_2[359:352]) ? 1 : 0;
assign detect_min[43][16] = (mid_1[359:352] < mid_2[367:360]) ? 1 : 0;
assign detect_min[43][17] = (mid_1[359:352] < btm_0[351:344]) ? 1 : 0;
assign detect_min[43][18] = (mid_1[359:352] < btm_0[359:352]) ? 1 : 0;
assign detect_min[43][19] = (mid_1[359:352] < btm_0[367:360]) ? 1 : 0;
assign detect_min[43][20] = (mid_1[359:352] < btm_1[351:344]) ? 1 : 0;
assign detect_min[43][21] = (mid_1[359:352] < btm_1[359:352]) ? 1 : 0;
assign detect_min[43][22] = (mid_1[359:352] < btm_1[367:360]) ? 1 : 0;
assign detect_min[43][23] = (mid_1[359:352] < btm_2[351:344]) ? 1 : 0;
assign detect_min[43][24] = (mid_1[359:352] < btm_2[359:352]) ? 1 : 0;
assign detect_min[43][25] = (mid_1[359:352] < btm_2[367:360]) ? 1 : 0;

assign detect_min[44][0] = (mid_1[367:360] < top_0[359:352]) ? 1 : 0;
assign detect_min[44][1] = (mid_1[367:360] < top_0[367:360]) ? 1 : 0;
assign detect_min[44][2] = (mid_1[367:360] < top_0[375:368]) ? 1 : 0;
assign detect_min[44][3] = (mid_1[367:360] < top_1[359:352]) ? 1 : 0;
assign detect_min[44][4] = (mid_1[367:360] < top_1[367:360]) ? 1 : 0;
assign detect_min[44][5] = (mid_1[367:360] < top_1[375:368]) ? 1 : 0;
assign detect_min[44][6] = (mid_1[367:360] < top_2[359:352]) ? 1 : 0;
assign detect_min[44][7] = (mid_1[367:360] < top_2[367:360]) ? 1 : 0;
assign detect_min[44][8] = (mid_1[367:360] < top_2[375:368]) ? 1 : 0;
assign detect_min[44][9] = (mid_1[367:360] < mid_0[359:352]) ? 1 : 0;
assign detect_min[44][10] = (mid_1[367:360] < mid_0[367:360]) ? 1 : 0;
assign detect_min[44][11] = (mid_1[367:360] < mid_0[375:368]) ? 1 : 0;
assign detect_min[44][12] = (mid_1[367:360] < mid_1[359:352]) ? 1 : 0;
assign detect_min[44][13] = (mid_1[367:360] < mid_1[375:368]) ? 1 : 0;
assign detect_min[44][14] = (mid_1[367:360] < mid_2[359:352]) ? 1 : 0;
assign detect_min[44][15] = (mid_1[367:360] < mid_2[367:360]) ? 1 : 0;
assign detect_min[44][16] = (mid_1[367:360] < mid_2[375:368]) ? 1 : 0;
assign detect_min[44][17] = (mid_1[367:360] < btm_0[359:352]) ? 1 : 0;
assign detect_min[44][18] = (mid_1[367:360] < btm_0[367:360]) ? 1 : 0;
assign detect_min[44][19] = (mid_1[367:360] < btm_0[375:368]) ? 1 : 0;
assign detect_min[44][20] = (mid_1[367:360] < btm_1[359:352]) ? 1 : 0;
assign detect_min[44][21] = (mid_1[367:360] < btm_1[367:360]) ? 1 : 0;
assign detect_min[44][22] = (mid_1[367:360] < btm_1[375:368]) ? 1 : 0;
assign detect_min[44][23] = (mid_1[367:360] < btm_2[359:352]) ? 1 : 0;
assign detect_min[44][24] = (mid_1[367:360] < btm_2[367:360]) ? 1 : 0;
assign detect_min[44][25] = (mid_1[367:360] < btm_2[375:368]) ? 1 : 0;

assign detect_min[45][0] = (mid_1[375:368] < top_0[367:360]) ? 1 : 0;
assign detect_min[45][1] = (mid_1[375:368] < top_0[375:368]) ? 1 : 0;
assign detect_min[45][2] = (mid_1[375:368] < top_0[383:376]) ? 1 : 0;
assign detect_min[45][3] = (mid_1[375:368] < top_1[367:360]) ? 1 : 0;
assign detect_min[45][4] = (mid_1[375:368] < top_1[375:368]) ? 1 : 0;
assign detect_min[45][5] = (mid_1[375:368] < top_1[383:376]) ? 1 : 0;
assign detect_min[45][6] = (mid_1[375:368] < top_2[367:360]) ? 1 : 0;
assign detect_min[45][7] = (mid_1[375:368] < top_2[375:368]) ? 1 : 0;
assign detect_min[45][8] = (mid_1[375:368] < top_2[383:376]) ? 1 : 0;
assign detect_min[45][9] = (mid_1[375:368] < mid_0[367:360]) ? 1 : 0;
assign detect_min[45][10] = (mid_1[375:368] < mid_0[375:368]) ? 1 : 0;
assign detect_min[45][11] = (mid_1[375:368] < mid_0[383:376]) ? 1 : 0;
assign detect_min[45][12] = (mid_1[375:368] < mid_1[367:360]) ? 1 : 0;
assign detect_min[45][13] = (mid_1[375:368] < mid_1[383:376]) ? 1 : 0;
assign detect_min[45][14] = (mid_1[375:368] < mid_2[367:360]) ? 1 : 0;
assign detect_min[45][15] = (mid_1[375:368] < mid_2[375:368]) ? 1 : 0;
assign detect_min[45][16] = (mid_1[375:368] < mid_2[383:376]) ? 1 : 0;
assign detect_min[45][17] = (mid_1[375:368] < btm_0[367:360]) ? 1 : 0;
assign detect_min[45][18] = (mid_1[375:368] < btm_0[375:368]) ? 1 : 0;
assign detect_min[45][19] = (mid_1[375:368] < btm_0[383:376]) ? 1 : 0;
assign detect_min[45][20] = (mid_1[375:368] < btm_1[367:360]) ? 1 : 0;
assign detect_min[45][21] = (mid_1[375:368] < btm_1[375:368]) ? 1 : 0;
assign detect_min[45][22] = (mid_1[375:368] < btm_1[383:376]) ? 1 : 0;
assign detect_min[45][23] = (mid_1[375:368] < btm_2[367:360]) ? 1 : 0;
assign detect_min[45][24] = (mid_1[375:368] < btm_2[375:368]) ? 1 : 0;
assign detect_min[45][25] = (mid_1[375:368] < btm_2[383:376]) ? 1 : 0;

assign detect_min[46][0] = (mid_1[383:376] < top_0[375:368]) ? 1 : 0;
assign detect_min[46][1] = (mid_1[383:376] < top_0[383:376]) ? 1 : 0;
assign detect_min[46][2] = (mid_1[383:376] < top_0[391:384]) ? 1 : 0;
assign detect_min[46][3] = (mid_1[383:376] < top_1[375:368]) ? 1 : 0;
assign detect_min[46][4] = (mid_1[383:376] < top_1[383:376]) ? 1 : 0;
assign detect_min[46][5] = (mid_1[383:376] < top_1[391:384]) ? 1 : 0;
assign detect_min[46][6] = (mid_1[383:376] < top_2[375:368]) ? 1 : 0;
assign detect_min[46][7] = (mid_1[383:376] < top_2[383:376]) ? 1 : 0;
assign detect_min[46][8] = (mid_1[383:376] < top_2[391:384]) ? 1 : 0;
assign detect_min[46][9] = (mid_1[383:376] < mid_0[375:368]) ? 1 : 0;
assign detect_min[46][10] = (mid_1[383:376] < mid_0[383:376]) ? 1 : 0;
assign detect_min[46][11] = (mid_1[383:376] < mid_0[391:384]) ? 1 : 0;
assign detect_min[46][12] = (mid_1[383:376] < mid_1[375:368]) ? 1 : 0;
assign detect_min[46][13] = (mid_1[383:376] < mid_1[391:384]) ? 1 : 0;
assign detect_min[46][14] = (mid_1[383:376] < mid_2[375:368]) ? 1 : 0;
assign detect_min[46][15] = (mid_1[383:376] < mid_2[383:376]) ? 1 : 0;
assign detect_min[46][16] = (mid_1[383:376] < mid_2[391:384]) ? 1 : 0;
assign detect_min[46][17] = (mid_1[383:376] < btm_0[375:368]) ? 1 : 0;
assign detect_min[46][18] = (mid_1[383:376] < btm_0[383:376]) ? 1 : 0;
assign detect_min[46][19] = (mid_1[383:376] < btm_0[391:384]) ? 1 : 0;
assign detect_min[46][20] = (mid_1[383:376] < btm_1[375:368]) ? 1 : 0;
assign detect_min[46][21] = (mid_1[383:376] < btm_1[383:376]) ? 1 : 0;
assign detect_min[46][22] = (mid_1[383:376] < btm_1[391:384]) ? 1 : 0;
assign detect_min[46][23] = (mid_1[383:376] < btm_2[375:368]) ? 1 : 0;
assign detect_min[46][24] = (mid_1[383:376] < btm_2[383:376]) ? 1 : 0;
assign detect_min[46][25] = (mid_1[383:376] < btm_2[391:384]) ? 1 : 0;

assign detect_min[47][0] = (mid_1[391:384] < top_0[383:376]) ? 1 : 0;
assign detect_min[47][1] = (mid_1[391:384] < top_0[391:384]) ? 1 : 0;
assign detect_min[47][2] = (mid_1[391:384] < top_0[399:392]) ? 1 : 0;
assign detect_min[47][3] = (mid_1[391:384] < top_1[383:376]) ? 1 : 0;
assign detect_min[47][4] = (mid_1[391:384] < top_1[391:384]) ? 1 : 0;
assign detect_min[47][5] = (mid_1[391:384] < top_1[399:392]) ? 1 : 0;
assign detect_min[47][6] = (mid_1[391:384] < top_2[383:376]) ? 1 : 0;
assign detect_min[47][7] = (mid_1[391:384] < top_2[391:384]) ? 1 : 0;
assign detect_min[47][8] = (mid_1[391:384] < top_2[399:392]) ? 1 : 0;
assign detect_min[47][9] = (mid_1[391:384] < mid_0[383:376]) ? 1 : 0;
assign detect_min[47][10] = (mid_1[391:384] < mid_0[391:384]) ? 1 : 0;
assign detect_min[47][11] = (mid_1[391:384] < mid_0[399:392]) ? 1 : 0;
assign detect_min[47][12] = (mid_1[391:384] < mid_1[383:376]) ? 1 : 0;
assign detect_min[47][13] = (mid_1[391:384] < mid_1[399:392]) ? 1 : 0;
assign detect_min[47][14] = (mid_1[391:384] < mid_2[383:376]) ? 1 : 0;
assign detect_min[47][15] = (mid_1[391:384] < mid_2[391:384]) ? 1 : 0;
assign detect_min[47][16] = (mid_1[391:384] < mid_2[399:392]) ? 1 : 0;
assign detect_min[47][17] = (mid_1[391:384] < btm_0[383:376]) ? 1 : 0;
assign detect_min[47][18] = (mid_1[391:384] < btm_0[391:384]) ? 1 : 0;
assign detect_min[47][19] = (mid_1[391:384] < btm_0[399:392]) ? 1 : 0;
assign detect_min[47][20] = (mid_1[391:384] < btm_1[383:376]) ? 1 : 0;
assign detect_min[47][21] = (mid_1[391:384] < btm_1[391:384]) ? 1 : 0;
assign detect_min[47][22] = (mid_1[391:384] < btm_1[399:392]) ? 1 : 0;
assign detect_min[47][23] = (mid_1[391:384] < btm_2[383:376]) ? 1 : 0;
assign detect_min[47][24] = (mid_1[391:384] < btm_2[391:384]) ? 1 : 0;
assign detect_min[47][25] = (mid_1[391:384] < btm_2[399:392]) ? 1 : 0;

assign detect_min[48][0] = (mid_1[399:392] < top_0[391:384]) ? 1 : 0;
assign detect_min[48][1] = (mid_1[399:392] < top_0[399:392]) ? 1 : 0;
assign detect_min[48][2] = (mid_1[399:392] < top_0[407:400]) ? 1 : 0;
assign detect_min[48][3] = (mid_1[399:392] < top_1[391:384]) ? 1 : 0;
assign detect_min[48][4] = (mid_1[399:392] < top_1[399:392]) ? 1 : 0;
assign detect_min[48][5] = (mid_1[399:392] < top_1[407:400]) ? 1 : 0;
assign detect_min[48][6] = (mid_1[399:392] < top_2[391:384]) ? 1 : 0;
assign detect_min[48][7] = (mid_1[399:392] < top_2[399:392]) ? 1 : 0;
assign detect_min[48][8] = (mid_1[399:392] < top_2[407:400]) ? 1 : 0;
assign detect_min[48][9] = (mid_1[399:392] < mid_0[391:384]) ? 1 : 0;
assign detect_min[48][10] = (mid_1[399:392] < mid_0[399:392]) ? 1 : 0;
assign detect_min[48][11] = (mid_1[399:392] < mid_0[407:400]) ? 1 : 0;
assign detect_min[48][12] = (mid_1[399:392] < mid_1[391:384]) ? 1 : 0;
assign detect_min[48][13] = (mid_1[399:392] < mid_1[407:400]) ? 1 : 0;
assign detect_min[48][14] = (mid_1[399:392] < mid_2[391:384]) ? 1 : 0;
assign detect_min[48][15] = (mid_1[399:392] < mid_2[399:392]) ? 1 : 0;
assign detect_min[48][16] = (mid_1[399:392] < mid_2[407:400]) ? 1 : 0;
assign detect_min[48][17] = (mid_1[399:392] < btm_0[391:384]) ? 1 : 0;
assign detect_min[48][18] = (mid_1[399:392] < btm_0[399:392]) ? 1 : 0;
assign detect_min[48][19] = (mid_1[399:392] < btm_0[407:400]) ? 1 : 0;
assign detect_min[48][20] = (mid_1[399:392] < btm_1[391:384]) ? 1 : 0;
assign detect_min[48][21] = (mid_1[399:392] < btm_1[399:392]) ? 1 : 0;
assign detect_min[48][22] = (mid_1[399:392] < btm_1[407:400]) ? 1 : 0;
assign detect_min[48][23] = (mid_1[399:392] < btm_2[391:384]) ? 1 : 0;
assign detect_min[48][24] = (mid_1[399:392] < btm_2[399:392]) ? 1 : 0;
assign detect_min[48][25] = (mid_1[399:392] < btm_2[407:400]) ? 1 : 0;

assign detect_min[49][0] = (mid_1[407:400] < top_0[399:392]) ? 1 : 0;
assign detect_min[49][1] = (mid_1[407:400] < top_0[407:400]) ? 1 : 0;
assign detect_min[49][2] = (mid_1[407:400] < top_0[415:408]) ? 1 : 0;
assign detect_min[49][3] = (mid_1[407:400] < top_1[399:392]) ? 1 : 0;
assign detect_min[49][4] = (mid_1[407:400] < top_1[407:400]) ? 1 : 0;
assign detect_min[49][5] = (mid_1[407:400] < top_1[415:408]) ? 1 : 0;
assign detect_min[49][6] = (mid_1[407:400] < top_2[399:392]) ? 1 : 0;
assign detect_min[49][7] = (mid_1[407:400] < top_2[407:400]) ? 1 : 0;
assign detect_min[49][8] = (mid_1[407:400] < top_2[415:408]) ? 1 : 0;
assign detect_min[49][9] = (mid_1[407:400] < mid_0[399:392]) ? 1 : 0;
assign detect_min[49][10] = (mid_1[407:400] < mid_0[407:400]) ? 1 : 0;
assign detect_min[49][11] = (mid_1[407:400] < mid_0[415:408]) ? 1 : 0;
assign detect_min[49][12] = (mid_1[407:400] < mid_1[399:392]) ? 1 : 0;
assign detect_min[49][13] = (mid_1[407:400] < mid_1[415:408]) ? 1 : 0;
assign detect_min[49][14] = (mid_1[407:400] < mid_2[399:392]) ? 1 : 0;
assign detect_min[49][15] = (mid_1[407:400] < mid_2[407:400]) ? 1 : 0;
assign detect_min[49][16] = (mid_1[407:400] < mid_2[415:408]) ? 1 : 0;
assign detect_min[49][17] = (mid_1[407:400] < btm_0[399:392]) ? 1 : 0;
assign detect_min[49][18] = (mid_1[407:400] < btm_0[407:400]) ? 1 : 0;
assign detect_min[49][19] = (mid_1[407:400] < btm_0[415:408]) ? 1 : 0;
assign detect_min[49][20] = (mid_1[407:400] < btm_1[399:392]) ? 1 : 0;
assign detect_min[49][21] = (mid_1[407:400] < btm_1[407:400]) ? 1 : 0;
assign detect_min[49][22] = (mid_1[407:400] < btm_1[415:408]) ? 1 : 0;
assign detect_min[49][23] = (mid_1[407:400] < btm_2[399:392]) ? 1 : 0;
assign detect_min[49][24] = (mid_1[407:400] < btm_2[407:400]) ? 1 : 0;
assign detect_min[49][25] = (mid_1[407:400] < btm_2[415:408]) ? 1 : 0;

assign detect_min[50][0] = (mid_1[415:408] < top_0[407:400]) ? 1 : 0;
assign detect_min[50][1] = (mid_1[415:408] < top_0[415:408]) ? 1 : 0;
assign detect_min[50][2] = (mid_1[415:408] < top_0[423:416]) ? 1 : 0;
assign detect_min[50][3] = (mid_1[415:408] < top_1[407:400]) ? 1 : 0;
assign detect_min[50][4] = (mid_1[415:408] < top_1[415:408]) ? 1 : 0;
assign detect_min[50][5] = (mid_1[415:408] < top_1[423:416]) ? 1 : 0;
assign detect_min[50][6] = (mid_1[415:408] < top_2[407:400]) ? 1 : 0;
assign detect_min[50][7] = (mid_1[415:408] < top_2[415:408]) ? 1 : 0;
assign detect_min[50][8] = (mid_1[415:408] < top_2[423:416]) ? 1 : 0;
assign detect_min[50][9] = (mid_1[415:408] < mid_0[407:400]) ? 1 : 0;
assign detect_min[50][10] = (mid_1[415:408] < mid_0[415:408]) ? 1 : 0;
assign detect_min[50][11] = (mid_1[415:408] < mid_0[423:416]) ? 1 : 0;
assign detect_min[50][12] = (mid_1[415:408] < mid_1[407:400]) ? 1 : 0;
assign detect_min[50][13] = (mid_1[415:408] < mid_1[423:416]) ? 1 : 0;
assign detect_min[50][14] = (mid_1[415:408] < mid_2[407:400]) ? 1 : 0;
assign detect_min[50][15] = (mid_1[415:408] < mid_2[415:408]) ? 1 : 0;
assign detect_min[50][16] = (mid_1[415:408] < mid_2[423:416]) ? 1 : 0;
assign detect_min[50][17] = (mid_1[415:408] < btm_0[407:400]) ? 1 : 0;
assign detect_min[50][18] = (mid_1[415:408] < btm_0[415:408]) ? 1 : 0;
assign detect_min[50][19] = (mid_1[415:408] < btm_0[423:416]) ? 1 : 0;
assign detect_min[50][20] = (mid_1[415:408] < btm_1[407:400]) ? 1 : 0;
assign detect_min[50][21] = (mid_1[415:408] < btm_1[415:408]) ? 1 : 0;
assign detect_min[50][22] = (mid_1[415:408] < btm_1[423:416]) ? 1 : 0;
assign detect_min[50][23] = (mid_1[415:408] < btm_2[407:400]) ? 1 : 0;
assign detect_min[50][24] = (mid_1[415:408] < btm_2[415:408]) ? 1 : 0;
assign detect_min[50][25] = (mid_1[415:408] < btm_2[423:416]) ? 1 : 0;

assign detect_min[51][0] = (mid_1[423:416] < top_0[415:408]) ? 1 : 0;
assign detect_min[51][1] = (mid_1[423:416] < top_0[423:416]) ? 1 : 0;
assign detect_min[51][2] = (mid_1[423:416] < top_0[431:424]) ? 1 : 0;
assign detect_min[51][3] = (mid_1[423:416] < top_1[415:408]) ? 1 : 0;
assign detect_min[51][4] = (mid_1[423:416] < top_1[423:416]) ? 1 : 0;
assign detect_min[51][5] = (mid_1[423:416] < top_1[431:424]) ? 1 : 0;
assign detect_min[51][6] = (mid_1[423:416] < top_2[415:408]) ? 1 : 0;
assign detect_min[51][7] = (mid_1[423:416] < top_2[423:416]) ? 1 : 0;
assign detect_min[51][8] = (mid_1[423:416] < top_2[431:424]) ? 1 : 0;
assign detect_min[51][9] = (mid_1[423:416] < mid_0[415:408]) ? 1 : 0;
assign detect_min[51][10] = (mid_1[423:416] < mid_0[423:416]) ? 1 : 0;
assign detect_min[51][11] = (mid_1[423:416] < mid_0[431:424]) ? 1 : 0;
assign detect_min[51][12] = (mid_1[423:416] < mid_1[415:408]) ? 1 : 0;
assign detect_min[51][13] = (mid_1[423:416] < mid_1[431:424]) ? 1 : 0;
assign detect_min[51][14] = (mid_1[423:416] < mid_2[415:408]) ? 1 : 0;
assign detect_min[51][15] = (mid_1[423:416] < mid_2[423:416]) ? 1 : 0;
assign detect_min[51][16] = (mid_1[423:416] < mid_2[431:424]) ? 1 : 0;
assign detect_min[51][17] = (mid_1[423:416] < btm_0[415:408]) ? 1 : 0;
assign detect_min[51][18] = (mid_1[423:416] < btm_0[423:416]) ? 1 : 0;
assign detect_min[51][19] = (mid_1[423:416] < btm_0[431:424]) ? 1 : 0;
assign detect_min[51][20] = (mid_1[423:416] < btm_1[415:408]) ? 1 : 0;
assign detect_min[51][21] = (mid_1[423:416] < btm_1[423:416]) ? 1 : 0;
assign detect_min[51][22] = (mid_1[423:416] < btm_1[431:424]) ? 1 : 0;
assign detect_min[51][23] = (mid_1[423:416] < btm_2[415:408]) ? 1 : 0;
assign detect_min[51][24] = (mid_1[423:416] < btm_2[423:416]) ? 1 : 0;
assign detect_min[51][25] = (mid_1[423:416] < btm_2[431:424]) ? 1 : 0;

assign detect_min[52][0] = (mid_1[431:424] < top_0[423:416]) ? 1 : 0;
assign detect_min[52][1] = (mid_1[431:424] < top_0[431:424]) ? 1 : 0;
assign detect_min[52][2] = (mid_1[431:424] < top_0[439:432]) ? 1 : 0;
assign detect_min[52][3] = (mid_1[431:424] < top_1[423:416]) ? 1 : 0;
assign detect_min[52][4] = (mid_1[431:424] < top_1[431:424]) ? 1 : 0;
assign detect_min[52][5] = (mid_1[431:424] < top_1[439:432]) ? 1 : 0;
assign detect_min[52][6] = (mid_1[431:424] < top_2[423:416]) ? 1 : 0;
assign detect_min[52][7] = (mid_1[431:424] < top_2[431:424]) ? 1 : 0;
assign detect_min[52][8] = (mid_1[431:424] < top_2[439:432]) ? 1 : 0;
assign detect_min[52][9] = (mid_1[431:424] < mid_0[423:416]) ? 1 : 0;
assign detect_min[52][10] = (mid_1[431:424] < mid_0[431:424]) ? 1 : 0;
assign detect_min[52][11] = (mid_1[431:424] < mid_0[439:432]) ? 1 : 0;
assign detect_min[52][12] = (mid_1[431:424] < mid_1[423:416]) ? 1 : 0;
assign detect_min[52][13] = (mid_1[431:424] < mid_1[439:432]) ? 1 : 0;
assign detect_min[52][14] = (mid_1[431:424] < mid_2[423:416]) ? 1 : 0;
assign detect_min[52][15] = (mid_1[431:424] < mid_2[431:424]) ? 1 : 0;
assign detect_min[52][16] = (mid_1[431:424] < mid_2[439:432]) ? 1 : 0;
assign detect_min[52][17] = (mid_1[431:424] < btm_0[423:416]) ? 1 : 0;
assign detect_min[52][18] = (mid_1[431:424] < btm_0[431:424]) ? 1 : 0;
assign detect_min[52][19] = (mid_1[431:424] < btm_0[439:432]) ? 1 : 0;
assign detect_min[52][20] = (mid_1[431:424] < btm_1[423:416]) ? 1 : 0;
assign detect_min[52][21] = (mid_1[431:424] < btm_1[431:424]) ? 1 : 0;
assign detect_min[52][22] = (mid_1[431:424] < btm_1[439:432]) ? 1 : 0;
assign detect_min[52][23] = (mid_1[431:424] < btm_2[423:416]) ? 1 : 0;
assign detect_min[52][24] = (mid_1[431:424] < btm_2[431:424]) ? 1 : 0;
assign detect_min[52][25] = (mid_1[431:424] < btm_2[439:432]) ? 1 : 0;

assign detect_min[53][0] = (mid_1[439:432] < top_0[431:424]) ? 1 : 0;
assign detect_min[53][1] = (mid_1[439:432] < top_0[439:432]) ? 1 : 0;
assign detect_min[53][2] = (mid_1[439:432] < top_0[447:440]) ? 1 : 0;
assign detect_min[53][3] = (mid_1[439:432] < top_1[431:424]) ? 1 : 0;
assign detect_min[53][4] = (mid_1[439:432] < top_1[439:432]) ? 1 : 0;
assign detect_min[53][5] = (mid_1[439:432] < top_1[447:440]) ? 1 : 0;
assign detect_min[53][6] = (mid_1[439:432] < top_2[431:424]) ? 1 : 0;
assign detect_min[53][7] = (mid_1[439:432] < top_2[439:432]) ? 1 : 0;
assign detect_min[53][8] = (mid_1[439:432] < top_2[447:440]) ? 1 : 0;
assign detect_min[53][9] = (mid_1[439:432] < mid_0[431:424]) ? 1 : 0;
assign detect_min[53][10] = (mid_1[439:432] < mid_0[439:432]) ? 1 : 0;
assign detect_min[53][11] = (mid_1[439:432] < mid_0[447:440]) ? 1 : 0;
assign detect_min[53][12] = (mid_1[439:432] < mid_1[431:424]) ? 1 : 0;
assign detect_min[53][13] = (mid_1[439:432] < mid_1[447:440]) ? 1 : 0;
assign detect_min[53][14] = (mid_1[439:432] < mid_2[431:424]) ? 1 : 0;
assign detect_min[53][15] = (mid_1[439:432] < mid_2[439:432]) ? 1 : 0;
assign detect_min[53][16] = (mid_1[439:432] < mid_2[447:440]) ? 1 : 0;
assign detect_min[53][17] = (mid_1[439:432] < btm_0[431:424]) ? 1 : 0;
assign detect_min[53][18] = (mid_1[439:432] < btm_0[439:432]) ? 1 : 0;
assign detect_min[53][19] = (mid_1[439:432] < btm_0[447:440]) ? 1 : 0;
assign detect_min[53][20] = (mid_1[439:432] < btm_1[431:424]) ? 1 : 0;
assign detect_min[53][21] = (mid_1[439:432] < btm_1[439:432]) ? 1 : 0;
assign detect_min[53][22] = (mid_1[439:432] < btm_1[447:440]) ? 1 : 0;
assign detect_min[53][23] = (mid_1[439:432] < btm_2[431:424]) ? 1 : 0;
assign detect_min[53][24] = (mid_1[439:432] < btm_2[439:432]) ? 1 : 0;
assign detect_min[53][25] = (mid_1[439:432] < btm_2[447:440]) ? 1 : 0;

assign detect_min[54][0] = (mid_1[447:440] < top_0[439:432]) ? 1 : 0;
assign detect_min[54][1] = (mid_1[447:440] < top_0[447:440]) ? 1 : 0;
assign detect_min[54][2] = (mid_1[447:440] < top_0[455:448]) ? 1 : 0;
assign detect_min[54][3] = (mid_1[447:440] < top_1[439:432]) ? 1 : 0;
assign detect_min[54][4] = (mid_1[447:440] < top_1[447:440]) ? 1 : 0;
assign detect_min[54][5] = (mid_1[447:440] < top_1[455:448]) ? 1 : 0;
assign detect_min[54][6] = (mid_1[447:440] < top_2[439:432]) ? 1 : 0;
assign detect_min[54][7] = (mid_1[447:440] < top_2[447:440]) ? 1 : 0;
assign detect_min[54][8] = (mid_1[447:440] < top_2[455:448]) ? 1 : 0;
assign detect_min[54][9] = (mid_1[447:440] < mid_0[439:432]) ? 1 : 0;
assign detect_min[54][10] = (mid_1[447:440] < mid_0[447:440]) ? 1 : 0;
assign detect_min[54][11] = (mid_1[447:440] < mid_0[455:448]) ? 1 : 0;
assign detect_min[54][12] = (mid_1[447:440] < mid_1[439:432]) ? 1 : 0;
assign detect_min[54][13] = (mid_1[447:440] < mid_1[455:448]) ? 1 : 0;
assign detect_min[54][14] = (mid_1[447:440] < mid_2[439:432]) ? 1 : 0;
assign detect_min[54][15] = (mid_1[447:440] < mid_2[447:440]) ? 1 : 0;
assign detect_min[54][16] = (mid_1[447:440] < mid_2[455:448]) ? 1 : 0;
assign detect_min[54][17] = (mid_1[447:440] < btm_0[439:432]) ? 1 : 0;
assign detect_min[54][18] = (mid_1[447:440] < btm_0[447:440]) ? 1 : 0;
assign detect_min[54][19] = (mid_1[447:440] < btm_0[455:448]) ? 1 : 0;
assign detect_min[54][20] = (mid_1[447:440] < btm_1[439:432]) ? 1 : 0;
assign detect_min[54][21] = (mid_1[447:440] < btm_1[447:440]) ? 1 : 0;
assign detect_min[54][22] = (mid_1[447:440] < btm_1[455:448]) ? 1 : 0;
assign detect_min[54][23] = (mid_1[447:440] < btm_2[439:432]) ? 1 : 0;
assign detect_min[54][24] = (mid_1[447:440] < btm_2[447:440]) ? 1 : 0;
assign detect_min[54][25] = (mid_1[447:440] < btm_2[455:448]) ? 1 : 0;

assign detect_min[55][0] = (mid_1[455:448] < top_0[447:440]) ? 1 : 0;
assign detect_min[55][1] = (mid_1[455:448] < top_0[455:448]) ? 1 : 0;
assign detect_min[55][2] = (mid_1[455:448] < top_0[463:456]) ? 1 : 0;
assign detect_min[55][3] = (mid_1[455:448] < top_1[447:440]) ? 1 : 0;
assign detect_min[55][4] = (mid_1[455:448] < top_1[455:448]) ? 1 : 0;
assign detect_min[55][5] = (mid_1[455:448] < top_1[463:456]) ? 1 : 0;
assign detect_min[55][6] = (mid_1[455:448] < top_2[447:440]) ? 1 : 0;
assign detect_min[55][7] = (mid_1[455:448] < top_2[455:448]) ? 1 : 0;
assign detect_min[55][8] = (mid_1[455:448] < top_2[463:456]) ? 1 : 0;
assign detect_min[55][9] = (mid_1[455:448] < mid_0[447:440]) ? 1 : 0;
assign detect_min[55][10] = (mid_1[455:448] < mid_0[455:448]) ? 1 : 0;
assign detect_min[55][11] = (mid_1[455:448] < mid_0[463:456]) ? 1 : 0;
assign detect_min[55][12] = (mid_1[455:448] < mid_1[447:440]) ? 1 : 0;
assign detect_min[55][13] = (mid_1[455:448] < mid_1[463:456]) ? 1 : 0;
assign detect_min[55][14] = (mid_1[455:448] < mid_2[447:440]) ? 1 : 0;
assign detect_min[55][15] = (mid_1[455:448] < mid_2[455:448]) ? 1 : 0;
assign detect_min[55][16] = (mid_1[455:448] < mid_2[463:456]) ? 1 : 0;
assign detect_min[55][17] = (mid_1[455:448] < btm_0[447:440]) ? 1 : 0;
assign detect_min[55][18] = (mid_1[455:448] < btm_0[455:448]) ? 1 : 0;
assign detect_min[55][19] = (mid_1[455:448] < btm_0[463:456]) ? 1 : 0;
assign detect_min[55][20] = (mid_1[455:448] < btm_1[447:440]) ? 1 : 0;
assign detect_min[55][21] = (mid_1[455:448] < btm_1[455:448]) ? 1 : 0;
assign detect_min[55][22] = (mid_1[455:448] < btm_1[463:456]) ? 1 : 0;
assign detect_min[55][23] = (mid_1[455:448] < btm_2[447:440]) ? 1 : 0;
assign detect_min[55][24] = (mid_1[455:448] < btm_2[455:448]) ? 1 : 0;
assign detect_min[55][25] = (mid_1[455:448] < btm_2[463:456]) ? 1 : 0;

assign detect_min[56][0] = (mid_1[463:456] < top_0[455:448]) ? 1 : 0;
assign detect_min[56][1] = (mid_1[463:456] < top_0[463:456]) ? 1 : 0;
assign detect_min[56][2] = (mid_1[463:456] < top_0[471:464]) ? 1 : 0;
assign detect_min[56][3] = (mid_1[463:456] < top_1[455:448]) ? 1 : 0;
assign detect_min[56][4] = (mid_1[463:456] < top_1[463:456]) ? 1 : 0;
assign detect_min[56][5] = (mid_1[463:456] < top_1[471:464]) ? 1 : 0;
assign detect_min[56][6] = (mid_1[463:456] < top_2[455:448]) ? 1 : 0;
assign detect_min[56][7] = (mid_1[463:456] < top_2[463:456]) ? 1 : 0;
assign detect_min[56][8] = (mid_1[463:456] < top_2[471:464]) ? 1 : 0;
assign detect_min[56][9] = (mid_1[463:456] < mid_0[455:448]) ? 1 : 0;
assign detect_min[56][10] = (mid_1[463:456] < mid_0[463:456]) ? 1 : 0;
assign detect_min[56][11] = (mid_1[463:456] < mid_0[471:464]) ? 1 : 0;
assign detect_min[56][12] = (mid_1[463:456] < mid_1[455:448]) ? 1 : 0;
assign detect_min[56][13] = (mid_1[463:456] < mid_1[471:464]) ? 1 : 0;
assign detect_min[56][14] = (mid_1[463:456] < mid_2[455:448]) ? 1 : 0;
assign detect_min[56][15] = (mid_1[463:456] < mid_2[463:456]) ? 1 : 0;
assign detect_min[56][16] = (mid_1[463:456] < mid_2[471:464]) ? 1 : 0;
assign detect_min[56][17] = (mid_1[463:456] < btm_0[455:448]) ? 1 : 0;
assign detect_min[56][18] = (mid_1[463:456] < btm_0[463:456]) ? 1 : 0;
assign detect_min[56][19] = (mid_1[463:456] < btm_0[471:464]) ? 1 : 0;
assign detect_min[56][20] = (mid_1[463:456] < btm_1[455:448]) ? 1 : 0;
assign detect_min[56][21] = (mid_1[463:456] < btm_1[463:456]) ? 1 : 0;
assign detect_min[56][22] = (mid_1[463:456] < btm_1[471:464]) ? 1 : 0;
assign detect_min[56][23] = (mid_1[463:456] < btm_2[455:448]) ? 1 : 0;
assign detect_min[56][24] = (mid_1[463:456] < btm_2[463:456]) ? 1 : 0;
assign detect_min[56][25] = (mid_1[463:456] < btm_2[471:464]) ? 1 : 0;

assign detect_min[57][0] = (mid_1[471:464] < top_0[463:456]) ? 1 : 0;
assign detect_min[57][1] = (mid_1[471:464] < top_0[471:464]) ? 1 : 0;
assign detect_min[57][2] = (mid_1[471:464] < top_0[479:472]) ? 1 : 0;
assign detect_min[57][3] = (mid_1[471:464] < top_1[463:456]) ? 1 : 0;
assign detect_min[57][4] = (mid_1[471:464] < top_1[471:464]) ? 1 : 0;
assign detect_min[57][5] = (mid_1[471:464] < top_1[479:472]) ? 1 : 0;
assign detect_min[57][6] = (mid_1[471:464] < top_2[463:456]) ? 1 : 0;
assign detect_min[57][7] = (mid_1[471:464] < top_2[471:464]) ? 1 : 0;
assign detect_min[57][8] = (mid_1[471:464] < top_2[479:472]) ? 1 : 0;
assign detect_min[57][9] = (mid_1[471:464] < mid_0[463:456]) ? 1 : 0;
assign detect_min[57][10] = (mid_1[471:464] < mid_0[471:464]) ? 1 : 0;
assign detect_min[57][11] = (mid_1[471:464] < mid_0[479:472]) ? 1 : 0;
assign detect_min[57][12] = (mid_1[471:464] < mid_1[463:456]) ? 1 : 0;
assign detect_min[57][13] = (mid_1[471:464] < mid_1[479:472]) ? 1 : 0;
assign detect_min[57][14] = (mid_1[471:464] < mid_2[463:456]) ? 1 : 0;
assign detect_min[57][15] = (mid_1[471:464] < mid_2[471:464]) ? 1 : 0;
assign detect_min[57][16] = (mid_1[471:464] < mid_2[479:472]) ? 1 : 0;
assign detect_min[57][17] = (mid_1[471:464] < btm_0[463:456]) ? 1 : 0;
assign detect_min[57][18] = (mid_1[471:464] < btm_0[471:464]) ? 1 : 0;
assign detect_min[57][19] = (mid_1[471:464] < btm_0[479:472]) ? 1 : 0;
assign detect_min[57][20] = (mid_1[471:464] < btm_1[463:456]) ? 1 : 0;
assign detect_min[57][21] = (mid_1[471:464] < btm_1[471:464]) ? 1 : 0;
assign detect_min[57][22] = (mid_1[471:464] < btm_1[479:472]) ? 1 : 0;
assign detect_min[57][23] = (mid_1[471:464] < btm_2[463:456]) ? 1 : 0;
assign detect_min[57][24] = (mid_1[471:464] < btm_2[471:464]) ? 1 : 0;
assign detect_min[57][25] = (mid_1[471:464] < btm_2[479:472]) ? 1 : 0;

assign detect_min[58][0] = (mid_1[479:472] < top_0[471:464]) ? 1 : 0;
assign detect_min[58][1] = (mid_1[479:472] < top_0[479:472]) ? 1 : 0;
assign detect_min[58][2] = (mid_1[479:472] < top_0[487:480]) ? 1 : 0;
assign detect_min[58][3] = (mid_1[479:472] < top_1[471:464]) ? 1 : 0;
assign detect_min[58][4] = (mid_1[479:472] < top_1[479:472]) ? 1 : 0;
assign detect_min[58][5] = (mid_1[479:472] < top_1[487:480]) ? 1 : 0;
assign detect_min[58][6] = (mid_1[479:472] < top_2[471:464]) ? 1 : 0;
assign detect_min[58][7] = (mid_1[479:472] < top_2[479:472]) ? 1 : 0;
assign detect_min[58][8] = (mid_1[479:472] < top_2[487:480]) ? 1 : 0;
assign detect_min[58][9] = (mid_1[479:472] < mid_0[471:464]) ? 1 : 0;
assign detect_min[58][10] = (mid_1[479:472] < mid_0[479:472]) ? 1 : 0;
assign detect_min[58][11] = (mid_1[479:472] < mid_0[487:480]) ? 1 : 0;
assign detect_min[58][12] = (mid_1[479:472] < mid_1[471:464]) ? 1 : 0;
assign detect_min[58][13] = (mid_1[479:472] < mid_1[487:480]) ? 1 : 0;
assign detect_min[58][14] = (mid_1[479:472] < mid_2[471:464]) ? 1 : 0;
assign detect_min[58][15] = (mid_1[479:472] < mid_2[479:472]) ? 1 : 0;
assign detect_min[58][16] = (mid_1[479:472] < mid_2[487:480]) ? 1 : 0;
assign detect_min[58][17] = (mid_1[479:472] < btm_0[471:464]) ? 1 : 0;
assign detect_min[58][18] = (mid_1[479:472] < btm_0[479:472]) ? 1 : 0;
assign detect_min[58][19] = (mid_1[479:472] < btm_0[487:480]) ? 1 : 0;
assign detect_min[58][20] = (mid_1[479:472] < btm_1[471:464]) ? 1 : 0;
assign detect_min[58][21] = (mid_1[479:472] < btm_1[479:472]) ? 1 : 0;
assign detect_min[58][22] = (mid_1[479:472] < btm_1[487:480]) ? 1 : 0;
assign detect_min[58][23] = (mid_1[479:472] < btm_2[471:464]) ? 1 : 0;
assign detect_min[58][24] = (mid_1[479:472] < btm_2[479:472]) ? 1 : 0;
assign detect_min[58][25] = (mid_1[479:472] < btm_2[487:480]) ? 1 : 0;

assign detect_min[59][0] = (mid_1[487:480] < top_0[479:472]) ? 1 : 0;
assign detect_min[59][1] = (mid_1[487:480] < top_0[487:480]) ? 1 : 0;
assign detect_min[59][2] = (mid_1[487:480] < top_0[495:488]) ? 1 : 0;
assign detect_min[59][3] = (mid_1[487:480] < top_1[479:472]) ? 1 : 0;
assign detect_min[59][4] = (mid_1[487:480] < top_1[487:480]) ? 1 : 0;
assign detect_min[59][5] = (mid_1[487:480] < top_1[495:488]) ? 1 : 0;
assign detect_min[59][6] = (mid_1[487:480] < top_2[479:472]) ? 1 : 0;
assign detect_min[59][7] = (mid_1[487:480] < top_2[487:480]) ? 1 : 0;
assign detect_min[59][8] = (mid_1[487:480] < top_2[495:488]) ? 1 : 0;
assign detect_min[59][9] = (mid_1[487:480] < mid_0[479:472]) ? 1 : 0;
assign detect_min[59][10] = (mid_1[487:480] < mid_0[487:480]) ? 1 : 0;
assign detect_min[59][11] = (mid_1[487:480] < mid_0[495:488]) ? 1 : 0;
assign detect_min[59][12] = (mid_1[487:480] < mid_1[479:472]) ? 1 : 0;
assign detect_min[59][13] = (mid_1[487:480] < mid_1[495:488]) ? 1 : 0;
assign detect_min[59][14] = (mid_1[487:480] < mid_2[479:472]) ? 1 : 0;
assign detect_min[59][15] = (mid_1[487:480] < mid_2[487:480]) ? 1 : 0;
assign detect_min[59][16] = (mid_1[487:480] < mid_2[495:488]) ? 1 : 0;
assign detect_min[59][17] = (mid_1[487:480] < btm_0[479:472]) ? 1 : 0;
assign detect_min[59][18] = (mid_1[487:480] < btm_0[487:480]) ? 1 : 0;
assign detect_min[59][19] = (mid_1[487:480] < btm_0[495:488]) ? 1 : 0;
assign detect_min[59][20] = (mid_1[487:480] < btm_1[479:472]) ? 1 : 0;
assign detect_min[59][21] = (mid_1[487:480] < btm_1[487:480]) ? 1 : 0;
assign detect_min[59][22] = (mid_1[487:480] < btm_1[495:488]) ? 1 : 0;
assign detect_min[59][23] = (mid_1[487:480] < btm_2[479:472]) ? 1 : 0;
assign detect_min[59][24] = (mid_1[487:480] < btm_2[487:480]) ? 1 : 0;
assign detect_min[59][25] = (mid_1[487:480] < btm_2[495:488]) ? 1 : 0;

assign detect_min[60][0] = (mid_1[495:488] < top_0[487:480]) ? 1 : 0;
assign detect_min[60][1] = (mid_1[495:488] < top_0[495:488]) ? 1 : 0;
assign detect_min[60][2] = (mid_1[495:488] < top_0[503:496]) ? 1 : 0;
assign detect_min[60][3] = (mid_1[495:488] < top_1[487:480]) ? 1 : 0;
assign detect_min[60][4] = (mid_1[495:488] < top_1[495:488]) ? 1 : 0;
assign detect_min[60][5] = (mid_1[495:488] < top_1[503:496]) ? 1 : 0;
assign detect_min[60][6] = (mid_1[495:488] < top_2[487:480]) ? 1 : 0;
assign detect_min[60][7] = (mid_1[495:488] < top_2[495:488]) ? 1 : 0;
assign detect_min[60][8] = (mid_1[495:488] < top_2[503:496]) ? 1 : 0;
assign detect_min[60][9] = (mid_1[495:488] < mid_0[487:480]) ? 1 : 0;
assign detect_min[60][10] = (mid_1[495:488] < mid_0[495:488]) ? 1 : 0;
assign detect_min[60][11] = (mid_1[495:488] < mid_0[503:496]) ? 1 : 0;
assign detect_min[60][12] = (mid_1[495:488] < mid_1[487:480]) ? 1 : 0;
assign detect_min[60][13] = (mid_1[495:488] < mid_1[503:496]) ? 1 : 0;
assign detect_min[60][14] = (mid_1[495:488] < mid_2[487:480]) ? 1 : 0;
assign detect_min[60][15] = (mid_1[495:488] < mid_2[495:488]) ? 1 : 0;
assign detect_min[60][16] = (mid_1[495:488] < mid_2[503:496]) ? 1 : 0;
assign detect_min[60][17] = (mid_1[495:488] < btm_0[487:480]) ? 1 : 0;
assign detect_min[60][18] = (mid_1[495:488] < btm_0[495:488]) ? 1 : 0;
assign detect_min[60][19] = (mid_1[495:488] < btm_0[503:496]) ? 1 : 0;
assign detect_min[60][20] = (mid_1[495:488] < btm_1[487:480]) ? 1 : 0;
assign detect_min[60][21] = (mid_1[495:488] < btm_1[495:488]) ? 1 : 0;
assign detect_min[60][22] = (mid_1[495:488] < btm_1[503:496]) ? 1 : 0;
assign detect_min[60][23] = (mid_1[495:488] < btm_2[487:480]) ? 1 : 0;
assign detect_min[60][24] = (mid_1[495:488] < btm_2[495:488]) ? 1 : 0;
assign detect_min[60][25] = (mid_1[495:488] < btm_2[503:496]) ? 1 : 0;

assign detect_min[61][0] = (mid_1[503:496] < top_0[495:488]) ? 1 : 0;
assign detect_min[61][1] = (mid_1[503:496] < top_0[503:496]) ? 1 : 0;
assign detect_min[61][2] = (mid_1[503:496] < top_0[511:504]) ? 1 : 0;
assign detect_min[61][3] = (mid_1[503:496] < top_1[495:488]) ? 1 : 0;
assign detect_min[61][4] = (mid_1[503:496] < top_1[503:496]) ? 1 : 0;
assign detect_min[61][5] = (mid_1[503:496] < top_1[511:504]) ? 1 : 0;
assign detect_min[61][6] = (mid_1[503:496] < top_2[495:488]) ? 1 : 0;
assign detect_min[61][7] = (mid_1[503:496] < top_2[503:496]) ? 1 : 0;
assign detect_min[61][8] = (mid_1[503:496] < top_2[511:504]) ? 1 : 0;
assign detect_min[61][9] = (mid_1[503:496] < mid_0[495:488]) ? 1 : 0;
assign detect_min[61][10] = (mid_1[503:496] < mid_0[503:496]) ? 1 : 0;
assign detect_min[61][11] = (mid_1[503:496] < mid_0[511:504]) ? 1 : 0;
assign detect_min[61][12] = (mid_1[503:496] < mid_1[495:488]) ? 1 : 0;
assign detect_min[61][13] = (mid_1[503:496] < mid_1[511:504]) ? 1 : 0;
assign detect_min[61][14] = (mid_1[503:496] < mid_2[495:488]) ? 1 : 0;
assign detect_min[61][15] = (mid_1[503:496] < mid_2[503:496]) ? 1 : 0;
assign detect_min[61][16] = (mid_1[503:496] < mid_2[511:504]) ? 1 : 0;
assign detect_min[61][17] = (mid_1[503:496] < btm_0[495:488]) ? 1 : 0;
assign detect_min[61][18] = (mid_1[503:496] < btm_0[503:496]) ? 1 : 0;
assign detect_min[61][19] = (mid_1[503:496] < btm_0[511:504]) ? 1 : 0;
assign detect_min[61][20] = (mid_1[503:496] < btm_1[495:488]) ? 1 : 0;
assign detect_min[61][21] = (mid_1[503:496] < btm_1[503:496]) ? 1 : 0;
assign detect_min[61][22] = (mid_1[503:496] < btm_1[511:504]) ? 1 : 0;
assign detect_min[61][23] = (mid_1[503:496] < btm_2[495:488]) ? 1 : 0;
assign detect_min[61][24] = (mid_1[503:496] < btm_2[503:496]) ? 1 : 0;
assign detect_min[61][25] = (mid_1[503:496] < btm_2[511:504]) ? 1 : 0;

assign detect_min[62][0] = (mid_1[511:504] < top_0[503:496]) ? 1 : 0;
assign detect_min[62][1] = (mid_1[511:504] < top_0[511:504]) ? 1 : 0;
assign detect_min[62][2] = (mid_1[511:504] < top_0[519:512]) ? 1 : 0;
assign detect_min[62][3] = (mid_1[511:504] < top_1[503:496]) ? 1 : 0;
assign detect_min[62][4] = (mid_1[511:504] < top_1[511:504]) ? 1 : 0;
assign detect_min[62][5] = (mid_1[511:504] < top_1[519:512]) ? 1 : 0;
assign detect_min[62][6] = (mid_1[511:504] < top_2[503:496]) ? 1 : 0;
assign detect_min[62][7] = (mid_1[511:504] < top_2[511:504]) ? 1 : 0;
assign detect_min[62][8] = (mid_1[511:504] < top_2[519:512]) ? 1 : 0;
assign detect_min[62][9] = (mid_1[511:504] < mid_0[503:496]) ? 1 : 0;
assign detect_min[62][10] = (mid_1[511:504] < mid_0[511:504]) ? 1 : 0;
assign detect_min[62][11] = (mid_1[511:504] < mid_0[519:512]) ? 1 : 0;
assign detect_min[62][12] = (mid_1[511:504] < mid_1[503:496]) ? 1 : 0;
assign detect_min[62][13] = (mid_1[511:504] < mid_1[519:512]) ? 1 : 0;
assign detect_min[62][14] = (mid_1[511:504] < mid_2[503:496]) ? 1 : 0;
assign detect_min[62][15] = (mid_1[511:504] < mid_2[511:504]) ? 1 : 0;
assign detect_min[62][16] = (mid_1[511:504] < mid_2[519:512]) ? 1 : 0;
assign detect_min[62][17] = (mid_1[511:504] < btm_0[503:496]) ? 1 : 0;
assign detect_min[62][18] = (mid_1[511:504] < btm_0[511:504]) ? 1 : 0;
assign detect_min[62][19] = (mid_1[511:504] < btm_0[519:512]) ? 1 : 0;
assign detect_min[62][20] = (mid_1[511:504] < btm_1[503:496]) ? 1 : 0;
assign detect_min[62][21] = (mid_1[511:504] < btm_1[511:504]) ? 1 : 0;
assign detect_min[62][22] = (mid_1[511:504] < btm_1[519:512]) ? 1 : 0;
assign detect_min[62][23] = (mid_1[511:504] < btm_2[503:496]) ? 1 : 0;
assign detect_min[62][24] = (mid_1[511:504] < btm_2[511:504]) ? 1 : 0;
assign detect_min[62][25] = (mid_1[511:504] < btm_2[519:512]) ? 1 : 0;

assign detect_min[63][0] = (mid_1[519:512] < top_0[511:504]) ? 1 : 0;
assign detect_min[63][1] = (mid_1[519:512] < top_0[519:512]) ? 1 : 0;
assign detect_min[63][2] = (mid_1[519:512] < top_0[527:520]) ? 1 : 0;
assign detect_min[63][3] = (mid_1[519:512] < top_1[511:504]) ? 1 : 0;
assign detect_min[63][4] = (mid_1[519:512] < top_1[519:512]) ? 1 : 0;
assign detect_min[63][5] = (mid_1[519:512] < top_1[527:520]) ? 1 : 0;
assign detect_min[63][6] = (mid_1[519:512] < top_2[511:504]) ? 1 : 0;
assign detect_min[63][7] = (mid_1[519:512] < top_2[519:512]) ? 1 : 0;
assign detect_min[63][8] = (mid_1[519:512] < top_2[527:520]) ? 1 : 0;
assign detect_min[63][9] = (mid_1[519:512] < mid_0[511:504]) ? 1 : 0;
assign detect_min[63][10] = (mid_1[519:512] < mid_0[519:512]) ? 1 : 0;
assign detect_min[63][11] = (mid_1[519:512] < mid_0[527:520]) ? 1 : 0;
assign detect_min[63][12] = (mid_1[519:512] < mid_1[511:504]) ? 1 : 0;
assign detect_min[63][13] = (mid_1[519:512] < mid_1[527:520]) ? 1 : 0;
assign detect_min[63][14] = (mid_1[519:512] < mid_2[511:504]) ? 1 : 0;
assign detect_min[63][15] = (mid_1[519:512] < mid_2[519:512]) ? 1 : 0;
assign detect_min[63][16] = (mid_1[519:512] < mid_2[527:520]) ? 1 : 0;
assign detect_min[63][17] = (mid_1[519:512] < btm_0[511:504]) ? 1 : 0;
assign detect_min[63][18] = (mid_1[519:512] < btm_0[519:512]) ? 1 : 0;
assign detect_min[63][19] = (mid_1[519:512] < btm_0[527:520]) ? 1 : 0;
assign detect_min[63][20] = (mid_1[519:512] < btm_1[511:504]) ? 1 : 0;
assign detect_min[63][21] = (mid_1[519:512] < btm_1[519:512]) ? 1 : 0;
assign detect_min[63][22] = (mid_1[519:512] < btm_1[527:520]) ? 1 : 0;
assign detect_min[63][23] = (mid_1[519:512] < btm_2[511:504]) ? 1 : 0;
assign detect_min[63][24] = (mid_1[519:512] < btm_2[519:512]) ? 1 : 0;
assign detect_min[63][25] = (mid_1[519:512] < btm_2[527:520]) ? 1 : 0;

assign detect_min[64][0] = (mid_1[527:520] < top_0[519:512]) ? 1 : 0;
assign detect_min[64][1] = (mid_1[527:520] < top_0[527:520]) ? 1 : 0;
assign detect_min[64][2] = (mid_1[527:520] < top_0[535:528]) ? 1 : 0;
assign detect_min[64][3] = (mid_1[527:520] < top_1[519:512]) ? 1 : 0;
assign detect_min[64][4] = (mid_1[527:520] < top_1[527:520]) ? 1 : 0;
assign detect_min[64][5] = (mid_1[527:520] < top_1[535:528]) ? 1 : 0;
assign detect_min[64][6] = (mid_1[527:520] < top_2[519:512]) ? 1 : 0;
assign detect_min[64][7] = (mid_1[527:520] < top_2[527:520]) ? 1 : 0;
assign detect_min[64][8] = (mid_1[527:520] < top_2[535:528]) ? 1 : 0;
assign detect_min[64][9] = (mid_1[527:520] < mid_0[519:512]) ? 1 : 0;
assign detect_min[64][10] = (mid_1[527:520] < mid_0[527:520]) ? 1 : 0;
assign detect_min[64][11] = (mid_1[527:520] < mid_0[535:528]) ? 1 : 0;
assign detect_min[64][12] = (mid_1[527:520] < mid_1[519:512]) ? 1 : 0;
assign detect_min[64][13] = (mid_1[527:520] < mid_1[535:528]) ? 1 : 0;
assign detect_min[64][14] = (mid_1[527:520] < mid_2[519:512]) ? 1 : 0;
assign detect_min[64][15] = (mid_1[527:520] < mid_2[527:520]) ? 1 : 0;
assign detect_min[64][16] = (mid_1[527:520] < mid_2[535:528]) ? 1 : 0;
assign detect_min[64][17] = (mid_1[527:520] < btm_0[519:512]) ? 1 : 0;
assign detect_min[64][18] = (mid_1[527:520] < btm_0[527:520]) ? 1 : 0;
assign detect_min[64][19] = (mid_1[527:520] < btm_0[535:528]) ? 1 : 0;
assign detect_min[64][20] = (mid_1[527:520] < btm_1[519:512]) ? 1 : 0;
assign detect_min[64][21] = (mid_1[527:520] < btm_1[527:520]) ? 1 : 0;
assign detect_min[64][22] = (mid_1[527:520] < btm_1[535:528]) ? 1 : 0;
assign detect_min[64][23] = (mid_1[527:520] < btm_2[519:512]) ? 1 : 0;
assign detect_min[64][24] = (mid_1[527:520] < btm_2[527:520]) ? 1 : 0;
assign detect_min[64][25] = (mid_1[527:520] < btm_2[535:528]) ? 1 : 0;

assign detect_min[65][0] = (mid_1[535:528] < top_0[527:520]) ? 1 : 0;
assign detect_min[65][1] = (mid_1[535:528] < top_0[535:528]) ? 1 : 0;
assign detect_min[65][2] = (mid_1[535:528] < top_0[543:536]) ? 1 : 0;
assign detect_min[65][3] = (mid_1[535:528] < top_1[527:520]) ? 1 : 0;
assign detect_min[65][4] = (mid_1[535:528] < top_1[535:528]) ? 1 : 0;
assign detect_min[65][5] = (mid_1[535:528] < top_1[543:536]) ? 1 : 0;
assign detect_min[65][6] = (mid_1[535:528] < top_2[527:520]) ? 1 : 0;
assign detect_min[65][7] = (mid_1[535:528] < top_2[535:528]) ? 1 : 0;
assign detect_min[65][8] = (mid_1[535:528] < top_2[543:536]) ? 1 : 0;
assign detect_min[65][9] = (mid_1[535:528] < mid_0[527:520]) ? 1 : 0;
assign detect_min[65][10] = (mid_1[535:528] < mid_0[535:528]) ? 1 : 0;
assign detect_min[65][11] = (mid_1[535:528] < mid_0[543:536]) ? 1 : 0;
assign detect_min[65][12] = (mid_1[535:528] < mid_1[527:520]) ? 1 : 0;
assign detect_min[65][13] = (mid_1[535:528] < mid_1[543:536]) ? 1 : 0;
assign detect_min[65][14] = (mid_1[535:528] < mid_2[527:520]) ? 1 : 0;
assign detect_min[65][15] = (mid_1[535:528] < mid_2[535:528]) ? 1 : 0;
assign detect_min[65][16] = (mid_1[535:528] < mid_2[543:536]) ? 1 : 0;
assign detect_min[65][17] = (mid_1[535:528] < btm_0[527:520]) ? 1 : 0;
assign detect_min[65][18] = (mid_1[535:528] < btm_0[535:528]) ? 1 : 0;
assign detect_min[65][19] = (mid_1[535:528] < btm_0[543:536]) ? 1 : 0;
assign detect_min[65][20] = (mid_1[535:528] < btm_1[527:520]) ? 1 : 0;
assign detect_min[65][21] = (mid_1[535:528] < btm_1[535:528]) ? 1 : 0;
assign detect_min[65][22] = (mid_1[535:528] < btm_1[543:536]) ? 1 : 0;
assign detect_min[65][23] = (mid_1[535:528] < btm_2[527:520]) ? 1 : 0;
assign detect_min[65][24] = (mid_1[535:528] < btm_2[535:528]) ? 1 : 0;
assign detect_min[65][25] = (mid_1[535:528] < btm_2[543:536]) ? 1 : 0;

assign detect_min[66][0] = (mid_1[543:536] < top_0[535:528]) ? 1 : 0;
assign detect_min[66][1] = (mid_1[543:536] < top_0[543:536]) ? 1 : 0;
assign detect_min[66][2] = (mid_1[543:536] < top_0[551:544]) ? 1 : 0;
assign detect_min[66][3] = (mid_1[543:536] < top_1[535:528]) ? 1 : 0;
assign detect_min[66][4] = (mid_1[543:536] < top_1[543:536]) ? 1 : 0;
assign detect_min[66][5] = (mid_1[543:536] < top_1[551:544]) ? 1 : 0;
assign detect_min[66][6] = (mid_1[543:536] < top_2[535:528]) ? 1 : 0;
assign detect_min[66][7] = (mid_1[543:536] < top_2[543:536]) ? 1 : 0;
assign detect_min[66][8] = (mid_1[543:536] < top_2[551:544]) ? 1 : 0;
assign detect_min[66][9] = (mid_1[543:536] < mid_0[535:528]) ? 1 : 0;
assign detect_min[66][10] = (mid_1[543:536] < mid_0[543:536]) ? 1 : 0;
assign detect_min[66][11] = (mid_1[543:536] < mid_0[551:544]) ? 1 : 0;
assign detect_min[66][12] = (mid_1[543:536] < mid_1[535:528]) ? 1 : 0;
assign detect_min[66][13] = (mid_1[543:536] < mid_1[551:544]) ? 1 : 0;
assign detect_min[66][14] = (mid_1[543:536] < mid_2[535:528]) ? 1 : 0;
assign detect_min[66][15] = (mid_1[543:536] < mid_2[543:536]) ? 1 : 0;
assign detect_min[66][16] = (mid_1[543:536] < mid_2[551:544]) ? 1 : 0;
assign detect_min[66][17] = (mid_1[543:536] < btm_0[535:528]) ? 1 : 0;
assign detect_min[66][18] = (mid_1[543:536] < btm_0[543:536]) ? 1 : 0;
assign detect_min[66][19] = (mid_1[543:536] < btm_0[551:544]) ? 1 : 0;
assign detect_min[66][20] = (mid_1[543:536] < btm_1[535:528]) ? 1 : 0;
assign detect_min[66][21] = (mid_1[543:536] < btm_1[543:536]) ? 1 : 0;
assign detect_min[66][22] = (mid_1[543:536] < btm_1[551:544]) ? 1 : 0;
assign detect_min[66][23] = (mid_1[543:536] < btm_2[535:528]) ? 1 : 0;
assign detect_min[66][24] = (mid_1[543:536] < btm_2[543:536]) ? 1 : 0;
assign detect_min[66][25] = (mid_1[543:536] < btm_2[551:544]) ? 1 : 0;

assign detect_min[67][0] = (mid_1[551:544] < top_0[543:536]) ? 1 : 0;
assign detect_min[67][1] = (mid_1[551:544] < top_0[551:544]) ? 1 : 0;
assign detect_min[67][2] = (mid_1[551:544] < top_0[559:552]) ? 1 : 0;
assign detect_min[67][3] = (mid_1[551:544] < top_1[543:536]) ? 1 : 0;
assign detect_min[67][4] = (mid_1[551:544] < top_1[551:544]) ? 1 : 0;
assign detect_min[67][5] = (mid_1[551:544] < top_1[559:552]) ? 1 : 0;
assign detect_min[67][6] = (mid_1[551:544] < top_2[543:536]) ? 1 : 0;
assign detect_min[67][7] = (mid_1[551:544] < top_2[551:544]) ? 1 : 0;
assign detect_min[67][8] = (mid_1[551:544] < top_2[559:552]) ? 1 : 0;
assign detect_min[67][9] = (mid_1[551:544] < mid_0[543:536]) ? 1 : 0;
assign detect_min[67][10] = (mid_1[551:544] < mid_0[551:544]) ? 1 : 0;
assign detect_min[67][11] = (mid_1[551:544] < mid_0[559:552]) ? 1 : 0;
assign detect_min[67][12] = (mid_1[551:544] < mid_1[543:536]) ? 1 : 0;
assign detect_min[67][13] = (mid_1[551:544] < mid_1[559:552]) ? 1 : 0;
assign detect_min[67][14] = (mid_1[551:544] < mid_2[543:536]) ? 1 : 0;
assign detect_min[67][15] = (mid_1[551:544] < mid_2[551:544]) ? 1 : 0;
assign detect_min[67][16] = (mid_1[551:544] < mid_2[559:552]) ? 1 : 0;
assign detect_min[67][17] = (mid_1[551:544] < btm_0[543:536]) ? 1 : 0;
assign detect_min[67][18] = (mid_1[551:544] < btm_0[551:544]) ? 1 : 0;
assign detect_min[67][19] = (mid_1[551:544] < btm_0[559:552]) ? 1 : 0;
assign detect_min[67][20] = (mid_1[551:544] < btm_1[543:536]) ? 1 : 0;
assign detect_min[67][21] = (mid_1[551:544] < btm_1[551:544]) ? 1 : 0;
assign detect_min[67][22] = (mid_1[551:544] < btm_1[559:552]) ? 1 : 0;
assign detect_min[67][23] = (mid_1[551:544] < btm_2[543:536]) ? 1 : 0;
assign detect_min[67][24] = (mid_1[551:544] < btm_2[551:544]) ? 1 : 0;
assign detect_min[67][25] = (mid_1[551:544] < btm_2[559:552]) ? 1 : 0;

assign detect_min[68][0] = (mid_1[559:552] < top_0[551:544]) ? 1 : 0;
assign detect_min[68][1] = (mid_1[559:552] < top_0[559:552]) ? 1 : 0;
assign detect_min[68][2] = (mid_1[559:552] < top_0[567:560]) ? 1 : 0;
assign detect_min[68][3] = (mid_1[559:552] < top_1[551:544]) ? 1 : 0;
assign detect_min[68][4] = (mid_1[559:552] < top_1[559:552]) ? 1 : 0;
assign detect_min[68][5] = (mid_1[559:552] < top_1[567:560]) ? 1 : 0;
assign detect_min[68][6] = (mid_1[559:552] < top_2[551:544]) ? 1 : 0;
assign detect_min[68][7] = (mid_1[559:552] < top_2[559:552]) ? 1 : 0;
assign detect_min[68][8] = (mid_1[559:552] < top_2[567:560]) ? 1 : 0;
assign detect_min[68][9] = (mid_1[559:552] < mid_0[551:544]) ? 1 : 0;
assign detect_min[68][10] = (mid_1[559:552] < mid_0[559:552]) ? 1 : 0;
assign detect_min[68][11] = (mid_1[559:552] < mid_0[567:560]) ? 1 : 0;
assign detect_min[68][12] = (mid_1[559:552] < mid_1[551:544]) ? 1 : 0;
assign detect_min[68][13] = (mid_1[559:552] < mid_1[567:560]) ? 1 : 0;
assign detect_min[68][14] = (mid_1[559:552] < mid_2[551:544]) ? 1 : 0;
assign detect_min[68][15] = (mid_1[559:552] < mid_2[559:552]) ? 1 : 0;
assign detect_min[68][16] = (mid_1[559:552] < mid_2[567:560]) ? 1 : 0;
assign detect_min[68][17] = (mid_1[559:552] < btm_0[551:544]) ? 1 : 0;
assign detect_min[68][18] = (mid_1[559:552] < btm_0[559:552]) ? 1 : 0;
assign detect_min[68][19] = (mid_1[559:552] < btm_0[567:560]) ? 1 : 0;
assign detect_min[68][20] = (mid_1[559:552] < btm_1[551:544]) ? 1 : 0;
assign detect_min[68][21] = (mid_1[559:552] < btm_1[559:552]) ? 1 : 0;
assign detect_min[68][22] = (mid_1[559:552] < btm_1[567:560]) ? 1 : 0;
assign detect_min[68][23] = (mid_1[559:552] < btm_2[551:544]) ? 1 : 0;
assign detect_min[68][24] = (mid_1[559:552] < btm_2[559:552]) ? 1 : 0;
assign detect_min[68][25] = (mid_1[559:552] < btm_2[567:560]) ? 1 : 0;

assign detect_min[69][0] = (mid_1[567:560] < top_0[559:552]) ? 1 : 0;
assign detect_min[69][1] = (mid_1[567:560] < top_0[567:560]) ? 1 : 0;
assign detect_min[69][2] = (mid_1[567:560] < top_0[575:568]) ? 1 : 0;
assign detect_min[69][3] = (mid_1[567:560] < top_1[559:552]) ? 1 : 0;
assign detect_min[69][4] = (mid_1[567:560] < top_1[567:560]) ? 1 : 0;
assign detect_min[69][5] = (mid_1[567:560] < top_1[575:568]) ? 1 : 0;
assign detect_min[69][6] = (mid_1[567:560] < top_2[559:552]) ? 1 : 0;
assign detect_min[69][7] = (mid_1[567:560] < top_2[567:560]) ? 1 : 0;
assign detect_min[69][8] = (mid_1[567:560] < top_2[575:568]) ? 1 : 0;
assign detect_min[69][9] = (mid_1[567:560] < mid_0[559:552]) ? 1 : 0;
assign detect_min[69][10] = (mid_1[567:560] < mid_0[567:560]) ? 1 : 0;
assign detect_min[69][11] = (mid_1[567:560] < mid_0[575:568]) ? 1 : 0;
assign detect_min[69][12] = (mid_1[567:560] < mid_1[559:552]) ? 1 : 0;
assign detect_min[69][13] = (mid_1[567:560] < mid_1[575:568]) ? 1 : 0;
assign detect_min[69][14] = (mid_1[567:560] < mid_2[559:552]) ? 1 : 0;
assign detect_min[69][15] = (mid_1[567:560] < mid_2[567:560]) ? 1 : 0;
assign detect_min[69][16] = (mid_1[567:560] < mid_2[575:568]) ? 1 : 0;
assign detect_min[69][17] = (mid_1[567:560] < btm_0[559:552]) ? 1 : 0;
assign detect_min[69][18] = (mid_1[567:560] < btm_0[567:560]) ? 1 : 0;
assign detect_min[69][19] = (mid_1[567:560] < btm_0[575:568]) ? 1 : 0;
assign detect_min[69][20] = (mid_1[567:560] < btm_1[559:552]) ? 1 : 0;
assign detect_min[69][21] = (mid_1[567:560] < btm_1[567:560]) ? 1 : 0;
assign detect_min[69][22] = (mid_1[567:560] < btm_1[575:568]) ? 1 : 0;
assign detect_min[69][23] = (mid_1[567:560] < btm_2[559:552]) ? 1 : 0;
assign detect_min[69][24] = (mid_1[567:560] < btm_2[567:560]) ? 1 : 0;
assign detect_min[69][25] = (mid_1[567:560] < btm_2[575:568]) ? 1 : 0;

assign detect_min[70][0] = (mid_1[575:568] < top_0[567:560]) ? 1 : 0;
assign detect_min[70][1] = (mid_1[575:568] < top_0[575:568]) ? 1 : 0;
assign detect_min[70][2] = (mid_1[575:568] < top_0[583:576]) ? 1 : 0;
assign detect_min[70][3] = (mid_1[575:568] < top_1[567:560]) ? 1 : 0;
assign detect_min[70][4] = (mid_1[575:568] < top_1[575:568]) ? 1 : 0;
assign detect_min[70][5] = (mid_1[575:568] < top_1[583:576]) ? 1 : 0;
assign detect_min[70][6] = (mid_1[575:568] < top_2[567:560]) ? 1 : 0;
assign detect_min[70][7] = (mid_1[575:568] < top_2[575:568]) ? 1 : 0;
assign detect_min[70][8] = (mid_1[575:568] < top_2[583:576]) ? 1 : 0;
assign detect_min[70][9] = (mid_1[575:568] < mid_0[567:560]) ? 1 : 0;
assign detect_min[70][10] = (mid_1[575:568] < mid_0[575:568]) ? 1 : 0;
assign detect_min[70][11] = (mid_1[575:568] < mid_0[583:576]) ? 1 : 0;
assign detect_min[70][12] = (mid_1[575:568] < mid_1[567:560]) ? 1 : 0;
assign detect_min[70][13] = (mid_1[575:568] < mid_1[583:576]) ? 1 : 0;
assign detect_min[70][14] = (mid_1[575:568] < mid_2[567:560]) ? 1 : 0;
assign detect_min[70][15] = (mid_1[575:568] < mid_2[575:568]) ? 1 : 0;
assign detect_min[70][16] = (mid_1[575:568] < mid_2[583:576]) ? 1 : 0;
assign detect_min[70][17] = (mid_1[575:568] < btm_0[567:560]) ? 1 : 0;
assign detect_min[70][18] = (mid_1[575:568] < btm_0[575:568]) ? 1 : 0;
assign detect_min[70][19] = (mid_1[575:568] < btm_0[583:576]) ? 1 : 0;
assign detect_min[70][20] = (mid_1[575:568] < btm_1[567:560]) ? 1 : 0;
assign detect_min[70][21] = (mid_1[575:568] < btm_1[575:568]) ? 1 : 0;
assign detect_min[70][22] = (mid_1[575:568] < btm_1[583:576]) ? 1 : 0;
assign detect_min[70][23] = (mid_1[575:568] < btm_2[567:560]) ? 1 : 0;
assign detect_min[70][24] = (mid_1[575:568] < btm_2[575:568]) ? 1 : 0;
assign detect_min[70][25] = (mid_1[575:568] < btm_2[583:576]) ? 1 : 0;

assign detect_min[71][0] = (mid_1[583:576] < top_0[575:568]) ? 1 : 0;
assign detect_min[71][1] = (mid_1[583:576] < top_0[583:576]) ? 1 : 0;
assign detect_min[71][2] = (mid_1[583:576] < top_0[591:584]) ? 1 : 0;
assign detect_min[71][3] = (mid_1[583:576] < top_1[575:568]) ? 1 : 0;
assign detect_min[71][4] = (mid_1[583:576] < top_1[583:576]) ? 1 : 0;
assign detect_min[71][5] = (mid_1[583:576] < top_1[591:584]) ? 1 : 0;
assign detect_min[71][6] = (mid_1[583:576] < top_2[575:568]) ? 1 : 0;
assign detect_min[71][7] = (mid_1[583:576] < top_2[583:576]) ? 1 : 0;
assign detect_min[71][8] = (mid_1[583:576] < top_2[591:584]) ? 1 : 0;
assign detect_min[71][9] = (mid_1[583:576] < mid_0[575:568]) ? 1 : 0;
assign detect_min[71][10] = (mid_1[583:576] < mid_0[583:576]) ? 1 : 0;
assign detect_min[71][11] = (mid_1[583:576] < mid_0[591:584]) ? 1 : 0;
assign detect_min[71][12] = (mid_1[583:576] < mid_1[575:568]) ? 1 : 0;
assign detect_min[71][13] = (mid_1[583:576] < mid_1[591:584]) ? 1 : 0;
assign detect_min[71][14] = (mid_1[583:576] < mid_2[575:568]) ? 1 : 0;
assign detect_min[71][15] = (mid_1[583:576] < mid_2[583:576]) ? 1 : 0;
assign detect_min[71][16] = (mid_1[583:576] < mid_2[591:584]) ? 1 : 0;
assign detect_min[71][17] = (mid_1[583:576] < btm_0[575:568]) ? 1 : 0;
assign detect_min[71][18] = (mid_1[583:576] < btm_0[583:576]) ? 1 : 0;
assign detect_min[71][19] = (mid_1[583:576] < btm_0[591:584]) ? 1 : 0;
assign detect_min[71][20] = (mid_1[583:576] < btm_1[575:568]) ? 1 : 0;
assign detect_min[71][21] = (mid_1[583:576] < btm_1[583:576]) ? 1 : 0;
assign detect_min[71][22] = (mid_1[583:576] < btm_1[591:584]) ? 1 : 0;
assign detect_min[71][23] = (mid_1[583:576] < btm_2[575:568]) ? 1 : 0;
assign detect_min[71][24] = (mid_1[583:576] < btm_2[583:576]) ? 1 : 0;
assign detect_min[71][25] = (mid_1[583:576] < btm_2[591:584]) ? 1 : 0;

assign detect_min[72][0] = (mid_1[591:584] < top_0[583:576]) ? 1 : 0;
assign detect_min[72][1] = (mid_1[591:584] < top_0[591:584]) ? 1 : 0;
assign detect_min[72][2] = (mid_1[591:584] < top_0[599:592]) ? 1 : 0;
assign detect_min[72][3] = (mid_1[591:584] < top_1[583:576]) ? 1 : 0;
assign detect_min[72][4] = (mid_1[591:584] < top_1[591:584]) ? 1 : 0;
assign detect_min[72][5] = (mid_1[591:584] < top_1[599:592]) ? 1 : 0;
assign detect_min[72][6] = (mid_1[591:584] < top_2[583:576]) ? 1 : 0;
assign detect_min[72][7] = (mid_1[591:584] < top_2[591:584]) ? 1 : 0;
assign detect_min[72][8] = (mid_1[591:584] < top_2[599:592]) ? 1 : 0;
assign detect_min[72][9] = (mid_1[591:584] < mid_0[583:576]) ? 1 : 0;
assign detect_min[72][10] = (mid_1[591:584] < mid_0[591:584]) ? 1 : 0;
assign detect_min[72][11] = (mid_1[591:584] < mid_0[599:592]) ? 1 : 0;
assign detect_min[72][12] = (mid_1[591:584] < mid_1[583:576]) ? 1 : 0;
assign detect_min[72][13] = (mid_1[591:584] < mid_1[599:592]) ? 1 : 0;
assign detect_min[72][14] = (mid_1[591:584] < mid_2[583:576]) ? 1 : 0;
assign detect_min[72][15] = (mid_1[591:584] < mid_2[591:584]) ? 1 : 0;
assign detect_min[72][16] = (mid_1[591:584] < mid_2[599:592]) ? 1 : 0;
assign detect_min[72][17] = (mid_1[591:584] < btm_0[583:576]) ? 1 : 0;
assign detect_min[72][18] = (mid_1[591:584] < btm_0[591:584]) ? 1 : 0;
assign detect_min[72][19] = (mid_1[591:584] < btm_0[599:592]) ? 1 : 0;
assign detect_min[72][20] = (mid_1[591:584] < btm_1[583:576]) ? 1 : 0;
assign detect_min[72][21] = (mid_1[591:584] < btm_1[591:584]) ? 1 : 0;
assign detect_min[72][22] = (mid_1[591:584] < btm_1[599:592]) ? 1 : 0;
assign detect_min[72][23] = (mid_1[591:584] < btm_2[583:576]) ? 1 : 0;
assign detect_min[72][24] = (mid_1[591:584] < btm_2[591:584]) ? 1 : 0;
assign detect_min[72][25] = (mid_1[591:584] < btm_2[599:592]) ? 1 : 0;

assign detect_min[73][0] = (mid_1[599:592] < top_0[591:584]) ? 1 : 0;
assign detect_min[73][1] = (mid_1[599:592] < top_0[599:592]) ? 1 : 0;
assign detect_min[73][2] = (mid_1[599:592] < top_0[607:600]) ? 1 : 0;
assign detect_min[73][3] = (mid_1[599:592] < top_1[591:584]) ? 1 : 0;
assign detect_min[73][4] = (mid_1[599:592] < top_1[599:592]) ? 1 : 0;
assign detect_min[73][5] = (mid_1[599:592] < top_1[607:600]) ? 1 : 0;
assign detect_min[73][6] = (mid_1[599:592] < top_2[591:584]) ? 1 : 0;
assign detect_min[73][7] = (mid_1[599:592] < top_2[599:592]) ? 1 : 0;
assign detect_min[73][8] = (mid_1[599:592] < top_2[607:600]) ? 1 : 0;
assign detect_min[73][9] = (mid_1[599:592] < mid_0[591:584]) ? 1 : 0;
assign detect_min[73][10] = (mid_1[599:592] < mid_0[599:592]) ? 1 : 0;
assign detect_min[73][11] = (mid_1[599:592] < mid_0[607:600]) ? 1 : 0;
assign detect_min[73][12] = (mid_1[599:592] < mid_1[591:584]) ? 1 : 0;
assign detect_min[73][13] = (mid_1[599:592] < mid_1[607:600]) ? 1 : 0;
assign detect_min[73][14] = (mid_1[599:592] < mid_2[591:584]) ? 1 : 0;
assign detect_min[73][15] = (mid_1[599:592] < mid_2[599:592]) ? 1 : 0;
assign detect_min[73][16] = (mid_1[599:592] < mid_2[607:600]) ? 1 : 0;
assign detect_min[73][17] = (mid_1[599:592] < btm_0[591:584]) ? 1 : 0;
assign detect_min[73][18] = (mid_1[599:592] < btm_0[599:592]) ? 1 : 0;
assign detect_min[73][19] = (mid_1[599:592] < btm_0[607:600]) ? 1 : 0;
assign detect_min[73][20] = (mid_1[599:592] < btm_1[591:584]) ? 1 : 0;
assign detect_min[73][21] = (mid_1[599:592] < btm_1[599:592]) ? 1 : 0;
assign detect_min[73][22] = (mid_1[599:592] < btm_1[607:600]) ? 1 : 0;
assign detect_min[73][23] = (mid_1[599:592] < btm_2[591:584]) ? 1 : 0;
assign detect_min[73][24] = (mid_1[599:592] < btm_2[599:592]) ? 1 : 0;
assign detect_min[73][25] = (mid_1[599:592] < btm_2[607:600]) ? 1 : 0;

assign detect_min[74][0] = (mid_1[607:600] < top_0[599:592]) ? 1 : 0;
assign detect_min[74][1] = (mid_1[607:600] < top_0[607:600]) ? 1 : 0;
assign detect_min[74][2] = (mid_1[607:600] < top_0[615:608]) ? 1 : 0;
assign detect_min[74][3] = (mid_1[607:600] < top_1[599:592]) ? 1 : 0;
assign detect_min[74][4] = (mid_1[607:600] < top_1[607:600]) ? 1 : 0;
assign detect_min[74][5] = (mid_1[607:600] < top_1[615:608]) ? 1 : 0;
assign detect_min[74][6] = (mid_1[607:600] < top_2[599:592]) ? 1 : 0;
assign detect_min[74][7] = (mid_1[607:600] < top_2[607:600]) ? 1 : 0;
assign detect_min[74][8] = (mid_1[607:600] < top_2[615:608]) ? 1 : 0;
assign detect_min[74][9] = (mid_1[607:600] < mid_0[599:592]) ? 1 : 0;
assign detect_min[74][10] = (mid_1[607:600] < mid_0[607:600]) ? 1 : 0;
assign detect_min[74][11] = (mid_1[607:600] < mid_0[615:608]) ? 1 : 0;
assign detect_min[74][12] = (mid_1[607:600] < mid_1[599:592]) ? 1 : 0;
assign detect_min[74][13] = (mid_1[607:600] < mid_1[615:608]) ? 1 : 0;
assign detect_min[74][14] = (mid_1[607:600] < mid_2[599:592]) ? 1 : 0;
assign detect_min[74][15] = (mid_1[607:600] < mid_2[607:600]) ? 1 : 0;
assign detect_min[74][16] = (mid_1[607:600] < mid_2[615:608]) ? 1 : 0;
assign detect_min[74][17] = (mid_1[607:600] < btm_0[599:592]) ? 1 : 0;
assign detect_min[74][18] = (mid_1[607:600] < btm_0[607:600]) ? 1 : 0;
assign detect_min[74][19] = (mid_1[607:600] < btm_0[615:608]) ? 1 : 0;
assign detect_min[74][20] = (mid_1[607:600] < btm_1[599:592]) ? 1 : 0;
assign detect_min[74][21] = (mid_1[607:600] < btm_1[607:600]) ? 1 : 0;
assign detect_min[74][22] = (mid_1[607:600] < btm_1[615:608]) ? 1 : 0;
assign detect_min[74][23] = (mid_1[607:600] < btm_2[599:592]) ? 1 : 0;
assign detect_min[74][24] = (mid_1[607:600] < btm_2[607:600]) ? 1 : 0;
assign detect_min[74][25] = (mid_1[607:600] < btm_2[615:608]) ? 1 : 0;

assign detect_min[75][0] = (mid_1[615:608] < top_0[607:600]) ? 1 : 0;
assign detect_min[75][1] = (mid_1[615:608] < top_0[615:608]) ? 1 : 0;
assign detect_min[75][2] = (mid_1[615:608] < top_0[623:616]) ? 1 : 0;
assign detect_min[75][3] = (mid_1[615:608] < top_1[607:600]) ? 1 : 0;
assign detect_min[75][4] = (mid_1[615:608] < top_1[615:608]) ? 1 : 0;
assign detect_min[75][5] = (mid_1[615:608] < top_1[623:616]) ? 1 : 0;
assign detect_min[75][6] = (mid_1[615:608] < top_2[607:600]) ? 1 : 0;
assign detect_min[75][7] = (mid_1[615:608] < top_2[615:608]) ? 1 : 0;
assign detect_min[75][8] = (mid_1[615:608] < top_2[623:616]) ? 1 : 0;
assign detect_min[75][9] = (mid_1[615:608] < mid_0[607:600]) ? 1 : 0;
assign detect_min[75][10] = (mid_1[615:608] < mid_0[615:608]) ? 1 : 0;
assign detect_min[75][11] = (mid_1[615:608] < mid_0[623:616]) ? 1 : 0;
assign detect_min[75][12] = (mid_1[615:608] < mid_1[607:600]) ? 1 : 0;
assign detect_min[75][13] = (mid_1[615:608] < mid_1[623:616]) ? 1 : 0;
assign detect_min[75][14] = (mid_1[615:608] < mid_2[607:600]) ? 1 : 0;
assign detect_min[75][15] = (mid_1[615:608] < mid_2[615:608]) ? 1 : 0;
assign detect_min[75][16] = (mid_1[615:608] < mid_2[623:616]) ? 1 : 0;
assign detect_min[75][17] = (mid_1[615:608] < btm_0[607:600]) ? 1 : 0;
assign detect_min[75][18] = (mid_1[615:608] < btm_0[615:608]) ? 1 : 0;
assign detect_min[75][19] = (mid_1[615:608] < btm_0[623:616]) ? 1 : 0;
assign detect_min[75][20] = (mid_1[615:608] < btm_1[607:600]) ? 1 : 0;
assign detect_min[75][21] = (mid_1[615:608] < btm_1[615:608]) ? 1 : 0;
assign detect_min[75][22] = (mid_1[615:608] < btm_1[623:616]) ? 1 : 0;
assign detect_min[75][23] = (mid_1[615:608] < btm_2[607:600]) ? 1 : 0;
assign detect_min[75][24] = (mid_1[615:608] < btm_2[615:608]) ? 1 : 0;
assign detect_min[75][25] = (mid_1[615:608] < btm_2[623:616]) ? 1 : 0;

assign detect_min[76][0] = (mid_1[623:616] < top_0[615:608]) ? 1 : 0;
assign detect_min[76][1] = (mid_1[623:616] < top_0[623:616]) ? 1 : 0;
assign detect_min[76][2] = (mid_1[623:616] < top_0[631:624]) ? 1 : 0;
assign detect_min[76][3] = (mid_1[623:616] < top_1[615:608]) ? 1 : 0;
assign detect_min[76][4] = (mid_1[623:616] < top_1[623:616]) ? 1 : 0;
assign detect_min[76][5] = (mid_1[623:616] < top_1[631:624]) ? 1 : 0;
assign detect_min[76][6] = (mid_1[623:616] < top_2[615:608]) ? 1 : 0;
assign detect_min[76][7] = (mid_1[623:616] < top_2[623:616]) ? 1 : 0;
assign detect_min[76][8] = (mid_1[623:616] < top_2[631:624]) ? 1 : 0;
assign detect_min[76][9] = (mid_1[623:616] < mid_0[615:608]) ? 1 : 0;
assign detect_min[76][10] = (mid_1[623:616] < mid_0[623:616]) ? 1 : 0;
assign detect_min[76][11] = (mid_1[623:616] < mid_0[631:624]) ? 1 : 0;
assign detect_min[76][12] = (mid_1[623:616] < mid_1[615:608]) ? 1 : 0;
assign detect_min[76][13] = (mid_1[623:616] < mid_1[631:624]) ? 1 : 0;
assign detect_min[76][14] = (mid_1[623:616] < mid_2[615:608]) ? 1 : 0;
assign detect_min[76][15] = (mid_1[623:616] < mid_2[623:616]) ? 1 : 0;
assign detect_min[76][16] = (mid_1[623:616] < mid_2[631:624]) ? 1 : 0;
assign detect_min[76][17] = (mid_1[623:616] < btm_0[615:608]) ? 1 : 0;
assign detect_min[76][18] = (mid_1[623:616] < btm_0[623:616]) ? 1 : 0;
assign detect_min[76][19] = (mid_1[623:616] < btm_0[631:624]) ? 1 : 0;
assign detect_min[76][20] = (mid_1[623:616] < btm_1[615:608]) ? 1 : 0;
assign detect_min[76][21] = (mid_1[623:616] < btm_1[623:616]) ? 1 : 0;
assign detect_min[76][22] = (mid_1[623:616] < btm_1[631:624]) ? 1 : 0;
assign detect_min[76][23] = (mid_1[623:616] < btm_2[615:608]) ? 1 : 0;
assign detect_min[76][24] = (mid_1[623:616] < btm_2[623:616]) ? 1 : 0;
assign detect_min[76][25] = (mid_1[623:616] < btm_2[631:624]) ? 1 : 0;

assign detect_min[77][0] = (mid_1[631:624] < top_0[623:616]) ? 1 : 0;
assign detect_min[77][1] = (mid_1[631:624] < top_0[631:624]) ? 1 : 0;
assign detect_min[77][2] = (mid_1[631:624] < top_0[639:632]) ? 1 : 0;
assign detect_min[77][3] = (mid_1[631:624] < top_1[623:616]) ? 1 : 0;
assign detect_min[77][4] = (mid_1[631:624] < top_1[631:624]) ? 1 : 0;
assign detect_min[77][5] = (mid_1[631:624] < top_1[639:632]) ? 1 : 0;
assign detect_min[77][6] = (mid_1[631:624] < top_2[623:616]) ? 1 : 0;
assign detect_min[77][7] = (mid_1[631:624] < top_2[631:624]) ? 1 : 0;
assign detect_min[77][8] = (mid_1[631:624] < top_2[639:632]) ? 1 : 0;
assign detect_min[77][9] = (mid_1[631:624] < mid_0[623:616]) ? 1 : 0;
assign detect_min[77][10] = (mid_1[631:624] < mid_0[631:624]) ? 1 : 0;
assign detect_min[77][11] = (mid_1[631:624] < mid_0[639:632]) ? 1 : 0;
assign detect_min[77][12] = (mid_1[631:624] < mid_1[623:616]) ? 1 : 0;
assign detect_min[77][13] = (mid_1[631:624] < mid_1[639:632]) ? 1 : 0;
assign detect_min[77][14] = (mid_1[631:624] < mid_2[623:616]) ? 1 : 0;
assign detect_min[77][15] = (mid_1[631:624] < mid_2[631:624]) ? 1 : 0;
assign detect_min[77][16] = (mid_1[631:624] < mid_2[639:632]) ? 1 : 0;
assign detect_min[77][17] = (mid_1[631:624] < btm_0[623:616]) ? 1 : 0;
assign detect_min[77][18] = (mid_1[631:624] < btm_0[631:624]) ? 1 : 0;
assign detect_min[77][19] = (mid_1[631:624] < btm_0[639:632]) ? 1 : 0;
assign detect_min[77][20] = (mid_1[631:624] < btm_1[623:616]) ? 1 : 0;
assign detect_min[77][21] = (mid_1[631:624] < btm_1[631:624]) ? 1 : 0;
assign detect_min[77][22] = (mid_1[631:624] < btm_1[639:632]) ? 1 : 0;
assign detect_min[77][23] = (mid_1[631:624] < btm_2[623:616]) ? 1 : 0;
assign detect_min[77][24] = (mid_1[631:624] < btm_2[631:624]) ? 1 : 0;
assign detect_min[77][25] = (mid_1[631:624] < btm_2[639:632]) ? 1 : 0;

assign detect_min[78][0] = (mid_1[639:632] < top_0[631:624]) ? 1 : 0;
assign detect_min[78][1] = (mid_1[639:632] < top_0[639:632]) ? 1 : 0;
assign detect_min[78][2] = (mid_1[639:632] < top_0[647:640]) ? 1 : 0;
assign detect_min[78][3] = (mid_1[639:632] < top_1[631:624]) ? 1 : 0;
assign detect_min[78][4] = (mid_1[639:632] < top_1[639:632]) ? 1 : 0;
assign detect_min[78][5] = (mid_1[639:632] < top_1[647:640]) ? 1 : 0;
assign detect_min[78][6] = (mid_1[639:632] < top_2[631:624]) ? 1 : 0;
assign detect_min[78][7] = (mid_1[639:632] < top_2[639:632]) ? 1 : 0;
assign detect_min[78][8] = (mid_1[639:632] < top_2[647:640]) ? 1 : 0;
assign detect_min[78][9] = (mid_1[639:632] < mid_0[631:624]) ? 1 : 0;
assign detect_min[78][10] = (mid_1[639:632] < mid_0[639:632]) ? 1 : 0;
assign detect_min[78][11] = (mid_1[639:632] < mid_0[647:640]) ? 1 : 0;
assign detect_min[78][12] = (mid_1[639:632] < mid_1[631:624]) ? 1 : 0;
assign detect_min[78][13] = (mid_1[639:632] < mid_1[647:640]) ? 1 : 0;
assign detect_min[78][14] = (mid_1[639:632] < mid_2[631:624]) ? 1 : 0;
assign detect_min[78][15] = (mid_1[639:632] < mid_2[639:632]) ? 1 : 0;
assign detect_min[78][16] = (mid_1[639:632] < mid_2[647:640]) ? 1 : 0;
assign detect_min[78][17] = (mid_1[639:632] < btm_0[631:624]) ? 1 : 0;
assign detect_min[78][18] = (mid_1[639:632] < btm_0[639:632]) ? 1 : 0;
assign detect_min[78][19] = (mid_1[639:632] < btm_0[647:640]) ? 1 : 0;
assign detect_min[78][20] = (mid_1[639:632] < btm_1[631:624]) ? 1 : 0;
assign detect_min[78][21] = (mid_1[639:632] < btm_1[639:632]) ? 1 : 0;
assign detect_min[78][22] = (mid_1[639:632] < btm_1[647:640]) ? 1 : 0;
assign detect_min[78][23] = (mid_1[639:632] < btm_2[631:624]) ? 1 : 0;
assign detect_min[78][24] = (mid_1[639:632] < btm_2[639:632]) ? 1 : 0;
assign detect_min[78][25] = (mid_1[639:632] < btm_2[647:640]) ? 1 : 0;

assign detect_min[79][0] = (mid_1[647:640] < top_0[639:632]) ? 1 : 0;
assign detect_min[79][1] = (mid_1[647:640] < top_0[647:640]) ? 1 : 0;
assign detect_min[79][2] = (mid_1[647:640] < top_0[655:648]) ? 1 : 0;
assign detect_min[79][3] = (mid_1[647:640] < top_1[639:632]) ? 1 : 0;
assign detect_min[79][4] = (mid_1[647:640] < top_1[647:640]) ? 1 : 0;
assign detect_min[79][5] = (mid_1[647:640] < top_1[655:648]) ? 1 : 0;
assign detect_min[79][6] = (mid_1[647:640] < top_2[639:632]) ? 1 : 0;
assign detect_min[79][7] = (mid_1[647:640] < top_2[647:640]) ? 1 : 0;
assign detect_min[79][8] = (mid_1[647:640] < top_2[655:648]) ? 1 : 0;
assign detect_min[79][9] = (mid_1[647:640] < mid_0[639:632]) ? 1 : 0;
assign detect_min[79][10] = (mid_1[647:640] < mid_0[647:640]) ? 1 : 0;
assign detect_min[79][11] = (mid_1[647:640] < mid_0[655:648]) ? 1 : 0;
assign detect_min[79][12] = (mid_1[647:640] < mid_1[639:632]) ? 1 : 0;
assign detect_min[79][13] = (mid_1[647:640] < mid_1[655:648]) ? 1 : 0;
assign detect_min[79][14] = (mid_1[647:640] < mid_2[639:632]) ? 1 : 0;
assign detect_min[79][15] = (mid_1[647:640] < mid_2[647:640]) ? 1 : 0;
assign detect_min[79][16] = (mid_1[647:640] < mid_2[655:648]) ? 1 : 0;
assign detect_min[79][17] = (mid_1[647:640] < btm_0[639:632]) ? 1 : 0;
assign detect_min[79][18] = (mid_1[647:640] < btm_0[647:640]) ? 1 : 0;
assign detect_min[79][19] = (mid_1[647:640] < btm_0[655:648]) ? 1 : 0;
assign detect_min[79][20] = (mid_1[647:640] < btm_1[639:632]) ? 1 : 0;
assign detect_min[79][21] = (mid_1[647:640] < btm_1[647:640]) ? 1 : 0;
assign detect_min[79][22] = (mid_1[647:640] < btm_1[655:648]) ? 1 : 0;
assign detect_min[79][23] = (mid_1[647:640] < btm_2[639:632]) ? 1 : 0;
assign detect_min[79][24] = (mid_1[647:640] < btm_2[647:640]) ? 1 : 0;
assign detect_min[79][25] = (mid_1[647:640] < btm_2[655:648]) ? 1 : 0;

assign detect_min[80][0] = (mid_1[655:648] < top_0[647:640]) ? 1 : 0;
assign detect_min[80][1] = (mid_1[655:648] < top_0[655:648]) ? 1 : 0;
assign detect_min[80][2] = (mid_1[655:648] < top_0[663:656]) ? 1 : 0;
assign detect_min[80][3] = (mid_1[655:648] < top_1[647:640]) ? 1 : 0;
assign detect_min[80][4] = (mid_1[655:648] < top_1[655:648]) ? 1 : 0;
assign detect_min[80][5] = (mid_1[655:648] < top_1[663:656]) ? 1 : 0;
assign detect_min[80][6] = (mid_1[655:648] < top_2[647:640]) ? 1 : 0;
assign detect_min[80][7] = (mid_1[655:648] < top_2[655:648]) ? 1 : 0;
assign detect_min[80][8] = (mid_1[655:648] < top_2[663:656]) ? 1 : 0;
assign detect_min[80][9] = (mid_1[655:648] < mid_0[647:640]) ? 1 : 0;
assign detect_min[80][10] = (mid_1[655:648] < mid_0[655:648]) ? 1 : 0;
assign detect_min[80][11] = (mid_1[655:648] < mid_0[663:656]) ? 1 : 0;
assign detect_min[80][12] = (mid_1[655:648] < mid_1[647:640]) ? 1 : 0;
assign detect_min[80][13] = (mid_1[655:648] < mid_1[663:656]) ? 1 : 0;
assign detect_min[80][14] = (mid_1[655:648] < mid_2[647:640]) ? 1 : 0;
assign detect_min[80][15] = (mid_1[655:648] < mid_2[655:648]) ? 1 : 0;
assign detect_min[80][16] = (mid_1[655:648] < mid_2[663:656]) ? 1 : 0;
assign detect_min[80][17] = (mid_1[655:648] < btm_0[647:640]) ? 1 : 0;
assign detect_min[80][18] = (mid_1[655:648] < btm_0[655:648]) ? 1 : 0;
assign detect_min[80][19] = (mid_1[655:648] < btm_0[663:656]) ? 1 : 0;
assign detect_min[80][20] = (mid_1[655:648] < btm_1[647:640]) ? 1 : 0;
assign detect_min[80][21] = (mid_1[655:648] < btm_1[655:648]) ? 1 : 0;
assign detect_min[80][22] = (mid_1[655:648] < btm_1[663:656]) ? 1 : 0;
assign detect_min[80][23] = (mid_1[655:648] < btm_2[647:640]) ? 1 : 0;
assign detect_min[80][24] = (mid_1[655:648] < btm_2[655:648]) ? 1 : 0;
assign detect_min[80][25] = (mid_1[655:648] < btm_2[663:656]) ? 1 : 0;

assign detect_min[81][0] = (mid_1[663:656] < top_0[655:648]) ? 1 : 0;
assign detect_min[81][1] = (mid_1[663:656] < top_0[663:656]) ? 1 : 0;
assign detect_min[81][2] = (mid_1[663:656] < top_0[671:664]) ? 1 : 0;
assign detect_min[81][3] = (mid_1[663:656] < top_1[655:648]) ? 1 : 0;
assign detect_min[81][4] = (mid_1[663:656] < top_1[663:656]) ? 1 : 0;
assign detect_min[81][5] = (mid_1[663:656] < top_1[671:664]) ? 1 : 0;
assign detect_min[81][6] = (mid_1[663:656] < top_2[655:648]) ? 1 : 0;
assign detect_min[81][7] = (mid_1[663:656] < top_2[663:656]) ? 1 : 0;
assign detect_min[81][8] = (mid_1[663:656] < top_2[671:664]) ? 1 : 0;
assign detect_min[81][9] = (mid_1[663:656] < mid_0[655:648]) ? 1 : 0;
assign detect_min[81][10] = (mid_1[663:656] < mid_0[663:656]) ? 1 : 0;
assign detect_min[81][11] = (mid_1[663:656] < mid_0[671:664]) ? 1 : 0;
assign detect_min[81][12] = (mid_1[663:656] < mid_1[655:648]) ? 1 : 0;
assign detect_min[81][13] = (mid_1[663:656] < mid_1[671:664]) ? 1 : 0;
assign detect_min[81][14] = (mid_1[663:656] < mid_2[655:648]) ? 1 : 0;
assign detect_min[81][15] = (mid_1[663:656] < mid_2[663:656]) ? 1 : 0;
assign detect_min[81][16] = (mid_1[663:656] < mid_2[671:664]) ? 1 : 0;
assign detect_min[81][17] = (mid_1[663:656] < btm_0[655:648]) ? 1 : 0;
assign detect_min[81][18] = (mid_1[663:656] < btm_0[663:656]) ? 1 : 0;
assign detect_min[81][19] = (mid_1[663:656] < btm_0[671:664]) ? 1 : 0;
assign detect_min[81][20] = (mid_1[663:656] < btm_1[655:648]) ? 1 : 0;
assign detect_min[81][21] = (mid_1[663:656] < btm_1[663:656]) ? 1 : 0;
assign detect_min[81][22] = (mid_1[663:656] < btm_1[671:664]) ? 1 : 0;
assign detect_min[81][23] = (mid_1[663:656] < btm_2[655:648]) ? 1 : 0;
assign detect_min[81][24] = (mid_1[663:656] < btm_2[663:656]) ? 1 : 0;
assign detect_min[81][25] = (mid_1[663:656] < btm_2[671:664]) ? 1 : 0;

assign detect_min[82][0] = (mid_1[671:664] < top_0[663:656]) ? 1 : 0;
assign detect_min[82][1] = (mid_1[671:664] < top_0[671:664]) ? 1 : 0;
assign detect_min[82][2] = (mid_1[671:664] < top_0[679:672]) ? 1 : 0;
assign detect_min[82][3] = (mid_1[671:664] < top_1[663:656]) ? 1 : 0;
assign detect_min[82][4] = (mid_1[671:664] < top_1[671:664]) ? 1 : 0;
assign detect_min[82][5] = (mid_1[671:664] < top_1[679:672]) ? 1 : 0;
assign detect_min[82][6] = (mid_1[671:664] < top_2[663:656]) ? 1 : 0;
assign detect_min[82][7] = (mid_1[671:664] < top_2[671:664]) ? 1 : 0;
assign detect_min[82][8] = (mid_1[671:664] < top_2[679:672]) ? 1 : 0;
assign detect_min[82][9] = (mid_1[671:664] < mid_0[663:656]) ? 1 : 0;
assign detect_min[82][10] = (mid_1[671:664] < mid_0[671:664]) ? 1 : 0;
assign detect_min[82][11] = (mid_1[671:664] < mid_0[679:672]) ? 1 : 0;
assign detect_min[82][12] = (mid_1[671:664] < mid_1[663:656]) ? 1 : 0;
assign detect_min[82][13] = (mid_1[671:664] < mid_1[679:672]) ? 1 : 0;
assign detect_min[82][14] = (mid_1[671:664] < mid_2[663:656]) ? 1 : 0;
assign detect_min[82][15] = (mid_1[671:664] < mid_2[671:664]) ? 1 : 0;
assign detect_min[82][16] = (mid_1[671:664] < mid_2[679:672]) ? 1 : 0;
assign detect_min[82][17] = (mid_1[671:664] < btm_0[663:656]) ? 1 : 0;
assign detect_min[82][18] = (mid_1[671:664] < btm_0[671:664]) ? 1 : 0;
assign detect_min[82][19] = (mid_1[671:664] < btm_0[679:672]) ? 1 : 0;
assign detect_min[82][20] = (mid_1[671:664] < btm_1[663:656]) ? 1 : 0;
assign detect_min[82][21] = (mid_1[671:664] < btm_1[671:664]) ? 1 : 0;
assign detect_min[82][22] = (mid_1[671:664] < btm_1[679:672]) ? 1 : 0;
assign detect_min[82][23] = (mid_1[671:664] < btm_2[663:656]) ? 1 : 0;
assign detect_min[82][24] = (mid_1[671:664] < btm_2[671:664]) ? 1 : 0;
assign detect_min[82][25] = (mid_1[671:664] < btm_2[679:672]) ? 1 : 0;

assign detect_min[83][0] = (mid_1[679:672] < top_0[671:664]) ? 1 : 0;
assign detect_min[83][1] = (mid_1[679:672] < top_0[679:672]) ? 1 : 0;
assign detect_min[83][2] = (mid_1[679:672] < top_0[687:680]) ? 1 : 0;
assign detect_min[83][3] = (mid_1[679:672] < top_1[671:664]) ? 1 : 0;
assign detect_min[83][4] = (mid_1[679:672] < top_1[679:672]) ? 1 : 0;
assign detect_min[83][5] = (mid_1[679:672] < top_1[687:680]) ? 1 : 0;
assign detect_min[83][6] = (mid_1[679:672] < top_2[671:664]) ? 1 : 0;
assign detect_min[83][7] = (mid_1[679:672] < top_2[679:672]) ? 1 : 0;
assign detect_min[83][8] = (mid_1[679:672] < top_2[687:680]) ? 1 : 0;
assign detect_min[83][9] = (mid_1[679:672] < mid_0[671:664]) ? 1 : 0;
assign detect_min[83][10] = (mid_1[679:672] < mid_0[679:672]) ? 1 : 0;
assign detect_min[83][11] = (mid_1[679:672] < mid_0[687:680]) ? 1 : 0;
assign detect_min[83][12] = (mid_1[679:672] < mid_1[671:664]) ? 1 : 0;
assign detect_min[83][13] = (mid_1[679:672] < mid_1[687:680]) ? 1 : 0;
assign detect_min[83][14] = (mid_1[679:672] < mid_2[671:664]) ? 1 : 0;
assign detect_min[83][15] = (mid_1[679:672] < mid_2[679:672]) ? 1 : 0;
assign detect_min[83][16] = (mid_1[679:672] < mid_2[687:680]) ? 1 : 0;
assign detect_min[83][17] = (mid_1[679:672] < btm_0[671:664]) ? 1 : 0;
assign detect_min[83][18] = (mid_1[679:672] < btm_0[679:672]) ? 1 : 0;
assign detect_min[83][19] = (mid_1[679:672] < btm_0[687:680]) ? 1 : 0;
assign detect_min[83][20] = (mid_1[679:672] < btm_1[671:664]) ? 1 : 0;
assign detect_min[83][21] = (mid_1[679:672] < btm_1[679:672]) ? 1 : 0;
assign detect_min[83][22] = (mid_1[679:672] < btm_1[687:680]) ? 1 : 0;
assign detect_min[83][23] = (mid_1[679:672] < btm_2[671:664]) ? 1 : 0;
assign detect_min[83][24] = (mid_1[679:672] < btm_2[679:672]) ? 1 : 0;
assign detect_min[83][25] = (mid_1[679:672] < btm_2[687:680]) ? 1 : 0;

assign detect_min[84][0] = (mid_1[687:680] < top_0[679:672]) ? 1 : 0;
assign detect_min[84][1] = (mid_1[687:680] < top_0[687:680]) ? 1 : 0;
assign detect_min[84][2] = (mid_1[687:680] < top_0[695:688]) ? 1 : 0;
assign detect_min[84][3] = (mid_1[687:680] < top_1[679:672]) ? 1 : 0;
assign detect_min[84][4] = (mid_1[687:680] < top_1[687:680]) ? 1 : 0;
assign detect_min[84][5] = (mid_1[687:680] < top_1[695:688]) ? 1 : 0;
assign detect_min[84][6] = (mid_1[687:680] < top_2[679:672]) ? 1 : 0;
assign detect_min[84][7] = (mid_1[687:680] < top_2[687:680]) ? 1 : 0;
assign detect_min[84][8] = (mid_1[687:680] < top_2[695:688]) ? 1 : 0;
assign detect_min[84][9] = (mid_1[687:680] < mid_0[679:672]) ? 1 : 0;
assign detect_min[84][10] = (mid_1[687:680] < mid_0[687:680]) ? 1 : 0;
assign detect_min[84][11] = (mid_1[687:680] < mid_0[695:688]) ? 1 : 0;
assign detect_min[84][12] = (mid_1[687:680] < mid_1[679:672]) ? 1 : 0;
assign detect_min[84][13] = (mid_1[687:680] < mid_1[695:688]) ? 1 : 0;
assign detect_min[84][14] = (mid_1[687:680] < mid_2[679:672]) ? 1 : 0;
assign detect_min[84][15] = (mid_1[687:680] < mid_2[687:680]) ? 1 : 0;
assign detect_min[84][16] = (mid_1[687:680] < mid_2[695:688]) ? 1 : 0;
assign detect_min[84][17] = (mid_1[687:680] < btm_0[679:672]) ? 1 : 0;
assign detect_min[84][18] = (mid_1[687:680] < btm_0[687:680]) ? 1 : 0;
assign detect_min[84][19] = (mid_1[687:680] < btm_0[695:688]) ? 1 : 0;
assign detect_min[84][20] = (mid_1[687:680] < btm_1[679:672]) ? 1 : 0;
assign detect_min[84][21] = (mid_1[687:680] < btm_1[687:680]) ? 1 : 0;
assign detect_min[84][22] = (mid_1[687:680] < btm_1[695:688]) ? 1 : 0;
assign detect_min[84][23] = (mid_1[687:680] < btm_2[679:672]) ? 1 : 0;
assign detect_min[84][24] = (mid_1[687:680] < btm_2[687:680]) ? 1 : 0;
assign detect_min[84][25] = (mid_1[687:680] < btm_2[695:688]) ? 1 : 0;

assign detect_min[85][0] = (mid_1[695:688] < top_0[687:680]) ? 1 : 0;
assign detect_min[85][1] = (mid_1[695:688] < top_0[695:688]) ? 1 : 0;
assign detect_min[85][2] = (mid_1[695:688] < top_0[703:696]) ? 1 : 0;
assign detect_min[85][3] = (mid_1[695:688] < top_1[687:680]) ? 1 : 0;
assign detect_min[85][4] = (mid_1[695:688] < top_1[695:688]) ? 1 : 0;
assign detect_min[85][5] = (mid_1[695:688] < top_1[703:696]) ? 1 : 0;
assign detect_min[85][6] = (mid_1[695:688] < top_2[687:680]) ? 1 : 0;
assign detect_min[85][7] = (mid_1[695:688] < top_2[695:688]) ? 1 : 0;
assign detect_min[85][8] = (mid_1[695:688] < top_2[703:696]) ? 1 : 0;
assign detect_min[85][9] = (mid_1[695:688] < mid_0[687:680]) ? 1 : 0;
assign detect_min[85][10] = (mid_1[695:688] < mid_0[695:688]) ? 1 : 0;
assign detect_min[85][11] = (mid_1[695:688] < mid_0[703:696]) ? 1 : 0;
assign detect_min[85][12] = (mid_1[695:688] < mid_1[687:680]) ? 1 : 0;
assign detect_min[85][13] = (mid_1[695:688] < mid_1[703:696]) ? 1 : 0;
assign detect_min[85][14] = (mid_1[695:688] < mid_2[687:680]) ? 1 : 0;
assign detect_min[85][15] = (mid_1[695:688] < mid_2[695:688]) ? 1 : 0;
assign detect_min[85][16] = (mid_1[695:688] < mid_2[703:696]) ? 1 : 0;
assign detect_min[85][17] = (mid_1[695:688] < btm_0[687:680]) ? 1 : 0;
assign detect_min[85][18] = (mid_1[695:688] < btm_0[695:688]) ? 1 : 0;
assign detect_min[85][19] = (mid_1[695:688] < btm_0[703:696]) ? 1 : 0;
assign detect_min[85][20] = (mid_1[695:688] < btm_1[687:680]) ? 1 : 0;
assign detect_min[85][21] = (mid_1[695:688] < btm_1[695:688]) ? 1 : 0;
assign detect_min[85][22] = (mid_1[695:688] < btm_1[703:696]) ? 1 : 0;
assign detect_min[85][23] = (mid_1[695:688] < btm_2[687:680]) ? 1 : 0;
assign detect_min[85][24] = (mid_1[695:688] < btm_2[695:688]) ? 1 : 0;
assign detect_min[85][25] = (mid_1[695:688] < btm_2[703:696]) ? 1 : 0;

assign detect_min[86][0] = (mid_1[703:696] < top_0[695:688]) ? 1 : 0;
assign detect_min[86][1] = (mid_1[703:696] < top_0[703:696]) ? 1 : 0;
assign detect_min[86][2] = (mid_1[703:696] < top_0[711:704]) ? 1 : 0;
assign detect_min[86][3] = (mid_1[703:696] < top_1[695:688]) ? 1 : 0;
assign detect_min[86][4] = (mid_1[703:696] < top_1[703:696]) ? 1 : 0;
assign detect_min[86][5] = (mid_1[703:696] < top_1[711:704]) ? 1 : 0;
assign detect_min[86][6] = (mid_1[703:696] < top_2[695:688]) ? 1 : 0;
assign detect_min[86][7] = (mid_1[703:696] < top_2[703:696]) ? 1 : 0;
assign detect_min[86][8] = (mid_1[703:696] < top_2[711:704]) ? 1 : 0;
assign detect_min[86][9] = (mid_1[703:696] < mid_0[695:688]) ? 1 : 0;
assign detect_min[86][10] = (mid_1[703:696] < mid_0[703:696]) ? 1 : 0;
assign detect_min[86][11] = (mid_1[703:696] < mid_0[711:704]) ? 1 : 0;
assign detect_min[86][12] = (mid_1[703:696] < mid_1[695:688]) ? 1 : 0;
assign detect_min[86][13] = (mid_1[703:696] < mid_1[711:704]) ? 1 : 0;
assign detect_min[86][14] = (mid_1[703:696] < mid_2[695:688]) ? 1 : 0;
assign detect_min[86][15] = (mid_1[703:696] < mid_2[703:696]) ? 1 : 0;
assign detect_min[86][16] = (mid_1[703:696] < mid_2[711:704]) ? 1 : 0;
assign detect_min[86][17] = (mid_1[703:696] < btm_0[695:688]) ? 1 : 0;
assign detect_min[86][18] = (mid_1[703:696] < btm_0[703:696]) ? 1 : 0;
assign detect_min[86][19] = (mid_1[703:696] < btm_0[711:704]) ? 1 : 0;
assign detect_min[86][20] = (mid_1[703:696] < btm_1[695:688]) ? 1 : 0;
assign detect_min[86][21] = (mid_1[703:696] < btm_1[703:696]) ? 1 : 0;
assign detect_min[86][22] = (mid_1[703:696] < btm_1[711:704]) ? 1 : 0;
assign detect_min[86][23] = (mid_1[703:696] < btm_2[695:688]) ? 1 : 0;
assign detect_min[86][24] = (mid_1[703:696] < btm_2[703:696]) ? 1 : 0;
assign detect_min[86][25] = (mid_1[703:696] < btm_2[711:704]) ? 1 : 0;

assign detect_min[87][0] = (mid_1[711:704] < top_0[703:696]) ? 1 : 0;
assign detect_min[87][1] = (mid_1[711:704] < top_0[711:704]) ? 1 : 0;
assign detect_min[87][2] = (mid_1[711:704] < top_0[719:712]) ? 1 : 0;
assign detect_min[87][3] = (mid_1[711:704] < top_1[703:696]) ? 1 : 0;
assign detect_min[87][4] = (mid_1[711:704] < top_1[711:704]) ? 1 : 0;
assign detect_min[87][5] = (mid_1[711:704] < top_1[719:712]) ? 1 : 0;
assign detect_min[87][6] = (mid_1[711:704] < top_2[703:696]) ? 1 : 0;
assign detect_min[87][7] = (mid_1[711:704] < top_2[711:704]) ? 1 : 0;
assign detect_min[87][8] = (mid_1[711:704] < top_2[719:712]) ? 1 : 0;
assign detect_min[87][9] = (mid_1[711:704] < mid_0[703:696]) ? 1 : 0;
assign detect_min[87][10] = (mid_1[711:704] < mid_0[711:704]) ? 1 : 0;
assign detect_min[87][11] = (mid_1[711:704] < mid_0[719:712]) ? 1 : 0;
assign detect_min[87][12] = (mid_1[711:704] < mid_1[703:696]) ? 1 : 0;
assign detect_min[87][13] = (mid_1[711:704] < mid_1[719:712]) ? 1 : 0;
assign detect_min[87][14] = (mid_1[711:704] < mid_2[703:696]) ? 1 : 0;
assign detect_min[87][15] = (mid_1[711:704] < mid_2[711:704]) ? 1 : 0;
assign detect_min[87][16] = (mid_1[711:704] < mid_2[719:712]) ? 1 : 0;
assign detect_min[87][17] = (mid_1[711:704] < btm_0[703:696]) ? 1 : 0;
assign detect_min[87][18] = (mid_1[711:704] < btm_0[711:704]) ? 1 : 0;
assign detect_min[87][19] = (mid_1[711:704] < btm_0[719:712]) ? 1 : 0;
assign detect_min[87][20] = (mid_1[711:704] < btm_1[703:696]) ? 1 : 0;
assign detect_min[87][21] = (mid_1[711:704] < btm_1[711:704]) ? 1 : 0;
assign detect_min[87][22] = (mid_1[711:704] < btm_1[719:712]) ? 1 : 0;
assign detect_min[87][23] = (mid_1[711:704] < btm_2[703:696]) ? 1 : 0;
assign detect_min[87][24] = (mid_1[711:704] < btm_2[711:704]) ? 1 : 0;
assign detect_min[87][25] = (mid_1[711:704] < btm_2[719:712]) ? 1 : 0;

assign detect_min[88][0] = (mid_1[719:712] < top_0[711:704]) ? 1 : 0;
assign detect_min[88][1] = (mid_1[719:712] < top_0[719:712]) ? 1 : 0;
assign detect_min[88][2] = (mid_1[719:712] < top_0[727:720]) ? 1 : 0;
assign detect_min[88][3] = (mid_1[719:712] < top_1[711:704]) ? 1 : 0;
assign detect_min[88][4] = (mid_1[719:712] < top_1[719:712]) ? 1 : 0;
assign detect_min[88][5] = (mid_1[719:712] < top_1[727:720]) ? 1 : 0;
assign detect_min[88][6] = (mid_1[719:712] < top_2[711:704]) ? 1 : 0;
assign detect_min[88][7] = (mid_1[719:712] < top_2[719:712]) ? 1 : 0;
assign detect_min[88][8] = (mid_1[719:712] < top_2[727:720]) ? 1 : 0;
assign detect_min[88][9] = (mid_1[719:712] < mid_0[711:704]) ? 1 : 0;
assign detect_min[88][10] = (mid_1[719:712] < mid_0[719:712]) ? 1 : 0;
assign detect_min[88][11] = (mid_1[719:712] < mid_0[727:720]) ? 1 : 0;
assign detect_min[88][12] = (mid_1[719:712] < mid_1[711:704]) ? 1 : 0;
assign detect_min[88][13] = (mid_1[719:712] < mid_1[727:720]) ? 1 : 0;
assign detect_min[88][14] = (mid_1[719:712] < mid_2[711:704]) ? 1 : 0;
assign detect_min[88][15] = (mid_1[719:712] < mid_2[719:712]) ? 1 : 0;
assign detect_min[88][16] = (mid_1[719:712] < mid_2[727:720]) ? 1 : 0;
assign detect_min[88][17] = (mid_1[719:712] < btm_0[711:704]) ? 1 : 0;
assign detect_min[88][18] = (mid_1[719:712] < btm_0[719:712]) ? 1 : 0;
assign detect_min[88][19] = (mid_1[719:712] < btm_0[727:720]) ? 1 : 0;
assign detect_min[88][20] = (mid_1[719:712] < btm_1[711:704]) ? 1 : 0;
assign detect_min[88][21] = (mid_1[719:712] < btm_1[719:712]) ? 1 : 0;
assign detect_min[88][22] = (mid_1[719:712] < btm_1[727:720]) ? 1 : 0;
assign detect_min[88][23] = (mid_1[719:712] < btm_2[711:704]) ? 1 : 0;
assign detect_min[88][24] = (mid_1[719:712] < btm_2[719:712]) ? 1 : 0;
assign detect_min[88][25] = (mid_1[719:712] < btm_2[727:720]) ? 1 : 0;

assign detect_min[89][0] = (mid_1[727:720] < top_0[719:712]) ? 1 : 0;
assign detect_min[89][1] = (mid_1[727:720] < top_0[727:720]) ? 1 : 0;
assign detect_min[89][2] = (mid_1[727:720] < top_0[735:728]) ? 1 : 0;
assign detect_min[89][3] = (mid_1[727:720] < top_1[719:712]) ? 1 : 0;
assign detect_min[89][4] = (mid_1[727:720] < top_1[727:720]) ? 1 : 0;
assign detect_min[89][5] = (mid_1[727:720] < top_1[735:728]) ? 1 : 0;
assign detect_min[89][6] = (mid_1[727:720] < top_2[719:712]) ? 1 : 0;
assign detect_min[89][7] = (mid_1[727:720] < top_2[727:720]) ? 1 : 0;
assign detect_min[89][8] = (mid_1[727:720] < top_2[735:728]) ? 1 : 0;
assign detect_min[89][9] = (mid_1[727:720] < mid_0[719:712]) ? 1 : 0;
assign detect_min[89][10] = (mid_1[727:720] < mid_0[727:720]) ? 1 : 0;
assign detect_min[89][11] = (mid_1[727:720] < mid_0[735:728]) ? 1 : 0;
assign detect_min[89][12] = (mid_1[727:720] < mid_1[719:712]) ? 1 : 0;
assign detect_min[89][13] = (mid_1[727:720] < mid_1[735:728]) ? 1 : 0;
assign detect_min[89][14] = (mid_1[727:720] < mid_2[719:712]) ? 1 : 0;
assign detect_min[89][15] = (mid_1[727:720] < mid_2[727:720]) ? 1 : 0;
assign detect_min[89][16] = (mid_1[727:720] < mid_2[735:728]) ? 1 : 0;
assign detect_min[89][17] = (mid_1[727:720] < btm_0[719:712]) ? 1 : 0;
assign detect_min[89][18] = (mid_1[727:720] < btm_0[727:720]) ? 1 : 0;
assign detect_min[89][19] = (mid_1[727:720] < btm_0[735:728]) ? 1 : 0;
assign detect_min[89][20] = (mid_1[727:720] < btm_1[719:712]) ? 1 : 0;
assign detect_min[89][21] = (mid_1[727:720] < btm_1[727:720]) ? 1 : 0;
assign detect_min[89][22] = (mid_1[727:720] < btm_1[735:728]) ? 1 : 0;
assign detect_min[89][23] = (mid_1[727:720] < btm_2[719:712]) ? 1 : 0;
assign detect_min[89][24] = (mid_1[727:720] < btm_2[727:720]) ? 1 : 0;
assign detect_min[89][25] = (mid_1[727:720] < btm_2[735:728]) ? 1 : 0;

assign detect_min[90][0] = (mid_1[735:728] < top_0[727:720]) ? 1 : 0;
assign detect_min[90][1] = (mid_1[735:728] < top_0[735:728]) ? 1 : 0;
assign detect_min[90][2] = (mid_1[735:728] < top_0[743:736]) ? 1 : 0;
assign detect_min[90][3] = (mid_1[735:728] < top_1[727:720]) ? 1 : 0;
assign detect_min[90][4] = (mid_1[735:728] < top_1[735:728]) ? 1 : 0;
assign detect_min[90][5] = (mid_1[735:728] < top_1[743:736]) ? 1 : 0;
assign detect_min[90][6] = (mid_1[735:728] < top_2[727:720]) ? 1 : 0;
assign detect_min[90][7] = (mid_1[735:728] < top_2[735:728]) ? 1 : 0;
assign detect_min[90][8] = (mid_1[735:728] < top_2[743:736]) ? 1 : 0;
assign detect_min[90][9] = (mid_1[735:728] < mid_0[727:720]) ? 1 : 0;
assign detect_min[90][10] = (mid_1[735:728] < mid_0[735:728]) ? 1 : 0;
assign detect_min[90][11] = (mid_1[735:728] < mid_0[743:736]) ? 1 : 0;
assign detect_min[90][12] = (mid_1[735:728] < mid_1[727:720]) ? 1 : 0;
assign detect_min[90][13] = (mid_1[735:728] < mid_1[743:736]) ? 1 : 0;
assign detect_min[90][14] = (mid_1[735:728] < mid_2[727:720]) ? 1 : 0;
assign detect_min[90][15] = (mid_1[735:728] < mid_2[735:728]) ? 1 : 0;
assign detect_min[90][16] = (mid_1[735:728] < mid_2[743:736]) ? 1 : 0;
assign detect_min[90][17] = (mid_1[735:728] < btm_0[727:720]) ? 1 : 0;
assign detect_min[90][18] = (mid_1[735:728] < btm_0[735:728]) ? 1 : 0;
assign detect_min[90][19] = (mid_1[735:728] < btm_0[743:736]) ? 1 : 0;
assign detect_min[90][20] = (mid_1[735:728] < btm_1[727:720]) ? 1 : 0;
assign detect_min[90][21] = (mid_1[735:728] < btm_1[735:728]) ? 1 : 0;
assign detect_min[90][22] = (mid_1[735:728] < btm_1[743:736]) ? 1 : 0;
assign detect_min[90][23] = (mid_1[735:728] < btm_2[727:720]) ? 1 : 0;
assign detect_min[90][24] = (mid_1[735:728] < btm_2[735:728]) ? 1 : 0;
assign detect_min[90][25] = (mid_1[735:728] < btm_2[743:736]) ? 1 : 0;

assign detect_min[91][0] = (mid_1[743:736] < top_0[735:728]) ? 1 : 0;
assign detect_min[91][1] = (mid_1[743:736] < top_0[743:736]) ? 1 : 0;
assign detect_min[91][2] = (mid_1[743:736] < top_0[751:744]) ? 1 : 0;
assign detect_min[91][3] = (mid_1[743:736] < top_1[735:728]) ? 1 : 0;
assign detect_min[91][4] = (mid_1[743:736] < top_1[743:736]) ? 1 : 0;
assign detect_min[91][5] = (mid_1[743:736] < top_1[751:744]) ? 1 : 0;
assign detect_min[91][6] = (mid_1[743:736] < top_2[735:728]) ? 1 : 0;
assign detect_min[91][7] = (mid_1[743:736] < top_2[743:736]) ? 1 : 0;
assign detect_min[91][8] = (mid_1[743:736] < top_2[751:744]) ? 1 : 0;
assign detect_min[91][9] = (mid_1[743:736] < mid_0[735:728]) ? 1 : 0;
assign detect_min[91][10] = (mid_1[743:736] < mid_0[743:736]) ? 1 : 0;
assign detect_min[91][11] = (mid_1[743:736] < mid_0[751:744]) ? 1 : 0;
assign detect_min[91][12] = (mid_1[743:736] < mid_1[735:728]) ? 1 : 0;
assign detect_min[91][13] = (mid_1[743:736] < mid_1[751:744]) ? 1 : 0;
assign detect_min[91][14] = (mid_1[743:736] < mid_2[735:728]) ? 1 : 0;
assign detect_min[91][15] = (mid_1[743:736] < mid_2[743:736]) ? 1 : 0;
assign detect_min[91][16] = (mid_1[743:736] < mid_2[751:744]) ? 1 : 0;
assign detect_min[91][17] = (mid_1[743:736] < btm_0[735:728]) ? 1 : 0;
assign detect_min[91][18] = (mid_1[743:736] < btm_0[743:736]) ? 1 : 0;
assign detect_min[91][19] = (mid_1[743:736] < btm_0[751:744]) ? 1 : 0;
assign detect_min[91][20] = (mid_1[743:736] < btm_1[735:728]) ? 1 : 0;
assign detect_min[91][21] = (mid_1[743:736] < btm_1[743:736]) ? 1 : 0;
assign detect_min[91][22] = (mid_1[743:736] < btm_1[751:744]) ? 1 : 0;
assign detect_min[91][23] = (mid_1[743:736] < btm_2[735:728]) ? 1 : 0;
assign detect_min[91][24] = (mid_1[743:736] < btm_2[743:736]) ? 1 : 0;
assign detect_min[91][25] = (mid_1[743:736] < btm_2[751:744]) ? 1 : 0;

assign detect_min[92][0] = (mid_1[751:744] < top_0[743:736]) ? 1 : 0;
assign detect_min[92][1] = (mid_1[751:744] < top_0[751:744]) ? 1 : 0;
assign detect_min[92][2] = (mid_1[751:744] < top_0[759:752]) ? 1 : 0;
assign detect_min[92][3] = (mid_1[751:744] < top_1[743:736]) ? 1 : 0;
assign detect_min[92][4] = (mid_1[751:744] < top_1[751:744]) ? 1 : 0;
assign detect_min[92][5] = (mid_1[751:744] < top_1[759:752]) ? 1 : 0;
assign detect_min[92][6] = (mid_1[751:744] < top_2[743:736]) ? 1 : 0;
assign detect_min[92][7] = (mid_1[751:744] < top_2[751:744]) ? 1 : 0;
assign detect_min[92][8] = (mid_1[751:744] < top_2[759:752]) ? 1 : 0;
assign detect_min[92][9] = (mid_1[751:744] < mid_0[743:736]) ? 1 : 0;
assign detect_min[92][10] = (mid_1[751:744] < mid_0[751:744]) ? 1 : 0;
assign detect_min[92][11] = (mid_1[751:744] < mid_0[759:752]) ? 1 : 0;
assign detect_min[92][12] = (mid_1[751:744] < mid_1[743:736]) ? 1 : 0;
assign detect_min[92][13] = (mid_1[751:744] < mid_1[759:752]) ? 1 : 0;
assign detect_min[92][14] = (mid_1[751:744] < mid_2[743:736]) ? 1 : 0;
assign detect_min[92][15] = (mid_1[751:744] < mid_2[751:744]) ? 1 : 0;
assign detect_min[92][16] = (mid_1[751:744] < mid_2[759:752]) ? 1 : 0;
assign detect_min[92][17] = (mid_1[751:744] < btm_0[743:736]) ? 1 : 0;
assign detect_min[92][18] = (mid_1[751:744] < btm_0[751:744]) ? 1 : 0;
assign detect_min[92][19] = (mid_1[751:744] < btm_0[759:752]) ? 1 : 0;
assign detect_min[92][20] = (mid_1[751:744] < btm_1[743:736]) ? 1 : 0;
assign detect_min[92][21] = (mid_1[751:744] < btm_1[751:744]) ? 1 : 0;
assign detect_min[92][22] = (mid_1[751:744] < btm_1[759:752]) ? 1 : 0;
assign detect_min[92][23] = (mid_1[751:744] < btm_2[743:736]) ? 1 : 0;
assign detect_min[92][24] = (mid_1[751:744] < btm_2[751:744]) ? 1 : 0;
assign detect_min[92][25] = (mid_1[751:744] < btm_2[759:752]) ? 1 : 0;

assign detect_min[93][0] = (mid_1[759:752] < top_0[751:744]) ? 1 : 0;
assign detect_min[93][1] = (mid_1[759:752] < top_0[759:752]) ? 1 : 0;
assign detect_min[93][2] = (mid_1[759:752] < top_0[767:760]) ? 1 : 0;
assign detect_min[93][3] = (mid_1[759:752] < top_1[751:744]) ? 1 : 0;
assign detect_min[93][4] = (mid_1[759:752] < top_1[759:752]) ? 1 : 0;
assign detect_min[93][5] = (mid_1[759:752] < top_1[767:760]) ? 1 : 0;
assign detect_min[93][6] = (mid_1[759:752] < top_2[751:744]) ? 1 : 0;
assign detect_min[93][7] = (mid_1[759:752] < top_2[759:752]) ? 1 : 0;
assign detect_min[93][8] = (mid_1[759:752] < top_2[767:760]) ? 1 : 0;
assign detect_min[93][9] = (mid_1[759:752] < mid_0[751:744]) ? 1 : 0;
assign detect_min[93][10] = (mid_1[759:752] < mid_0[759:752]) ? 1 : 0;
assign detect_min[93][11] = (mid_1[759:752] < mid_0[767:760]) ? 1 : 0;
assign detect_min[93][12] = (mid_1[759:752] < mid_1[751:744]) ? 1 : 0;
assign detect_min[93][13] = (mid_1[759:752] < mid_1[767:760]) ? 1 : 0;
assign detect_min[93][14] = (mid_1[759:752] < mid_2[751:744]) ? 1 : 0;
assign detect_min[93][15] = (mid_1[759:752] < mid_2[759:752]) ? 1 : 0;
assign detect_min[93][16] = (mid_1[759:752] < mid_2[767:760]) ? 1 : 0;
assign detect_min[93][17] = (mid_1[759:752] < btm_0[751:744]) ? 1 : 0;
assign detect_min[93][18] = (mid_1[759:752] < btm_0[759:752]) ? 1 : 0;
assign detect_min[93][19] = (mid_1[759:752] < btm_0[767:760]) ? 1 : 0;
assign detect_min[93][20] = (mid_1[759:752] < btm_1[751:744]) ? 1 : 0;
assign detect_min[93][21] = (mid_1[759:752] < btm_1[759:752]) ? 1 : 0;
assign detect_min[93][22] = (mid_1[759:752] < btm_1[767:760]) ? 1 : 0;
assign detect_min[93][23] = (mid_1[759:752] < btm_2[751:744]) ? 1 : 0;
assign detect_min[93][24] = (mid_1[759:752] < btm_2[759:752]) ? 1 : 0;
assign detect_min[93][25] = (mid_1[759:752] < btm_2[767:760]) ? 1 : 0;

assign detect_min[94][0] = (mid_1[767:760] < top_0[759:752]) ? 1 : 0;
assign detect_min[94][1] = (mid_1[767:760] < top_0[767:760]) ? 1 : 0;
assign detect_min[94][2] = (mid_1[767:760] < top_0[775:768]) ? 1 : 0;
assign detect_min[94][3] = (mid_1[767:760] < top_1[759:752]) ? 1 : 0;
assign detect_min[94][4] = (mid_1[767:760] < top_1[767:760]) ? 1 : 0;
assign detect_min[94][5] = (mid_1[767:760] < top_1[775:768]) ? 1 : 0;
assign detect_min[94][6] = (mid_1[767:760] < top_2[759:752]) ? 1 : 0;
assign detect_min[94][7] = (mid_1[767:760] < top_2[767:760]) ? 1 : 0;
assign detect_min[94][8] = (mid_1[767:760] < top_2[775:768]) ? 1 : 0;
assign detect_min[94][9] = (mid_1[767:760] < mid_0[759:752]) ? 1 : 0;
assign detect_min[94][10] = (mid_1[767:760] < mid_0[767:760]) ? 1 : 0;
assign detect_min[94][11] = (mid_1[767:760] < mid_0[775:768]) ? 1 : 0;
assign detect_min[94][12] = (mid_1[767:760] < mid_1[759:752]) ? 1 : 0;
assign detect_min[94][13] = (mid_1[767:760] < mid_1[775:768]) ? 1 : 0;
assign detect_min[94][14] = (mid_1[767:760] < mid_2[759:752]) ? 1 : 0;
assign detect_min[94][15] = (mid_1[767:760] < mid_2[767:760]) ? 1 : 0;
assign detect_min[94][16] = (mid_1[767:760] < mid_2[775:768]) ? 1 : 0;
assign detect_min[94][17] = (mid_1[767:760] < btm_0[759:752]) ? 1 : 0;
assign detect_min[94][18] = (mid_1[767:760] < btm_0[767:760]) ? 1 : 0;
assign detect_min[94][19] = (mid_1[767:760] < btm_0[775:768]) ? 1 : 0;
assign detect_min[94][20] = (mid_1[767:760] < btm_1[759:752]) ? 1 : 0;
assign detect_min[94][21] = (mid_1[767:760] < btm_1[767:760]) ? 1 : 0;
assign detect_min[94][22] = (mid_1[767:760] < btm_1[775:768]) ? 1 : 0;
assign detect_min[94][23] = (mid_1[767:760] < btm_2[759:752]) ? 1 : 0;
assign detect_min[94][24] = (mid_1[767:760] < btm_2[767:760]) ? 1 : 0;
assign detect_min[94][25] = (mid_1[767:760] < btm_2[775:768]) ? 1 : 0;

assign detect_min[95][0] = (mid_1[775:768] < top_0[767:760]) ? 1 : 0;
assign detect_min[95][1] = (mid_1[775:768] < top_0[775:768]) ? 1 : 0;
assign detect_min[95][2] = (mid_1[775:768] < top_0[783:776]) ? 1 : 0;
assign detect_min[95][3] = (mid_1[775:768] < top_1[767:760]) ? 1 : 0;
assign detect_min[95][4] = (mid_1[775:768] < top_1[775:768]) ? 1 : 0;
assign detect_min[95][5] = (mid_1[775:768] < top_1[783:776]) ? 1 : 0;
assign detect_min[95][6] = (mid_1[775:768] < top_2[767:760]) ? 1 : 0;
assign detect_min[95][7] = (mid_1[775:768] < top_2[775:768]) ? 1 : 0;
assign detect_min[95][8] = (mid_1[775:768] < top_2[783:776]) ? 1 : 0;
assign detect_min[95][9] = (mid_1[775:768] < mid_0[767:760]) ? 1 : 0;
assign detect_min[95][10] = (mid_1[775:768] < mid_0[775:768]) ? 1 : 0;
assign detect_min[95][11] = (mid_1[775:768] < mid_0[783:776]) ? 1 : 0;
assign detect_min[95][12] = (mid_1[775:768] < mid_1[767:760]) ? 1 : 0;
assign detect_min[95][13] = (mid_1[775:768] < mid_1[783:776]) ? 1 : 0;
assign detect_min[95][14] = (mid_1[775:768] < mid_2[767:760]) ? 1 : 0;
assign detect_min[95][15] = (mid_1[775:768] < mid_2[775:768]) ? 1 : 0;
assign detect_min[95][16] = (mid_1[775:768] < mid_2[783:776]) ? 1 : 0;
assign detect_min[95][17] = (mid_1[775:768] < btm_0[767:760]) ? 1 : 0;
assign detect_min[95][18] = (mid_1[775:768] < btm_0[775:768]) ? 1 : 0;
assign detect_min[95][19] = (mid_1[775:768] < btm_0[783:776]) ? 1 : 0;
assign detect_min[95][20] = (mid_1[775:768] < btm_1[767:760]) ? 1 : 0;
assign detect_min[95][21] = (mid_1[775:768] < btm_1[775:768]) ? 1 : 0;
assign detect_min[95][22] = (mid_1[775:768] < btm_1[783:776]) ? 1 : 0;
assign detect_min[95][23] = (mid_1[775:768] < btm_2[767:760]) ? 1 : 0;
assign detect_min[95][24] = (mid_1[775:768] < btm_2[775:768]) ? 1 : 0;
assign detect_min[95][25] = (mid_1[775:768] < btm_2[783:776]) ? 1 : 0;

assign detect_min[96][0] = (mid_1[783:776] < top_0[775:768]) ? 1 : 0;
assign detect_min[96][1] = (mid_1[783:776] < top_0[783:776]) ? 1 : 0;
assign detect_min[96][2] = (mid_1[783:776] < top_0[791:784]) ? 1 : 0;
assign detect_min[96][3] = (mid_1[783:776] < top_1[775:768]) ? 1 : 0;
assign detect_min[96][4] = (mid_1[783:776] < top_1[783:776]) ? 1 : 0;
assign detect_min[96][5] = (mid_1[783:776] < top_1[791:784]) ? 1 : 0;
assign detect_min[96][6] = (mid_1[783:776] < top_2[775:768]) ? 1 : 0;
assign detect_min[96][7] = (mid_1[783:776] < top_2[783:776]) ? 1 : 0;
assign detect_min[96][8] = (mid_1[783:776] < top_2[791:784]) ? 1 : 0;
assign detect_min[96][9] = (mid_1[783:776] < mid_0[775:768]) ? 1 : 0;
assign detect_min[96][10] = (mid_1[783:776] < mid_0[783:776]) ? 1 : 0;
assign detect_min[96][11] = (mid_1[783:776] < mid_0[791:784]) ? 1 : 0;
assign detect_min[96][12] = (mid_1[783:776] < mid_1[775:768]) ? 1 : 0;
assign detect_min[96][13] = (mid_1[783:776] < mid_1[791:784]) ? 1 : 0;
assign detect_min[96][14] = (mid_1[783:776] < mid_2[775:768]) ? 1 : 0;
assign detect_min[96][15] = (mid_1[783:776] < mid_2[783:776]) ? 1 : 0;
assign detect_min[96][16] = (mid_1[783:776] < mid_2[791:784]) ? 1 : 0;
assign detect_min[96][17] = (mid_1[783:776] < btm_0[775:768]) ? 1 : 0;
assign detect_min[96][18] = (mid_1[783:776] < btm_0[783:776]) ? 1 : 0;
assign detect_min[96][19] = (mid_1[783:776] < btm_0[791:784]) ? 1 : 0;
assign detect_min[96][20] = (mid_1[783:776] < btm_1[775:768]) ? 1 : 0;
assign detect_min[96][21] = (mid_1[783:776] < btm_1[783:776]) ? 1 : 0;
assign detect_min[96][22] = (mid_1[783:776] < btm_1[791:784]) ? 1 : 0;
assign detect_min[96][23] = (mid_1[783:776] < btm_2[775:768]) ? 1 : 0;
assign detect_min[96][24] = (mid_1[783:776] < btm_2[783:776]) ? 1 : 0;
assign detect_min[96][25] = (mid_1[783:776] < btm_2[791:784]) ? 1 : 0;

assign detect_min[97][0] = (mid_1[791:784] < top_0[783:776]) ? 1 : 0;
assign detect_min[97][1] = (mid_1[791:784] < top_0[791:784]) ? 1 : 0;
assign detect_min[97][2] = (mid_1[791:784] < top_0[799:792]) ? 1 : 0;
assign detect_min[97][3] = (mid_1[791:784] < top_1[783:776]) ? 1 : 0;
assign detect_min[97][4] = (mid_1[791:784] < top_1[791:784]) ? 1 : 0;
assign detect_min[97][5] = (mid_1[791:784] < top_1[799:792]) ? 1 : 0;
assign detect_min[97][6] = (mid_1[791:784] < top_2[783:776]) ? 1 : 0;
assign detect_min[97][7] = (mid_1[791:784] < top_2[791:784]) ? 1 : 0;
assign detect_min[97][8] = (mid_1[791:784] < top_2[799:792]) ? 1 : 0;
assign detect_min[97][9] = (mid_1[791:784] < mid_0[783:776]) ? 1 : 0;
assign detect_min[97][10] = (mid_1[791:784] < mid_0[791:784]) ? 1 : 0;
assign detect_min[97][11] = (mid_1[791:784] < mid_0[799:792]) ? 1 : 0;
assign detect_min[97][12] = (mid_1[791:784] < mid_1[783:776]) ? 1 : 0;
assign detect_min[97][13] = (mid_1[791:784] < mid_1[799:792]) ? 1 : 0;
assign detect_min[97][14] = (mid_1[791:784] < mid_2[783:776]) ? 1 : 0;
assign detect_min[97][15] = (mid_1[791:784] < mid_2[791:784]) ? 1 : 0;
assign detect_min[97][16] = (mid_1[791:784] < mid_2[799:792]) ? 1 : 0;
assign detect_min[97][17] = (mid_1[791:784] < btm_0[783:776]) ? 1 : 0;
assign detect_min[97][18] = (mid_1[791:784] < btm_0[791:784]) ? 1 : 0;
assign detect_min[97][19] = (mid_1[791:784] < btm_0[799:792]) ? 1 : 0;
assign detect_min[97][20] = (mid_1[791:784] < btm_1[783:776]) ? 1 : 0;
assign detect_min[97][21] = (mid_1[791:784] < btm_1[791:784]) ? 1 : 0;
assign detect_min[97][22] = (mid_1[791:784] < btm_1[799:792]) ? 1 : 0;
assign detect_min[97][23] = (mid_1[791:784] < btm_2[783:776]) ? 1 : 0;
assign detect_min[97][24] = (mid_1[791:784] < btm_2[791:784]) ? 1 : 0;
assign detect_min[97][25] = (mid_1[791:784] < btm_2[799:792]) ? 1 : 0;

assign detect_min[98][0] = (mid_1[799:792] < top_0[791:784]) ? 1 : 0;
assign detect_min[98][1] = (mid_1[799:792] < top_0[799:792]) ? 1 : 0;
assign detect_min[98][2] = (mid_1[799:792] < top_0[807:800]) ? 1 : 0;
assign detect_min[98][3] = (mid_1[799:792] < top_1[791:784]) ? 1 : 0;
assign detect_min[98][4] = (mid_1[799:792] < top_1[799:792]) ? 1 : 0;
assign detect_min[98][5] = (mid_1[799:792] < top_1[807:800]) ? 1 : 0;
assign detect_min[98][6] = (mid_1[799:792] < top_2[791:784]) ? 1 : 0;
assign detect_min[98][7] = (mid_1[799:792] < top_2[799:792]) ? 1 : 0;
assign detect_min[98][8] = (mid_1[799:792] < top_2[807:800]) ? 1 : 0;
assign detect_min[98][9] = (mid_1[799:792] < mid_0[791:784]) ? 1 : 0;
assign detect_min[98][10] = (mid_1[799:792] < mid_0[799:792]) ? 1 : 0;
assign detect_min[98][11] = (mid_1[799:792] < mid_0[807:800]) ? 1 : 0;
assign detect_min[98][12] = (mid_1[799:792] < mid_1[791:784]) ? 1 : 0;
assign detect_min[98][13] = (mid_1[799:792] < mid_1[807:800]) ? 1 : 0;
assign detect_min[98][14] = (mid_1[799:792] < mid_2[791:784]) ? 1 : 0;
assign detect_min[98][15] = (mid_1[799:792] < mid_2[799:792]) ? 1 : 0;
assign detect_min[98][16] = (mid_1[799:792] < mid_2[807:800]) ? 1 : 0;
assign detect_min[98][17] = (mid_1[799:792] < btm_0[791:784]) ? 1 : 0;
assign detect_min[98][18] = (mid_1[799:792] < btm_0[799:792]) ? 1 : 0;
assign detect_min[98][19] = (mid_1[799:792] < btm_0[807:800]) ? 1 : 0;
assign detect_min[98][20] = (mid_1[799:792] < btm_1[791:784]) ? 1 : 0;
assign detect_min[98][21] = (mid_1[799:792] < btm_1[799:792]) ? 1 : 0;
assign detect_min[98][22] = (mid_1[799:792] < btm_1[807:800]) ? 1 : 0;
assign detect_min[98][23] = (mid_1[799:792] < btm_2[791:784]) ? 1 : 0;
assign detect_min[98][24] = (mid_1[799:792] < btm_2[799:792]) ? 1 : 0;
assign detect_min[98][25] = (mid_1[799:792] < btm_2[807:800]) ? 1 : 0;

assign detect_min[99][0] = (mid_1[807:800] < top_0[799:792]) ? 1 : 0;
assign detect_min[99][1] = (mid_1[807:800] < top_0[807:800]) ? 1 : 0;
assign detect_min[99][2] = (mid_1[807:800] < top_0[815:808]) ? 1 : 0;
assign detect_min[99][3] = (mid_1[807:800] < top_1[799:792]) ? 1 : 0;
assign detect_min[99][4] = (mid_1[807:800] < top_1[807:800]) ? 1 : 0;
assign detect_min[99][5] = (mid_1[807:800] < top_1[815:808]) ? 1 : 0;
assign detect_min[99][6] = (mid_1[807:800] < top_2[799:792]) ? 1 : 0;
assign detect_min[99][7] = (mid_1[807:800] < top_2[807:800]) ? 1 : 0;
assign detect_min[99][8] = (mid_1[807:800] < top_2[815:808]) ? 1 : 0;
assign detect_min[99][9] = (mid_1[807:800] < mid_0[799:792]) ? 1 : 0;
assign detect_min[99][10] = (mid_1[807:800] < mid_0[807:800]) ? 1 : 0;
assign detect_min[99][11] = (mid_1[807:800] < mid_0[815:808]) ? 1 : 0;
assign detect_min[99][12] = (mid_1[807:800] < mid_1[799:792]) ? 1 : 0;
assign detect_min[99][13] = (mid_1[807:800] < mid_1[815:808]) ? 1 : 0;
assign detect_min[99][14] = (mid_1[807:800] < mid_2[799:792]) ? 1 : 0;
assign detect_min[99][15] = (mid_1[807:800] < mid_2[807:800]) ? 1 : 0;
assign detect_min[99][16] = (mid_1[807:800] < mid_2[815:808]) ? 1 : 0;
assign detect_min[99][17] = (mid_1[807:800] < btm_0[799:792]) ? 1 : 0;
assign detect_min[99][18] = (mid_1[807:800] < btm_0[807:800]) ? 1 : 0;
assign detect_min[99][19] = (mid_1[807:800] < btm_0[815:808]) ? 1 : 0;
assign detect_min[99][20] = (mid_1[807:800] < btm_1[799:792]) ? 1 : 0;
assign detect_min[99][21] = (mid_1[807:800] < btm_1[807:800]) ? 1 : 0;
assign detect_min[99][22] = (mid_1[807:800] < btm_1[815:808]) ? 1 : 0;
assign detect_min[99][23] = (mid_1[807:800] < btm_2[799:792]) ? 1 : 0;
assign detect_min[99][24] = (mid_1[807:800] < btm_2[807:800]) ? 1 : 0;
assign detect_min[99][25] = (mid_1[807:800] < btm_2[815:808]) ? 1 : 0;

assign detect_min[100][0] = (mid_1[815:808] < top_0[807:800]) ? 1 : 0;
assign detect_min[100][1] = (mid_1[815:808] < top_0[815:808]) ? 1 : 0;
assign detect_min[100][2] = (mid_1[815:808] < top_0[823:816]) ? 1 : 0;
assign detect_min[100][3] = (mid_1[815:808] < top_1[807:800]) ? 1 : 0;
assign detect_min[100][4] = (mid_1[815:808] < top_1[815:808]) ? 1 : 0;
assign detect_min[100][5] = (mid_1[815:808] < top_1[823:816]) ? 1 : 0;
assign detect_min[100][6] = (mid_1[815:808] < top_2[807:800]) ? 1 : 0;
assign detect_min[100][7] = (mid_1[815:808] < top_2[815:808]) ? 1 : 0;
assign detect_min[100][8] = (mid_1[815:808] < top_2[823:816]) ? 1 : 0;
assign detect_min[100][9] = (mid_1[815:808] < mid_0[807:800]) ? 1 : 0;
assign detect_min[100][10] = (mid_1[815:808] < mid_0[815:808]) ? 1 : 0;
assign detect_min[100][11] = (mid_1[815:808] < mid_0[823:816]) ? 1 : 0;
assign detect_min[100][12] = (mid_1[815:808] < mid_1[807:800]) ? 1 : 0;
assign detect_min[100][13] = (mid_1[815:808] < mid_1[823:816]) ? 1 : 0;
assign detect_min[100][14] = (mid_1[815:808] < mid_2[807:800]) ? 1 : 0;
assign detect_min[100][15] = (mid_1[815:808] < mid_2[815:808]) ? 1 : 0;
assign detect_min[100][16] = (mid_1[815:808] < mid_2[823:816]) ? 1 : 0;
assign detect_min[100][17] = (mid_1[815:808] < btm_0[807:800]) ? 1 : 0;
assign detect_min[100][18] = (mid_1[815:808] < btm_0[815:808]) ? 1 : 0;
assign detect_min[100][19] = (mid_1[815:808] < btm_0[823:816]) ? 1 : 0;
assign detect_min[100][20] = (mid_1[815:808] < btm_1[807:800]) ? 1 : 0;
assign detect_min[100][21] = (mid_1[815:808] < btm_1[815:808]) ? 1 : 0;
assign detect_min[100][22] = (mid_1[815:808] < btm_1[823:816]) ? 1 : 0;
assign detect_min[100][23] = (mid_1[815:808] < btm_2[807:800]) ? 1 : 0;
assign detect_min[100][24] = (mid_1[815:808] < btm_2[815:808]) ? 1 : 0;
assign detect_min[100][25] = (mid_1[815:808] < btm_2[823:816]) ? 1 : 0;

assign detect_min[101][0] = (mid_1[823:816] < top_0[815:808]) ? 1 : 0;
assign detect_min[101][1] = (mid_1[823:816] < top_0[823:816]) ? 1 : 0;
assign detect_min[101][2] = (mid_1[823:816] < top_0[831:824]) ? 1 : 0;
assign detect_min[101][3] = (mid_1[823:816] < top_1[815:808]) ? 1 : 0;
assign detect_min[101][4] = (mid_1[823:816] < top_1[823:816]) ? 1 : 0;
assign detect_min[101][5] = (mid_1[823:816] < top_1[831:824]) ? 1 : 0;
assign detect_min[101][6] = (mid_1[823:816] < top_2[815:808]) ? 1 : 0;
assign detect_min[101][7] = (mid_1[823:816] < top_2[823:816]) ? 1 : 0;
assign detect_min[101][8] = (mid_1[823:816] < top_2[831:824]) ? 1 : 0;
assign detect_min[101][9] = (mid_1[823:816] < mid_0[815:808]) ? 1 : 0;
assign detect_min[101][10] = (mid_1[823:816] < mid_0[823:816]) ? 1 : 0;
assign detect_min[101][11] = (mid_1[823:816] < mid_0[831:824]) ? 1 : 0;
assign detect_min[101][12] = (mid_1[823:816] < mid_1[815:808]) ? 1 : 0;
assign detect_min[101][13] = (mid_1[823:816] < mid_1[831:824]) ? 1 : 0;
assign detect_min[101][14] = (mid_1[823:816] < mid_2[815:808]) ? 1 : 0;
assign detect_min[101][15] = (mid_1[823:816] < mid_2[823:816]) ? 1 : 0;
assign detect_min[101][16] = (mid_1[823:816] < mid_2[831:824]) ? 1 : 0;
assign detect_min[101][17] = (mid_1[823:816] < btm_0[815:808]) ? 1 : 0;
assign detect_min[101][18] = (mid_1[823:816] < btm_0[823:816]) ? 1 : 0;
assign detect_min[101][19] = (mid_1[823:816] < btm_0[831:824]) ? 1 : 0;
assign detect_min[101][20] = (mid_1[823:816] < btm_1[815:808]) ? 1 : 0;
assign detect_min[101][21] = (mid_1[823:816] < btm_1[823:816]) ? 1 : 0;
assign detect_min[101][22] = (mid_1[823:816] < btm_1[831:824]) ? 1 : 0;
assign detect_min[101][23] = (mid_1[823:816] < btm_2[815:808]) ? 1 : 0;
assign detect_min[101][24] = (mid_1[823:816] < btm_2[823:816]) ? 1 : 0;
assign detect_min[101][25] = (mid_1[823:816] < btm_2[831:824]) ? 1 : 0;

assign detect_min[102][0] = (mid_1[831:824] < top_0[823:816]) ? 1 : 0;
assign detect_min[102][1] = (mid_1[831:824] < top_0[831:824]) ? 1 : 0;
assign detect_min[102][2] = (mid_1[831:824] < top_0[839:832]) ? 1 : 0;
assign detect_min[102][3] = (mid_1[831:824] < top_1[823:816]) ? 1 : 0;
assign detect_min[102][4] = (mid_1[831:824] < top_1[831:824]) ? 1 : 0;
assign detect_min[102][5] = (mid_1[831:824] < top_1[839:832]) ? 1 : 0;
assign detect_min[102][6] = (mid_1[831:824] < top_2[823:816]) ? 1 : 0;
assign detect_min[102][7] = (mid_1[831:824] < top_2[831:824]) ? 1 : 0;
assign detect_min[102][8] = (mid_1[831:824] < top_2[839:832]) ? 1 : 0;
assign detect_min[102][9] = (mid_1[831:824] < mid_0[823:816]) ? 1 : 0;
assign detect_min[102][10] = (mid_1[831:824] < mid_0[831:824]) ? 1 : 0;
assign detect_min[102][11] = (mid_1[831:824] < mid_0[839:832]) ? 1 : 0;
assign detect_min[102][12] = (mid_1[831:824] < mid_1[823:816]) ? 1 : 0;
assign detect_min[102][13] = (mid_1[831:824] < mid_1[839:832]) ? 1 : 0;
assign detect_min[102][14] = (mid_1[831:824] < mid_2[823:816]) ? 1 : 0;
assign detect_min[102][15] = (mid_1[831:824] < mid_2[831:824]) ? 1 : 0;
assign detect_min[102][16] = (mid_1[831:824] < mid_2[839:832]) ? 1 : 0;
assign detect_min[102][17] = (mid_1[831:824] < btm_0[823:816]) ? 1 : 0;
assign detect_min[102][18] = (mid_1[831:824] < btm_0[831:824]) ? 1 : 0;
assign detect_min[102][19] = (mid_1[831:824] < btm_0[839:832]) ? 1 : 0;
assign detect_min[102][20] = (mid_1[831:824] < btm_1[823:816]) ? 1 : 0;
assign detect_min[102][21] = (mid_1[831:824] < btm_1[831:824]) ? 1 : 0;
assign detect_min[102][22] = (mid_1[831:824] < btm_1[839:832]) ? 1 : 0;
assign detect_min[102][23] = (mid_1[831:824] < btm_2[823:816]) ? 1 : 0;
assign detect_min[102][24] = (mid_1[831:824] < btm_2[831:824]) ? 1 : 0;
assign detect_min[102][25] = (mid_1[831:824] < btm_2[839:832]) ? 1 : 0;

assign detect_min[103][0] = (mid_1[839:832] < top_0[831:824]) ? 1 : 0;
assign detect_min[103][1] = (mid_1[839:832] < top_0[839:832]) ? 1 : 0;
assign detect_min[103][2] = (mid_1[839:832] < top_0[847:840]) ? 1 : 0;
assign detect_min[103][3] = (mid_1[839:832] < top_1[831:824]) ? 1 : 0;
assign detect_min[103][4] = (mid_1[839:832] < top_1[839:832]) ? 1 : 0;
assign detect_min[103][5] = (mid_1[839:832] < top_1[847:840]) ? 1 : 0;
assign detect_min[103][6] = (mid_1[839:832] < top_2[831:824]) ? 1 : 0;
assign detect_min[103][7] = (mid_1[839:832] < top_2[839:832]) ? 1 : 0;
assign detect_min[103][8] = (mid_1[839:832] < top_2[847:840]) ? 1 : 0;
assign detect_min[103][9] = (mid_1[839:832] < mid_0[831:824]) ? 1 : 0;
assign detect_min[103][10] = (mid_1[839:832] < mid_0[839:832]) ? 1 : 0;
assign detect_min[103][11] = (mid_1[839:832] < mid_0[847:840]) ? 1 : 0;
assign detect_min[103][12] = (mid_1[839:832] < mid_1[831:824]) ? 1 : 0;
assign detect_min[103][13] = (mid_1[839:832] < mid_1[847:840]) ? 1 : 0;
assign detect_min[103][14] = (mid_1[839:832] < mid_2[831:824]) ? 1 : 0;
assign detect_min[103][15] = (mid_1[839:832] < mid_2[839:832]) ? 1 : 0;
assign detect_min[103][16] = (mid_1[839:832] < mid_2[847:840]) ? 1 : 0;
assign detect_min[103][17] = (mid_1[839:832] < btm_0[831:824]) ? 1 : 0;
assign detect_min[103][18] = (mid_1[839:832] < btm_0[839:832]) ? 1 : 0;
assign detect_min[103][19] = (mid_1[839:832] < btm_0[847:840]) ? 1 : 0;
assign detect_min[103][20] = (mid_1[839:832] < btm_1[831:824]) ? 1 : 0;
assign detect_min[103][21] = (mid_1[839:832] < btm_1[839:832]) ? 1 : 0;
assign detect_min[103][22] = (mid_1[839:832] < btm_1[847:840]) ? 1 : 0;
assign detect_min[103][23] = (mid_1[839:832] < btm_2[831:824]) ? 1 : 0;
assign detect_min[103][24] = (mid_1[839:832] < btm_2[839:832]) ? 1 : 0;
assign detect_min[103][25] = (mid_1[839:832] < btm_2[847:840]) ? 1 : 0;

assign detect_min[104][0] = (mid_1[847:840] < top_0[839:832]) ? 1 : 0;
assign detect_min[104][1] = (mid_1[847:840] < top_0[847:840]) ? 1 : 0;
assign detect_min[104][2] = (mid_1[847:840] < top_0[855:848]) ? 1 : 0;
assign detect_min[104][3] = (mid_1[847:840] < top_1[839:832]) ? 1 : 0;
assign detect_min[104][4] = (mid_1[847:840] < top_1[847:840]) ? 1 : 0;
assign detect_min[104][5] = (mid_1[847:840] < top_1[855:848]) ? 1 : 0;
assign detect_min[104][6] = (mid_1[847:840] < top_2[839:832]) ? 1 : 0;
assign detect_min[104][7] = (mid_1[847:840] < top_2[847:840]) ? 1 : 0;
assign detect_min[104][8] = (mid_1[847:840] < top_2[855:848]) ? 1 : 0;
assign detect_min[104][9] = (mid_1[847:840] < mid_0[839:832]) ? 1 : 0;
assign detect_min[104][10] = (mid_1[847:840] < mid_0[847:840]) ? 1 : 0;
assign detect_min[104][11] = (mid_1[847:840] < mid_0[855:848]) ? 1 : 0;
assign detect_min[104][12] = (mid_1[847:840] < mid_1[839:832]) ? 1 : 0;
assign detect_min[104][13] = (mid_1[847:840] < mid_1[855:848]) ? 1 : 0;
assign detect_min[104][14] = (mid_1[847:840] < mid_2[839:832]) ? 1 : 0;
assign detect_min[104][15] = (mid_1[847:840] < mid_2[847:840]) ? 1 : 0;
assign detect_min[104][16] = (mid_1[847:840] < mid_2[855:848]) ? 1 : 0;
assign detect_min[104][17] = (mid_1[847:840] < btm_0[839:832]) ? 1 : 0;
assign detect_min[104][18] = (mid_1[847:840] < btm_0[847:840]) ? 1 : 0;
assign detect_min[104][19] = (mid_1[847:840] < btm_0[855:848]) ? 1 : 0;
assign detect_min[104][20] = (mid_1[847:840] < btm_1[839:832]) ? 1 : 0;
assign detect_min[104][21] = (mid_1[847:840] < btm_1[847:840]) ? 1 : 0;
assign detect_min[104][22] = (mid_1[847:840] < btm_1[855:848]) ? 1 : 0;
assign detect_min[104][23] = (mid_1[847:840] < btm_2[839:832]) ? 1 : 0;
assign detect_min[104][24] = (mid_1[847:840] < btm_2[847:840]) ? 1 : 0;
assign detect_min[104][25] = (mid_1[847:840] < btm_2[855:848]) ? 1 : 0;

assign detect_min[105][0] = (mid_1[855:848] < top_0[847:840]) ? 1 : 0;
assign detect_min[105][1] = (mid_1[855:848] < top_0[855:848]) ? 1 : 0;
assign detect_min[105][2] = (mid_1[855:848] < top_0[863:856]) ? 1 : 0;
assign detect_min[105][3] = (mid_1[855:848] < top_1[847:840]) ? 1 : 0;
assign detect_min[105][4] = (mid_1[855:848] < top_1[855:848]) ? 1 : 0;
assign detect_min[105][5] = (mid_1[855:848] < top_1[863:856]) ? 1 : 0;
assign detect_min[105][6] = (mid_1[855:848] < top_2[847:840]) ? 1 : 0;
assign detect_min[105][7] = (mid_1[855:848] < top_2[855:848]) ? 1 : 0;
assign detect_min[105][8] = (mid_1[855:848] < top_2[863:856]) ? 1 : 0;
assign detect_min[105][9] = (mid_1[855:848] < mid_0[847:840]) ? 1 : 0;
assign detect_min[105][10] = (mid_1[855:848] < mid_0[855:848]) ? 1 : 0;
assign detect_min[105][11] = (mid_1[855:848] < mid_0[863:856]) ? 1 : 0;
assign detect_min[105][12] = (mid_1[855:848] < mid_1[847:840]) ? 1 : 0;
assign detect_min[105][13] = (mid_1[855:848] < mid_1[863:856]) ? 1 : 0;
assign detect_min[105][14] = (mid_1[855:848] < mid_2[847:840]) ? 1 : 0;
assign detect_min[105][15] = (mid_1[855:848] < mid_2[855:848]) ? 1 : 0;
assign detect_min[105][16] = (mid_1[855:848] < mid_2[863:856]) ? 1 : 0;
assign detect_min[105][17] = (mid_1[855:848] < btm_0[847:840]) ? 1 : 0;
assign detect_min[105][18] = (mid_1[855:848] < btm_0[855:848]) ? 1 : 0;
assign detect_min[105][19] = (mid_1[855:848] < btm_0[863:856]) ? 1 : 0;
assign detect_min[105][20] = (mid_1[855:848] < btm_1[847:840]) ? 1 : 0;
assign detect_min[105][21] = (mid_1[855:848] < btm_1[855:848]) ? 1 : 0;
assign detect_min[105][22] = (mid_1[855:848] < btm_1[863:856]) ? 1 : 0;
assign detect_min[105][23] = (mid_1[855:848] < btm_2[847:840]) ? 1 : 0;
assign detect_min[105][24] = (mid_1[855:848] < btm_2[855:848]) ? 1 : 0;
assign detect_min[105][25] = (mid_1[855:848] < btm_2[863:856]) ? 1 : 0;

assign detect_min[106][0] = (mid_1[863:856] < top_0[855:848]) ? 1 : 0;
assign detect_min[106][1] = (mid_1[863:856] < top_0[863:856]) ? 1 : 0;
assign detect_min[106][2] = (mid_1[863:856] < top_0[871:864]) ? 1 : 0;
assign detect_min[106][3] = (mid_1[863:856] < top_1[855:848]) ? 1 : 0;
assign detect_min[106][4] = (mid_1[863:856] < top_1[863:856]) ? 1 : 0;
assign detect_min[106][5] = (mid_1[863:856] < top_1[871:864]) ? 1 : 0;
assign detect_min[106][6] = (mid_1[863:856] < top_2[855:848]) ? 1 : 0;
assign detect_min[106][7] = (mid_1[863:856] < top_2[863:856]) ? 1 : 0;
assign detect_min[106][8] = (mid_1[863:856] < top_2[871:864]) ? 1 : 0;
assign detect_min[106][9] = (mid_1[863:856] < mid_0[855:848]) ? 1 : 0;
assign detect_min[106][10] = (mid_1[863:856] < mid_0[863:856]) ? 1 : 0;
assign detect_min[106][11] = (mid_1[863:856] < mid_0[871:864]) ? 1 : 0;
assign detect_min[106][12] = (mid_1[863:856] < mid_1[855:848]) ? 1 : 0;
assign detect_min[106][13] = (mid_1[863:856] < mid_1[871:864]) ? 1 : 0;
assign detect_min[106][14] = (mid_1[863:856] < mid_2[855:848]) ? 1 : 0;
assign detect_min[106][15] = (mid_1[863:856] < mid_2[863:856]) ? 1 : 0;
assign detect_min[106][16] = (mid_1[863:856] < mid_2[871:864]) ? 1 : 0;
assign detect_min[106][17] = (mid_1[863:856] < btm_0[855:848]) ? 1 : 0;
assign detect_min[106][18] = (mid_1[863:856] < btm_0[863:856]) ? 1 : 0;
assign detect_min[106][19] = (mid_1[863:856] < btm_0[871:864]) ? 1 : 0;
assign detect_min[106][20] = (mid_1[863:856] < btm_1[855:848]) ? 1 : 0;
assign detect_min[106][21] = (mid_1[863:856] < btm_1[863:856]) ? 1 : 0;
assign detect_min[106][22] = (mid_1[863:856] < btm_1[871:864]) ? 1 : 0;
assign detect_min[106][23] = (mid_1[863:856] < btm_2[855:848]) ? 1 : 0;
assign detect_min[106][24] = (mid_1[863:856] < btm_2[863:856]) ? 1 : 0;
assign detect_min[106][25] = (mid_1[863:856] < btm_2[871:864]) ? 1 : 0;

assign detect_min[107][0] = (mid_1[871:864] < top_0[863:856]) ? 1 : 0;
assign detect_min[107][1] = (mid_1[871:864] < top_0[871:864]) ? 1 : 0;
assign detect_min[107][2] = (mid_1[871:864] < top_0[879:872]) ? 1 : 0;
assign detect_min[107][3] = (mid_1[871:864] < top_1[863:856]) ? 1 : 0;
assign detect_min[107][4] = (mid_1[871:864] < top_1[871:864]) ? 1 : 0;
assign detect_min[107][5] = (mid_1[871:864] < top_1[879:872]) ? 1 : 0;
assign detect_min[107][6] = (mid_1[871:864] < top_2[863:856]) ? 1 : 0;
assign detect_min[107][7] = (mid_1[871:864] < top_2[871:864]) ? 1 : 0;
assign detect_min[107][8] = (mid_1[871:864] < top_2[879:872]) ? 1 : 0;
assign detect_min[107][9] = (mid_1[871:864] < mid_0[863:856]) ? 1 : 0;
assign detect_min[107][10] = (mid_1[871:864] < mid_0[871:864]) ? 1 : 0;
assign detect_min[107][11] = (mid_1[871:864] < mid_0[879:872]) ? 1 : 0;
assign detect_min[107][12] = (mid_1[871:864] < mid_1[863:856]) ? 1 : 0;
assign detect_min[107][13] = (mid_1[871:864] < mid_1[879:872]) ? 1 : 0;
assign detect_min[107][14] = (mid_1[871:864] < mid_2[863:856]) ? 1 : 0;
assign detect_min[107][15] = (mid_1[871:864] < mid_2[871:864]) ? 1 : 0;
assign detect_min[107][16] = (mid_1[871:864] < mid_2[879:872]) ? 1 : 0;
assign detect_min[107][17] = (mid_1[871:864] < btm_0[863:856]) ? 1 : 0;
assign detect_min[107][18] = (mid_1[871:864] < btm_0[871:864]) ? 1 : 0;
assign detect_min[107][19] = (mid_1[871:864] < btm_0[879:872]) ? 1 : 0;
assign detect_min[107][20] = (mid_1[871:864] < btm_1[863:856]) ? 1 : 0;
assign detect_min[107][21] = (mid_1[871:864] < btm_1[871:864]) ? 1 : 0;
assign detect_min[107][22] = (mid_1[871:864] < btm_1[879:872]) ? 1 : 0;
assign detect_min[107][23] = (mid_1[871:864] < btm_2[863:856]) ? 1 : 0;
assign detect_min[107][24] = (mid_1[871:864] < btm_2[871:864]) ? 1 : 0;
assign detect_min[107][25] = (mid_1[871:864] < btm_2[879:872]) ? 1 : 0;

assign detect_min[108][0] = (mid_1[879:872] < top_0[871:864]) ? 1 : 0;
assign detect_min[108][1] = (mid_1[879:872] < top_0[879:872]) ? 1 : 0;
assign detect_min[108][2] = (mid_1[879:872] < top_0[887:880]) ? 1 : 0;
assign detect_min[108][3] = (mid_1[879:872] < top_1[871:864]) ? 1 : 0;
assign detect_min[108][4] = (mid_1[879:872] < top_1[879:872]) ? 1 : 0;
assign detect_min[108][5] = (mid_1[879:872] < top_1[887:880]) ? 1 : 0;
assign detect_min[108][6] = (mid_1[879:872] < top_2[871:864]) ? 1 : 0;
assign detect_min[108][7] = (mid_1[879:872] < top_2[879:872]) ? 1 : 0;
assign detect_min[108][8] = (mid_1[879:872] < top_2[887:880]) ? 1 : 0;
assign detect_min[108][9] = (mid_1[879:872] < mid_0[871:864]) ? 1 : 0;
assign detect_min[108][10] = (mid_1[879:872] < mid_0[879:872]) ? 1 : 0;
assign detect_min[108][11] = (mid_1[879:872] < mid_0[887:880]) ? 1 : 0;
assign detect_min[108][12] = (mid_1[879:872] < mid_1[871:864]) ? 1 : 0;
assign detect_min[108][13] = (mid_1[879:872] < mid_1[887:880]) ? 1 : 0;
assign detect_min[108][14] = (mid_1[879:872] < mid_2[871:864]) ? 1 : 0;
assign detect_min[108][15] = (mid_1[879:872] < mid_2[879:872]) ? 1 : 0;
assign detect_min[108][16] = (mid_1[879:872] < mid_2[887:880]) ? 1 : 0;
assign detect_min[108][17] = (mid_1[879:872] < btm_0[871:864]) ? 1 : 0;
assign detect_min[108][18] = (mid_1[879:872] < btm_0[879:872]) ? 1 : 0;
assign detect_min[108][19] = (mid_1[879:872] < btm_0[887:880]) ? 1 : 0;
assign detect_min[108][20] = (mid_1[879:872] < btm_1[871:864]) ? 1 : 0;
assign detect_min[108][21] = (mid_1[879:872] < btm_1[879:872]) ? 1 : 0;
assign detect_min[108][22] = (mid_1[879:872] < btm_1[887:880]) ? 1 : 0;
assign detect_min[108][23] = (mid_1[879:872] < btm_2[871:864]) ? 1 : 0;
assign detect_min[108][24] = (mid_1[879:872] < btm_2[879:872]) ? 1 : 0;
assign detect_min[108][25] = (mid_1[879:872] < btm_2[887:880]) ? 1 : 0;

assign detect_min[109][0] = (mid_1[887:880] < top_0[879:872]) ? 1 : 0;
assign detect_min[109][1] = (mid_1[887:880] < top_0[887:880]) ? 1 : 0;
assign detect_min[109][2] = (mid_1[887:880] < top_0[895:888]) ? 1 : 0;
assign detect_min[109][3] = (mid_1[887:880] < top_1[879:872]) ? 1 : 0;
assign detect_min[109][4] = (mid_1[887:880] < top_1[887:880]) ? 1 : 0;
assign detect_min[109][5] = (mid_1[887:880] < top_1[895:888]) ? 1 : 0;
assign detect_min[109][6] = (mid_1[887:880] < top_2[879:872]) ? 1 : 0;
assign detect_min[109][7] = (mid_1[887:880] < top_2[887:880]) ? 1 : 0;
assign detect_min[109][8] = (mid_1[887:880] < top_2[895:888]) ? 1 : 0;
assign detect_min[109][9] = (mid_1[887:880] < mid_0[879:872]) ? 1 : 0;
assign detect_min[109][10] = (mid_1[887:880] < mid_0[887:880]) ? 1 : 0;
assign detect_min[109][11] = (mid_1[887:880] < mid_0[895:888]) ? 1 : 0;
assign detect_min[109][12] = (mid_1[887:880] < mid_1[879:872]) ? 1 : 0;
assign detect_min[109][13] = (mid_1[887:880] < mid_1[895:888]) ? 1 : 0;
assign detect_min[109][14] = (mid_1[887:880] < mid_2[879:872]) ? 1 : 0;
assign detect_min[109][15] = (mid_1[887:880] < mid_2[887:880]) ? 1 : 0;
assign detect_min[109][16] = (mid_1[887:880] < mid_2[895:888]) ? 1 : 0;
assign detect_min[109][17] = (mid_1[887:880] < btm_0[879:872]) ? 1 : 0;
assign detect_min[109][18] = (mid_1[887:880] < btm_0[887:880]) ? 1 : 0;
assign detect_min[109][19] = (mid_1[887:880] < btm_0[895:888]) ? 1 : 0;
assign detect_min[109][20] = (mid_1[887:880] < btm_1[879:872]) ? 1 : 0;
assign detect_min[109][21] = (mid_1[887:880] < btm_1[887:880]) ? 1 : 0;
assign detect_min[109][22] = (mid_1[887:880] < btm_1[895:888]) ? 1 : 0;
assign detect_min[109][23] = (mid_1[887:880] < btm_2[879:872]) ? 1 : 0;
assign detect_min[109][24] = (mid_1[887:880] < btm_2[887:880]) ? 1 : 0;
assign detect_min[109][25] = (mid_1[887:880] < btm_2[895:888]) ? 1 : 0;

assign detect_min[110][0] = (mid_1[895:888] < top_0[887:880]) ? 1 : 0;
assign detect_min[110][1] = (mid_1[895:888] < top_0[895:888]) ? 1 : 0;
assign detect_min[110][2] = (mid_1[895:888] < top_0[903:896]) ? 1 : 0;
assign detect_min[110][3] = (mid_1[895:888] < top_1[887:880]) ? 1 : 0;
assign detect_min[110][4] = (mid_1[895:888] < top_1[895:888]) ? 1 : 0;
assign detect_min[110][5] = (mid_1[895:888] < top_1[903:896]) ? 1 : 0;
assign detect_min[110][6] = (mid_1[895:888] < top_2[887:880]) ? 1 : 0;
assign detect_min[110][7] = (mid_1[895:888] < top_2[895:888]) ? 1 : 0;
assign detect_min[110][8] = (mid_1[895:888] < top_2[903:896]) ? 1 : 0;
assign detect_min[110][9] = (mid_1[895:888] < mid_0[887:880]) ? 1 : 0;
assign detect_min[110][10] = (mid_1[895:888] < mid_0[895:888]) ? 1 : 0;
assign detect_min[110][11] = (mid_1[895:888] < mid_0[903:896]) ? 1 : 0;
assign detect_min[110][12] = (mid_1[895:888] < mid_1[887:880]) ? 1 : 0;
assign detect_min[110][13] = (mid_1[895:888] < mid_1[903:896]) ? 1 : 0;
assign detect_min[110][14] = (mid_1[895:888] < mid_2[887:880]) ? 1 : 0;
assign detect_min[110][15] = (mid_1[895:888] < mid_2[895:888]) ? 1 : 0;
assign detect_min[110][16] = (mid_1[895:888] < mid_2[903:896]) ? 1 : 0;
assign detect_min[110][17] = (mid_1[895:888] < btm_0[887:880]) ? 1 : 0;
assign detect_min[110][18] = (mid_1[895:888] < btm_0[895:888]) ? 1 : 0;
assign detect_min[110][19] = (mid_1[895:888] < btm_0[903:896]) ? 1 : 0;
assign detect_min[110][20] = (mid_1[895:888] < btm_1[887:880]) ? 1 : 0;
assign detect_min[110][21] = (mid_1[895:888] < btm_1[895:888]) ? 1 : 0;
assign detect_min[110][22] = (mid_1[895:888] < btm_1[903:896]) ? 1 : 0;
assign detect_min[110][23] = (mid_1[895:888] < btm_2[887:880]) ? 1 : 0;
assign detect_min[110][24] = (mid_1[895:888] < btm_2[895:888]) ? 1 : 0;
assign detect_min[110][25] = (mid_1[895:888] < btm_2[903:896]) ? 1 : 0;

assign detect_min[111][0] = (mid_1[903:896] < top_0[895:888]) ? 1 : 0;
assign detect_min[111][1] = (mid_1[903:896] < top_0[903:896]) ? 1 : 0;
assign detect_min[111][2] = (mid_1[903:896] < top_0[911:904]) ? 1 : 0;
assign detect_min[111][3] = (mid_1[903:896] < top_1[895:888]) ? 1 : 0;
assign detect_min[111][4] = (mid_1[903:896] < top_1[903:896]) ? 1 : 0;
assign detect_min[111][5] = (mid_1[903:896] < top_1[911:904]) ? 1 : 0;
assign detect_min[111][6] = (mid_1[903:896] < top_2[895:888]) ? 1 : 0;
assign detect_min[111][7] = (mid_1[903:896] < top_2[903:896]) ? 1 : 0;
assign detect_min[111][8] = (mid_1[903:896] < top_2[911:904]) ? 1 : 0;
assign detect_min[111][9] = (mid_1[903:896] < mid_0[895:888]) ? 1 : 0;
assign detect_min[111][10] = (mid_1[903:896] < mid_0[903:896]) ? 1 : 0;
assign detect_min[111][11] = (mid_1[903:896] < mid_0[911:904]) ? 1 : 0;
assign detect_min[111][12] = (mid_1[903:896] < mid_1[895:888]) ? 1 : 0;
assign detect_min[111][13] = (mid_1[903:896] < mid_1[911:904]) ? 1 : 0;
assign detect_min[111][14] = (mid_1[903:896] < mid_2[895:888]) ? 1 : 0;
assign detect_min[111][15] = (mid_1[903:896] < mid_2[903:896]) ? 1 : 0;
assign detect_min[111][16] = (mid_1[903:896] < mid_2[911:904]) ? 1 : 0;
assign detect_min[111][17] = (mid_1[903:896] < btm_0[895:888]) ? 1 : 0;
assign detect_min[111][18] = (mid_1[903:896] < btm_0[903:896]) ? 1 : 0;
assign detect_min[111][19] = (mid_1[903:896] < btm_0[911:904]) ? 1 : 0;
assign detect_min[111][20] = (mid_1[903:896] < btm_1[895:888]) ? 1 : 0;
assign detect_min[111][21] = (mid_1[903:896] < btm_1[903:896]) ? 1 : 0;
assign detect_min[111][22] = (mid_1[903:896] < btm_1[911:904]) ? 1 : 0;
assign detect_min[111][23] = (mid_1[903:896] < btm_2[895:888]) ? 1 : 0;
assign detect_min[111][24] = (mid_1[903:896] < btm_2[903:896]) ? 1 : 0;
assign detect_min[111][25] = (mid_1[903:896] < btm_2[911:904]) ? 1 : 0;

assign detect_min[112][0] = (mid_1[911:904] < top_0[903:896]) ? 1 : 0;
assign detect_min[112][1] = (mid_1[911:904] < top_0[911:904]) ? 1 : 0;
assign detect_min[112][2] = (mid_1[911:904] < top_0[919:912]) ? 1 : 0;
assign detect_min[112][3] = (mid_1[911:904] < top_1[903:896]) ? 1 : 0;
assign detect_min[112][4] = (mid_1[911:904] < top_1[911:904]) ? 1 : 0;
assign detect_min[112][5] = (mid_1[911:904] < top_1[919:912]) ? 1 : 0;
assign detect_min[112][6] = (mid_1[911:904] < top_2[903:896]) ? 1 : 0;
assign detect_min[112][7] = (mid_1[911:904] < top_2[911:904]) ? 1 : 0;
assign detect_min[112][8] = (mid_1[911:904] < top_2[919:912]) ? 1 : 0;
assign detect_min[112][9] = (mid_1[911:904] < mid_0[903:896]) ? 1 : 0;
assign detect_min[112][10] = (mid_1[911:904] < mid_0[911:904]) ? 1 : 0;
assign detect_min[112][11] = (mid_1[911:904] < mid_0[919:912]) ? 1 : 0;
assign detect_min[112][12] = (mid_1[911:904] < mid_1[903:896]) ? 1 : 0;
assign detect_min[112][13] = (mid_1[911:904] < mid_1[919:912]) ? 1 : 0;
assign detect_min[112][14] = (mid_1[911:904] < mid_2[903:896]) ? 1 : 0;
assign detect_min[112][15] = (mid_1[911:904] < mid_2[911:904]) ? 1 : 0;
assign detect_min[112][16] = (mid_1[911:904] < mid_2[919:912]) ? 1 : 0;
assign detect_min[112][17] = (mid_1[911:904] < btm_0[903:896]) ? 1 : 0;
assign detect_min[112][18] = (mid_1[911:904] < btm_0[911:904]) ? 1 : 0;
assign detect_min[112][19] = (mid_1[911:904] < btm_0[919:912]) ? 1 : 0;
assign detect_min[112][20] = (mid_1[911:904] < btm_1[903:896]) ? 1 : 0;
assign detect_min[112][21] = (mid_1[911:904] < btm_1[911:904]) ? 1 : 0;
assign detect_min[112][22] = (mid_1[911:904] < btm_1[919:912]) ? 1 : 0;
assign detect_min[112][23] = (mid_1[911:904] < btm_2[903:896]) ? 1 : 0;
assign detect_min[112][24] = (mid_1[911:904] < btm_2[911:904]) ? 1 : 0;
assign detect_min[112][25] = (mid_1[911:904] < btm_2[919:912]) ? 1 : 0;

assign detect_min[113][0] = (mid_1[919:912] < top_0[911:904]) ? 1 : 0;
assign detect_min[113][1] = (mid_1[919:912] < top_0[919:912]) ? 1 : 0;
assign detect_min[113][2] = (mid_1[919:912] < top_0[927:920]) ? 1 : 0;
assign detect_min[113][3] = (mid_1[919:912] < top_1[911:904]) ? 1 : 0;
assign detect_min[113][4] = (mid_1[919:912] < top_1[919:912]) ? 1 : 0;
assign detect_min[113][5] = (mid_1[919:912] < top_1[927:920]) ? 1 : 0;
assign detect_min[113][6] = (mid_1[919:912] < top_2[911:904]) ? 1 : 0;
assign detect_min[113][7] = (mid_1[919:912] < top_2[919:912]) ? 1 : 0;
assign detect_min[113][8] = (mid_1[919:912] < top_2[927:920]) ? 1 : 0;
assign detect_min[113][9] = (mid_1[919:912] < mid_0[911:904]) ? 1 : 0;
assign detect_min[113][10] = (mid_1[919:912] < mid_0[919:912]) ? 1 : 0;
assign detect_min[113][11] = (mid_1[919:912] < mid_0[927:920]) ? 1 : 0;
assign detect_min[113][12] = (mid_1[919:912] < mid_1[911:904]) ? 1 : 0;
assign detect_min[113][13] = (mid_1[919:912] < mid_1[927:920]) ? 1 : 0;
assign detect_min[113][14] = (mid_1[919:912] < mid_2[911:904]) ? 1 : 0;
assign detect_min[113][15] = (mid_1[919:912] < mid_2[919:912]) ? 1 : 0;
assign detect_min[113][16] = (mid_1[919:912] < mid_2[927:920]) ? 1 : 0;
assign detect_min[113][17] = (mid_1[919:912] < btm_0[911:904]) ? 1 : 0;
assign detect_min[113][18] = (mid_1[919:912] < btm_0[919:912]) ? 1 : 0;
assign detect_min[113][19] = (mid_1[919:912] < btm_0[927:920]) ? 1 : 0;
assign detect_min[113][20] = (mid_1[919:912] < btm_1[911:904]) ? 1 : 0;
assign detect_min[113][21] = (mid_1[919:912] < btm_1[919:912]) ? 1 : 0;
assign detect_min[113][22] = (mid_1[919:912] < btm_1[927:920]) ? 1 : 0;
assign detect_min[113][23] = (mid_1[919:912] < btm_2[911:904]) ? 1 : 0;
assign detect_min[113][24] = (mid_1[919:912] < btm_2[919:912]) ? 1 : 0;
assign detect_min[113][25] = (mid_1[919:912] < btm_2[927:920]) ? 1 : 0;

assign detect_min[114][0] = (mid_1[927:920] < top_0[919:912]) ? 1 : 0;
assign detect_min[114][1] = (mid_1[927:920] < top_0[927:920]) ? 1 : 0;
assign detect_min[114][2] = (mid_1[927:920] < top_0[935:928]) ? 1 : 0;
assign detect_min[114][3] = (mid_1[927:920] < top_1[919:912]) ? 1 : 0;
assign detect_min[114][4] = (mid_1[927:920] < top_1[927:920]) ? 1 : 0;
assign detect_min[114][5] = (mid_1[927:920] < top_1[935:928]) ? 1 : 0;
assign detect_min[114][6] = (mid_1[927:920] < top_2[919:912]) ? 1 : 0;
assign detect_min[114][7] = (mid_1[927:920] < top_2[927:920]) ? 1 : 0;
assign detect_min[114][8] = (mid_1[927:920] < top_2[935:928]) ? 1 : 0;
assign detect_min[114][9] = (mid_1[927:920] < mid_0[919:912]) ? 1 : 0;
assign detect_min[114][10] = (mid_1[927:920] < mid_0[927:920]) ? 1 : 0;
assign detect_min[114][11] = (mid_1[927:920] < mid_0[935:928]) ? 1 : 0;
assign detect_min[114][12] = (mid_1[927:920] < mid_1[919:912]) ? 1 : 0;
assign detect_min[114][13] = (mid_1[927:920] < mid_1[935:928]) ? 1 : 0;
assign detect_min[114][14] = (mid_1[927:920] < mid_2[919:912]) ? 1 : 0;
assign detect_min[114][15] = (mid_1[927:920] < mid_2[927:920]) ? 1 : 0;
assign detect_min[114][16] = (mid_1[927:920] < mid_2[935:928]) ? 1 : 0;
assign detect_min[114][17] = (mid_1[927:920] < btm_0[919:912]) ? 1 : 0;
assign detect_min[114][18] = (mid_1[927:920] < btm_0[927:920]) ? 1 : 0;
assign detect_min[114][19] = (mid_1[927:920] < btm_0[935:928]) ? 1 : 0;
assign detect_min[114][20] = (mid_1[927:920] < btm_1[919:912]) ? 1 : 0;
assign detect_min[114][21] = (mid_1[927:920] < btm_1[927:920]) ? 1 : 0;
assign detect_min[114][22] = (mid_1[927:920] < btm_1[935:928]) ? 1 : 0;
assign detect_min[114][23] = (mid_1[927:920] < btm_2[919:912]) ? 1 : 0;
assign detect_min[114][24] = (mid_1[927:920] < btm_2[927:920]) ? 1 : 0;
assign detect_min[114][25] = (mid_1[927:920] < btm_2[935:928]) ? 1 : 0;

assign detect_min[115][0] = (mid_1[935:928] < top_0[927:920]) ? 1 : 0;
assign detect_min[115][1] = (mid_1[935:928] < top_0[935:928]) ? 1 : 0;
assign detect_min[115][2] = (mid_1[935:928] < top_0[943:936]) ? 1 : 0;
assign detect_min[115][3] = (mid_1[935:928] < top_1[927:920]) ? 1 : 0;
assign detect_min[115][4] = (mid_1[935:928] < top_1[935:928]) ? 1 : 0;
assign detect_min[115][5] = (mid_1[935:928] < top_1[943:936]) ? 1 : 0;
assign detect_min[115][6] = (mid_1[935:928] < top_2[927:920]) ? 1 : 0;
assign detect_min[115][7] = (mid_1[935:928] < top_2[935:928]) ? 1 : 0;
assign detect_min[115][8] = (mid_1[935:928] < top_2[943:936]) ? 1 : 0;
assign detect_min[115][9] = (mid_1[935:928] < mid_0[927:920]) ? 1 : 0;
assign detect_min[115][10] = (mid_1[935:928] < mid_0[935:928]) ? 1 : 0;
assign detect_min[115][11] = (mid_1[935:928] < mid_0[943:936]) ? 1 : 0;
assign detect_min[115][12] = (mid_1[935:928] < mid_1[927:920]) ? 1 : 0;
assign detect_min[115][13] = (mid_1[935:928] < mid_1[943:936]) ? 1 : 0;
assign detect_min[115][14] = (mid_1[935:928] < mid_2[927:920]) ? 1 : 0;
assign detect_min[115][15] = (mid_1[935:928] < mid_2[935:928]) ? 1 : 0;
assign detect_min[115][16] = (mid_1[935:928] < mid_2[943:936]) ? 1 : 0;
assign detect_min[115][17] = (mid_1[935:928] < btm_0[927:920]) ? 1 : 0;
assign detect_min[115][18] = (mid_1[935:928] < btm_0[935:928]) ? 1 : 0;
assign detect_min[115][19] = (mid_1[935:928] < btm_0[943:936]) ? 1 : 0;
assign detect_min[115][20] = (mid_1[935:928] < btm_1[927:920]) ? 1 : 0;
assign detect_min[115][21] = (mid_1[935:928] < btm_1[935:928]) ? 1 : 0;
assign detect_min[115][22] = (mid_1[935:928] < btm_1[943:936]) ? 1 : 0;
assign detect_min[115][23] = (mid_1[935:928] < btm_2[927:920]) ? 1 : 0;
assign detect_min[115][24] = (mid_1[935:928] < btm_2[935:928]) ? 1 : 0;
assign detect_min[115][25] = (mid_1[935:928] < btm_2[943:936]) ? 1 : 0;

assign detect_min[116][0] = (mid_1[943:936] < top_0[935:928]) ? 1 : 0;
assign detect_min[116][1] = (mid_1[943:936] < top_0[943:936]) ? 1 : 0;
assign detect_min[116][2] = (mid_1[943:936] < top_0[951:944]) ? 1 : 0;
assign detect_min[116][3] = (mid_1[943:936] < top_1[935:928]) ? 1 : 0;
assign detect_min[116][4] = (mid_1[943:936] < top_1[943:936]) ? 1 : 0;
assign detect_min[116][5] = (mid_1[943:936] < top_1[951:944]) ? 1 : 0;
assign detect_min[116][6] = (mid_1[943:936] < top_2[935:928]) ? 1 : 0;
assign detect_min[116][7] = (mid_1[943:936] < top_2[943:936]) ? 1 : 0;
assign detect_min[116][8] = (mid_1[943:936] < top_2[951:944]) ? 1 : 0;
assign detect_min[116][9] = (mid_1[943:936] < mid_0[935:928]) ? 1 : 0;
assign detect_min[116][10] = (mid_1[943:936] < mid_0[943:936]) ? 1 : 0;
assign detect_min[116][11] = (mid_1[943:936] < mid_0[951:944]) ? 1 : 0;
assign detect_min[116][12] = (mid_1[943:936] < mid_1[935:928]) ? 1 : 0;
assign detect_min[116][13] = (mid_1[943:936] < mid_1[951:944]) ? 1 : 0;
assign detect_min[116][14] = (mid_1[943:936] < mid_2[935:928]) ? 1 : 0;
assign detect_min[116][15] = (mid_1[943:936] < mid_2[943:936]) ? 1 : 0;
assign detect_min[116][16] = (mid_1[943:936] < mid_2[951:944]) ? 1 : 0;
assign detect_min[116][17] = (mid_1[943:936] < btm_0[935:928]) ? 1 : 0;
assign detect_min[116][18] = (mid_1[943:936] < btm_0[943:936]) ? 1 : 0;
assign detect_min[116][19] = (mid_1[943:936] < btm_0[951:944]) ? 1 : 0;
assign detect_min[116][20] = (mid_1[943:936] < btm_1[935:928]) ? 1 : 0;
assign detect_min[116][21] = (mid_1[943:936] < btm_1[943:936]) ? 1 : 0;
assign detect_min[116][22] = (mid_1[943:936] < btm_1[951:944]) ? 1 : 0;
assign detect_min[116][23] = (mid_1[943:936] < btm_2[935:928]) ? 1 : 0;
assign detect_min[116][24] = (mid_1[943:936] < btm_2[943:936]) ? 1 : 0;
assign detect_min[116][25] = (mid_1[943:936] < btm_2[951:944]) ? 1 : 0;

assign detect_min[117][0] = (mid_1[951:944] < top_0[943:936]) ? 1 : 0;
assign detect_min[117][1] = (mid_1[951:944] < top_0[951:944]) ? 1 : 0;
assign detect_min[117][2] = (mid_1[951:944] < top_0[959:952]) ? 1 : 0;
assign detect_min[117][3] = (mid_1[951:944] < top_1[943:936]) ? 1 : 0;
assign detect_min[117][4] = (mid_1[951:944] < top_1[951:944]) ? 1 : 0;
assign detect_min[117][5] = (mid_1[951:944] < top_1[959:952]) ? 1 : 0;
assign detect_min[117][6] = (mid_1[951:944] < top_2[943:936]) ? 1 : 0;
assign detect_min[117][7] = (mid_1[951:944] < top_2[951:944]) ? 1 : 0;
assign detect_min[117][8] = (mid_1[951:944] < top_2[959:952]) ? 1 : 0;
assign detect_min[117][9] = (mid_1[951:944] < mid_0[943:936]) ? 1 : 0;
assign detect_min[117][10] = (mid_1[951:944] < mid_0[951:944]) ? 1 : 0;
assign detect_min[117][11] = (mid_1[951:944] < mid_0[959:952]) ? 1 : 0;
assign detect_min[117][12] = (mid_1[951:944] < mid_1[943:936]) ? 1 : 0;
assign detect_min[117][13] = (mid_1[951:944] < mid_1[959:952]) ? 1 : 0;
assign detect_min[117][14] = (mid_1[951:944] < mid_2[943:936]) ? 1 : 0;
assign detect_min[117][15] = (mid_1[951:944] < mid_2[951:944]) ? 1 : 0;
assign detect_min[117][16] = (mid_1[951:944] < mid_2[959:952]) ? 1 : 0;
assign detect_min[117][17] = (mid_1[951:944] < btm_0[943:936]) ? 1 : 0;
assign detect_min[117][18] = (mid_1[951:944] < btm_0[951:944]) ? 1 : 0;
assign detect_min[117][19] = (mid_1[951:944] < btm_0[959:952]) ? 1 : 0;
assign detect_min[117][20] = (mid_1[951:944] < btm_1[943:936]) ? 1 : 0;
assign detect_min[117][21] = (mid_1[951:944] < btm_1[951:944]) ? 1 : 0;
assign detect_min[117][22] = (mid_1[951:944] < btm_1[959:952]) ? 1 : 0;
assign detect_min[117][23] = (mid_1[951:944] < btm_2[943:936]) ? 1 : 0;
assign detect_min[117][24] = (mid_1[951:944] < btm_2[951:944]) ? 1 : 0;
assign detect_min[117][25] = (mid_1[951:944] < btm_2[959:952]) ? 1 : 0;

assign detect_min[118][0] = (mid_1[959:952] < top_0[951:944]) ? 1 : 0;
assign detect_min[118][1] = (mid_1[959:952] < top_0[959:952]) ? 1 : 0;
assign detect_min[118][2] = (mid_1[959:952] < top_0[967:960]) ? 1 : 0;
assign detect_min[118][3] = (mid_1[959:952] < top_1[951:944]) ? 1 : 0;
assign detect_min[118][4] = (mid_1[959:952] < top_1[959:952]) ? 1 : 0;
assign detect_min[118][5] = (mid_1[959:952] < top_1[967:960]) ? 1 : 0;
assign detect_min[118][6] = (mid_1[959:952] < top_2[951:944]) ? 1 : 0;
assign detect_min[118][7] = (mid_1[959:952] < top_2[959:952]) ? 1 : 0;
assign detect_min[118][8] = (mid_1[959:952] < top_2[967:960]) ? 1 : 0;
assign detect_min[118][9] = (mid_1[959:952] < mid_0[951:944]) ? 1 : 0;
assign detect_min[118][10] = (mid_1[959:952] < mid_0[959:952]) ? 1 : 0;
assign detect_min[118][11] = (mid_1[959:952] < mid_0[967:960]) ? 1 : 0;
assign detect_min[118][12] = (mid_1[959:952] < mid_1[951:944]) ? 1 : 0;
assign detect_min[118][13] = (mid_1[959:952] < mid_1[967:960]) ? 1 : 0;
assign detect_min[118][14] = (mid_1[959:952] < mid_2[951:944]) ? 1 : 0;
assign detect_min[118][15] = (mid_1[959:952] < mid_2[959:952]) ? 1 : 0;
assign detect_min[118][16] = (mid_1[959:952] < mid_2[967:960]) ? 1 : 0;
assign detect_min[118][17] = (mid_1[959:952] < btm_0[951:944]) ? 1 : 0;
assign detect_min[118][18] = (mid_1[959:952] < btm_0[959:952]) ? 1 : 0;
assign detect_min[118][19] = (mid_1[959:952] < btm_0[967:960]) ? 1 : 0;
assign detect_min[118][20] = (mid_1[959:952] < btm_1[951:944]) ? 1 : 0;
assign detect_min[118][21] = (mid_1[959:952] < btm_1[959:952]) ? 1 : 0;
assign detect_min[118][22] = (mid_1[959:952] < btm_1[967:960]) ? 1 : 0;
assign detect_min[118][23] = (mid_1[959:952] < btm_2[951:944]) ? 1 : 0;
assign detect_min[118][24] = (mid_1[959:952] < btm_2[959:952]) ? 1 : 0;
assign detect_min[118][25] = (mid_1[959:952] < btm_2[967:960]) ? 1 : 0;

assign detect_min[119][0] = (mid_1[967:960] < top_0[959:952]) ? 1 : 0;
assign detect_min[119][1] = (mid_1[967:960] < top_0[967:960]) ? 1 : 0;
assign detect_min[119][2] = (mid_1[967:960] < top_0[975:968]) ? 1 : 0;
assign detect_min[119][3] = (mid_1[967:960] < top_1[959:952]) ? 1 : 0;
assign detect_min[119][4] = (mid_1[967:960] < top_1[967:960]) ? 1 : 0;
assign detect_min[119][5] = (mid_1[967:960] < top_1[975:968]) ? 1 : 0;
assign detect_min[119][6] = (mid_1[967:960] < top_2[959:952]) ? 1 : 0;
assign detect_min[119][7] = (mid_1[967:960] < top_2[967:960]) ? 1 : 0;
assign detect_min[119][8] = (mid_1[967:960] < top_2[975:968]) ? 1 : 0;
assign detect_min[119][9] = (mid_1[967:960] < mid_0[959:952]) ? 1 : 0;
assign detect_min[119][10] = (mid_1[967:960] < mid_0[967:960]) ? 1 : 0;
assign detect_min[119][11] = (mid_1[967:960] < mid_0[975:968]) ? 1 : 0;
assign detect_min[119][12] = (mid_1[967:960] < mid_1[959:952]) ? 1 : 0;
assign detect_min[119][13] = (mid_1[967:960] < mid_1[975:968]) ? 1 : 0;
assign detect_min[119][14] = (mid_1[967:960] < mid_2[959:952]) ? 1 : 0;
assign detect_min[119][15] = (mid_1[967:960] < mid_2[967:960]) ? 1 : 0;
assign detect_min[119][16] = (mid_1[967:960] < mid_2[975:968]) ? 1 : 0;
assign detect_min[119][17] = (mid_1[967:960] < btm_0[959:952]) ? 1 : 0;
assign detect_min[119][18] = (mid_1[967:960] < btm_0[967:960]) ? 1 : 0;
assign detect_min[119][19] = (mid_1[967:960] < btm_0[975:968]) ? 1 : 0;
assign detect_min[119][20] = (mid_1[967:960] < btm_1[959:952]) ? 1 : 0;
assign detect_min[119][21] = (mid_1[967:960] < btm_1[967:960]) ? 1 : 0;
assign detect_min[119][22] = (mid_1[967:960] < btm_1[975:968]) ? 1 : 0;
assign detect_min[119][23] = (mid_1[967:960] < btm_2[959:952]) ? 1 : 0;
assign detect_min[119][24] = (mid_1[967:960] < btm_2[967:960]) ? 1 : 0;
assign detect_min[119][25] = (mid_1[967:960] < btm_2[975:968]) ? 1 : 0;

assign detect_min[120][0] = (mid_1[975:968] < top_0[967:960]) ? 1 : 0;
assign detect_min[120][1] = (mid_1[975:968] < top_0[975:968]) ? 1 : 0;
assign detect_min[120][2] = (mid_1[975:968] < top_0[983:976]) ? 1 : 0;
assign detect_min[120][3] = (mid_1[975:968] < top_1[967:960]) ? 1 : 0;
assign detect_min[120][4] = (mid_1[975:968] < top_1[975:968]) ? 1 : 0;
assign detect_min[120][5] = (mid_1[975:968] < top_1[983:976]) ? 1 : 0;
assign detect_min[120][6] = (mid_1[975:968] < top_2[967:960]) ? 1 : 0;
assign detect_min[120][7] = (mid_1[975:968] < top_2[975:968]) ? 1 : 0;
assign detect_min[120][8] = (mid_1[975:968] < top_2[983:976]) ? 1 : 0;
assign detect_min[120][9] = (mid_1[975:968] < mid_0[967:960]) ? 1 : 0;
assign detect_min[120][10] = (mid_1[975:968] < mid_0[975:968]) ? 1 : 0;
assign detect_min[120][11] = (mid_1[975:968] < mid_0[983:976]) ? 1 : 0;
assign detect_min[120][12] = (mid_1[975:968] < mid_1[967:960]) ? 1 : 0;
assign detect_min[120][13] = (mid_1[975:968] < mid_1[983:976]) ? 1 : 0;
assign detect_min[120][14] = (mid_1[975:968] < mid_2[967:960]) ? 1 : 0;
assign detect_min[120][15] = (mid_1[975:968] < mid_2[975:968]) ? 1 : 0;
assign detect_min[120][16] = (mid_1[975:968] < mid_2[983:976]) ? 1 : 0;
assign detect_min[120][17] = (mid_1[975:968] < btm_0[967:960]) ? 1 : 0;
assign detect_min[120][18] = (mid_1[975:968] < btm_0[975:968]) ? 1 : 0;
assign detect_min[120][19] = (mid_1[975:968] < btm_0[983:976]) ? 1 : 0;
assign detect_min[120][20] = (mid_1[975:968] < btm_1[967:960]) ? 1 : 0;
assign detect_min[120][21] = (mid_1[975:968] < btm_1[975:968]) ? 1 : 0;
assign detect_min[120][22] = (mid_1[975:968] < btm_1[983:976]) ? 1 : 0;
assign detect_min[120][23] = (mid_1[975:968] < btm_2[967:960]) ? 1 : 0;
assign detect_min[120][24] = (mid_1[975:968] < btm_2[975:968]) ? 1 : 0;
assign detect_min[120][25] = (mid_1[975:968] < btm_2[983:976]) ? 1 : 0;

assign detect_min[121][0] = (mid_1[983:976] < top_0[975:968]) ? 1 : 0;
assign detect_min[121][1] = (mid_1[983:976] < top_0[983:976]) ? 1 : 0;
assign detect_min[121][2] = (mid_1[983:976] < top_0[991:984]) ? 1 : 0;
assign detect_min[121][3] = (mid_1[983:976] < top_1[975:968]) ? 1 : 0;
assign detect_min[121][4] = (mid_1[983:976] < top_1[983:976]) ? 1 : 0;
assign detect_min[121][5] = (mid_1[983:976] < top_1[991:984]) ? 1 : 0;
assign detect_min[121][6] = (mid_1[983:976] < top_2[975:968]) ? 1 : 0;
assign detect_min[121][7] = (mid_1[983:976] < top_2[983:976]) ? 1 : 0;
assign detect_min[121][8] = (mid_1[983:976] < top_2[991:984]) ? 1 : 0;
assign detect_min[121][9] = (mid_1[983:976] < mid_0[975:968]) ? 1 : 0;
assign detect_min[121][10] = (mid_1[983:976] < mid_0[983:976]) ? 1 : 0;
assign detect_min[121][11] = (mid_1[983:976] < mid_0[991:984]) ? 1 : 0;
assign detect_min[121][12] = (mid_1[983:976] < mid_1[975:968]) ? 1 : 0;
assign detect_min[121][13] = (mid_1[983:976] < mid_1[991:984]) ? 1 : 0;
assign detect_min[121][14] = (mid_1[983:976] < mid_2[975:968]) ? 1 : 0;
assign detect_min[121][15] = (mid_1[983:976] < mid_2[983:976]) ? 1 : 0;
assign detect_min[121][16] = (mid_1[983:976] < mid_2[991:984]) ? 1 : 0;
assign detect_min[121][17] = (mid_1[983:976] < btm_0[975:968]) ? 1 : 0;
assign detect_min[121][18] = (mid_1[983:976] < btm_0[983:976]) ? 1 : 0;
assign detect_min[121][19] = (mid_1[983:976] < btm_0[991:984]) ? 1 : 0;
assign detect_min[121][20] = (mid_1[983:976] < btm_1[975:968]) ? 1 : 0;
assign detect_min[121][21] = (mid_1[983:976] < btm_1[983:976]) ? 1 : 0;
assign detect_min[121][22] = (mid_1[983:976] < btm_1[991:984]) ? 1 : 0;
assign detect_min[121][23] = (mid_1[983:976] < btm_2[975:968]) ? 1 : 0;
assign detect_min[121][24] = (mid_1[983:976] < btm_2[983:976]) ? 1 : 0;
assign detect_min[121][25] = (mid_1[983:976] < btm_2[991:984]) ? 1 : 0;

assign detect_min[122][0] = (mid_1[991:984] < top_0[983:976]) ? 1 : 0;
assign detect_min[122][1] = (mid_1[991:984] < top_0[991:984]) ? 1 : 0;
assign detect_min[122][2] = (mid_1[991:984] < top_0[999:992]) ? 1 : 0;
assign detect_min[122][3] = (mid_1[991:984] < top_1[983:976]) ? 1 : 0;
assign detect_min[122][4] = (mid_1[991:984] < top_1[991:984]) ? 1 : 0;
assign detect_min[122][5] = (mid_1[991:984] < top_1[999:992]) ? 1 : 0;
assign detect_min[122][6] = (mid_1[991:984] < top_2[983:976]) ? 1 : 0;
assign detect_min[122][7] = (mid_1[991:984] < top_2[991:984]) ? 1 : 0;
assign detect_min[122][8] = (mid_1[991:984] < top_2[999:992]) ? 1 : 0;
assign detect_min[122][9] = (mid_1[991:984] < mid_0[983:976]) ? 1 : 0;
assign detect_min[122][10] = (mid_1[991:984] < mid_0[991:984]) ? 1 : 0;
assign detect_min[122][11] = (mid_1[991:984] < mid_0[999:992]) ? 1 : 0;
assign detect_min[122][12] = (mid_1[991:984] < mid_1[983:976]) ? 1 : 0;
assign detect_min[122][13] = (mid_1[991:984] < mid_1[999:992]) ? 1 : 0;
assign detect_min[122][14] = (mid_1[991:984] < mid_2[983:976]) ? 1 : 0;
assign detect_min[122][15] = (mid_1[991:984] < mid_2[991:984]) ? 1 : 0;
assign detect_min[122][16] = (mid_1[991:984] < mid_2[999:992]) ? 1 : 0;
assign detect_min[122][17] = (mid_1[991:984] < btm_0[983:976]) ? 1 : 0;
assign detect_min[122][18] = (mid_1[991:984] < btm_0[991:984]) ? 1 : 0;
assign detect_min[122][19] = (mid_1[991:984] < btm_0[999:992]) ? 1 : 0;
assign detect_min[122][20] = (mid_1[991:984] < btm_1[983:976]) ? 1 : 0;
assign detect_min[122][21] = (mid_1[991:984] < btm_1[991:984]) ? 1 : 0;
assign detect_min[122][22] = (mid_1[991:984] < btm_1[999:992]) ? 1 : 0;
assign detect_min[122][23] = (mid_1[991:984] < btm_2[983:976]) ? 1 : 0;
assign detect_min[122][24] = (mid_1[991:984] < btm_2[991:984]) ? 1 : 0;
assign detect_min[122][25] = (mid_1[991:984] < btm_2[999:992]) ? 1 : 0;

assign detect_min[123][0] = (mid_1[999:992] < top_0[991:984]) ? 1 : 0;
assign detect_min[123][1] = (mid_1[999:992] < top_0[999:992]) ? 1 : 0;
assign detect_min[123][2] = (mid_1[999:992] < top_0[1007:1000]) ? 1 : 0;
assign detect_min[123][3] = (mid_1[999:992] < top_1[991:984]) ? 1 : 0;
assign detect_min[123][4] = (mid_1[999:992] < top_1[999:992]) ? 1 : 0;
assign detect_min[123][5] = (mid_1[999:992] < top_1[1007:1000]) ? 1 : 0;
assign detect_min[123][6] = (mid_1[999:992] < top_2[991:984]) ? 1 : 0;
assign detect_min[123][7] = (mid_1[999:992] < top_2[999:992]) ? 1 : 0;
assign detect_min[123][8] = (mid_1[999:992] < top_2[1007:1000]) ? 1 : 0;
assign detect_min[123][9] = (mid_1[999:992] < mid_0[991:984]) ? 1 : 0;
assign detect_min[123][10] = (mid_1[999:992] < mid_0[999:992]) ? 1 : 0;
assign detect_min[123][11] = (mid_1[999:992] < mid_0[1007:1000]) ? 1 : 0;
assign detect_min[123][12] = (mid_1[999:992] < mid_1[991:984]) ? 1 : 0;
assign detect_min[123][13] = (mid_1[999:992] < mid_1[1007:1000]) ? 1 : 0;
assign detect_min[123][14] = (mid_1[999:992] < mid_2[991:984]) ? 1 : 0;
assign detect_min[123][15] = (mid_1[999:992] < mid_2[999:992]) ? 1 : 0;
assign detect_min[123][16] = (mid_1[999:992] < mid_2[1007:1000]) ? 1 : 0;
assign detect_min[123][17] = (mid_1[999:992] < btm_0[991:984]) ? 1 : 0;
assign detect_min[123][18] = (mid_1[999:992] < btm_0[999:992]) ? 1 : 0;
assign detect_min[123][19] = (mid_1[999:992] < btm_0[1007:1000]) ? 1 : 0;
assign detect_min[123][20] = (mid_1[999:992] < btm_1[991:984]) ? 1 : 0;
assign detect_min[123][21] = (mid_1[999:992] < btm_1[999:992]) ? 1 : 0;
assign detect_min[123][22] = (mid_1[999:992] < btm_1[1007:1000]) ? 1 : 0;
assign detect_min[123][23] = (mid_1[999:992] < btm_2[991:984]) ? 1 : 0;
assign detect_min[123][24] = (mid_1[999:992] < btm_2[999:992]) ? 1 : 0;
assign detect_min[123][25] = (mid_1[999:992] < btm_2[1007:1000]) ? 1 : 0;

assign detect_min[124][0] = (mid_1[1007:1000] < top_0[999:992]) ? 1 : 0;
assign detect_min[124][1] = (mid_1[1007:1000] < top_0[1007:1000]) ? 1 : 0;
assign detect_min[124][2] = (mid_1[1007:1000] < top_0[1015:1008]) ? 1 : 0;
assign detect_min[124][3] = (mid_1[1007:1000] < top_1[999:992]) ? 1 : 0;
assign detect_min[124][4] = (mid_1[1007:1000] < top_1[1007:1000]) ? 1 : 0;
assign detect_min[124][5] = (mid_1[1007:1000] < top_1[1015:1008]) ? 1 : 0;
assign detect_min[124][6] = (mid_1[1007:1000] < top_2[999:992]) ? 1 : 0;
assign detect_min[124][7] = (mid_1[1007:1000] < top_2[1007:1000]) ? 1 : 0;
assign detect_min[124][8] = (mid_1[1007:1000] < top_2[1015:1008]) ? 1 : 0;
assign detect_min[124][9] = (mid_1[1007:1000] < mid_0[999:992]) ? 1 : 0;
assign detect_min[124][10] = (mid_1[1007:1000] < mid_0[1007:1000]) ? 1 : 0;
assign detect_min[124][11] = (mid_1[1007:1000] < mid_0[1015:1008]) ? 1 : 0;
assign detect_min[124][12] = (mid_1[1007:1000] < mid_1[999:992]) ? 1 : 0;
assign detect_min[124][13] = (mid_1[1007:1000] < mid_1[1015:1008]) ? 1 : 0;
assign detect_min[124][14] = (mid_1[1007:1000] < mid_2[999:992]) ? 1 : 0;
assign detect_min[124][15] = (mid_1[1007:1000] < mid_2[1007:1000]) ? 1 : 0;
assign detect_min[124][16] = (mid_1[1007:1000] < mid_2[1015:1008]) ? 1 : 0;
assign detect_min[124][17] = (mid_1[1007:1000] < btm_0[999:992]) ? 1 : 0;
assign detect_min[124][18] = (mid_1[1007:1000] < btm_0[1007:1000]) ? 1 : 0;
assign detect_min[124][19] = (mid_1[1007:1000] < btm_0[1015:1008]) ? 1 : 0;
assign detect_min[124][20] = (mid_1[1007:1000] < btm_1[999:992]) ? 1 : 0;
assign detect_min[124][21] = (mid_1[1007:1000] < btm_1[1007:1000]) ? 1 : 0;
assign detect_min[124][22] = (mid_1[1007:1000] < btm_1[1015:1008]) ? 1 : 0;
assign detect_min[124][23] = (mid_1[1007:1000] < btm_2[999:992]) ? 1 : 0;
assign detect_min[124][24] = (mid_1[1007:1000] < btm_2[1007:1000]) ? 1 : 0;
assign detect_min[124][25] = (mid_1[1007:1000] < btm_2[1015:1008]) ? 1 : 0;

assign detect_min[125][0] = (mid_1[1015:1008] < top_0[1007:1000]) ? 1 : 0;
assign detect_min[125][1] = (mid_1[1015:1008] < top_0[1015:1008]) ? 1 : 0;
assign detect_min[125][2] = (mid_1[1015:1008] < top_0[1023:1016]) ? 1 : 0;
assign detect_min[125][3] = (mid_1[1015:1008] < top_1[1007:1000]) ? 1 : 0;
assign detect_min[125][4] = (mid_1[1015:1008] < top_1[1015:1008]) ? 1 : 0;
assign detect_min[125][5] = (mid_1[1015:1008] < top_1[1023:1016]) ? 1 : 0;
assign detect_min[125][6] = (mid_1[1015:1008] < top_2[1007:1000]) ? 1 : 0;
assign detect_min[125][7] = (mid_1[1015:1008] < top_2[1015:1008]) ? 1 : 0;
assign detect_min[125][8] = (mid_1[1015:1008] < top_2[1023:1016]) ? 1 : 0;
assign detect_min[125][9] = (mid_1[1015:1008] < mid_0[1007:1000]) ? 1 : 0;
assign detect_min[125][10] = (mid_1[1015:1008] < mid_0[1015:1008]) ? 1 : 0;
assign detect_min[125][11] = (mid_1[1015:1008] < mid_0[1023:1016]) ? 1 : 0;
assign detect_min[125][12] = (mid_1[1015:1008] < mid_1[1007:1000]) ? 1 : 0;
assign detect_min[125][13] = (mid_1[1015:1008] < mid_1[1023:1016]) ? 1 : 0;
assign detect_min[125][14] = (mid_1[1015:1008] < mid_2[1007:1000]) ? 1 : 0;
assign detect_min[125][15] = (mid_1[1015:1008] < mid_2[1015:1008]) ? 1 : 0;
assign detect_min[125][16] = (mid_1[1015:1008] < mid_2[1023:1016]) ? 1 : 0;
assign detect_min[125][17] = (mid_1[1015:1008] < btm_0[1007:1000]) ? 1 : 0;
assign detect_min[125][18] = (mid_1[1015:1008] < btm_0[1015:1008]) ? 1 : 0;
assign detect_min[125][19] = (mid_1[1015:1008] < btm_0[1023:1016]) ? 1 : 0;
assign detect_min[125][20] = (mid_1[1015:1008] < btm_1[1007:1000]) ? 1 : 0;
assign detect_min[125][21] = (mid_1[1015:1008] < btm_1[1015:1008]) ? 1 : 0;
assign detect_min[125][22] = (mid_1[1015:1008] < btm_1[1023:1016]) ? 1 : 0;
assign detect_min[125][23] = (mid_1[1015:1008] < btm_2[1007:1000]) ? 1 : 0;
assign detect_min[125][24] = (mid_1[1015:1008] < btm_2[1015:1008]) ? 1 : 0;
assign detect_min[125][25] = (mid_1[1015:1008] < btm_2[1023:1016]) ? 1 : 0;

assign detect_min[126][0] = (mid_1[1023:1016] < top_0[1015:1008]) ? 1 : 0;
assign detect_min[126][1] = (mid_1[1023:1016] < top_0[1023:1016]) ? 1 : 0;
assign detect_min[126][2] = (mid_1[1023:1016] < top_0[1031:1024]) ? 1 : 0;
assign detect_min[126][3] = (mid_1[1023:1016] < top_1[1015:1008]) ? 1 : 0;
assign detect_min[126][4] = (mid_1[1023:1016] < top_1[1023:1016]) ? 1 : 0;
assign detect_min[126][5] = (mid_1[1023:1016] < top_1[1031:1024]) ? 1 : 0;
assign detect_min[126][6] = (mid_1[1023:1016] < top_2[1015:1008]) ? 1 : 0;
assign detect_min[126][7] = (mid_1[1023:1016] < top_2[1023:1016]) ? 1 : 0;
assign detect_min[126][8] = (mid_1[1023:1016] < top_2[1031:1024]) ? 1 : 0;
assign detect_min[126][9] = (mid_1[1023:1016] < mid_0[1015:1008]) ? 1 : 0;
assign detect_min[126][10] = (mid_1[1023:1016] < mid_0[1023:1016]) ? 1 : 0;
assign detect_min[126][11] = (mid_1[1023:1016] < mid_0[1031:1024]) ? 1 : 0;
assign detect_min[126][12] = (mid_1[1023:1016] < mid_1[1015:1008]) ? 1 : 0;
assign detect_min[126][13] = (mid_1[1023:1016] < mid_1[1031:1024]) ? 1 : 0;
assign detect_min[126][14] = (mid_1[1023:1016] < mid_2[1015:1008]) ? 1 : 0;
assign detect_min[126][15] = (mid_1[1023:1016] < mid_2[1023:1016]) ? 1 : 0;
assign detect_min[126][16] = (mid_1[1023:1016] < mid_2[1031:1024]) ? 1 : 0;
assign detect_min[126][17] = (mid_1[1023:1016] < btm_0[1015:1008]) ? 1 : 0;
assign detect_min[126][18] = (mid_1[1023:1016] < btm_0[1023:1016]) ? 1 : 0;
assign detect_min[126][19] = (mid_1[1023:1016] < btm_0[1031:1024]) ? 1 : 0;
assign detect_min[126][20] = (mid_1[1023:1016] < btm_1[1015:1008]) ? 1 : 0;
assign detect_min[126][21] = (mid_1[1023:1016] < btm_1[1023:1016]) ? 1 : 0;
assign detect_min[126][22] = (mid_1[1023:1016] < btm_1[1031:1024]) ? 1 : 0;
assign detect_min[126][23] = (mid_1[1023:1016] < btm_2[1015:1008]) ? 1 : 0;
assign detect_min[126][24] = (mid_1[1023:1016] < btm_2[1023:1016]) ? 1 : 0;
assign detect_min[126][25] = (mid_1[1023:1016] < btm_2[1031:1024]) ? 1 : 0;

assign detect_min[127][0] = (mid_1[1031:1024] < top_0[1023:1016]) ? 1 : 0;
assign detect_min[127][1] = (mid_1[1031:1024] < top_0[1031:1024]) ? 1 : 0;
assign detect_min[127][2] = (mid_1[1031:1024] < top_0[1039:1032]) ? 1 : 0;
assign detect_min[127][3] = (mid_1[1031:1024] < top_1[1023:1016]) ? 1 : 0;
assign detect_min[127][4] = (mid_1[1031:1024] < top_1[1031:1024]) ? 1 : 0;
assign detect_min[127][5] = (mid_1[1031:1024] < top_1[1039:1032]) ? 1 : 0;
assign detect_min[127][6] = (mid_1[1031:1024] < top_2[1023:1016]) ? 1 : 0;
assign detect_min[127][7] = (mid_1[1031:1024] < top_2[1031:1024]) ? 1 : 0;
assign detect_min[127][8] = (mid_1[1031:1024] < top_2[1039:1032]) ? 1 : 0;
assign detect_min[127][9] = (mid_1[1031:1024] < mid_0[1023:1016]) ? 1 : 0;
assign detect_min[127][10] = (mid_1[1031:1024] < mid_0[1031:1024]) ? 1 : 0;
assign detect_min[127][11] = (mid_1[1031:1024] < mid_0[1039:1032]) ? 1 : 0;
assign detect_min[127][12] = (mid_1[1031:1024] < mid_1[1023:1016]) ? 1 : 0;
assign detect_min[127][13] = (mid_1[1031:1024] < mid_1[1039:1032]) ? 1 : 0;
assign detect_min[127][14] = (mid_1[1031:1024] < mid_2[1023:1016]) ? 1 : 0;
assign detect_min[127][15] = (mid_1[1031:1024] < mid_2[1031:1024]) ? 1 : 0;
assign detect_min[127][16] = (mid_1[1031:1024] < mid_2[1039:1032]) ? 1 : 0;
assign detect_min[127][17] = (mid_1[1031:1024] < btm_0[1023:1016]) ? 1 : 0;
assign detect_min[127][18] = (mid_1[1031:1024] < btm_0[1031:1024]) ? 1 : 0;
assign detect_min[127][19] = (mid_1[1031:1024] < btm_0[1039:1032]) ? 1 : 0;
assign detect_min[127][20] = (mid_1[1031:1024] < btm_1[1023:1016]) ? 1 : 0;
assign detect_min[127][21] = (mid_1[1031:1024] < btm_1[1031:1024]) ? 1 : 0;
assign detect_min[127][22] = (mid_1[1031:1024] < btm_1[1039:1032]) ? 1 : 0;
assign detect_min[127][23] = (mid_1[1031:1024] < btm_2[1023:1016]) ? 1 : 0;
assign detect_min[127][24] = (mid_1[1031:1024] < btm_2[1031:1024]) ? 1 : 0;
assign detect_min[127][25] = (mid_1[1031:1024] < btm_2[1039:1032]) ? 1 : 0;

assign detect_min[128][0] = (mid_1[1039:1032] < top_0[1031:1024]) ? 1 : 0;
assign detect_min[128][1] = (mid_1[1039:1032] < top_0[1039:1032]) ? 1 : 0;
assign detect_min[128][2] = (mid_1[1039:1032] < top_0[1047:1040]) ? 1 : 0;
assign detect_min[128][3] = (mid_1[1039:1032] < top_1[1031:1024]) ? 1 : 0;
assign detect_min[128][4] = (mid_1[1039:1032] < top_1[1039:1032]) ? 1 : 0;
assign detect_min[128][5] = (mid_1[1039:1032] < top_1[1047:1040]) ? 1 : 0;
assign detect_min[128][6] = (mid_1[1039:1032] < top_2[1031:1024]) ? 1 : 0;
assign detect_min[128][7] = (mid_1[1039:1032] < top_2[1039:1032]) ? 1 : 0;
assign detect_min[128][8] = (mid_1[1039:1032] < top_2[1047:1040]) ? 1 : 0;
assign detect_min[128][9] = (mid_1[1039:1032] < mid_0[1031:1024]) ? 1 : 0;
assign detect_min[128][10] = (mid_1[1039:1032] < mid_0[1039:1032]) ? 1 : 0;
assign detect_min[128][11] = (mid_1[1039:1032] < mid_0[1047:1040]) ? 1 : 0;
assign detect_min[128][12] = (mid_1[1039:1032] < mid_1[1031:1024]) ? 1 : 0;
assign detect_min[128][13] = (mid_1[1039:1032] < mid_1[1047:1040]) ? 1 : 0;
assign detect_min[128][14] = (mid_1[1039:1032] < mid_2[1031:1024]) ? 1 : 0;
assign detect_min[128][15] = (mid_1[1039:1032] < mid_2[1039:1032]) ? 1 : 0;
assign detect_min[128][16] = (mid_1[1039:1032] < mid_2[1047:1040]) ? 1 : 0;
assign detect_min[128][17] = (mid_1[1039:1032] < btm_0[1031:1024]) ? 1 : 0;
assign detect_min[128][18] = (mid_1[1039:1032] < btm_0[1039:1032]) ? 1 : 0;
assign detect_min[128][19] = (mid_1[1039:1032] < btm_0[1047:1040]) ? 1 : 0;
assign detect_min[128][20] = (mid_1[1039:1032] < btm_1[1031:1024]) ? 1 : 0;
assign detect_min[128][21] = (mid_1[1039:1032] < btm_1[1039:1032]) ? 1 : 0;
assign detect_min[128][22] = (mid_1[1039:1032] < btm_1[1047:1040]) ? 1 : 0;
assign detect_min[128][23] = (mid_1[1039:1032] < btm_2[1031:1024]) ? 1 : 0;
assign detect_min[128][24] = (mid_1[1039:1032] < btm_2[1039:1032]) ? 1 : 0;
assign detect_min[128][25] = (mid_1[1039:1032] < btm_2[1047:1040]) ? 1 : 0;

assign detect_min[129][0] = (mid_1[1047:1040] < top_0[1039:1032]) ? 1 : 0;
assign detect_min[129][1] = (mid_1[1047:1040] < top_0[1047:1040]) ? 1 : 0;
assign detect_min[129][2] = (mid_1[1047:1040] < top_0[1055:1048]) ? 1 : 0;
assign detect_min[129][3] = (mid_1[1047:1040] < top_1[1039:1032]) ? 1 : 0;
assign detect_min[129][4] = (mid_1[1047:1040] < top_1[1047:1040]) ? 1 : 0;
assign detect_min[129][5] = (mid_1[1047:1040] < top_1[1055:1048]) ? 1 : 0;
assign detect_min[129][6] = (mid_1[1047:1040] < top_2[1039:1032]) ? 1 : 0;
assign detect_min[129][7] = (mid_1[1047:1040] < top_2[1047:1040]) ? 1 : 0;
assign detect_min[129][8] = (mid_1[1047:1040] < top_2[1055:1048]) ? 1 : 0;
assign detect_min[129][9] = (mid_1[1047:1040] < mid_0[1039:1032]) ? 1 : 0;
assign detect_min[129][10] = (mid_1[1047:1040] < mid_0[1047:1040]) ? 1 : 0;
assign detect_min[129][11] = (mid_1[1047:1040] < mid_0[1055:1048]) ? 1 : 0;
assign detect_min[129][12] = (mid_1[1047:1040] < mid_1[1039:1032]) ? 1 : 0;
assign detect_min[129][13] = (mid_1[1047:1040] < mid_1[1055:1048]) ? 1 : 0;
assign detect_min[129][14] = (mid_1[1047:1040] < mid_2[1039:1032]) ? 1 : 0;
assign detect_min[129][15] = (mid_1[1047:1040] < mid_2[1047:1040]) ? 1 : 0;
assign detect_min[129][16] = (mid_1[1047:1040] < mid_2[1055:1048]) ? 1 : 0;
assign detect_min[129][17] = (mid_1[1047:1040] < btm_0[1039:1032]) ? 1 : 0;
assign detect_min[129][18] = (mid_1[1047:1040] < btm_0[1047:1040]) ? 1 : 0;
assign detect_min[129][19] = (mid_1[1047:1040] < btm_0[1055:1048]) ? 1 : 0;
assign detect_min[129][20] = (mid_1[1047:1040] < btm_1[1039:1032]) ? 1 : 0;
assign detect_min[129][21] = (mid_1[1047:1040] < btm_1[1047:1040]) ? 1 : 0;
assign detect_min[129][22] = (mid_1[1047:1040] < btm_1[1055:1048]) ? 1 : 0;
assign detect_min[129][23] = (mid_1[1047:1040] < btm_2[1039:1032]) ? 1 : 0;
assign detect_min[129][24] = (mid_1[1047:1040] < btm_2[1047:1040]) ? 1 : 0;
assign detect_min[129][25] = (mid_1[1047:1040] < btm_2[1055:1048]) ? 1 : 0;

assign detect_min[130][0] = (mid_1[1055:1048] < top_0[1047:1040]) ? 1 : 0;
assign detect_min[130][1] = (mid_1[1055:1048] < top_0[1055:1048]) ? 1 : 0;
assign detect_min[130][2] = (mid_1[1055:1048] < top_0[1063:1056]) ? 1 : 0;
assign detect_min[130][3] = (mid_1[1055:1048] < top_1[1047:1040]) ? 1 : 0;
assign detect_min[130][4] = (mid_1[1055:1048] < top_1[1055:1048]) ? 1 : 0;
assign detect_min[130][5] = (mid_1[1055:1048] < top_1[1063:1056]) ? 1 : 0;
assign detect_min[130][6] = (mid_1[1055:1048] < top_2[1047:1040]) ? 1 : 0;
assign detect_min[130][7] = (mid_1[1055:1048] < top_2[1055:1048]) ? 1 : 0;
assign detect_min[130][8] = (mid_1[1055:1048] < top_2[1063:1056]) ? 1 : 0;
assign detect_min[130][9] = (mid_1[1055:1048] < mid_0[1047:1040]) ? 1 : 0;
assign detect_min[130][10] = (mid_1[1055:1048] < mid_0[1055:1048]) ? 1 : 0;
assign detect_min[130][11] = (mid_1[1055:1048] < mid_0[1063:1056]) ? 1 : 0;
assign detect_min[130][12] = (mid_1[1055:1048] < mid_1[1047:1040]) ? 1 : 0;
assign detect_min[130][13] = (mid_1[1055:1048] < mid_1[1063:1056]) ? 1 : 0;
assign detect_min[130][14] = (mid_1[1055:1048] < mid_2[1047:1040]) ? 1 : 0;
assign detect_min[130][15] = (mid_1[1055:1048] < mid_2[1055:1048]) ? 1 : 0;
assign detect_min[130][16] = (mid_1[1055:1048] < mid_2[1063:1056]) ? 1 : 0;
assign detect_min[130][17] = (mid_1[1055:1048] < btm_0[1047:1040]) ? 1 : 0;
assign detect_min[130][18] = (mid_1[1055:1048] < btm_0[1055:1048]) ? 1 : 0;
assign detect_min[130][19] = (mid_1[1055:1048] < btm_0[1063:1056]) ? 1 : 0;
assign detect_min[130][20] = (mid_1[1055:1048] < btm_1[1047:1040]) ? 1 : 0;
assign detect_min[130][21] = (mid_1[1055:1048] < btm_1[1055:1048]) ? 1 : 0;
assign detect_min[130][22] = (mid_1[1055:1048] < btm_1[1063:1056]) ? 1 : 0;
assign detect_min[130][23] = (mid_1[1055:1048] < btm_2[1047:1040]) ? 1 : 0;
assign detect_min[130][24] = (mid_1[1055:1048] < btm_2[1055:1048]) ? 1 : 0;
assign detect_min[130][25] = (mid_1[1055:1048] < btm_2[1063:1056]) ? 1 : 0;

assign detect_min[131][0] = (mid_1[1063:1056] < top_0[1055:1048]) ? 1 : 0;
assign detect_min[131][1] = (mid_1[1063:1056] < top_0[1063:1056]) ? 1 : 0;
assign detect_min[131][2] = (mid_1[1063:1056] < top_0[1071:1064]) ? 1 : 0;
assign detect_min[131][3] = (mid_1[1063:1056] < top_1[1055:1048]) ? 1 : 0;
assign detect_min[131][4] = (mid_1[1063:1056] < top_1[1063:1056]) ? 1 : 0;
assign detect_min[131][5] = (mid_1[1063:1056] < top_1[1071:1064]) ? 1 : 0;
assign detect_min[131][6] = (mid_1[1063:1056] < top_2[1055:1048]) ? 1 : 0;
assign detect_min[131][7] = (mid_1[1063:1056] < top_2[1063:1056]) ? 1 : 0;
assign detect_min[131][8] = (mid_1[1063:1056] < top_2[1071:1064]) ? 1 : 0;
assign detect_min[131][9] = (mid_1[1063:1056] < mid_0[1055:1048]) ? 1 : 0;
assign detect_min[131][10] = (mid_1[1063:1056] < mid_0[1063:1056]) ? 1 : 0;
assign detect_min[131][11] = (mid_1[1063:1056] < mid_0[1071:1064]) ? 1 : 0;
assign detect_min[131][12] = (mid_1[1063:1056] < mid_1[1055:1048]) ? 1 : 0;
assign detect_min[131][13] = (mid_1[1063:1056] < mid_1[1071:1064]) ? 1 : 0;
assign detect_min[131][14] = (mid_1[1063:1056] < mid_2[1055:1048]) ? 1 : 0;
assign detect_min[131][15] = (mid_1[1063:1056] < mid_2[1063:1056]) ? 1 : 0;
assign detect_min[131][16] = (mid_1[1063:1056] < mid_2[1071:1064]) ? 1 : 0;
assign detect_min[131][17] = (mid_1[1063:1056] < btm_0[1055:1048]) ? 1 : 0;
assign detect_min[131][18] = (mid_1[1063:1056] < btm_0[1063:1056]) ? 1 : 0;
assign detect_min[131][19] = (mid_1[1063:1056] < btm_0[1071:1064]) ? 1 : 0;
assign detect_min[131][20] = (mid_1[1063:1056] < btm_1[1055:1048]) ? 1 : 0;
assign detect_min[131][21] = (mid_1[1063:1056] < btm_1[1063:1056]) ? 1 : 0;
assign detect_min[131][22] = (mid_1[1063:1056] < btm_1[1071:1064]) ? 1 : 0;
assign detect_min[131][23] = (mid_1[1063:1056] < btm_2[1055:1048]) ? 1 : 0;
assign detect_min[131][24] = (mid_1[1063:1056] < btm_2[1063:1056]) ? 1 : 0;
assign detect_min[131][25] = (mid_1[1063:1056] < btm_2[1071:1064]) ? 1 : 0;

assign detect_min[132][0] = (mid_1[1071:1064] < top_0[1063:1056]) ? 1 : 0;
assign detect_min[132][1] = (mid_1[1071:1064] < top_0[1071:1064]) ? 1 : 0;
assign detect_min[132][2] = (mid_1[1071:1064] < top_0[1079:1072]) ? 1 : 0;
assign detect_min[132][3] = (mid_1[1071:1064] < top_1[1063:1056]) ? 1 : 0;
assign detect_min[132][4] = (mid_1[1071:1064] < top_1[1071:1064]) ? 1 : 0;
assign detect_min[132][5] = (mid_1[1071:1064] < top_1[1079:1072]) ? 1 : 0;
assign detect_min[132][6] = (mid_1[1071:1064] < top_2[1063:1056]) ? 1 : 0;
assign detect_min[132][7] = (mid_1[1071:1064] < top_2[1071:1064]) ? 1 : 0;
assign detect_min[132][8] = (mid_1[1071:1064] < top_2[1079:1072]) ? 1 : 0;
assign detect_min[132][9] = (mid_1[1071:1064] < mid_0[1063:1056]) ? 1 : 0;
assign detect_min[132][10] = (mid_1[1071:1064] < mid_0[1071:1064]) ? 1 : 0;
assign detect_min[132][11] = (mid_1[1071:1064] < mid_0[1079:1072]) ? 1 : 0;
assign detect_min[132][12] = (mid_1[1071:1064] < mid_1[1063:1056]) ? 1 : 0;
assign detect_min[132][13] = (mid_1[1071:1064] < mid_1[1079:1072]) ? 1 : 0;
assign detect_min[132][14] = (mid_1[1071:1064] < mid_2[1063:1056]) ? 1 : 0;
assign detect_min[132][15] = (mid_1[1071:1064] < mid_2[1071:1064]) ? 1 : 0;
assign detect_min[132][16] = (mid_1[1071:1064] < mid_2[1079:1072]) ? 1 : 0;
assign detect_min[132][17] = (mid_1[1071:1064] < btm_0[1063:1056]) ? 1 : 0;
assign detect_min[132][18] = (mid_1[1071:1064] < btm_0[1071:1064]) ? 1 : 0;
assign detect_min[132][19] = (mid_1[1071:1064] < btm_0[1079:1072]) ? 1 : 0;
assign detect_min[132][20] = (mid_1[1071:1064] < btm_1[1063:1056]) ? 1 : 0;
assign detect_min[132][21] = (mid_1[1071:1064] < btm_1[1071:1064]) ? 1 : 0;
assign detect_min[132][22] = (mid_1[1071:1064] < btm_1[1079:1072]) ? 1 : 0;
assign detect_min[132][23] = (mid_1[1071:1064] < btm_2[1063:1056]) ? 1 : 0;
assign detect_min[132][24] = (mid_1[1071:1064] < btm_2[1071:1064]) ? 1 : 0;
assign detect_min[132][25] = (mid_1[1071:1064] < btm_2[1079:1072]) ? 1 : 0;

assign detect_min[133][0] = (mid_1[1079:1072] < top_0[1071:1064]) ? 1 : 0;
assign detect_min[133][1] = (mid_1[1079:1072] < top_0[1079:1072]) ? 1 : 0;
assign detect_min[133][2] = (mid_1[1079:1072] < top_0[1087:1080]) ? 1 : 0;
assign detect_min[133][3] = (mid_1[1079:1072] < top_1[1071:1064]) ? 1 : 0;
assign detect_min[133][4] = (mid_1[1079:1072] < top_1[1079:1072]) ? 1 : 0;
assign detect_min[133][5] = (mid_1[1079:1072] < top_1[1087:1080]) ? 1 : 0;
assign detect_min[133][6] = (mid_1[1079:1072] < top_2[1071:1064]) ? 1 : 0;
assign detect_min[133][7] = (mid_1[1079:1072] < top_2[1079:1072]) ? 1 : 0;
assign detect_min[133][8] = (mid_1[1079:1072] < top_2[1087:1080]) ? 1 : 0;
assign detect_min[133][9] = (mid_1[1079:1072] < mid_0[1071:1064]) ? 1 : 0;
assign detect_min[133][10] = (mid_1[1079:1072] < mid_0[1079:1072]) ? 1 : 0;
assign detect_min[133][11] = (mid_1[1079:1072] < mid_0[1087:1080]) ? 1 : 0;
assign detect_min[133][12] = (mid_1[1079:1072] < mid_1[1071:1064]) ? 1 : 0;
assign detect_min[133][13] = (mid_1[1079:1072] < mid_1[1087:1080]) ? 1 : 0;
assign detect_min[133][14] = (mid_1[1079:1072] < mid_2[1071:1064]) ? 1 : 0;
assign detect_min[133][15] = (mid_1[1079:1072] < mid_2[1079:1072]) ? 1 : 0;
assign detect_min[133][16] = (mid_1[1079:1072] < mid_2[1087:1080]) ? 1 : 0;
assign detect_min[133][17] = (mid_1[1079:1072] < btm_0[1071:1064]) ? 1 : 0;
assign detect_min[133][18] = (mid_1[1079:1072] < btm_0[1079:1072]) ? 1 : 0;
assign detect_min[133][19] = (mid_1[1079:1072] < btm_0[1087:1080]) ? 1 : 0;
assign detect_min[133][20] = (mid_1[1079:1072] < btm_1[1071:1064]) ? 1 : 0;
assign detect_min[133][21] = (mid_1[1079:1072] < btm_1[1079:1072]) ? 1 : 0;
assign detect_min[133][22] = (mid_1[1079:1072] < btm_1[1087:1080]) ? 1 : 0;
assign detect_min[133][23] = (mid_1[1079:1072] < btm_2[1071:1064]) ? 1 : 0;
assign detect_min[133][24] = (mid_1[1079:1072] < btm_2[1079:1072]) ? 1 : 0;
assign detect_min[133][25] = (mid_1[1079:1072] < btm_2[1087:1080]) ? 1 : 0;

assign detect_min[134][0] = (mid_1[1087:1080] < top_0[1079:1072]) ? 1 : 0;
assign detect_min[134][1] = (mid_1[1087:1080] < top_0[1087:1080]) ? 1 : 0;
assign detect_min[134][2] = (mid_1[1087:1080] < top_0[1095:1088]) ? 1 : 0;
assign detect_min[134][3] = (mid_1[1087:1080] < top_1[1079:1072]) ? 1 : 0;
assign detect_min[134][4] = (mid_1[1087:1080] < top_1[1087:1080]) ? 1 : 0;
assign detect_min[134][5] = (mid_1[1087:1080] < top_1[1095:1088]) ? 1 : 0;
assign detect_min[134][6] = (mid_1[1087:1080] < top_2[1079:1072]) ? 1 : 0;
assign detect_min[134][7] = (mid_1[1087:1080] < top_2[1087:1080]) ? 1 : 0;
assign detect_min[134][8] = (mid_1[1087:1080] < top_2[1095:1088]) ? 1 : 0;
assign detect_min[134][9] = (mid_1[1087:1080] < mid_0[1079:1072]) ? 1 : 0;
assign detect_min[134][10] = (mid_1[1087:1080] < mid_0[1087:1080]) ? 1 : 0;
assign detect_min[134][11] = (mid_1[1087:1080] < mid_0[1095:1088]) ? 1 : 0;
assign detect_min[134][12] = (mid_1[1087:1080] < mid_1[1079:1072]) ? 1 : 0;
assign detect_min[134][13] = (mid_1[1087:1080] < mid_1[1095:1088]) ? 1 : 0;
assign detect_min[134][14] = (mid_1[1087:1080] < mid_2[1079:1072]) ? 1 : 0;
assign detect_min[134][15] = (mid_1[1087:1080] < mid_2[1087:1080]) ? 1 : 0;
assign detect_min[134][16] = (mid_1[1087:1080] < mid_2[1095:1088]) ? 1 : 0;
assign detect_min[134][17] = (mid_1[1087:1080] < btm_0[1079:1072]) ? 1 : 0;
assign detect_min[134][18] = (mid_1[1087:1080] < btm_0[1087:1080]) ? 1 : 0;
assign detect_min[134][19] = (mid_1[1087:1080] < btm_0[1095:1088]) ? 1 : 0;
assign detect_min[134][20] = (mid_1[1087:1080] < btm_1[1079:1072]) ? 1 : 0;
assign detect_min[134][21] = (mid_1[1087:1080] < btm_1[1087:1080]) ? 1 : 0;
assign detect_min[134][22] = (mid_1[1087:1080] < btm_1[1095:1088]) ? 1 : 0;
assign detect_min[134][23] = (mid_1[1087:1080] < btm_2[1079:1072]) ? 1 : 0;
assign detect_min[134][24] = (mid_1[1087:1080] < btm_2[1087:1080]) ? 1 : 0;
assign detect_min[134][25] = (mid_1[1087:1080] < btm_2[1095:1088]) ? 1 : 0;

assign detect_min[135][0] = (mid_1[1095:1088] < top_0[1087:1080]) ? 1 : 0;
assign detect_min[135][1] = (mid_1[1095:1088] < top_0[1095:1088]) ? 1 : 0;
assign detect_min[135][2] = (mid_1[1095:1088] < top_0[1103:1096]) ? 1 : 0;
assign detect_min[135][3] = (mid_1[1095:1088] < top_1[1087:1080]) ? 1 : 0;
assign detect_min[135][4] = (mid_1[1095:1088] < top_1[1095:1088]) ? 1 : 0;
assign detect_min[135][5] = (mid_1[1095:1088] < top_1[1103:1096]) ? 1 : 0;
assign detect_min[135][6] = (mid_1[1095:1088] < top_2[1087:1080]) ? 1 : 0;
assign detect_min[135][7] = (mid_1[1095:1088] < top_2[1095:1088]) ? 1 : 0;
assign detect_min[135][8] = (mid_1[1095:1088] < top_2[1103:1096]) ? 1 : 0;
assign detect_min[135][9] = (mid_1[1095:1088] < mid_0[1087:1080]) ? 1 : 0;
assign detect_min[135][10] = (mid_1[1095:1088] < mid_0[1095:1088]) ? 1 : 0;
assign detect_min[135][11] = (mid_1[1095:1088] < mid_0[1103:1096]) ? 1 : 0;
assign detect_min[135][12] = (mid_1[1095:1088] < mid_1[1087:1080]) ? 1 : 0;
assign detect_min[135][13] = (mid_1[1095:1088] < mid_1[1103:1096]) ? 1 : 0;
assign detect_min[135][14] = (mid_1[1095:1088] < mid_2[1087:1080]) ? 1 : 0;
assign detect_min[135][15] = (mid_1[1095:1088] < mid_2[1095:1088]) ? 1 : 0;
assign detect_min[135][16] = (mid_1[1095:1088] < mid_2[1103:1096]) ? 1 : 0;
assign detect_min[135][17] = (mid_1[1095:1088] < btm_0[1087:1080]) ? 1 : 0;
assign detect_min[135][18] = (mid_1[1095:1088] < btm_0[1095:1088]) ? 1 : 0;
assign detect_min[135][19] = (mid_1[1095:1088] < btm_0[1103:1096]) ? 1 : 0;
assign detect_min[135][20] = (mid_1[1095:1088] < btm_1[1087:1080]) ? 1 : 0;
assign detect_min[135][21] = (mid_1[1095:1088] < btm_1[1095:1088]) ? 1 : 0;
assign detect_min[135][22] = (mid_1[1095:1088] < btm_1[1103:1096]) ? 1 : 0;
assign detect_min[135][23] = (mid_1[1095:1088] < btm_2[1087:1080]) ? 1 : 0;
assign detect_min[135][24] = (mid_1[1095:1088] < btm_2[1095:1088]) ? 1 : 0;
assign detect_min[135][25] = (mid_1[1095:1088] < btm_2[1103:1096]) ? 1 : 0;

assign detect_min[136][0] = (mid_1[1103:1096] < top_0[1095:1088]) ? 1 : 0;
assign detect_min[136][1] = (mid_1[1103:1096] < top_0[1103:1096]) ? 1 : 0;
assign detect_min[136][2] = (mid_1[1103:1096] < top_0[1111:1104]) ? 1 : 0;
assign detect_min[136][3] = (mid_1[1103:1096] < top_1[1095:1088]) ? 1 : 0;
assign detect_min[136][4] = (mid_1[1103:1096] < top_1[1103:1096]) ? 1 : 0;
assign detect_min[136][5] = (mid_1[1103:1096] < top_1[1111:1104]) ? 1 : 0;
assign detect_min[136][6] = (mid_1[1103:1096] < top_2[1095:1088]) ? 1 : 0;
assign detect_min[136][7] = (mid_1[1103:1096] < top_2[1103:1096]) ? 1 : 0;
assign detect_min[136][8] = (mid_1[1103:1096] < top_2[1111:1104]) ? 1 : 0;
assign detect_min[136][9] = (mid_1[1103:1096] < mid_0[1095:1088]) ? 1 : 0;
assign detect_min[136][10] = (mid_1[1103:1096] < mid_0[1103:1096]) ? 1 : 0;
assign detect_min[136][11] = (mid_1[1103:1096] < mid_0[1111:1104]) ? 1 : 0;
assign detect_min[136][12] = (mid_1[1103:1096] < mid_1[1095:1088]) ? 1 : 0;
assign detect_min[136][13] = (mid_1[1103:1096] < mid_1[1111:1104]) ? 1 : 0;
assign detect_min[136][14] = (mid_1[1103:1096] < mid_2[1095:1088]) ? 1 : 0;
assign detect_min[136][15] = (mid_1[1103:1096] < mid_2[1103:1096]) ? 1 : 0;
assign detect_min[136][16] = (mid_1[1103:1096] < mid_2[1111:1104]) ? 1 : 0;
assign detect_min[136][17] = (mid_1[1103:1096] < btm_0[1095:1088]) ? 1 : 0;
assign detect_min[136][18] = (mid_1[1103:1096] < btm_0[1103:1096]) ? 1 : 0;
assign detect_min[136][19] = (mid_1[1103:1096] < btm_0[1111:1104]) ? 1 : 0;
assign detect_min[136][20] = (mid_1[1103:1096] < btm_1[1095:1088]) ? 1 : 0;
assign detect_min[136][21] = (mid_1[1103:1096] < btm_1[1103:1096]) ? 1 : 0;
assign detect_min[136][22] = (mid_1[1103:1096] < btm_1[1111:1104]) ? 1 : 0;
assign detect_min[136][23] = (mid_1[1103:1096] < btm_2[1095:1088]) ? 1 : 0;
assign detect_min[136][24] = (mid_1[1103:1096] < btm_2[1103:1096]) ? 1 : 0;
assign detect_min[136][25] = (mid_1[1103:1096] < btm_2[1111:1104]) ? 1 : 0;

assign detect_min[137][0] = (mid_1[1111:1104] < top_0[1103:1096]) ? 1 : 0;
assign detect_min[137][1] = (mid_1[1111:1104] < top_0[1111:1104]) ? 1 : 0;
assign detect_min[137][2] = (mid_1[1111:1104] < top_0[1119:1112]) ? 1 : 0;
assign detect_min[137][3] = (mid_1[1111:1104] < top_1[1103:1096]) ? 1 : 0;
assign detect_min[137][4] = (mid_1[1111:1104] < top_1[1111:1104]) ? 1 : 0;
assign detect_min[137][5] = (mid_1[1111:1104] < top_1[1119:1112]) ? 1 : 0;
assign detect_min[137][6] = (mid_1[1111:1104] < top_2[1103:1096]) ? 1 : 0;
assign detect_min[137][7] = (mid_1[1111:1104] < top_2[1111:1104]) ? 1 : 0;
assign detect_min[137][8] = (mid_1[1111:1104] < top_2[1119:1112]) ? 1 : 0;
assign detect_min[137][9] = (mid_1[1111:1104] < mid_0[1103:1096]) ? 1 : 0;
assign detect_min[137][10] = (mid_1[1111:1104] < mid_0[1111:1104]) ? 1 : 0;
assign detect_min[137][11] = (mid_1[1111:1104] < mid_0[1119:1112]) ? 1 : 0;
assign detect_min[137][12] = (mid_1[1111:1104] < mid_1[1103:1096]) ? 1 : 0;
assign detect_min[137][13] = (mid_1[1111:1104] < mid_1[1119:1112]) ? 1 : 0;
assign detect_min[137][14] = (mid_1[1111:1104] < mid_2[1103:1096]) ? 1 : 0;
assign detect_min[137][15] = (mid_1[1111:1104] < mid_2[1111:1104]) ? 1 : 0;
assign detect_min[137][16] = (mid_1[1111:1104] < mid_2[1119:1112]) ? 1 : 0;
assign detect_min[137][17] = (mid_1[1111:1104] < btm_0[1103:1096]) ? 1 : 0;
assign detect_min[137][18] = (mid_1[1111:1104] < btm_0[1111:1104]) ? 1 : 0;
assign detect_min[137][19] = (mid_1[1111:1104] < btm_0[1119:1112]) ? 1 : 0;
assign detect_min[137][20] = (mid_1[1111:1104] < btm_1[1103:1096]) ? 1 : 0;
assign detect_min[137][21] = (mid_1[1111:1104] < btm_1[1111:1104]) ? 1 : 0;
assign detect_min[137][22] = (mid_1[1111:1104] < btm_1[1119:1112]) ? 1 : 0;
assign detect_min[137][23] = (mid_1[1111:1104] < btm_2[1103:1096]) ? 1 : 0;
assign detect_min[137][24] = (mid_1[1111:1104] < btm_2[1111:1104]) ? 1 : 0;
assign detect_min[137][25] = (mid_1[1111:1104] < btm_2[1119:1112]) ? 1 : 0;

assign detect_min[138][0] = (mid_1[1119:1112] < top_0[1111:1104]) ? 1 : 0;
assign detect_min[138][1] = (mid_1[1119:1112] < top_0[1119:1112]) ? 1 : 0;
assign detect_min[138][2] = (mid_1[1119:1112] < top_0[1127:1120]) ? 1 : 0;
assign detect_min[138][3] = (mid_1[1119:1112] < top_1[1111:1104]) ? 1 : 0;
assign detect_min[138][4] = (mid_1[1119:1112] < top_1[1119:1112]) ? 1 : 0;
assign detect_min[138][5] = (mid_1[1119:1112] < top_1[1127:1120]) ? 1 : 0;
assign detect_min[138][6] = (mid_1[1119:1112] < top_2[1111:1104]) ? 1 : 0;
assign detect_min[138][7] = (mid_1[1119:1112] < top_2[1119:1112]) ? 1 : 0;
assign detect_min[138][8] = (mid_1[1119:1112] < top_2[1127:1120]) ? 1 : 0;
assign detect_min[138][9] = (mid_1[1119:1112] < mid_0[1111:1104]) ? 1 : 0;
assign detect_min[138][10] = (mid_1[1119:1112] < mid_0[1119:1112]) ? 1 : 0;
assign detect_min[138][11] = (mid_1[1119:1112] < mid_0[1127:1120]) ? 1 : 0;
assign detect_min[138][12] = (mid_1[1119:1112] < mid_1[1111:1104]) ? 1 : 0;
assign detect_min[138][13] = (mid_1[1119:1112] < mid_1[1127:1120]) ? 1 : 0;
assign detect_min[138][14] = (mid_1[1119:1112] < mid_2[1111:1104]) ? 1 : 0;
assign detect_min[138][15] = (mid_1[1119:1112] < mid_2[1119:1112]) ? 1 : 0;
assign detect_min[138][16] = (mid_1[1119:1112] < mid_2[1127:1120]) ? 1 : 0;
assign detect_min[138][17] = (mid_1[1119:1112] < btm_0[1111:1104]) ? 1 : 0;
assign detect_min[138][18] = (mid_1[1119:1112] < btm_0[1119:1112]) ? 1 : 0;
assign detect_min[138][19] = (mid_1[1119:1112] < btm_0[1127:1120]) ? 1 : 0;
assign detect_min[138][20] = (mid_1[1119:1112] < btm_1[1111:1104]) ? 1 : 0;
assign detect_min[138][21] = (mid_1[1119:1112] < btm_1[1119:1112]) ? 1 : 0;
assign detect_min[138][22] = (mid_1[1119:1112] < btm_1[1127:1120]) ? 1 : 0;
assign detect_min[138][23] = (mid_1[1119:1112] < btm_2[1111:1104]) ? 1 : 0;
assign detect_min[138][24] = (mid_1[1119:1112] < btm_2[1119:1112]) ? 1 : 0;
assign detect_min[138][25] = (mid_1[1119:1112] < btm_2[1127:1120]) ? 1 : 0;

assign detect_min[139][0] = (mid_1[1127:1120] < top_0[1119:1112]) ? 1 : 0;
assign detect_min[139][1] = (mid_1[1127:1120] < top_0[1127:1120]) ? 1 : 0;
assign detect_min[139][2] = (mid_1[1127:1120] < top_0[1135:1128]) ? 1 : 0;
assign detect_min[139][3] = (mid_1[1127:1120] < top_1[1119:1112]) ? 1 : 0;
assign detect_min[139][4] = (mid_1[1127:1120] < top_1[1127:1120]) ? 1 : 0;
assign detect_min[139][5] = (mid_1[1127:1120] < top_1[1135:1128]) ? 1 : 0;
assign detect_min[139][6] = (mid_1[1127:1120] < top_2[1119:1112]) ? 1 : 0;
assign detect_min[139][7] = (mid_1[1127:1120] < top_2[1127:1120]) ? 1 : 0;
assign detect_min[139][8] = (mid_1[1127:1120] < top_2[1135:1128]) ? 1 : 0;
assign detect_min[139][9] = (mid_1[1127:1120] < mid_0[1119:1112]) ? 1 : 0;
assign detect_min[139][10] = (mid_1[1127:1120] < mid_0[1127:1120]) ? 1 : 0;
assign detect_min[139][11] = (mid_1[1127:1120] < mid_0[1135:1128]) ? 1 : 0;
assign detect_min[139][12] = (mid_1[1127:1120] < mid_1[1119:1112]) ? 1 : 0;
assign detect_min[139][13] = (mid_1[1127:1120] < mid_1[1135:1128]) ? 1 : 0;
assign detect_min[139][14] = (mid_1[1127:1120] < mid_2[1119:1112]) ? 1 : 0;
assign detect_min[139][15] = (mid_1[1127:1120] < mid_2[1127:1120]) ? 1 : 0;
assign detect_min[139][16] = (mid_1[1127:1120] < mid_2[1135:1128]) ? 1 : 0;
assign detect_min[139][17] = (mid_1[1127:1120] < btm_0[1119:1112]) ? 1 : 0;
assign detect_min[139][18] = (mid_1[1127:1120] < btm_0[1127:1120]) ? 1 : 0;
assign detect_min[139][19] = (mid_1[1127:1120] < btm_0[1135:1128]) ? 1 : 0;
assign detect_min[139][20] = (mid_1[1127:1120] < btm_1[1119:1112]) ? 1 : 0;
assign detect_min[139][21] = (mid_1[1127:1120] < btm_1[1127:1120]) ? 1 : 0;
assign detect_min[139][22] = (mid_1[1127:1120] < btm_1[1135:1128]) ? 1 : 0;
assign detect_min[139][23] = (mid_1[1127:1120] < btm_2[1119:1112]) ? 1 : 0;
assign detect_min[139][24] = (mid_1[1127:1120] < btm_2[1127:1120]) ? 1 : 0;
assign detect_min[139][25] = (mid_1[1127:1120] < btm_2[1135:1128]) ? 1 : 0;

assign detect_min[140][0] = (mid_1[1135:1128] < top_0[1127:1120]) ? 1 : 0;
assign detect_min[140][1] = (mid_1[1135:1128] < top_0[1135:1128]) ? 1 : 0;
assign detect_min[140][2] = (mid_1[1135:1128] < top_0[1143:1136]) ? 1 : 0;
assign detect_min[140][3] = (mid_1[1135:1128] < top_1[1127:1120]) ? 1 : 0;
assign detect_min[140][4] = (mid_1[1135:1128] < top_1[1135:1128]) ? 1 : 0;
assign detect_min[140][5] = (mid_1[1135:1128] < top_1[1143:1136]) ? 1 : 0;
assign detect_min[140][6] = (mid_1[1135:1128] < top_2[1127:1120]) ? 1 : 0;
assign detect_min[140][7] = (mid_1[1135:1128] < top_2[1135:1128]) ? 1 : 0;
assign detect_min[140][8] = (mid_1[1135:1128] < top_2[1143:1136]) ? 1 : 0;
assign detect_min[140][9] = (mid_1[1135:1128] < mid_0[1127:1120]) ? 1 : 0;
assign detect_min[140][10] = (mid_1[1135:1128] < mid_0[1135:1128]) ? 1 : 0;
assign detect_min[140][11] = (mid_1[1135:1128] < mid_0[1143:1136]) ? 1 : 0;
assign detect_min[140][12] = (mid_1[1135:1128] < mid_1[1127:1120]) ? 1 : 0;
assign detect_min[140][13] = (mid_1[1135:1128] < mid_1[1143:1136]) ? 1 : 0;
assign detect_min[140][14] = (mid_1[1135:1128] < mid_2[1127:1120]) ? 1 : 0;
assign detect_min[140][15] = (mid_1[1135:1128] < mid_2[1135:1128]) ? 1 : 0;
assign detect_min[140][16] = (mid_1[1135:1128] < mid_2[1143:1136]) ? 1 : 0;
assign detect_min[140][17] = (mid_1[1135:1128] < btm_0[1127:1120]) ? 1 : 0;
assign detect_min[140][18] = (mid_1[1135:1128] < btm_0[1135:1128]) ? 1 : 0;
assign detect_min[140][19] = (mid_1[1135:1128] < btm_0[1143:1136]) ? 1 : 0;
assign detect_min[140][20] = (mid_1[1135:1128] < btm_1[1127:1120]) ? 1 : 0;
assign detect_min[140][21] = (mid_1[1135:1128] < btm_1[1135:1128]) ? 1 : 0;
assign detect_min[140][22] = (mid_1[1135:1128] < btm_1[1143:1136]) ? 1 : 0;
assign detect_min[140][23] = (mid_1[1135:1128] < btm_2[1127:1120]) ? 1 : 0;
assign detect_min[140][24] = (mid_1[1135:1128] < btm_2[1135:1128]) ? 1 : 0;
assign detect_min[140][25] = (mid_1[1135:1128] < btm_2[1143:1136]) ? 1 : 0;

assign detect_min[141][0] = (mid_1[1143:1136] < top_0[1135:1128]) ? 1 : 0;
assign detect_min[141][1] = (mid_1[1143:1136] < top_0[1143:1136]) ? 1 : 0;
assign detect_min[141][2] = (mid_1[1143:1136] < top_0[1151:1144]) ? 1 : 0;
assign detect_min[141][3] = (mid_1[1143:1136] < top_1[1135:1128]) ? 1 : 0;
assign detect_min[141][4] = (mid_1[1143:1136] < top_1[1143:1136]) ? 1 : 0;
assign detect_min[141][5] = (mid_1[1143:1136] < top_1[1151:1144]) ? 1 : 0;
assign detect_min[141][6] = (mid_1[1143:1136] < top_2[1135:1128]) ? 1 : 0;
assign detect_min[141][7] = (mid_1[1143:1136] < top_2[1143:1136]) ? 1 : 0;
assign detect_min[141][8] = (mid_1[1143:1136] < top_2[1151:1144]) ? 1 : 0;
assign detect_min[141][9] = (mid_1[1143:1136] < mid_0[1135:1128]) ? 1 : 0;
assign detect_min[141][10] = (mid_1[1143:1136] < mid_0[1143:1136]) ? 1 : 0;
assign detect_min[141][11] = (mid_1[1143:1136] < mid_0[1151:1144]) ? 1 : 0;
assign detect_min[141][12] = (mid_1[1143:1136] < mid_1[1135:1128]) ? 1 : 0;
assign detect_min[141][13] = (mid_1[1143:1136] < mid_1[1151:1144]) ? 1 : 0;
assign detect_min[141][14] = (mid_1[1143:1136] < mid_2[1135:1128]) ? 1 : 0;
assign detect_min[141][15] = (mid_1[1143:1136] < mid_2[1143:1136]) ? 1 : 0;
assign detect_min[141][16] = (mid_1[1143:1136] < mid_2[1151:1144]) ? 1 : 0;
assign detect_min[141][17] = (mid_1[1143:1136] < btm_0[1135:1128]) ? 1 : 0;
assign detect_min[141][18] = (mid_1[1143:1136] < btm_0[1143:1136]) ? 1 : 0;
assign detect_min[141][19] = (mid_1[1143:1136] < btm_0[1151:1144]) ? 1 : 0;
assign detect_min[141][20] = (mid_1[1143:1136] < btm_1[1135:1128]) ? 1 : 0;
assign detect_min[141][21] = (mid_1[1143:1136] < btm_1[1143:1136]) ? 1 : 0;
assign detect_min[141][22] = (mid_1[1143:1136] < btm_1[1151:1144]) ? 1 : 0;
assign detect_min[141][23] = (mid_1[1143:1136] < btm_2[1135:1128]) ? 1 : 0;
assign detect_min[141][24] = (mid_1[1143:1136] < btm_2[1143:1136]) ? 1 : 0;
assign detect_min[141][25] = (mid_1[1143:1136] < btm_2[1151:1144]) ? 1 : 0;

assign detect_min[142][0] = (mid_1[1151:1144] < top_0[1143:1136]) ? 1 : 0;
assign detect_min[142][1] = (mid_1[1151:1144] < top_0[1151:1144]) ? 1 : 0;
assign detect_min[142][2] = (mid_1[1151:1144] < top_0[1159:1152]) ? 1 : 0;
assign detect_min[142][3] = (mid_1[1151:1144] < top_1[1143:1136]) ? 1 : 0;
assign detect_min[142][4] = (mid_1[1151:1144] < top_1[1151:1144]) ? 1 : 0;
assign detect_min[142][5] = (mid_1[1151:1144] < top_1[1159:1152]) ? 1 : 0;
assign detect_min[142][6] = (mid_1[1151:1144] < top_2[1143:1136]) ? 1 : 0;
assign detect_min[142][7] = (mid_1[1151:1144] < top_2[1151:1144]) ? 1 : 0;
assign detect_min[142][8] = (mid_1[1151:1144] < top_2[1159:1152]) ? 1 : 0;
assign detect_min[142][9] = (mid_1[1151:1144] < mid_0[1143:1136]) ? 1 : 0;
assign detect_min[142][10] = (mid_1[1151:1144] < mid_0[1151:1144]) ? 1 : 0;
assign detect_min[142][11] = (mid_1[1151:1144] < mid_0[1159:1152]) ? 1 : 0;
assign detect_min[142][12] = (mid_1[1151:1144] < mid_1[1143:1136]) ? 1 : 0;
assign detect_min[142][13] = (mid_1[1151:1144] < mid_1[1159:1152]) ? 1 : 0;
assign detect_min[142][14] = (mid_1[1151:1144] < mid_2[1143:1136]) ? 1 : 0;
assign detect_min[142][15] = (mid_1[1151:1144] < mid_2[1151:1144]) ? 1 : 0;
assign detect_min[142][16] = (mid_1[1151:1144] < mid_2[1159:1152]) ? 1 : 0;
assign detect_min[142][17] = (mid_1[1151:1144] < btm_0[1143:1136]) ? 1 : 0;
assign detect_min[142][18] = (mid_1[1151:1144] < btm_0[1151:1144]) ? 1 : 0;
assign detect_min[142][19] = (mid_1[1151:1144] < btm_0[1159:1152]) ? 1 : 0;
assign detect_min[142][20] = (mid_1[1151:1144] < btm_1[1143:1136]) ? 1 : 0;
assign detect_min[142][21] = (mid_1[1151:1144] < btm_1[1151:1144]) ? 1 : 0;
assign detect_min[142][22] = (mid_1[1151:1144] < btm_1[1159:1152]) ? 1 : 0;
assign detect_min[142][23] = (mid_1[1151:1144] < btm_2[1143:1136]) ? 1 : 0;
assign detect_min[142][24] = (mid_1[1151:1144] < btm_2[1151:1144]) ? 1 : 0;
assign detect_min[142][25] = (mid_1[1151:1144] < btm_2[1159:1152]) ? 1 : 0;

assign detect_min[143][0] = (mid_1[1159:1152] < top_0[1151:1144]) ? 1 : 0;
assign detect_min[143][1] = (mid_1[1159:1152] < top_0[1159:1152]) ? 1 : 0;
assign detect_min[143][2] = (mid_1[1159:1152] < top_0[1167:1160]) ? 1 : 0;
assign detect_min[143][3] = (mid_1[1159:1152] < top_1[1151:1144]) ? 1 : 0;
assign detect_min[143][4] = (mid_1[1159:1152] < top_1[1159:1152]) ? 1 : 0;
assign detect_min[143][5] = (mid_1[1159:1152] < top_1[1167:1160]) ? 1 : 0;
assign detect_min[143][6] = (mid_1[1159:1152] < top_2[1151:1144]) ? 1 : 0;
assign detect_min[143][7] = (mid_1[1159:1152] < top_2[1159:1152]) ? 1 : 0;
assign detect_min[143][8] = (mid_1[1159:1152] < top_2[1167:1160]) ? 1 : 0;
assign detect_min[143][9] = (mid_1[1159:1152] < mid_0[1151:1144]) ? 1 : 0;
assign detect_min[143][10] = (mid_1[1159:1152] < mid_0[1159:1152]) ? 1 : 0;
assign detect_min[143][11] = (mid_1[1159:1152] < mid_0[1167:1160]) ? 1 : 0;
assign detect_min[143][12] = (mid_1[1159:1152] < mid_1[1151:1144]) ? 1 : 0;
assign detect_min[143][13] = (mid_1[1159:1152] < mid_1[1167:1160]) ? 1 : 0;
assign detect_min[143][14] = (mid_1[1159:1152] < mid_2[1151:1144]) ? 1 : 0;
assign detect_min[143][15] = (mid_1[1159:1152] < mid_2[1159:1152]) ? 1 : 0;
assign detect_min[143][16] = (mid_1[1159:1152] < mid_2[1167:1160]) ? 1 : 0;
assign detect_min[143][17] = (mid_1[1159:1152] < btm_0[1151:1144]) ? 1 : 0;
assign detect_min[143][18] = (mid_1[1159:1152] < btm_0[1159:1152]) ? 1 : 0;
assign detect_min[143][19] = (mid_1[1159:1152] < btm_0[1167:1160]) ? 1 : 0;
assign detect_min[143][20] = (mid_1[1159:1152] < btm_1[1151:1144]) ? 1 : 0;
assign detect_min[143][21] = (mid_1[1159:1152] < btm_1[1159:1152]) ? 1 : 0;
assign detect_min[143][22] = (mid_1[1159:1152] < btm_1[1167:1160]) ? 1 : 0;
assign detect_min[143][23] = (mid_1[1159:1152] < btm_2[1151:1144]) ? 1 : 0;
assign detect_min[143][24] = (mid_1[1159:1152] < btm_2[1159:1152]) ? 1 : 0;
assign detect_min[143][25] = (mid_1[1159:1152] < btm_2[1167:1160]) ? 1 : 0;

assign detect_min[144][0] = (mid_1[1167:1160] < top_0[1159:1152]) ? 1 : 0;
assign detect_min[144][1] = (mid_1[1167:1160] < top_0[1167:1160]) ? 1 : 0;
assign detect_min[144][2] = (mid_1[1167:1160] < top_0[1175:1168]) ? 1 : 0;
assign detect_min[144][3] = (mid_1[1167:1160] < top_1[1159:1152]) ? 1 : 0;
assign detect_min[144][4] = (mid_1[1167:1160] < top_1[1167:1160]) ? 1 : 0;
assign detect_min[144][5] = (mid_1[1167:1160] < top_1[1175:1168]) ? 1 : 0;
assign detect_min[144][6] = (mid_1[1167:1160] < top_2[1159:1152]) ? 1 : 0;
assign detect_min[144][7] = (mid_1[1167:1160] < top_2[1167:1160]) ? 1 : 0;
assign detect_min[144][8] = (mid_1[1167:1160] < top_2[1175:1168]) ? 1 : 0;
assign detect_min[144][9] = (mid_1[1167:1160] < mid_0[1159:1152]) ? 1 : 0;
assign detect_min[144][10] = (mid_1[1167:1160] < mid_0[1167:1160]) ? 1 : 0;
assign detect_min[144][11] = (mid_1[1167:1160] < mid_0[1175:1168]) ? 1 : 0;
assign detect_min[144][12] = (mid_1[1167:1160] < mid_1[1159:1152]) ? 1 : 0;
assign detect_min[144][13] = (mid_1[1167:1160] < mid_1[1175:1168]) ? 1 : 0;
assign detect_min[144][14] = (mid_1[1167:1160] < mid_2[1159:1152]) ? 1 : 0;
assign detect_min[144][15] = (mid_1[1167:1160] < mid_2[1167:1160]) ? 1 : 0;
assign detect_min[144][16] = (mid_1[1167:1160] < mid_2[1175:1168]) ? 1 : 0;
assign detect_min[144][17] = (mid_1[1167:1160] < btm_0[1159:1152]) ? 1 : 0;
assign detect_min[144][18] = (mid_1[1167:1160] < btm_0[1167:1160]) ? 1 : 0;
assign detect_min[144][19] = (mid_1[1167:1160] < btm_0[1175:1168]) ? 1 : 0;
assign detect_min[144][20] = (mid_1[1167:1160] < btm_1[1159:1152]) ? 1 : 0;
assign detect_min[144][21] = (mid_1[1167:1160] < btm_1[1167:1160]) ? 1 : 0;
assign detect_min[144][22] = (mid_1[1167:1160] < btm_1[1175:1168]) ? 1 : 0;
assign detect_min[144][23] = (mid_1[1167:1160] < btm_2[1159:1152]) ? 1 : 0;
assign detect_min[144][24] = (mid_1[1167:1160] < btm_2[1167:1160]) ? 1 : 0;
assign detect_min[144][25] = (mid_1[1167:1160] < btm_2[1175:1168]) ? 1 : 0;

assign detect_min[145][0] = (mid_1[1175:1168] < top_0[1167:1160]) ? 1 : 0;
assign detect_min[145][1] = (mid_1[1175:1168] < top_0[1175:1168]) ? 1 : 0;
assign detect_min[145][2] = (mid_1[1175:1168] < top_0[1183:1176]) ? 1 : 0;
assign detect_min[145][3] = (mid_1[1175:1168] < top_1[1167:1160]) ? 1 : 0;
assign detect_min[145][4] = (mid_1[1175:1168] < top_1[1175:1168]) ? 1 : 0;
assign detect_min[145][5] = (mid_1[1175:1168] < top_1[1183:1176]) ? 1 : 0;
assign detect_min[145][6] = (mid_1[1175:1168] < top_2[1167:1160]) ? 1 : 0;
assign detect_min[145][7] = (mid_1[1175:1168] < top_2[1175:1168]) ? 1 : 0;
assign detect_min[145][8] = (mid_1[1175:1168] < top_2[1183:1176]) ? 1 : 0;
assign detect_min[145][9] = (mid_1[1175:1168] < mid_0[1167:1160]) ? 1 : 0;
assign detect_min[145][10] = (mid_1[1175:1168] < mid_0[1175:1168]) ? 1 : 0;
assign detect_min[145][11] = (mid_1[1175:1168] < mid_0[1183:1176]) ? 1 : 0;
assign detect_min[145][12] = (mid_1[1175:1168] < mid_1[1167:1160]) ? 1 : 0;
assign detect_min[145][13] = (mid_1[1175:1168] < mid_1[1183:1176]) ? 1 : 0;
assign detect_min[145][14] = (mid_1[1175:1168] < mid_2[1167:1160]) ? 1 : 0;
assign detect_min[145][15] = (mid_1[1175:1168] < mid_2[1175:1168]) ? 1 : 0;
assign detect_min[145][16] = (mid_1[1175:1168] < mid_2[1183:1176]) ? 1 : 0;
assign detect_min[145][17] = (mid_1[1175:1168] < btm_0[1167:1160]) ? 1 : 0;
assign detect_min[145][18] = (mid_1[1175:1168] < btm_0[1175:1168]) ? 1 : 0;
assign detect_min[145][19] = (mid_1[1175:1168] < btm_0[1183:1176]) ? 1 : 0;
assign detect_min[145][20] = (mid_1[1175:1168] < btm_1[1167:1160]) ? 1 : 0;
assign detect_min[145][21] = (mid_1[1175:1168] < btm_1[1175:1168]) ? 1 : 0;
assign detect_min[145][22] = (mid_1[1175:1168] < btm_1[1183:1176]) ? 1 : 0;
assign detect_min[145][23] = (mid_1[1175:1168] < btm_2[1167:1160]) ? 1 : 0;
assign detect_min[145][24] = (mid_1[1175:1168] < btm_2[1175:1168]) ? 1 : 0;
assign detect_min[145][25] = (mid_1[1175:1168] < btm_2[1183:1176]) ? 1 : 0;

assign detect_min[146][0] = (mid_1[1183:1176] < top_0[1175:1168]) ? 1 : 0;
assign detect_min[146][1] = (mid_1[1183:1176] < top_0[1183:1176]) ? 1 : 0;
assign detect_min[146][2] = (mid_1[1183:1176] < top_0[1191:1184]) ? 1 : 0;
assign detect_min[146][3] = (mid_1[1183:1176] < top_1[1175:1168]) ? 1 : 0;
assign detect_min[146][4] = (mid_1[1183:1176] < top_1[1183:1176]) ? 1 : 0;
assign detect_min[146][5] = (mid_1[1183:1176] < top_1[1191:1184]) ? 1 : 0;
assign detect_min[146][6] = (mid_1[1183:1176] < top_2[1175:1168]) ? 1 : 0;
assign detect_min[146][7] = (mid_1[1183:1176] < top_2[1183:1176]) ? 1 : 0;
assign detect_min[146][8] = (mid_1[1183:1176] < top_2[1191:1184]) ? 1 : 0;
assign detect_min[146][9] = (mid_1[1183:1176] < mid_0[1175:1168]) ? 1 : 0;
assign detect_min[146][10] = (mid_1[1183:1176] < mid_0[1183:1176]) ? 1 : 0;
assign detect_min[146][11] = (mid_1[1183:1176] < mid_0[1191:1184]) ? 1 : 0;
assign detect_min[146][12] = (mid_1[1183:1176] < mid_1[1175:1168]) ? 1 : 0;
assign detect_min[146][13] = (mid_1[1183:1176] < mid_1[1191:1184]) ? 1 : 0;
assign detect_min[146][14] = (mid_1[1183:1176] < mid_2[1175:1168]) ? 1 : 0;
assign detect_min[146][15] = (mid_1[1183:1176] < mid_2[1183:1176]) ? 1 : 0;
assign detect_min[146][16] = (mid_1[1183:1176] < mid_2[1191:1184]) ? 1 : 0;
assign detect_min[146][17] = (mid_1[1183:1176] < btm_0[1175:1168]) ? 1 : 0;
assign detect_min[146][18] = (mid_1[1183:1176] < btm_0[1183:1176]) ? 1 : 0;
assign detect_min[146][19] = (mid_1[1183:1176] < btm_0[1191:1184]) ? 1 : 0;
assign detect_min[146][20] = (mid_1[1183:1176] < btm_1[1175:1168]) ? 1 : 0;
assign detect_min[146][21] = (mid_1[1183:1176] < btm_1[1183:1176]) ? 1 : 0;
assign detect_min[146][22] = (mid_1[1183:1176] < btm_1[1191:1184]) ? 1 : 0;
assign detect_min[146][23] = (mid_1[1183:1176] < btm_2[1175:1168]) ? 1 : 0;
assign detect_min[146][24] = (mid_1[1183:1176] < btm_2[1183:1176]) ? 1 : 0;
assign detect_min[146][25] = (mid_1[1183:1176] < btm_2[1191:1184]) ? 1 : 0;

assign detect_min[147][0] = (mid_1[1191:1184] < top_0[1183:1176]) ? 1 : 0;
assign detect_min[147][1] = (mid_1[1191:1184] < top_0[1191:1184]) ? 1 : 0;
assign detect_min[147][2] = (mid_1[1191:1184] < top_0[1199:1192]) ? 1 : 0;
assign detect_min[147][3] = (mid_1[1191:1184] < top_1[1183:1176]) ? 1 : 0;
assign detect_min[147][4] = (mid_1[1191:1184] < top_1[1191:1184]) ? 1 : 0;
assign detect_min[147][5] = (mid_1[1191:1184] < top_1[1199:1192]) ? 1 : 0;
assign detect_min[147][6] = (mid_1[1191:1184] < top_2[1183:1176]) ? 1 : 0;
assign detect_min[147][7] = (mid_1[1191:1184] < top_2[1191:1184]) ? 1 : 0;
assign detect_min[147][8] = (mid_1[1191:1184] < top_2[1199:1192]) ? 1 : 0;
assign detect_min[147][9] = (mid_1[1191:1184] < mid_0[1183:1176]) ? 1 : 0;
assign detect_min[147][10] = (mid_1[1191:1184] < mid_0[1191:1184]) ? 1 : 0;
assign detect_min[147][11] = (mid_1[1191:1184] < mid_0[1199:1192]) ? 1 : 0;
assign detect_min[147][12] = (mid_1[1191:1184] < mid_1[1183:1176]) ? 1 : 0;
assign detect_min[147][13] = (mid_1[1191:1184] < mid_1[1199:1192]) ? 1 : 0;
assign detect_min[147][14] = (mid_1[1191:1184] < mid_2[1183:1176]) ? 1 : 0;
assign detect_min[147][15] = (mid_1[1191:1184] < mid_2[1191:1184]) ? 1 : 0;
assign detect_min[147][16] = (mid_1[1191:1184] < mid_2[1199:1192]) ? 1 : 0;
assign detect_min[147][17] = (mid_1[1191:1184] < btm_0[1183:1176]) ? 1 : 0;
assign detect_min[147][18] = (mid_1[1191:1184] < btm_0[1191:1184]) ? 1 : 0;
assign detect_min[147][19] = (mid_1[1191:1184] < btm_0[1199:1192]) ? 1 : 0;
assign detect_min[147][20] = (mid_1[1191:1184] < btm_1[1183:1176]) ? 1 : 0;
assign detect_min[147][21] = (mid_1[1191:1184] < btm_1[1191:1184]) ? 1 : 0;
assign detect_min[147][22] = (mid_1[1191:1184] < btm_1[1199:1192]) ? 1 : 0;
assign detect_min[147][23] = (mid_1[1191:1184] < btm_2[1183:1176]) ? 1 : 0;
assign detect_min[147][24] = (mid_1[1191:1184] < btm_2[1191:1184]) ? 1 : 0;
assign detect_min[147][25] = (mid_1[1191:1184] < btm_2[1199:1192]) ? 1 : 0;

assign detect_min[148][0] = (mid_1[1199:1192] < top_0[1191:1184]) ? 1 : 0;
assign detect_min[148][1] = (mid_1[1199:1192] < top_0[1199:1192]) ? 1 : 0;
assign detect_min[148][2] = (mid_1[1199:1192] < top_0[1207:1200]) ? 1 : 0;
assign detect_min[148][3] = (mid_1[1199:1192] < top_1[1191:1184]) ? 1 : 0;
assign detect_min[148][4] = (mid_1[1199:1192] < top_1[1199:1192]) ? 1 : 0;
assign detect_min[148][5] = (mid_1[1199:1192] < top_1[1207:1200]) ? 1 : 0;
assign detect_min[148][6] = (mid_1[1199:1192] < top_2[1191:1184]) ? 1 : 0;
assign detect_min[148][7] = (mid_1[1199:1192] < top_2[1199:1192]) ? 1 : 0;
assign detect_min[148][8] = (mid_1[1199:1192] < top_2[1207:1200]) ? 1 : 0;
assign detect_min[148][9] = (mid_1[1199:1192] < mid_0[1191:1184]) ? 1 : 0;
assign detect_min[148][10] = (mid_1[1199:1192] < mid_0[1199:1192]) ? 1 : 0;
assign detect_min[148][11] = (mid_1[1199:1192] < mid_0[1207:1200]) ? 1 : 0;
assign detect_min[148][12] = (mid_1[1199:1192] < mid_1[1191:1184]) ? 1 : 0;
assign detect_min[148][13] = (mid_1[1199:1192] < mid_1[1207:1200]) ? 1 : 0;
assign detect_min[148][14] = (mid_1[1199:1192] < mid_2[1191:1184]) ? 1 : 0;
assign detect_min[148][15] = (mid_1[1199:1192] < mid_2[1199:1192]) ? 1 : 0;
assign detect_min[148][16] = (mid_1[1199:1192] < mid_2[1207:1200]) ? 1 : 0;
assign detect_min[148][17] = (mid_1[1199:1192] < btm_0[1191:1184]) ? 1 : 0;
assign detect_min[148][18] = (mid_1[1199:1192] < btm_0[1199:1192]) ? 1 : 0;
assign detect_min[148][19] = (mid_1[1199:1192] < btm_0[1207:1200]) ? 1 : 0;
assign detect_min[148][20] = (mid_1[1199:1192] < btm_1[1191:1184]) ? 1 : 0;
assign detect_min[148][21] = (mid_1[1199:1192] < btm_1[1199:1192]) ? 1 : 0;
assign detect_min[148][22] = (mid_1[1199:1192] < btm_1[1207:1200]) ? 1 : 0;
assign detect_min[148][23] = (mid_1[1199:1192] < btm_2[1191:1184]) ? 1 : 0;
assign detect_min[148][24] = (mid_1[1199:1192] < btm_2[1199:1192]) ? 1 : 0;
assign detect_min[148][25] = (mid_1[1199:1192] < btm_2[1207:1200]) ? 1 : 0;

assign detect_min[149][0] = (mid_1[1207:1200] < top_0[1199:1192]) ? 1 : 0;
assign detect_min[149][1] = (mid_1[1207:1200] < top_0[1207:1200]) ? 1 : 0;
assign detect_min[149][2] = (mid_1[1207:1200] < top_0[1215:1208]) ? 1 : 0;
assign detect_min[149][3] = (mid_1[1207:1200] < top_1[1199:1192]) ? 1 : 0;
assign detect_min[149][4] = (mid_1[1207:1200] < top_1[1207:1200]) ? 1 : 0;
assign detect_min[149][5] = (mid_1[1207:1200] < top_1[1215:1208]) ? 1 : 0;
assign detect_min[149][6] = (mid_1[1207:1200] < top_2[1199:1192]) ? 1 : 0;
assign detect_min[149][7] = (mid_1[1207:1200] < top_2[1207:1200]) ? 1 : 0;
assign detect_min[149][8] = (mid_1[1207:1200] < top_2[1215:1208]) ? 1 : 0;
assign detect_min[149][9] = (mid_1[1207:1200] < mid_0[1199:1192]) ? 1 : 0;
assign detect_min[149][10] = (mid_1[1207:1200] < mid_0[1207:1200]) ? 1 : 0;
assign detect_min[149][11] = (mid_1[1207:1200] < mid_0[1215:1208]) ? 1 : 0;
assign detect_min[149][12] = (mid_1[1207:1200] < mid_1[1199:1192]) ? 1 : 0;
assign detect_min[149][13] = (mid_1[1207:1200] < mid_1[1215:1208]) ? 1 : 0;
assign detect_min[149][14] = (mid_1[1207:1200] < mid_2[1199:1192]) ? 1 : 0;
assign detect_min[149][15] = (mid_1[1207:1200] < mid_2[1207:1200]) ? 1 : 0;
assign detect_min[149][16] = (mid_1[1207:1200] < mid_2[1215:1208]) ? 1 : 0;
assign detect_min[149][17] = (mid_1[1207:1200] < btm_0[1199:1192]) ? 1 : 0;
assign detect_min[149][18] = (mid_1[1207:1200] < btm_0[1207:1200]) ? 1 : 0;
assign detect_min[149][19] = (mid_1[1207:1200] < btm_0[1215:1208]) ? 1 : 0;
assign detect_min[149][20] = (mid_1[1207:1200] < btm_1[1199:1192]) ? 1 : 0;
assign detect_min[149][21] = (mid_1[1207:1200] < btm_1[1207:1200]) ? 1 : 0;
assign detect_min[149][22] = (mid_1[1207:1200] < btm_1[1215:1208]) ? 1 : 0;
assign detect_min[149][23] = (mid_1[1207:1200] < btm_2[1199:1192]) ? 1 : 0;
assign detect_min[149][24] = (mid_1[1207:1200] < btm_2[1207:1200]) ? 1 : 0;
assign detect_min[149][25] = (mid_1[1207:1200] < btm_2[1215:1208]) ? 1 : 0;

assign detect_min[150][0] = (mid_1[1215:1208] < top_0[1207:1200]) ? 1 : 0;
assign detect_min[150][1] = (mid_1[1215:1208] < top_0[1215:1208]) ? 1 : 0;
assign detect_min[150][2] = (mid_1[1215:1208] < top_0[1223:1216]) ? 1 : 0;
assign detect_min[150][3] = (mid_1[1215:1208] < top_1[1207:1200]) ? 1 : 0;
assign detect_min[150][4] = (mid_1[1215:1208] < top_1[1215:1208]) ? 1 : 0;
assign detect_min[150][5] = (mid_1[1215:1208] < top_1[1223:1216]) ? 1 : 0;
assign detect_min[150][6] = (mid_1[1215:1208] < top_2[1207:1200]) ? 1 : 0;
assign detect_min[150][7] = (mid_1[1215:1208] < top_2[1215:1208]) ? 1 : 0;
assign detect_min[150][8] = (mid_1[1215:1208] < top_2[1223:1216]) ? 1 : 0;
assign detect_min[150][9] = (mid_1[1215:1208] < mid_0[1207:1200]) ? 1 : 0;
assign detect_min[150][10] = (mid_1[1215:1208] < mid_0[1215:1208]) ? 1 : 0;
assign detect_min[150][11] = (mid_1[1215:1208] < mid_0[1223:1216]) ? 1 : 0;
assign detect_min[150][12] = (mid_1[1215:1208] < mid_1[1207:1200]) ? 1 : 0;
assign detect_min[150][13] = (mid_1[1215:1208] < mid_1[1223:1216]) ? 1 : 0;
assign detect_min[150][14] = (mid_1[1215:1208] < mid_2[1207:1200]) ? 1 : 0;
assign detect_min[150][15] = (mid_1[1215:1208] < mid_2[1215:1208]) ? 1 : 0;
assign detect_min[150][16] = (mid_1[1215:1208] < mid_2[1223:1216]) ? 1 : 0;
assign detect_min[150][17] = (mid_1[1215:1208] < btm_0[1207:1200]) ? 1 : 0;
assign detect_min[150][18] = (mid_1[1215:1208] < btm_0[1215:1208]) ? 1 : 0;
assign detect_min[150][19] = (mid_1[1215:1208] < btm_0[1223:1216]) ? 1 : 0;
assign detect_min[150][20] = (mid_1[1215:1208] < btm_1[1207:1200]) ? 1 : 0;
assign detect_min[150][21] = (mid_1[1215:1208] < btm_1[1215:1208]) ? 1 : 0;
assign detect_min[150][22] = (mid_1[1215:1208] < btm_1[1223:1216]) ? 1 : 0;
assign detect_min[150][23] = (mid_1[1215:1208] < btm_2[1207:1200]) ? 1 : 0;
assign detect_min[150][24] = (mid_1[1215:1208] < btm_2[1215:1208]) ? 1 : 0;
assign detect_min[150][25] = (mid_1[1215:1208] < btm_2[1223:1216]) ? 1 : 0;

assign detect_min[151][0] = (mid_1[1223:1216] < top_0[1215:1208]) ? 1 : 0;
assign detect_min[151][1] = (mid_1[1223:1216] < top_0[1223:1216]) ? 1 : 0;
assign detect_min[151][2] = (mid_1[1223:1216] < top_0[1231:1224]) ? 1 : 0;
assign detect_min[151][3] = (mid_1[1223:1216] < top_1[1215:1208]) ? 1 : 0;
assign detect_min[151][4] = (mid_1[1223:1216] < top_1[1223:1216]) ? 1 : 0;
assign detect_min[151][5] = (mid_1[1223:1216] < top_1[1231:1224]) ? 1 : 0;
assign detect_min[151][6] = (mid_1[1223:1216] < top_2[1215:1208]) ? 1 : 0;
assign detect_min[151][7] = (mid_1[1223:1216] < top_2[1223:1216]) ? 1 : 0;
assign detect_min[151][8] = (mid_1[1223:1216] < top_2[1231:1224]) ? 1 : 0;
assign detect_min[151][9] = (mid_1[1223:1216] < mid_0[1215:1208]) ? 1 : 0;
assign detect_min[151][10] = (mid_1[1223:1216] < mid_0[1223:1216]) ? 1 : 0;
assign detect_min[151][11] = (mid_1[1223:1216] < mid_0[1231:1224]) ? 1 : 0;
assign detect_min[151][12] = (mid_1[1223:1216] < mid_1[1215:1208]) ? 1 : 0;
assign detect_min[151][13] = (mid_1[1223:1216] < mid_1[1231:1224]) ? 1 : 0;
assign detect_min[151][14] = (mid_1[1223:1216] < mid_2[1215:1208]) ? 1 : 0;
assign detect_min[151][15] = (mid_1[1223:1216] < mid_2[1223:1216]) ? 1 : 0;
assign detect_min[151][16] = (mid_1[1223:1216] < mid_2[1231:1224]) ? 1 : 0;
assign detect_min[151][17] = (mid_1[1223:1216] < btm_0[1215:1208]) ? 1 : 0;
assign detect_min[151][18] = (mid_1[1223:1216] < btm_0[1223:1216]) ? 1 : 0;
assign detect_min[151][19] = (mid_1[1223:1216] < btm_0[1231:1224]) ? 1 : 0;
assign detect_min[151][20] = (mid_1[1223:1216] < btm_1[1215:1208]) ? 1 : 0;
assign detect_min[151][21] = (mid_1[1223:1216] < btm_1[1223:1216]) ? 1 : 0;
assign detect_min[151][22] = (mid_1[1223:1216] < btm_1[1231:1224]) ? 1 : 0;
assign detect_min[151][23] = (mid_1[1223:1216] < btm_2[1215:1208]) ? 1 : 0;
assign detect_min[151][24] = (mid_1[1223:1216] < btm_2[1223:1216]) ? 1 : 0;
assign detect_min[151][25] = (mid_1[1223:1216] < btm_2[1231:1224]) ? 1 : 0;

assign detect_min[152][0] = (mid_1[1231:1224] < top_0[1223:1216]) ? 1 : 0;
assign detect_min[152][1] = (mid_1[1231:1224] < top_0[1231:1224]) ? 1 : 0;
assign detect_min[152][2] = (mid_1[1231:1224] < top_0[1239:1232]) ? 1 : 0;
assign detect_min[152][3] = (mid_1[1231:1224] < top_1[1223:1216]) ? 1 : 0;
assign detect_min[152][4] = (mid_1[1231:1224] < top_1[1231:1224]) ? 1 : 0;
assign detect_min[152][5] = (mid_1[1231:1224] < top_1[1239:1232]) ? 1 : 0;
assign detect_min[152][6] = (mid_1[1231:1224] < top_2[1223:1216]) ? 1 : 0;
assign detect_min[152][7] = (mid_1[1231:1224] < top_2[1231:1224]) ? 1 : 0;
assign detect_min[152][8] = (mid_1[1231:1224] < top_2[1239:1232]) ? 1 : 0;
assign detect_min[152][9] = (mid_1[1231:1224] < mid_0[1223:1216]) ? 1 : 0;
assign detect_min[152][10] = (mid_1[1231:1224] < mid_0[1231:1224]) ? 1 : 0;
assign detect_min[152][11] = (mid_1[1231:1224] < mid_0[1239:1232]) ? 1 : 0;
assign detect_min[152][12] = (mid_1[1231:1224] < mid_1[1223:1216]) ? 1 : 0;
assign detect_min[152][13] = (mid_1[1231:1224] < mid_1[1239:1232]) ? 1 : 0;
assign detect_min[152][14] = (mid_1[1231:1224] < mid_2[1223:1216]) ? 1 : 0;
assign detect_min[152][15] = (mid_1[1231:1224] < mid_2[1231:1224]) ? 1 : 0;
assign detect_min[152][16] = (mid_1[1231:1224] < mid_2[1239:1232]) ? 1 : 0;
assign detect_min[152][17] = (mid_1[1231:1224] < btm_0[1223:1216]) ? 1 : 0;
assign detect_min[152][18] = (mid_1[1231:1224] < btm_0[1231:1224]) ? 1 : 0;
assign detect_min[152][19] = (mid_1[1231:1224] < btm_0[1239:1232]) ? 1 : 0;
assign detect_min[152][20] = (mid_1[1231:1224] < btm_1[1223:1216]) ? 1 : 0;
assign detect_min[152][21] = (mid_1[1231:1224] < btm_1[1231:1224]) ? 1 : 0;
assign detect_min[152][22] = (mid_1[1231:1224] < btm_1[1239:1232]) ? 1 : 0;
assign detect_min[152][23] = (mid_1[1231:1224] < btm_2[1223:1216]) ? 1 : 0;
assign detect_min[152][24] = (mid_1[1231:1224] < btm_2[1231:1224]) ? 1 : 0;
assign detect_min[152][25] = (mid_1[1231:1224] < btm_2[1239:1232]) ? 1 : 0;

assign detect_min[153][0] = (mid_1[1239:1232] < top_0[1231:1224]) ? 1 : 0;
assign detect_min[153][1] = (mid_1[1239:1232] < top_0[1239:1232]) ? 1 : 0;
assign detect_min[153][2] = (mid_1[1239:1232] < top_0[1247:1240]) ? 1 : 0;
assign detect_min[153][3] = (mid_1[1239:1232] < top_1[1231:1224]) ? 1 : 0;
assign detect_min[153][4] = (mid_1[1239:1232] < top_1[1239:1232]) ? 1 : 0;
assign detect_min[153][5] = (mid_1[1239:1232] < top_1[1247:1240]) ? 1 : 0;
assign detect_min[153][6] = (mid_1[1239:1232] < top_2[1231:1224]) ? 1 : 0;
assign detect_min[153][7] = (mid_1[1239:1232] < top_2[1239:1232]) ? 1 : 0;
assign detect_min[153][8] = (mid_1[1239:1232] < top_2[1247:1240]) ? 1 : 0;
assign detect_min[153][9] = (mid_1[1239:1232] < mid_0[1231:1224]) ? 1 : 0;
assign detect_min[153][10] = (mid_1[1239:1232] < mid_0[1239:1232]) ? 1 : 0;
assign detect_min[153][11] = (mid_1[1239:1232] < mid_0[1247:1240]) ? 1 : 0;
assign detect_min[153][12] = (mid_1[1239:1232] < mid_1[1231:1224]) ? 1 : 0;
assign detect_min[153][13] = (mid_1[1239:1232] < mid_1[1247:1240]) ? 1 : 0;
assign detect_min[153][14] = (mid_1[1239:1232] < mid_2[1231:1224]) ? 1 : 0;
assign detect_min[153][15] = (mid_1[1239:1232] < mid_2[1239:1232]) ? 1 : 0;
assign detect_min[153][16] = (mid_1[1239:1232] < mid_2[1247:1240]) ? 1 : 0;
assign detect_min[153][17] = (mid_1[1239:1232] < btm_0[1231:1224]) ? 1 : 0;
assign detect_min[153][18] = (mid_1[1239:1232] < btm_0[1239:1232]) ? 1 : 0;
assign detect_min[153][19] = (mid_1[1239:1232] < btm_0[1247:1240]) ? 1 : 0;
assign detect_min[153][20] = (mid_1[1239:1232] < btm_1[1231:1224]) ? 1 : 0;
assign detect_min[153][21] = (mid_1[1239:1232] < btm_1[1239:1232]) ? 1 : 0;
assign detect_min[153][22] = (mid_1[1239:1232] < btm_1[1247:1240]) ? 1 : 0;
assign detect_min[153][23] = (mid_1[1239:1232] < btm_2[1231:1224]) ? 1 : 0;
assign detect_min[153][24] = (mid_1[1239:1232] < btm_2[1239:1232]) ? 1 : 0;
assign detect_min[153][25] = (mid_1[1239:1232] < btm_2[1247:1240]) ? 1 : 0;

assign detect_min[154][0] = (mid_1[1247:1240] < top_0[1239:1232]) ? 1 : 0;
assign detect_min[154][1] = (mid_1[1247:1240] < top_0[1247:1240]) ? 1 : 0;
assign detect_min[154][2] = (mid_1[1247:1240] < top_0[1255:1248]) ? 1 : 0;
assign detect_min[154][3] = (mid_1[1247:1240] < top_1[1239:1232]) ? 1 : 0;
assign detect_min[154][4] = (mid_1[1247:1240] < top_1[1247:1240]) ? 1 : 0;
assign detect_min[154][5] = (mid_1[1247:1240] < top_1[1255:1248]) ? 1 : 0;
assign detect_min[154][6] = (mid_1[1247:1240] < top_2[1239:1232]) ? 1 : 0;
assign detect_min[154][7] = (mid_1[1247:1240] < top_2[1247:1240]) ? 1 : 0;
assign detect_min[154][8] = (mid_1[1247:1240] < top_2[1255:1248]) ? 1 : 0;
assign detect_min[154][9] = (mid_1[1247:1240] < mid_0[1239:1232]) ? 1 : 0;
assign detect_min[154][10] = (mid_1[1247:1240] < mid_0[1247:1240]) ? 1 : 0;
assign detect_min[154][11] = (mid_1[1247:1240] < mid_0[1255:1248]) ? 1 : 0;
assign detect_min[154][12] = (mid_1[1247:1240] < mid_1[1239:1232]) ? 1 : 0;
assign detect_min[154][13] = (mid_1[1247:1240] < mid_1[1255:1248]) ? 1 : 0;
assign detect_min[154][14] = (mid_1[1247:1240] < mid_2[1239:1232]) ? 1 : 0;
assign detect_min[154][15] = (mid_1[1247:1240] < mid_2[1247:1240]) ? 1 : 0;
assign detect_min[154][16] = (mid_1[1247:1240] < mid_2[1255:1248]) ? 1 : 0;
assign detect_min[154][17] = (mid_1[1247:1240] < btm_0[1239:1232]) ? 1 : 0;
assign detect_min[154][18] = (mid_1[1247:1240] < btm_0[1247:1240]) ? 1 : 0;
assign detect_min[154][19] = (mid_1[1247:1240] < btm_0[1255:1248]) ? 1 : 0;
assign detect_min[154][20] = (mid_1[1247:1240] < btm_1[1239:1232]) ? 1 : 0;
assign detect_min[154][21] = (mid_1[1247:1240] < btm_1[1247:1240]) ? 1 : 0;
assign detect_min[154][22] = (mid_1[1247:1240] < btm_1[1255:1248]) ? 1 : 0;
assign detect_min[154][23] = (mid_1[1247:1240] < btm_2[1239:1232]) ? 1 : 0;
assign detect_min[154][24] = (mid_1[1247:1240] < btm_2[1247:1240]) ? 1 : 0;
assign detect_min[154][25] = (mid_1[1247:1240] < btm_2[1255:1248]) ? 1 : 0;

assign detect_min[155][0] = (mid_1[1255:1248] < top_0[1247:1240]) ? 1 : 0;
assign detect_min[155][1] = (mid_1[1255:1248] < top_0[1255:1248]) ? 1 : 0;
assign detect_min[155][2] = (mid_1[1255:1248] < top_0[1263:1256]) ? 1 : 0;
assign detect_min[155][3] = (mid_1[1255:1248] < top_1[1247:1240]) ? 1 : 0;
assign detect_min[155][4] = (mid_1[1255:1248] < top_1[1255:1248]) ? 1 : 0;
assign detect_min[155][5] = (mid_1[1255:1248] < top_1[1263:1256]) ? 1 : 0;
assign detect_min[155][6] = (mid_1[1255:1248] < top_2[1247:1240]) ? 1 : 0;
assign detect_min[155][7] = (mid_1[1255:1248] < top_2[1255:1248]) ? 1 : 0;
assign detect_min[155][8] = (mid_1[1255:1248] < top_2[1263:1256]) ? 1 : 0;
assign detect_min[155][9] = (mid_1[1255:1248] < mid_0[1247:1240]) ? 1 : 0;
assign detect_min[155][10] = (mid_1[1255:1248] < mid_0[1255:1248]) ? 1 : 0;
assign detect_min[155][11] = (mid_1[1255:1248] < mid_0[1263:1256]) ? 1 : 0;
assign detect_min[155][12] = (mid_1[1255:1248] < mid_1[1247:1240]) ? 1 : 0;
assign detect_min[155][13] = (mid_1[1255:1248] < mid_1[1263:1256]) ? 1 : 0;
assign detect_min[155][14] = (mid_1[1255:1248] < mid_2[1247:1240]) ? 1 : 0;
assign detect_min[155][15] = (mid_1[1255:1248] < mid_2[1255:1248]) ? 1 : 0;
assign detect_min[155][16] = (mid_1[1255:1248] < mid_2[1263:1256]) ? 1 : 0;
assign detect_min[155][17] = (mid_1[1255:1248] < btm_0[1247:1240]) ? 1 : 0;
assign detect_min[155][18] = (mid_1[1255:1248] < btm_0[1255:1248]) ? 1 : 0;
assign detect_min[155][19] = (mid_1[1255:1248] < btm_0[1263:1256]) ? 1 : 0;
assign detect_min[155][20] = (mid_1[1255:1248] < btm_1[1247:1240]) ? 1 : 0;
assign detect_min[155][21] = (mid_1[1255:1248] < btm_1[1255:1248]) ? 1 : 0;
assign detect_min[155][22] = (mid_1[1255:1248] < btm_1[1263:1256]) ? 1 : 0;
assign detect_min[155][23] = (mid_1[1255:1248] < btm_2[1247:1240]) ? 1 : 0;
assign detect_min[155][24] = (mid_1[1255:1248] < btm_2[1255:1248]) ? 1 : 0;
assign detect_min[155][25] = (mid_1[1255:1248] < btm_2[1263:1256]) ? 1 : 0;

assign detect_min[156][0] = (mid_1[1263:1256] < top_0[1255:1248]) ? 1 : 0;
assign detect_min[156][1] = (mid_1[1263:1256] < top_0[1263:1256]) ? 1 : 0;
assign detect_min[156][2] = (mid_1[1263:1256] < top_0[1271:1264]) ? 1 : 0;
assign detect_min[156][3] = (mid_1[1263:1256] < top_1[1255:1248]) ? 1 : 0;
assign detect_min[156][4] = (mid_1[1263:1256] < top_1[1263:1256]) ? 1 : 0;
assign detect_min[156][5] = (mid_1[1263:1256] < top_1[1271:1264]) ? 1 : 0;
assign detect_min[156][6] = (mid_1[1263:1256] < top_2[1255:1248]) ? 1 : 0;
assign detect_min[156][7] = (mid_1[1263:1256] < top_2[1263:1256]) ? 1 : 0;
assign detect_min[156][8] = (mid_1[1263:1256] < top_2[1271:1264]) ? 1 : 0;
assign detect_min[156][9] = (mid_1[1263:1256] < mid_0[1255:1248]) ? 1 : 0;
assign detect_min[156][10] = (mid_1[1263:1256] < mid_0[1263:1256]) ? 1 : 0;
assign detect_min[156][11] = (mid_1[1263:1256] < mid_0[1271:1264]) ? 1 : 0;
assign detect_min[156][12] = (mid_1[1263:1256] < mid_1[1255:1248]) ? 1 : 0;
assign detect_min[156][13] = (mid_1[1263:1256] < mid_1[1271:1264]) ? 1 : 0;
assign detect_min[156][14] = (mid_1[1263:1256] < mid_2[1255:1248]) ? 1 : 0;
assign detect_min[156][15] = (mid_1[1263:1256] < mid_2[1263:1256]) ? 1 : 0;
assign detect_min[156][16] = (mid_1[1263:1256] < mid_2[1271:1264]) ? 1 : 0;
assign detect_min[156][17] = (mid_1[1263:1256] < btm_0[1255:1248]) ? 1 : 0;
assign detect_min[156][18] = (mid_1[1263:1256] < btm_0[1263:1256]) ? 1 : 0;
assign detect_min[156][19] = (mid_1[1263:1256] < btm_0[1271:1264]) ? 1 : 0;
assign detect_min[156][20] = (mid_1[1263:1256] < btm_1[1255:1248]) ? 1 : 0;
assign detect_min[156][21] = (mid_1[1263:1256] < btm_1[1263:1256]) ? 1 : 0;
assign detect_min[156][22] = (mid_1[1263:1256] < btm_1[1271:1264]) ? 1 : 0;
assign detect_min[156][23] = (mid_1[1263:1256] < btm_2[1255:1248]) ? 1 : 0;
assign detect_min[156][24] = (mid_1[1263:1256] < btm_2[1263:1256]) ? 1 : 0;
assign detect_min[156][25] = (mid_1[1263:1256] < btm_2[1271:1264]) ? 1 : 0;

assign detect_min[157][0] = (mid_1[1271:1264] < top_0[1263:1256]) ? 1 : 0;
assign detect_min[157][1] = (mid_1[1271:1264] < top_0[1271:1264]) ? 1 : 0;
assign detect_min[157][2] = (mid_1[1271:1264] < top_0[1279:1272]) ? 1 : 0;
assign detect_min[157][3] = (mid_1[1271:1264] < top_1[1263:1256]) ? 1 : 0;
assign detect_min[157][4] = (mid_1[1271:1264] < top_1[1271:1264]) ? 1 : 0;
assign detect_min[157][5] = (mid_1[1271:1264] < top_1[1279:1272]) ? 1 : 0;
assign detect_min[157][6] = (mid_1[1271:1264] < top_2[1263:1256]) ? 1 : 0;
assign detect_min[157][7] = (mid_1[1271:1264] < top_2[1271:1264]) ? 1 : 0;
assign detect_min[157][8] = (mid_1[1271:1264] < top_2[1279:1272]) ? 1 : 0;
assign detect_min[157][9] = (mid_1[1271:1264] < mid_0[1263:1256]) ? 1 : 0;
assign detect_min[157][10] = (mid_1[1271:1264] < mid_0[1271:1264]) ? 1 : 0;
assign detect_min[157][11] = (mid_1[1271:1264] < mid_0[1279:1272]) ? 1 : 0;
assign detect_min[157][12] = (mid_1[1271:1264] < mid_1[1263:1256]) ? 1 : 0;
assign detect_min[157][13] = (mid_1[1271:1264] < mid_1[1279:1272]) ? 1 : 0;
assign detect_min[157][14] = (mid_1[1271:1264] < mid_2[1263:1256]) ? 1 : 0;
assign detect_min[157][15] = (mid_1[1271:1264] < mid_2[1271:1264]) ? 1 : 0;
assign detect_min[157][16] = (mid_1[1271:1264] < mid_2[1279:1272]) ? 1 : 0;
assign detect_min[157][17] = (mid_1[1271:1264] < btm_0[1263:1256]) ? 1 : 0;
assign detect_min[157][18] = (mid_1[1271:1264] < btm_0[1271:1264]) ? 1 : 0;
assign detect_min[157][19] = (mid_1[1271:1264] < btm_0[1279:1272]) ? 1 : 0;
assign detect_min[157][20] = (mid_1[1271:1264] < btm_1[1263:1256]) ? 1 : 0;
assign detect_min[157][21] = (mid_1[1271:1264] < btm_1[1271:1264]) ? 1 : 0;
assign detect_min[157][22] = (mid_1[1271:1264] < btm_1[1279:1272]) ? 1 : 0;
assign detect_min[157][23] = (mid_1[1271:1264] < btm_2[1263:1256]) ? 1 : 0;
assign detect_min[157][24] = (mid_1[1271:1264] < btm_2[1271:1264]) ? 1 : 0;
assign detect_min[157][25] = (mid_1[1271:1264] < btm_2[1279:1272]) ? 1 : 0;

assign detect_min[158][0] = (mid_1[1279:1272] < top_0[1271:1264]) ? 1 : 0;
assign detect_min[158][1] = (mid_1[1279:1272] < top_0[1279:1272]) ? 1 : 0;
assign detect_min[158][2] = (mid_1[1279:1272] < top_0[1287:1280]) ? 1 : 0;
assign detect_min[158][3] = (mid_1[1279:1272] < top_1[1271:1264]) ? 1 : 0;
assign detect_min[158][4] = (mid_1[1279:1272] < top_1[1279:1272]) ? 1 : 0;
assign detect_min[158][5] = (mid_1[1279:1272] < top_1[1287:1280]) ? 1 : 0;
assign detect_min[158][6] = (mid_1[1279:1272] < top_2[1271:1264]) ? 1 : 0;
assign detect_min[158][7] = (mid_1[1279:1272] < top_2[1279:1272]) ? 1 : 0;
assign detect_min[158][8] = (mid_1[1279:1272] < top_2[1287:1280]) ? 1 : 0;
assign detect_min[158][9] = (mid_1[1279:1272] < mid_0[1271:1264]) ? 1 : 0;
assign detect_min[158][10] = (mid_1[1279:1272] < mid_0[1279:1272]) ? 1 : 0;
assign detect_min[158][11] = (mid_1[1279:1272] < mid_0[1287:1280]) ? 1 : 0;
assign detect_min[158][12] = (mid_1[1279:1272] < mid_1[1271:1264]) ? 1 : 0;
assign detect_min[158][13] = (mid_1[1279:1272] < mid_1[1287:1280]) ? 1 : 0;
assign detect_min[158][14] = (mid_1[1279:1272] < mid_2[1271:1264]) ? 1 : 0;
assign detect_min[158][15] = (mid_1[1279:1272] < mid_2[1279:1272]) ? 1 : 0;
assign detect_min[158][16] = (mid_1[1279:1272] < mid_2[1287:1280]) ? 1 : 0;
assign detect_min[158][17] = (mid_1[1279:1272] < btm_0[1271:1264]) ? 1 : 0;
assign detect_min[158][18] = (mid_1[1279:1272] < btm_0[1279:1272]) ? 1 : 0;
assign detect_min[158][19] = (mid_1[1279:1272] < btm_0[1287:1280]) ? 1 : 0;
assign detect_min[158][20] = (mid_1[1279:1272] < btm_1[1271:1264]) ? 1 : 0;
assign detect_min[158][21] = (mid_1[1279:1272] < btm_1[1279:1272]) ? 1 : 0;
assign detect_min[158][22] = (mid_1[1279:1272] < btm_1[1287:1280]) ? 1 : 0;
assign detect_min[158][23] = (mid_1[1279:1272] < btm_2[1271:1264]) ? 1 : 0;
assign detect_min[158][24] = (mid_1[1279:1272] < btm_2[1279:1272]) ? 1 : 0;
assign detect_min[158][25] = (mid_1[1279:1272] < btm_2[1287:1280]) ? 1 : 0;

assign detect_min[159][0] = (mid_1[1287:1280] < top_0[1279:1272]) ? 1 : 0;
assign detect_min[159][1] = (mid_1[1287:1280] < top_0[1287:1280]) ? 1 : 0;
assign detect_min[159][2] = (mid_1[1287:1280] < top_0[1295:1288]) ? 1 : 0;
assign detect_min[159][3] = (mid_1[1287:1280] < top_1[1279:1272]) ? 1 : 0;
assign detect_min[159][4] = (mid_1[1287:1280] < top_1[1287:1280]) ? 1 : 0;
assign detect_min[159][5] = (mid_1[1287:1280] < top_1[1295:1288]) ? 1 : 0;
assign detect_min[159][6] = (mid_1[1287:1280] < top_2[1279:1272]) ? 1 : 0;
assign detect_min[159][7] = (mid_1[1287:1280] < top_2[1287:1280]) ? 1 : 0;
assign detect_min[159][8] = (mid_1[1287:1280] < top_2[1295:1288]) ? 1 : 0;
assign detect_min[159][9] = (mid_1[1287:1280] < mid_0[1279:1272]) ? 1 : 0;
assign detect_min[159][10] = (mid_1[1287:1280] < mid_0[1287:1280]) ? 1 : 0;
assign detect_min[159][11] = (mid_1[1287:1280] < mid_0[1295:1288]) ? 1 : 0;
assign detect_min[159][12] = (mid_1[1287:1280] < mid_1[1279:1272]) ? 1 : 0;
assign detect_min[159][13] = (mid_1[1287:1280] < mid_1[1295:1288]) ? 1 : 0;
assign detect_min[159][14] = (mid_1[1287:1280] < mid_2[1279:1272]) ? 1 : 0;
assign detect_min[159][15] = (mid_1[1287:1280] < mid_2[1287:1280]) ? 1 : 0;
assign detect_min[159][16] = (mid_1[1287:1280] < mid_2[1295:1288]) ? 1 : 0;
assign detect_min[159][17] = (mid_1[1287:1280] < btm_0[1279:1272]) ? 1 : 0;
assign detect_min[159][18] = (mid_1[1287:1280] < btm_0[1287:1280]) ? 1 : 0;
assign detect_min[159][19] = (mid_1[1287:1280] < btm_0[1295:1288]) ? 1 : 0;
assign detect_min[159][20] = (mid_1[1287:1280] < btm_1[1279:1272]) ? 1 : 0;
assign detect_min[159][21] = (mid_1[1287:1280] < btm_1[1287:1280]) ? 1 : 0;
assign detect_min[159][22] = (mid_1[1287:1280] < btm_1[1295:1288]) ? 1 : 0;
assign detect_min[159][23] = (mid_1[1287:1280] < btm_2[1279:1272]) ? 1 : 0;
assign detect_min[159][24] = (mid_1[1287:1280] < btm_2[1287:1280]) ? 1 : 0;
assign detect_min[159][25] = (mid_1[1287:1280] < btm_2[1295:1288]) ? 1 : 0;

assign detect_min[160][0] = (mid_1[1295:1288] < top_0[1287:1280]) ? 1 : 0;
assign detect_min[160][1] = (mid_1[1295:1288] < top_0[1295:1288]) ? 1 : 0;
assign detect_min[160][2] = (mid_1[1295:1288] < top_0[1303:1296]) ? 1 : 0;
assign detect_min[160][3] = (mid_1[1295:1288] < top_1[1287:1280]) ? 1 : 0;
assign detect_min[160][4] = (mid_1[1295:1288] < top_1[1295:1288]) ? 1 : 0;
assign detect_min[160][5] = (mid_1[1295:1288] < top_1[1303:1296]) ? 1 : 0;
assign detect_min[160][6] = (mid_1[1295:1288] < top_2[1287:1280]) ? 1 : 0;
assign detect_min[160][7] = (mid_1[1295:1288] < top_2[1295:1288]) ? 1 : 0;
assign detect_min[160][8] = (mid_1[1295:1288] < top_2[1303:1296]) ? 1 : 0;
assign detect_min[160][9] = (mid_1[1295:1288] < mid_0[1287:1280]) ? 1 : 0;
assign detect_min[160][10] = (mid_1[1295:1288] < mid_0[1295:1288]) ? 1 : 0;
assign detect_min[160][11] = (mid_1[1295:1288] < mid_0[1303:1296]) ? 1 : 0;
assign detect_min[160][12] = (mid_1[1295:1288] < mid_1[1287:1280]) ? 1 : 0;
assign detect_min[160][13] = (mid_1[1295:1288] < mid_1[1303:1296]) ? 1 : 0;
assign detect_min[160][14] = (mid_1[1295:1288] < mid_2[1287:1280]) ? 1 : 0;
assign detect_min[160][15] = (mid_1[1295:1288] < mid_2[1295:1288]) ? 1 : 0;
assign detect_min[160][16] = (mid_1[1295:1288] < mid_2[1303:1296]) ? 1 : 0;
assign detect_min[160][17] = (mid_1[1295:1288] < btm_0[1287:1280]) ? 1 : 0;
assign detect_min[160][18] = (mid_1[1295:1288] < btm_0[1295:1288]) ? 1 : 0;
assign detect_min[160][19] = (mid_1[1295:1288] < btm_0[1303:1296]) ? 1 : 0;
assign detect_min[160][20] = (mid_1[1295:1288] < btm_1[1287:1280]) ? 1 : 0;
assign detect_min[160][21] = (mid_1[1295:1288] < btm_1[1295:1288]) ? 1 : 0;
assign detect_min[160][22] = (mid_1[1295:1288] < btm_1[1303:1296]) ? 1 : 0;
assign detect_min[160][23] = (mid_1[1295:1288] < btm_2[1287:1280]) ? 1 : 0;
assign detect_min[160][24] = (mid_1[1295:1288] < btm_2[1295:1288]) ? 1 : 0;
assign detect_min[160][25] = (mid_1[1295:1288] < btm_2[1303:1296]) ? 1 : 0;

assign detect_min[161][0] = (mid_1[1303:1296] < top_0[1295:1288]) ? 1 : 0;
assign detect_min[161][1] = (mid_1[1303:1296] < top_0[1303:1296]) ? 1 : 0;
assign detect_min[161][2] = (mid_1[1303:1296] < top_0[1311:1304]) ? 1 : 0;
assign detect_min[161][3] = (mid_1[1303:1296] < top_1[1295:1288]) ? 1 : 0;
assign detect_min[161][4] = (mid_1[1303:1296] < top_1[1303:1296]) ? 1 : 0;
assign detect_min[161][5] = (mid_1[1303:1296] < top_1[1311:1304]) ? 1 : 0;
assign detect_min[161][6] = (mid_1[1303:1296] < top_2[1295:1288]) ? 1 : 0;
assign detect_min[161][7] = (mid_1[1303:1296] < top_2[1303:1296]) ? 1 : 0;
assign detect_min[161][8] = (mid_1[1303:1296] < top_2[1311:1304]) ? 1 : 0;
assign detect_min[161][9] = (mid_1[1303:1296] < mid_0[1295:1288]) ? 1 : 0;
assign detect_min[161][10] = (mid_1[1303:1296] < mid_0[1303:1296]) ? 1 : 0;
assign detect_min[161][11] = (mid_1[1303:1296] < mid_0[1311:1304]) ? 1 : 0;
assign detect_min[161][12] = (mid_1[1303:1296] < mid_1[1295:1288]) ? 1 : 0;
assign detect_min[161][13] = (mid_1[1303:1296] < mid_1[1311:1304]) ? 1 : 0;
assign detect_min[161][14] = (mid_1[1303:1296] < mid_2[1295:1288]) ? 1 : 0;
assign detect_min[161][15] = (mid_1[1303:1296] < mid_2[1303:1296]) ? 1 : 0;
assign detect_min[161][16] = (mid_1[1303:1296] < mid_2[1311:1304]) ? 1 : 0;
assign detect_min[161][17] = (mid_1[1303:1296] < btm_0[1295:1288]) ? 1 : 0;
assign detect_min[161][18] = (mid_1[1303:1296] < btm_0[1303:1296]) ? 1 : 0;
assign detect_min[161][19] = (mid_1[1303:1296] < btm_0[1311:1304]) ? 1 : 0;
assign detect_min[161][20] = (mid_1[1303:1296] < btm_1[1295:1288]) ? 1 : 0;
assign detect_min[161][21] = (mid_1[1303:1296] < btm_1[1303:1296]) ? 1 : 0;
assign detect_min[161][22] = (mid_1[1303:1296] < btm_1[1311:1304]) ? 1 : 0;
assign detect_min[161][23] = (mid_1[1303:1296] < btm_2[1295:1288]) ? 1 : 0;
assign detect_min[161][24] = (mid_1[1303:1296] < btm_2[1303:1296]) ? 1 : 0;
assign detect_min[161][25] = (mid_1[1303:1296] < btm_2[1311:1304]) ? 1 : 0;

assign detect_min[162][0] = (mid_1[1311:1304] < top_0[1303:1296]) ? 1 : 0;
assign detect_min[162][1] = (mid_1[1311:1304] < top_0[1311:1304]) ? 1 : 0;
assign detect_min[162][2] = (mid_1[1311:1304] < top_0[1319:1312]) ? 1 : 0;
assign detect_min[162][3] = (mid_1[1311:1304] < top_1[1303:1296]) ? 1 : 0;
assign detect_min[162][4] = (mid_1[1311:1304] < top_1[1311:1304]) ? 1 : 0;
assign detect_min[162][5] = (mid_1[1311:1304] < top_1[1319:1312]) ? 1 : 0;
assign detect_min[162][6] = (mid_1[1311:1304] < top_2[1303:1296]) ? 1 : 0;
assign detect_min[162][7] = (mid_1[1311:1304] < top_2[1311:1304]) ? 1 : 0;
assign detect_min[162][8] = (mid_1[1311:1304] < top_2[1319:1312]) ? 1 : 0;
assign detect_min[162][9] = (mid_1[1311:1304] < mid_0[1303:1296]) ? 1 : 0;
assign detect_min[162][10] = (mid_1[1311:1304] < mid_0[1311:1304]) ? 1 : 0;
assign detect_min[162][11] = (mid_1[1311:1304] < mid_0[1319:1312]) ? 1 : 0;
assign detect_min[162][12] = (mid_1[1311:1304] < mid_1[1303:1296]) ? 1 : 0;
assign detect_min[162][13] = (mid_1[1311:1304] < mid_1[1319:1312]) ? 1 : 0;
assign detect_min[162][14] = (mid_1[1311:1304] < mid_2[1303:1296]) ? 1 : 0;
assign detect_min[162][15] = (mid_1[1311:1304] < mid_2[1311:1304]) ? 1 : 0;
assign detect_min[162][16] = (mid_1[1311:1304] < mid_2[1319:1312]) ? 1 : 0;
assign detect_min[162][17] = (mid_1[1311:1304] < btm_0[1303:1296]) ? 1 : 0;
assign detect_min[162][18] = (mid_1[1311:1304] < btm_0[1311:1304]) ? 1 : 0;
assign detect_min[162][19] = (mid_1[1311:1304] < btm_0[1319:1312]) ? 1 : 0;
assign detect_min[162][20] = (mid_1[1311:1304] < btm_1[1303:1296]) ? 1 : 0;
assign detect_min[162][21] = (mid_1[1311:1304] < btm_1[1311:1304]) ? 1 : 0;
assign detect_min[162][22] = (mid_1[1311:1304] < btm_1[1319:1312]) ? 1 : 0;
assign detect_min[162][23] = (mid_1[1311:1304] < btm_2[1303:1296]) ? 1 : 0;
assign detect_min[162][24] = (mid_1[1311:1304] < btm_2[1311:1304]) ? 1 : 0;
assign detect_min[162][25] = (mid_1[1311:1304] < btm_2[1319:1312]) ? 1 : 0;

assign detect_min[163][0] = (mid_1[1319:1312] < top_0[1311:1304]) ? 1 : 0;
assign detect_min[163][1] = (mid_1[1319:1312] < top_0[1319:1312]) ? 1 : 0;
assign detect_min[163][2] = (mid_1[1319:1312] < top_0[1327:1320]) ? 1 : 0;
assign detect_min[163][3] = (mid_1[1319:1312] < top_1[1311:1304]) ? 1 : 0;
assign detect_min[163][4] = (mid_1[1319:1312] < top_1[1319:1312]) ? 1 : 0;
assign detect_min[163][5] = (mid_1[1319:1312] < top_1[1327:1320]) ? 1 : 0;
assign detect_min[163][6] = (mid_1[1319:1312] < top_2[1311:1304]) ? 1 : 0;
assign detect_min[163][7] = (mid_1[1319:1312] < top_2[1319:1312]) ? 1 : 0;
assign detect_min[163][8] = (mid_1[1319:1312] < top_2[1327:1320]) ? 1 : 0;
assign detect_min[163][9] = (mid_1[1319:1312] < mid_0[1311:1304]) ? 1 : 0;
assign detect_min[163][10] = (mid_1[1319:1312] < mid_0[1319:1312]) ? 1 : 0;
assign detect_min[163][11] = (mid_1[1319:1312] < mid_0[1327:1320]) ? 1 : 0;
assign detect_min[163][12] = (mid_1[1319:1312] < mid_1[1311:1304]) ? 1 : 0;
assign detect_min[163][13] = (mid_1[1319:1312] < mid_1[1327:1320]) ? 1 : 0;
assign detect_min[163][14] = (mid_1[1319:1312] < mid_2[1311:1304]) ? 1 : 0;
assign detect_min[163][15] = (mid_1[1319:1312] < mid_2[1319:1312]) ? 1 : 0;
assign detect_min[163][16] = (mid_1[1319:1312] < mid_2[1327:1320]) ? 1 : 0;
assign detect_min[163][17] = (mid_1[1319:1312] < btm_0[1311:1304]) ? 1 : 0;
assign detect_min[163][18] = (mid_1[1319:1312] < btm_0[1319:1312]) ? 1 : 0;
assign detect_min[163][19] = (mid_1[1319:1312] < btm_0[1327:1320]) ? 1 : 0;
assign detect_min[163][20] = (mid_1[1319:1312] < btm_1[1311:1304]) ? 1 : 0;
assign detect_min[163][21] = (mid_1[1319:1312] < btm_1[1319:1312]) ? 1 : 0;
assign detect_min[163][22] = (mid_1[1319:1312] < btm_1[1327:1320]) ? 1 : 0;
assign detect_min[163][23] = (mid_1[1319:1312] < btm_2[1311:1304]) ? 1 : 0;
assign detect_min[163][24] = (mid_1[1319:1312] < btm_2[1319:1312]) ? 1 : 0;
assign detect_min[163][25] = (mid_1[1319:1312] < btm_2[1327:1320]) ? 1 : 0;

assign detect_min[164][0] = (mid_1[1327:1320] < top_0[1319:1312]) ? 1 : 0;
assign detect_min[164][1] = (mid_1[1327:1320] < top_0[1327:1320]) ? 1 : 0;
assign detect_min[164][2] = (mid_1[1327:1320] < top_0[1335:1328]) ? 1 : 0;
assign detect_min[164][3] = (mid_1[1327:1320] < top_1[1319:1312]) ? 1 : 0;
assign detect_min[164][4] = (mid_1[1327:1320] < top_1[1327:1320]) ? 1 : 0;
assign detect_min[164][5] = (mid_1[1327:1320] < top_1[1335:1328]) ? 1 : 0;
assign detect_min[164][6] = (mid_1[1327:1320] < top_2[1319:1312]) ? 1 : 0;
assign detect_min[164][7] = (mid_1[1327:1320] < top_2[1327:1320]) ? 1 : 0;
assign detect_min[164][8] = (mid_1[1327:1320] < top_2[1335:1328]) ? 1 : 0;
assign detect_min[164][9] = (mid_1[1327:1320] < mid_0[1319:1312]) ? 1 : 0;
assign detect_min[164][10] = (mid_1[1327:1320] < mid_0[1327:1320]) ? 1 : 0;
assign detect_min[164][11] = (mid_1[1327:1320] < mid_0[1335:1328]) ? 1 : 0;
assign detect_min[164][12] = (mid_1[1327:1320] < mid_1[1319:1312]) ? 1 : 0;
assign detect_min[164][13] = (mid_1[1327:1320] < mid_1[1335:1328]) ? 1 : 0;
assign detect_min[164][14] = (mid_1[1327:1320] < mid_2[1319:1312]) ? 1 : 0;
assign detect_min[164][15] = (mid_1[1327:1320] < mid_2[1327:1320]) ? 1 : 0;
assign detect_min[164][16] = (mid_1[1327:1320] < mid_2[1335:1328]) ? 1 : 0;
assign detect_min[164][17] = (mid_1[1327:1320] < btm_0[1319:1312]) ? 1 : 0;
assign detect_min[164][18] = (mid_1[1327:1320] < btm_0[1327:1320]) ? 1 : 0;
assign detect_min[164][19] = (mid_1[1327:1320] < btm_0[1335:1328]) ? 1 : 0;
assign detect_min[164][20] = (mid_1[1327:1320] < btm_1[1319:1312]) ? 1 : 0;
assign detect_min[164][21] = (mid_1[1327:1320] < btm_1[1327:1320]) ? 1 : 0;
assign detect_min[164][22] = (mid_1[1327:1320] < btm_1[1335:1328]) ? 1 : 0;
assign detect_min[164][23] = (mid_1[1327:1320] < btm_2[1319:1312]) ? 1 : 0;
assign detect_min[164][24] = (mid_1[1327:1320] < btm_2[1327:1320]) ? 1 : 0;
assign detect_min[164][25] = (mid_1[1327:1320] < btm_2[1335:1328]) ? 1 : 0;

assign detect_min[165][0] = (mid_1[1335:1328] < top_0[1327:1320]) ? 1 : 0;
assign detect_min[165][1] = (mid_1[1335:1328] < top_0[1335:1328]) ? 1 : 0;
assign detect_min[165][2] = (mid_1[1335:1328] < top_0[1343:1336]) ? 1 : 0;
assign detect_min[165][3] = (mid_1[1335:1328] < top_1[1327:1320]) ? 1 : 0;
assign detect_min[165][4] = (mid_1[1335:1328] < top_1[1335:1328]) ? 1 : 0;
assign detect_min[165][5] = (mid_1[1335:1328] < top_1[1343:1336]) ? 1 : 0;
assign detect_min[165][6] = (mid_1[1335:1328] < top_2[1327:1320]) ? 1 : 0;
assign detect_min[165][7] = (mid_1[1335:1328] < top_2[1335:1328]) ? 1 : 0;
assign detect_min[165][8] = (mid_1[1335:1328] < top_2[1343:1336]) ? 1 : 0;
assign detect_min[165][9] = (mid_1[1335:1328] < mid_0[1327:1320]) ? 1 : 0;
assign detect_min[165][10] = (mid_1[1335:1328] < mid_0[1335:1328]) ? 1 : 0;
assign detect_min[165][11] = (mid_1[1335:1328] < mid_0[1343:1336]) ? 1 : 0;
assign detect_min[165][12] = (mid_1[1335:1328] < mid_1[1327:1320]) ? 1 : 0;
assign detect_min[165][13] = (mid_1[1335:1328] < mid_1[1343:1336]) ? 1 : 0;
assign detect_min[165][14] = (mid_1[1335:1328] < mid_2[1327:1320]) ? 1 : 0;
assign detect_min[165][15] = (mid_1[1335:1328] < mid_2[1335:1328]) ? 1 : 0;
assign detect_min[165][16] = (mid_1[1335:1328] < mid_2[1343:1336]) ? 1 : 0;
assign detect_min[165][17] = (mid_1[1335:1328] < btm_0[1327:1320]) ? 1 : 0;
assign detect_min[165][18] = (mid_1[1335:1328] < btm_0[1335:1328]) ? 1 : 0;
assign detect_min[165][19] = (mid_1[1335:1328] < btm_0[1343:1336]) ? 1 : 0;
assign detect_min[165][20] = (mid_1[1335:1328] < btm_1[1327:1320]) ? 1 : 0;
assign detect_min[165][21] = (mid_1[1335:1328] < btm_1[1335:1328]) ? 1 : 0;
assign detect_min[165][22] = (mid_1[1335:1328] < btm_1[1343:1336]) ? 1 : 0;
assign detect_min[165][23] = (mid_1[1335:1328] < btm_2[1327:1320]) ? 1 : 0;
assign detect_min[165][24] = (mid_1[1335:1328] < btm_2[1335:1328]) ? 1 : 0;
assign detect_min[165][25] = (mid_1[1335:1328] < btm_2[1343:1336]) ? 1 : 0;

assign detect_min[166][0] = (mid_1[1343:1336] < top_0[1335:1328]) ? 1 : 0;
assign detect_min[166][1] = (mid_1[1343:1336] < top_0[1343:1336]) ? 1 : 0;
assign detect_min[166][2] = (mid_1[1343:1336] < top_0[1351:1344]) ? 1 : 0;
assign detect_min[166][3] = (mid_1[1343:1336] < top_1[1335:1328]) ? 1 : 0;
assign detect_min[166][4] = (mid_1[1343:1336] < top_1[1343:1336]) ? 1 : 0;
assign detect_min[166][5] = (mid_1[1343:1336] < top_1[1351:1344]) ? 1 : 0;
assign detect_min[166][6] = (mid_1[1343:1336] < top_2[1335:1328]) ? 1 : 0;
assign detect_min[166][7] = (mid_1[1343:1336] < top_2[1343:1336]) ? 1 : 0;
assign detect_min[166][8] = (mid_1[1343:1336] < top_2[1351:1344]) ? 1 : 0;
assign detect_min[166][9] = (mid_1[1343:1336] < mid_0[1335:1328]) ? 1 : 0;
assign detect_min[166][10] = (mid_1[1343:1336] < mid_0[1343:1336]) ? 1 : 0;
assign detect_min[166][11] = (mid_1[1343:1336] < mid_0[1351:1344]) ? 1 : 0;
assign detect_min[166][12] = (mid_1[1343:1336] < mid_1[1335:1328]) ? 1 : 0;
assign detect_min[166][13] = (mid_1[1343:1336] < mid_1[1351:1344]) ? 1 : 0;
assign detect_min[166][14] = (mid_1[1343:1336] < mid_2[1335:1328]) ? 1 : 0;
assign detect_min[166][15] = (mid_1[1343:1336] < mid_2[1343:1336]) ? 1 : 0;
assign detect_min[166][16] = (mid_1[1343:1336] < mid_2[1351:1344]) ? 1 : 0;
assign detect_min[166][17] = (mid_1[1343:1336] < btm_0[1335:1328]) ? 1 : 0;
assign detect_min[166][18] = (mid_1[1343:1336] < btm_0[1343:1336]) ? 1 : 0;
assign detect_min[166][19] = (mid_1[1343:1336] < btm_0[1351:1344]) ? 1 : 0;
assign detect_min[166][20] = (mid_1[1343:1336] < btm_1[1335:1328]) ? 1 : 0;
assign detect_min[166][21] = (mid_1[1343:1336] < btm_1[1343:1336]) ? 1 : 0;
assign detect_min[166][22] = (mid_1[1343:1336] < btm_1[1351:1344]) ? 1 : 0;
assign detect_min[166][23] = (mid_1[1343:1336] < btm_2[1335:1328]) ? 1 : 0;
assign detect_min[166][24] = (mid_1[1343:1336] < btm_2[1343:1336]) ? 1 : 0;
assign detect_min[166][25] = (mid_1[1343:1336] < btm_2[1351:1344]) ? 1 : 0;

assign detect_min[167][0] = (mid_1[1351:1344] < top_0[1343:1336]) ? 1 : 0;
assign detect_min[167][1] = (mid_1[1351:1344] < top_0[1351:1344]) ? 1 : 0;
assign detect_min[167][2] = (mid_1[1351:1344] < top_0[1359:1352]) ? 1 : 0;
assign detect_min[167][3] = (mid_1[1351:1344] < top_1[1343:1336]) ? 1 : 0;
assign detect_min[167][4] = (mid_1[1351:1344] < top_1[1351:1344]) ? 1 : 0;
assign detect_min[167][5] = (mid_1[1351:1344] < top_1[1359:1352]) ? 1 : 0;
assign detect_min[167][6] = (mid_1[1351:1344] < top_2[1343:1336]) ? 1 : 0;
assign detect_min[167][7] = (mid_1[1351:1344] < top_2[1351:1344]) ? 1 : 0;
assign detect_min[167][8] = (mid_1[1351:1344] < top_2[1359:1352]) ? 1 : 0;
assign detect_min[167][9] = (mid_1[1351:1344] < mid_0[1343:1336]) ? 1 : 0;
assign detect_min[167][10] = (mid_1[1351:1344] < mid_0[1351:1344]) ? 1 : 0;
assign detect_min[167][11] = (mid_1[1351:1344] < mid_0[1359:1352]) ? 1 : 0;
assign detect_min[167][12] = (mid_1[1351:1344] < mid_1[1343:1336]) ? 1 : 0;
assign detect_min[167][13] = (mid_1[1351:1344] < mid_1[1359:1352]) ? 1 : 0;
assign detect_min[167][14] = (mid_1[1351:1344] < mid_2[1343:1336]) ? 1 : 0;
assign detect_min[167][15] = (mid_1[1351:1344] < mid_2[1351:1344]) ? 1 : 0;
assign detect_min[167][16] = (mid_1[1351:1344] < mid_2[1359:1352]) ? 1 : 0;
assign detect_min[167][17] = (mid_1[1351:1344] < btm_0[1343:1336]) ? 1 : 0;
assign detect_min[167][18] = (mid_1[1351:1344] < btm_0[1351:1344]) ? 1 : 0;
assign detect_min[167][19] = (mid_1[1351:1344] < btm_0[1359:1352]) ? 1 : 0;
assign detect_min[167][20] = (mid_1[1351:1344] < btm_1[1343:1336]) ? 1 : 0;
assign detect_min[167][21] = (mid_1[1351:1344] < btm_1[1351:1344]) ? 1 : 0;
assign detect_min[167][22] = (mid_1[1351:1344] < btm_1[1359:1352]) ? 1 : 0;
assign detect_min[167][23] = (mid_1[1351:1344] < btm_2[1343:1336]) ? 1 : 0;
assign detect_min[167][24] = (mid_1[1351:1344] < btm_2[1351:1344]) ? 1 : 0;
assign detect_min[167][25] = (mid_1[1351:1344] < btm_2[1359:1352]) ? 1 : 0;

assign detect_min[168][0] = (mid_1[1359:1352] < top_0[1351:1344]) ? 1 : 0;
assign detect_min[168][1] = (mid_1[1359:1352] < top_0[1359:1352]) ? 1 : 0;
assign detect_min[168][2] = (mid_1[1359:1352] < top_0[1367:1360]) ? 1 : 0;
assign detect_min[168][3] = (mid_1[1359:1352] < top_1[1351:1344]) ? 1 : 0;
assign detect_min[168][4] = (mid_1[1359:1352] < top_1[1359:1352]) ? 1 : 0;
assign detect_min[168][5] = (mid_1[1359:1352] < top_1[1367:1360]) ? 1 : 0;
assign detect_min[168][6] = (mid_1[1359:1352] < top_2[1351:1344]) ? 1 : 0;
assign detect_min[168][7] = (mid_1[1359:1352] < top_2[1359:1352]) ? 1 : 0;
assign detect_min[168][8] = (mid_1[1359:1352] < top_2[1367:1360]) ? 1 : 0;
assign detect_min[168][9] = (mid_1[1359:1352] < mid_0[1351:1344]) ? 1 : 0;
assign detect_min[168][10] = (mid_1[1359:1352] < mid_0[1359:1352]) ? 1 : 0;
assign detect_min[168][11] = (mid_1[1359:1352] < mid_0[1367:1360]) ? 1 : 0;
assign detect_min[168][12] = (mid_1[1359:1352] < mid_1[1351:1344]) ? 1 : 0;
assign detect_min[168][13] = (mid_1[1359:1352] < mid_1[1367:1360]) ? 1 : 0;
assign detect_min[168][14] = (mid_1[1359:1352] < mid_2[1351:1344]) ? 1 : 0;
assign detect_min[168][15] = (mid_1[1359:1352] < mid_2[1359:1352]) ? 1 : 0;
assign detect_min[168][16] = (mid_1[1359:1352] < mid_2[1367:1360]) ? 1 : 0;
assign detect_min[168][17] = (mid_1[1359:1352] < btm_0[1351:1344]) ? 1 : 0;
assign detect_min[168][18] = (mid_1[1359:1352] < btm_0[1359:1352]) ? 1 : 0;
assign detect_min[168][19] = (mid_1[1359:1352] < btm_0[1367:1360]) ? 1 : 0;
assign detect_min[168][20] = (mid_1[1359:1352] < btm_1[1351:1344]) ? 1 : 0;
assign detect_min[168][21] = (mid_1[1359:1352] < btm_1[1359:1352]) ? 1 : 0;
assign detect_min[168][22] = (mid_1[1359:1352] < btm_1[1367:1360]) ? 1 : 0;
assign detect_min[168][23] = (mid_1[1359:1352] < btm_2[1351:1344]) ? 1 : 0;
assign detect_min[168][24] = (mid_1[1359:1352] < btm_2[1359:1352]) ? 1 : 0;
assign detect_min[168][25] = (mid_1[1359:1352] < btm_2[1367:1360]) ? 1 : 0;

assign detect_min[169][0] = (mid_1[1367:1360] < top_0[1359:1352]) ? 1 : 0;
assign detect_min[169][1] = (mid_1[1367:1360] < top_0[1367:1360]) ? 1 : 0;
assign detect_min[169][2] = (mid_1[1367:1360] < top_0[1375:1368]) ? 1 : 0;
assign detect_min[169][3] = (mid_1[1367:1360] < top_1[1359:1352]) ? 1 : 0;
assign detect_min[169][4] = (mid_1[1367:1360] < top_1[1367:1360]) ? 1 : 0;
assign detect_min[169][5] = (mid_1[1367:1360] < top_1[1375:1368]) ? 1 : 0;
assign detect_min[169][6] = (mid_1[1367:1360] < top_2[1359:1352]) ? 1 : 0;
assign detect_min[169][7] = (mid_1[1367:1360] < top_2[1367:1360]) ? 1 : 0;
assign detect_min[169][8] = (mid_1[1367:1360] < top_2[1375:1368]) ? 1 : 0;
assign detect_min[169][9] = (mid_1[1367:1360] < mid_0[1359:1352]) ? 1 : 0;
assign detect_min[169][10] = (mid_1[1367:1360] < mid_0[1367:1360]) ? 1 : 0;
assign detect_min[169][11] = (mid_1[1367:1360] < mid_0[1375:1368]) ? 1 : 0;
assign detect_min[169][12] = (mid_1[1367:1360] < mid_1[1359:1352]) ? 1 : 0;
assign detect_min[169][13] = (mid_1[1367:1360] < mid_1[1375:1368]) ? 1 : 0;
assign detect_min[169][14] = (mid_1[1367:1360] < mid_2[1359:1352]) ? 1 : 0;
assign detect_min[169][15] = (mid_1[1367:1360] < mid_2[1367:1360]) ? 1 : 0;
assign detect_min[169][16] = (mid_1[1367:1360] < mid_2[1375:1368]) ? 1 : 0;
assign detect_min[169][17] = (mid_1[1367:1360] < btm_0[1359:1352]) ? 1 : 0;
assign detect_min[169][18] = (mid_1[1367:1360] < btm_0[1367:1360]) ? 1 : 0;
assign detect_min[169][19] = (mid_1[1367:1360] < btm_0[1375:1368]) ? 1 : 0;
assign detect_min[169][20] = (mid_1[1367:1360] < btm_1[1359:1352]) ? 1 : 0;
assign detect_min[169][21] = (mid_1[1367:1360] < btm_1[1367:1360]) ? 1 : 0;
assign detect_min[169][22] = (mid_1[1367:1360] < btm_1[1375:1368]) ? 1 : 0;
assign detect_min[169][23] = (mid_1[1367:1360] < btm_2[1359:1352]) ? 1 : 0;
assign detect_min[169][24] = (mid_1[1367:1360] < btm_2[1367:1360]) ? 1 : 0;
assign detect_min[169][25] = (mid_1[1367:1360] < btm_2[1375:1368]) ? 1 : 0;

assign detect_min[170][0] = (mid_1[1375:1368] < top_0[1367:1360]) ? 1 : 0;
assign detect_min[170][1] = (mid_1[1375:1368] < top_0[1375:1368]) ? 1 : 0;
assign detect_min[170][2] = (mid_1[1375:1368] < top_0[1383:1376]) ? 1 : 0;
assign detect_min[170][3] = (mid_1[1375:1368] < top_1[1367:1360]) ? 1 : 0;
assign detect_min[170][4] = (mid_1[1375:1368] < top_1[1375:1368]) ? 1 : 0;
assign detect_min[170][5] = (mid_1[1375:1368] < top_1[1383:1376]) ? 1 : 0;
assign detect_min[170][6] = (mid_1[1375:1368] < top_2[1367:1360]) ? 1 : 0;
assign detect_min[170][7] = (mid_1[1375:1368] < top_2[1375:1368]) ? 1 : 0;
assign detect_min[170][8] = (mid_1[1375:1368] < top_2[1383:1376]) ? 1 : 0;
assign detect_min[170][9] = (mid_1[1375:1368] < mid_0[1367:1360]) ? 1 : 0;
assign detect_min[170][10] = (mid_1[1375:1368] < mid_0[1375:1368]) ? 1 : 0;
assign detect_min[170][11] = (mid_1[1375:1368] < mid_0[1383:1376]) ? 1 : 0;
assign detect_min[170][12] = (mid_1[1375:1368] < mid_1[1367:1360]) ? 1 : 0;
assign detect_min[170][13] = (mid_1[1375:1368] < mid_1[1383:1376]) ? 1 : 0;
assign detect_min[170][14] = (mid_1[1375:1368] < mid_2[1367:1360]) ? 1 : 0;
assign detect_min[170][15] = (mid_1[1375:1368] < mid_2[1375:1368]) ? 1 : 0;
assign detect_min[170][16] = (mid_1[1375:1368] < mid_2[1383:1376]) ? 1 : 0;
assign detect_min[170][17] = (mid_1[1375:1368] < btm_0[1367:1360]) ? 1 : 0;
assign detect_min[170][18] = (mid_1[1375:1368] < btm_0[1375:1368]) ? 1 : 0;
assign detect_min[170][19] = (mid_1[1375:1368] < btm_0[1383:1376]) ? 1 : 0;
assign detect_min[170][20] = (mid_1[1375:1368] < btm_1[1367:1360]) ? 1 : 0;
assign detect_min[170][21] = (mid_1[1375:1368] < btm_1[1375:1368]) ? 1 : 0;
assign detect_min[170][22] = (mid_1[1375:1368] < btm_1[1383:1376]) ? 1 : 0;
assign detect_min[170][23] = (mid_1[1375:1368] < btm_2[1367:1360]) ? 1 : 0;
assign detect_min[170][24] = (mid_1[1375:1368] < btm_2[1375:1368]) ? 1 : 0;
assign detect_min[170][25] = (mid_1[1375:1368] < btm_2[1383:1376]) ? 1 : 0;

assign detect_min[171][0] = (mid_1[1383:1376] < top_0[1375:1368]) ? 1 : 0;
assign detect_min[171][1] = (mid_1[1383:1376] < top_0[1383:1376]) ? 1 : 0;
assign detect_min[171][2] = (mid_1[1383:1376] < top_0[1391:1384]) ? 1 : 0;
assign detect_min[171][3] = (mid_1[1383:1376] < top_1[1375:1368]) ? 1 : 0;
assign detect_min[171][4] = (mid_1[1383:1376] < top_1[1383:1376]) ? 1 : 0;
assign detect_min[171][5] = (mid_1[1383:1376] < top_1[1391:1384]) ? 1 : 0;
assign detect_min[171][6] = (mid_1[1383:1376] < top_2[1375:1368]) ? 1 : 0;
assign detect_min[171][7] = (mid_1[1383:1376] < top_2[1383:1376]) ? 1 : 0;
assign detect_min[171][8] = (mid_1[1383:1376] < top_2[1391:1384]) ? 1 : 0;
assign detect_min[171][9] = (mid_1[1383:1376] < mid_0[1375:1368]) ? 1 : 0;
assign detect_min[171][10] = (mid_1[1383:1376] < mid_0[1383:1376]) ? 1 : 0;
assign detect_min[171][11] = (mid_1[1383:1376] < mid_0[1391:1384]) ? 1 : 0;
assign detect_min[171][12] = (mid_1[1383:1376] < mid_1[1375:1368]) ? 1 : 0;
assign detect_min[171][13] = (mid_1[1383:1376] < mid_1[1391:1384]) ? 1 : 0;
assign detect_min[171][14] = (mid_1[1383:1376] < mid_2[1375:1368]) ? 1 : 0;
assign detect_min[171][15] = (mid_1[1383:1376] < mid_2[1383:1376]) ? 1 : 0;
assign detect_min[171][16] = (mid_1[1383:1376] < mid_2[1391:1384]) ? 1 : 0;
assign detect_min[171][17] = (mid_1[1383:1376] < btm_0[1375:1368]) ? 1 : 0;
assign detect_min[171][18] = (mid_1[1383:1376] < btm_0[1383:1376]) ? 1 : 0;
assign detect_min[171][19] = (mid_1[1383:1376] < btm_0[1391:1384]) ? 1 : 0;
assign detect_min[171][20] = (mid_1[1383:1376] < btm_1[1375:1368]) ? 1 : 0;
assign detect_min[171][21] = (mid_1[1383:1376] < btm_1[1383:1376]) ? 1 : 0;
assign detect_min[171][22] = (mid_1[1383:1376] < btm_1[1391:1384]) ? 1 : 0;
assign detect_min[171][23] = (mid_1[1383:1376] < btm_2[1375:1368]) ? 1 : 0;
assign detect_min[171][24] = (mid_1[1383:1376] < btm_2[1383:1376]) ? 1 : 0;
assign detect_min[171][25] = (mid_1[1383:1376] < btm_2[1391:1384]) ? 1 : 0;

assign detect_min[172][0] = (mid_1[1391:1384] < top_0[1383:1376]) ? 1 : 0;
assign detect_min[172][1] = (mid_1[1391:1384] < top_0[1391:1384]) ? 1 : 0;
assign detect_min[172][2] = (mid_1[1391:1384] < top_0[1399:1392]) ? 1 : 0;
assign detect_min[172][3] = (mid_1[1391:1384] < top_1[1383:1376]) ? 1 : 0;
assign detect_min[172][4] = (mid_1[1391:1384] < top_1[1391:1384]) ? 1 : 0;
assign detect_min[172][5] = (mid_1[1391:1384] < top_1[1399:1392]) ? 1 : 0;
assign detect_min[172][6] = (mid_1[1391:1384] < top_2[1383:1376]) ? 1 : 0;
assign detect_min[172][7] = (mid_1[1391:1384] < top_2[1391:1384]) ? 1 : 0;
assign detect_min[172][8] = (mid_1[1391:1384] < top_2[1399:1392]) ? 1 : 0;
assign detect_min[172][9] = (mid_1[1391:1384] < mid_0[1383:1376]) ? 1 : 0;
assign detect_min[172][10] = (mid_1[1391:1384] < mid_0[1391:1384]) ? 1 : 0;
assign detect_min[172][11] = (mid_1[1391:1384] < mid_0[1399:1392]) ? 1 : 0;
assign detect_min[172][12] = (mid_1[1391:1384] < mid_1[1383:1376]) ? 1 : 0;
assign detect_min[172][13] = (mid_1[1391:1384] < mid_1[1399:1392]) ? 1 : 0;
assign detect_min[172][14] = (mid_1[1391:1384] < mid_2[1383:1376]) ? 1 : 0;
assign detect_min[172][15] = (mid_1[1391:1384] < mid_2[1391:1384]) ? 1 : 0;
assign detect_min[172][16] = (mid_1[1391:1384] < mid_2[1399:1392]) ? 1 : 0;
assign detect_min[172][17] = (mid_1[1391:1384] < btm_0[1383:1376]) ? 1 : 0;
assign detect_min[172][18] = (mid_1[1391:1384] < btm_0[1391:1384]) ? 1 : 0;
assign detect_min[172][19] = (mid_1[1391:1384] < btm_0[1399:1392]) ? 1 : 0;
assign detect_min[172][20] = (mid_1[1391:1384] < btm_1[1383:1376]) ? 1 : 0;
assign detect_min[172][21] = (mid_1[1391:1384] < btm_1[1391:1384]) ? 1 : 0;
assign detect_min[172][22] = (mid_1[1391:1384] < btm_1[1399:1392]) ? 1 : 0;
assign detect_min[172][23] = (mid_1[1391:1384] < btm_2[1383:1376]) ? 1 : 0;
assign detect_min[172][24] = (mid_1[1391:1384] < btm_2[1391:1384]) ? 1 : 0;
assign detect_min[172][25] = (mid_1[1391:1384] < btm_2[1399:1392]) ? 1 : 0;

assign detect_min[173][0] = (mid_1[1399:1392] < top_0[1391:1384]) ? 1 : 0;
assign detect_min[173][1] = (mid_1[1399:1392] < top_0[1399:1392]) ? 1 : 0;
assign detect_min[173][2] = (mid_1[1399:1392] < top_0[1407:1400]) ? 1 : 0;
assign detect_min[173][3] = (mid_1[1399:1392] < top_1[1391:1384]) ? 1 : 0;
assign detect_min[173][4] = (mid_1[1399:1392] < top_1[1399:1392]) ? 1 : 0;
assign detect_min[173][5] = (mid_1[1399:1392] < top_1[1407:1400]) ? 1 : 0;
assign detect_min[173][6] = (mid_1[1399:1392] < top_2[1391:1384]) ? 1 : 0;
assign detect_min[173][7] = (mid_1[1399:1392] < top_2[1399:1392]) ? 1 : 0;
assign detect_min[173][8] = (mid_1[1399:1392] < top_2[1407:1400]) ? 1 : 0;
assign detect_min[173][9] = (mid_1[1399:1392] < mid_0[1391:1384]) ? 1 : 0;
assign detect_min[173][10] = (mid_1[1399:1392] < mid_0[1399:1392]) ? 1 : 0;
assign detect_min[173][11] = (mid_1[1399:1392] < mid_0[1407:1400]) ? 1 : 0;
assign detect_min[173][12] = (mid_1[1399:1392] < mid_1[1391:1384]) ? 1 : 0;
assign detect_min[173][13] = (mid_1[1399:1392] < mid_1[1407:1400]) ? 1 : 0;
assign detect_min[173][14] = (mid_1[1399:1392] < mid_2[1391:1384]) ? 1 : 0;
assign detect_min[173][15] = (mid_1[1399:1392] < mid_2[1399:1392]) ? 1 : 0;
assign detect_min[173][16] = (mid_1[1399:1392] < mid_2[1407:1400]) ? 1 : 0;
assign detect_min[173][17] = (mid_1[1399:1392] < btm_0[1391:1384]) ? 1 : 0;
assign detect_min[173][18] = (mid_1[1399:1392] < btm_0[1399:1392]) ? 1 : 0;
assign detect_min[173][19] = (mid_1[1399:1392] < btm_0[1407:1400]) ? 1 : 0;
assign detect_min[173][20] = (mid_1[1399:1392] < btm_1[1391:1384]) ? 1 : 0;
assign detect_min[173][21] = (mid_1[1399:1392] < btm_1[1399:1392]) ? 1 : 0;
assign detect_min[173][22] = (mid_1[1399:1392] < btm_1[1407:1400]) ? 1 : 0;
assign detect_min[173][23] = (mid_1[1399:1392] < btm_2[1391:1384]) ? 1 : 0;
assign detect_min[173][24] = (mid_1[1399:1392] < btm_2[1399:1392]) ? 1 : 0;
assign detect_min[173][25] = (mid_1[1399:1392] < btm_2[1407:1400]) ? 1 : 0;

assign detect_min[174][0] = (mid_1[1407:1400] < top_0[1399:1392]) ? 1 : 0;
assign detect_min[174][1] = (mid_1[1407:1400] < top_0[1407:1400]) ? 1 : 0;
assign detect_min[174][2] = (mid_1[1407:1400] < top_0[1415:1408]) ? 1 : 0;
assign detect_min[174][3] = (mid_1[1407:1400] < top_1[1399:1392]) ? 1 : 0;
assign detect_min[174][4] = (mid_1[1407:1400] < top_1[1407:1400]) ? 1 : 0;
assign detect_min[174][5] = (mid_1[1407:1400] < top_1[1415:1408]) ? 1 : 0;
assign detect_min[174][6] = (mid_1[1407:1400] < top_2[1399:1392]) ? 1 : 0;
assign detect_min[174][7] = (mid_1[1407:1400] < top_2[1407:1400]) ? 1 : 0;
assign detect_min[174][8] = (mid_1[1407:1400] < top_2[1415:1408]) ? 1 : 0;
assign detect_min[174][9] = (mid_1[1407:1400] < mid_0[1399:1392]) ? 1 : 0;
assign detect_min[174][10] = (mid_1[1407:1400] < mid_0[1407:1400]) ? 1 : 0;
assign detect_min[174][11] = (mid_1[1407:1400] < mid_0[1415:1408]) ? 1 : 0;
assign detect_min[174][12] = (mid_1[1407:1400] < mid_1[1399:1392]) ? 1 : 0;
assign detect_min[174][13] = (mid_1[1407:1400] < mid_1[1415:1408]) ? 1 : 0;
assign detect_min[174][14] = (mid_1[1407:1400] < mid_2[1399:1392]) ? 1 : 0;
assign detect_min[174][15] = (mid_1[1407:1400] < mid_2[1407:1400]) ? 1 : 0;
assign detect_min[174][16] = (mid_1[1407:1400] < mid_2[1415:1408]) ? 1 : 0;
assign detect_min[174][17] = (mid_1[1407:1400] < btm_0[1399:1392]) ? 1 : 0;
assign detect_min[174][18] = (mid_1[1407:1400] < btm_0[1407:1400]) ? 1 : 0;
assign detect_min[174][19] = (mid_1[1407:1400] < btm_0[1415:1408]) ? 1 : 0;
assign detect_min[174][20] = (mid_1[1407:1400] < btm_1[1399:1392]) ? 1 : 0;
assign detect_min[174][21] = (mid_1[1407:1400] < btm_1[1407:1400]) ? 1 : 0;
assign detect_min[174][22] = (mid_1[1407:1400] < btm_1[1415:1408]) ? 1 : 0;
assign detect_min[174][23] = (mid_1[1407:1400] < btm_2[1399:1392]) ? 1 : 0;
assign detect_min[174][24] = (mid_1[1407:1400] < btm_2[1407:1400]) ? 1 : 0;
assign detect_min[174][25] = (mid_1[1407:1400] < btm_2[1415:1408]) ? 1 : 0;

assign detect_min[175][0] = (mid_1[1415:1408] < top_0[1407:1400]) ? 1 : 0;
assign detect_min[175][1] = (mid_1[1415:1408] < top_0[1415:1408]) ? 1 : 0;
assign detect_min[175][2] = (mid_1[1415:1408] < top_0[1423:1416]) ? 1 : 0;
assign detect_min[175][3] = (mid_1[1415:1408] < top_1[1407:1400]) ? 1 : 0;
assign detect_min[175][4] = (mid_1[1415:1408] < top_1[1415:1408]) ? 1 : 0;
assign detect_min[175][5] = (mid_1[1415:1408] < top_1[1423:1416]) ? 1 : 0;
assign detect_min[175][6] = (mid_1[1415:1408] < top_2[1407:1400]) ? 1 : 0;
assign detect_min[175][7] = (mid_1[1415:1408] < top_2[1415:1408]) ? 1 : 0;
assign detect_min[175][8] = (mid_1[1415:1408] < top_2[1423:1416]) ? 1 : 0;
assign detect_min[175][9] = (mid_1[1415:1408] < mid_0[1407:1400]) ? 1 : 0;
assign detect_min[175][10] = (mid_1[1415:1408] < mid_0[1415:1408]) ? 1 : 0;
assign detect_min[175][11] = (mid_1[1415:1408] < mid_0[1423:1416]) ? 1 : 0;
assign detect_min[175][12] = (mid_1[1415:1408] < mid_1[1407:1400]) ? 1 : 0;
assign detect_min[175][13] = (mid_1[1415:1408] < mid_1[1423:1416]) ? 1 : 0;
assign detect_min[175][14] = (mid_1[1415:1408] < mid_2[1407:1400]) ? 1 : 0;
assign detect_min[175][15] = (mid_1[1415:1408] < mid_2[1415:1408]) ? 1 : 0;
assign detect_min[175][16] = (mid_1[1415:1408] < mid_2[1423:1416]) ? 1 : 0;
assign detect_min[175][17] = (mid_1[1415:1408] < btm_0[1407:1400]) ? 1 : 0;
assign detect_min[175][18] = (mid_1[1415:1408] < btm_0[1415:1408]) ? 1 : 0;
assign detect_min[175][19] = (mid_1[1415:1408] < btm_0[1423:1416]) ? 1 : 0;
assign detect_min[175][20] = (mid_1[1415:1408] < btm_1[1407:1400]) ? 1 : 0;
assign detect_min[175][21] = (mid_1[1415:1408] < btm_1[1415:1408]) ? 1 : 0;
assign detect_min[175][22] = (mid_1[1415:1408] < btm_1[1423:1416]) ? 1 : 0;
assign detect_min[175][23] = (mid_1[1415:1408] < btm_2[1407:1400]) ? 1 : 0;
assign detect_min[175][24] = (mid_1[1415:1408] < btm_2[1415:1408]) ? 1 : 0;
assign detect_min[175][25] = (mid_1[1415:1408] < btm_2[1423:1416]) ? 1 : 0;

assign detect_min[176][0] = (mid_1[1423:1416] < top_0[1415:1408]) ? 1 : 0;
assign detect_min[176][1] = (mid_1[1423:1416] < top_0[1423:1416]) ? 1 : 0;
assign detect_min[176][2] = (mid_1[1423:1416] < top_0[1431:1424]) ? 1 : 0;
assign detect_min[176][3] = (mid_1[1423:1416] < top_1[1415:1408]) ? 1 : 0;
assign detect_min[176][4] = (mid_1[1423:1416] < top_1[1423:1416]) ? 1 : 0;
assign detect_min[176][5] = (mid_1[1423:1416] < top_1[1431:1424]) ? 1 : 0;
assign detect_min[176][6] = (mid_1[1423:1416] < top_2[1415:1408]) ? 1 : 0;
assign detect_min[176][7] = (mid_1[1423:1416] < top_2[1423:1416]) ? 1 : 0;
assign detect_min[176][8] = (mid_1[1423:1416] < top_2[1431:1424]) ? 1 : 0;
assign detect_min[176][9] = (mid_1[1423:1416] < mid_0[1415:1408]) ? 1 : 0;
assign detect_min[176][10] = (mid_1[1423:1416] < mid_0[1423:1416]) ? 1 : 0;
assign detect_min[176][11] = (mid_1[1423:1416] < mid_0[1431:1424]) ? 1 : 0;
assign detect_min[176][12] = (mid_1[1423:1416] < mid_1[1415:1408]) ? 1 : 0;
assign detect_min[176][13] = (mid_1[1423:1416] < mid_1[1431:1424]) ? 1 : 0;
assign detect_min[176][14] = (mid_1[1423:1416] < mid_2[1415:1408]) ? 1 : 0;
assign detect_min[176][15] = (mid_1[1423:1416] < mid_2[1423:1416]) ? 1 : 0;
assign detect_min[176][16] = (mid_1[1423:1416] < mid_2[1431:1424]) ? 1 : 0;
assign detect_min[176][17] = (mid_1[1423:1416] < btm_0[1415:1408]) ? 1 : 0;
assign detect_min[176][18] = (mid_1[1423:1416] < btm_0[1423:1416]) ? 1 : 0;
assign detect_min[176][19] = (mid_1[1423:1416] < btm_0[1431:1424]) ? 1 : 0;
assign detect_min[176][20] = (mid_1[1423:1416] < btm_1[1415:1408]) ? 1 : 0;
assign detect_min[176][21] = (mid_1[1423:1416] < btm_1[1423:1416]) ? 1 : 0;
assign detect_min[176][22] = (mid_1[1423:1416] < btm_1[1431:1424]) ? 1 : 0;
assign detect_min[176][23] = (mid_1[1423:1416] < btm_2[1415:1408]) ? 1 : 0;
assign detect_min[176][24] = (mid_1[1423:1416] < btm_2[1423:1416]) ? 1 : 0;
assign detect_min[176][25] = (mid_1[1423:1416] < btm_2[1431:1424]) ? 1 : 0;

assign detect_min[177][0] = (mid_1[1431:1424] < top_0[1423:1416]) ? 1 : 0;
assign detect_min[177][1] = (mid_1[1431:1424] < top_0[1431:1424]) ? 1 : 0;
assign detect_min[177][2] = (mid_1[1431:1424] < top_0[1439:1432]) ? 1 : 0;
assign detect_min[177][3] = (mid_1[1431:1424] < top_1[1423:1416]) ? 1 : 0;
assign detect_min[177][4] = (mid_1[1431:1424] < top_1[1431:1424]) ? 1 : 0;
assign detect_min[177][5] = (mid_1[1431:1424] < top_1[1439:1432]) ? 1 : 0;
assign detect_min[177][6] = (mid_1[1431:1424] < top_2[1423:1416]) ? 1 : 0;
assign detect_min[177][7] = (mid_1[1431:1424] < top_2[1431:1424]) ? 1 : 0;
assign detect_min[177][8] = (mid_1[1431:1424] < top_2[1439:1432]) ? 1 : 0;
assign detect_min[177][9] = (mid_1[1431:1424] < mid_0[1423:1416]) ? 1 : 0;
assign detect_min[177][10] = (mid_1[1431:1424] < mid_0[1431:1424]) ? 1 : 0;
assign detect_min[177][11] = (mid_1[1431:1424] < mid_0[1439:1432]) ? 1 : 0;
assign detect_min[177][12] = (mid_1[1431:1424] < mid_1[1423:1416]) ? 1 : 0;
assign detect_min[177][13] = (mid_1[1431:1424] < mid_1[1439:1432]) ? 1 : 0;
assign detect_min[177][14] = (mid_1[1431:1424] < mid_2[1423:1416]) ? 1 : 0;
assign detect_min[177][15] = (mid_1[1431:1424] < mid_2[1431:1424]) ? 1 : 0;
assign detect_min[177][16] = (mid_1[1431:1424] < mid_2[1439:1432]) ? 1 : 0;
assign detect_min[177][17] = (mid_1[1431:1424] < btm_0[1423:1416]) ? 1 : 0;
assign detect_min[177][18] = (mid_1[1431:1424] < btm_0[1431:1424]) ? 1 : 0;
assign detect_min[177][19] = (mid_1[1431:1424] < btm_0[1439:1432]) ? 1 : 0;
assign detect_min[177][20] = (mid_1[1431:1424] < btm_1[1423:1416]) ? 1 : 0;
assign detect_min[177][21] = (mid_1[1431:1424] < btm_1[1431:1424]) ? 1 : 0;
assign detect_min[177][22] = (mid_1[1431:1424] < btm_1[1439:1432]) ? 1 : 0;
assign detect_min[177][23] = (mid_1[1431:1424] < btm_2[1423:1416]) ? 1 : 0;
assign detect_min[177][24] = (mid_1[1431:1424] < btm_2[1431:1424]) ? 1 : 0;
assign detect_min[177][25] = (mid_1[1431:1424] < btm_2[1439:1432]) ? 1 : 0;

assign detect_min[178][0] = (mid_1[1439:1432] < top_0[1431:1424]) ? 1 : 0;
assign detect_min[178][1] = (mid_1[1439:1432] < top_0[1439:1432]) ? 1 : 0;
assign detect_min[178][2] = (mid_1[1439:1432] < top_0[1447:1440]) ? 1 : 0;
assign detect_min[178][3] = (mid_1[1439:1432] < top_1[1431:1424]) ? 1 : 0;
assign detect_min[178][4] = (mid_1[1439:1432] < top_1[1439:1432]) ? 1 : 0;
assign detect_min[178][5] = (mid_1[1439:1432] < top_1[1447:1440]) ? 1 : 0;
assign detect_min[178][6] = (mid_1[1439:1432] < top_2[1431:1424]) ? 1 : 0;
assign detect_min[178][7] = (mid_1[1439:1432] < top_2[1439:1432]) ? 1 : 0;
assign detect_min[178][8] = (mid_1[1439:1432] < top_2[1447:1440]) ? 1 : 0;
assign detect_min[178][9] = (mid_1[1439:1432] < mid_0[1431:1424]) ? 1 : 0;
assign detect_min[178][10] = (mid_1[1439:1432] < mid_0[1439:1432]) ? 1 : 0;
assign detect_min[178][11] = (mid_1[1439:1432] < mid_0[1447:1440]) ? 1 : 0;
assign detect_min[178][12] = (mid_1[1439:1432] < mid_1[1431:1424]) ? 1 : 0;
assign detect_min[178][13] = (mid_1[1439:1432] < mid_1[1447:1440]) ? 1 : 0;
assign detect_min[178][14] = (mid_1[1439:1432] < mid_2[1431:1424]) ? 1 : 0;
assign detect_min[178][15] = (mid_1[1439:1432] < mid_2[1439:1432]) ? 1 : 0;
assign detect_min[178][16] = (mid_1[1439:1432] < mid_2[1447:1440]) ? 1 : 0;
assign detect_min[178][17] = (mid_1[1439:1432] < btm_0[1431:1424]) ? 1 : 0;
assign detect_min[178][18] = (mid_1[1439:1432] < btm_0[1439:1432]) ? 1 : 0;
assign detect_min[178][19] = (mid_1[1439:1432] < btm_0[1447:1440]) ? 1 : 0;
assign detect_min[178][20] = (mid_1[1439:1432] < btm_1[1431:1424]) ? 1 : 0;
assign detect_min[178][21] = (mid_1[1439:1432] < btm_1[1439:1432]) ? 1 : 0;
assign detect_min[178][22] = (mid_1[1439:1432] < btm_1[1447:1440]) ? 1 : 0;
assign detect_min[178][23] = (mid_1[1439:1432] < btm_2[1431:1424]) ? 1 : 0;
assign detect_min[178][24] = (mid_1[1439:1432] < btm_2[1439:1432]) ? 1 : 0;
assign detect_min[178][25] = (mid_1[1439:1432] < btm_2[1447:1440]) ? 1 : 0;

assign detect_min[179][0] = (mid_1[1447:1440] < top_0[1439:1432]) ? 1 : 0;
assign detect_min[179][1] = (mid_1[1447:1440] < top_0[1447:1440]) ? 1 : 0;
assign detect_min[179][2] = (mid_1[1447:1440] < top_0[1455:1448]) ? 1 : 0;
assign detect_min[179][3] = (mid_1[1447:1440] < top_1[1439:1432]) ? 1 : 0;
assign detect_min[179][4] = (mid_1[1447:1440] < top_1[1447:1440]) ? 1 : 0;
assign detect_min[179][5] = (mid_1[1447:1440] < top_1[1455:1448]) ? 1 : 0;
assign detect_min[179][6] = (mid_1[1447:1440] < top_2[1439:1432]) ? 1 : 0;
assign detect_min[179][7] = (mid_1[1447:1440] < top_2[1447:1440]) ? 1 : 0;
assign detect_min[179][8] = (mid_1[1447:1440] < top_2[1455:1448]) ? 1 : 0;
assign detect_min[179][9] = (mid_1[1447:1440] < mid_0[1439:1432]) ? 1 : 0;
assign detect_min[179][10] = (mid_1[1447:1440] < mid_0[1447:1440]) ? 1 : 0;
assign detect_min[179][11] = (mid_1[1447:1440] < mid_0[1455:1448]) ? 1 : 0;
assign detect_min[179][12] = (mid_1[1447:1440] < mid_1[1439:1432]) ? 1 : 0;
assign detect_min[179][13] = (mid_1[1447:1440] < mid_1[1455:1448]) ? 1 : 0;
assign detect_min[179][14] = (mid_1[1447:1440] < mid_2[1439:1432]) ? 1 : 0;
assign detect_min[179][15] = (mid_1[1447:1440] < mid_2[1447:1440]) ? 1 : 0;
assign detect_min[179][16] = (mid_1[1447:1440] < mid_2[1455:1448]) ? 1 : 0;
assign detect_min[179][17] = (mid_1[1447:1440] < btm_0[1439:1432]) ? 1 : 0;
assign detect_min[179][18] = (mid_1[1447:1440] < btm_0[1447:1440]) ? 1 : 0;
assign detect_min[179][19] = (mid_1[1447:1440] < btm_0[1455:1448]) ? 1 : 0;
assign detect_min[179][20] = (mid_1[1447:1440] < btm_1[1439:1432]) ? 1 : 0;
assign detect_min[179][21] = (mid_1[1447:1440] < btm_1[1447:1440]) ? 1 : 0;
assign detect_min[179][22] = (mid_1[1447:1440] < btm_1[1455:1448]) ? 1 : 0;
assign detect_min[179][23] = (mid_1[1447:1440] < btm_2[1439:1432]) ? 1 : 0;
assign detect_min[179][24] = (mid_1[1447:1440] < btm_2[1447:1440]) ? 1 : 0;
assign detect_min[179][25] = (mid_1[1447:1440] < btm_2[1455:1448]) ? 1 : 0;

assign detect_min[180][0] = (mid_1[1455:1448] < top_0[1447:1440]) ? 1 : 0;
assign detect_min[180][1] = (mid_1[1455:1448] < top_0[1455:1448]) ? 1 : 0;
assign detect_min[180][2] = (mid_1[1455:1448] < top_0[1463:1456]) ? 1 : 0;
assign detect_min[180][3] = (mid_1[1455:1448] < top_1[1447:1440]) ? 1 : 0;
assign detect_min[180][4] = (mid_1[1455:1448] < top_1[1455:1448]) ? 1 : 0;
assign detect_min[180][5] = (mid_1[1455:1448] < top_1[1463:1456]) ? 1 : 0;
assign detect_min[180][6] = (mid_1[1455:1448] < top_2[1447:1440]) ? 1 : 0;
assign detect_min[180][7] = (mid_1[1455:1448] < top_2[1455:1448]) ? 1 : 0;
assign detect_min[180][8] = (mid_1[1455:1448] < top_2[1463:1456]) ? 1 : 0;
assign detect_min[180][9] = (mid_1[1455:1448] < mid_0[1447:1440]) ? 1 : 0;
assign detect_min[180][10] = (mid_1[1455:1448] < mid_0[1455:1448]) ? 1 : 0;
assign detect_min[180][11] = (mid_1[1455:1448] < mid_0[1463:1456]) ? 1 : 0;
assign detect_min[180][12] = (mid_1[1455:1448] < mid_1[1447:1440]) ? 1 : 0;
assign detect_min[180][13] = (mid_1[1455:1448] < mid_1[1463:1456]) ? 1 : 0;
assign detect_min[180][14] = (mid_1[1455:1448] < mid_2[1447:1440]) ? 1 : 0;
assign detect_min[180][15] = (mid_1[1455:1448] < mid_2[1455:1448]) ? 1 : 0;
assign detect_min[180][16] = (mid_1[1455:1448] < mid_2[1463:1456]) ? 1 : 0;
assign detect_min[180][17] = (mid_1[1455:1448] < btm_0[1447:1440]) ? 1 : 0;
assign detect_min[180][18] = (mid_1[1455:1448] < btm_0[1455:1448]) ? 1 : 0;
assign detect_min[180][19] = (mid_1[1455:1448] < btm_0[1463:1456]) ? 1 : 0;
assign detect_min[180][20] = (mid_1[1455:1448] < btm_1[1447:1440]) ? 1 : 0;
assign detect_min[180][21] = (mid_1[1455:1448] < btm_1[1455:1448]) ? 1 : 0;
assign detect_min[180][22] = (mid_1[1455:1448] < btm_1[1463:1456]) ? 1 : 0;
assign detect_min[180][23] = (mid_1[1455:1448] < btm_2[1447:1440]) ? 1 : 0;
assign detect_min[180][24] = (mid_1[1455:1448] < btm_2[1455:1448]) ? 1 : 0;
assign detect_min[180][25] = (mid_1[1455:1448] < btm_2[1463:1456]) ? 1 : 0;

assign detect_min[181][0] = (mid_1[1463:1456] < top_0[1455:1448]) ? 1 : 0;
assign detect_min[181][1] = (mid_1[1463:1456] < top_0[1463:1456]) ? 1 : 0;
assign detect_min[181][2] = (mid_1[1463:1456] < top_0[1471:1464]) ? 1 : 0;
assign detect_min[181][3] = (mid_1[1463:1456] < top_1[1455:1448]) ? 1 : 0;
assign detect_min[181][4] = (mid_1[1463:1456] < top_1[1463:1456]) ? 1 : 0;
assign detect_min[181][5] = (mid_1[1463:1456] < top_1[1471:1464]) ? 1 : 0;
assign detect_min[181][6] = (mid_1[1463:1456] < top_2[1455:1448]) ? 1 : 0;
assign detect_min[181][7] = (mid_1[1463:1456] < top_2[1463:1456]) ? 1 : 0;
assign detect_min[181][8] = (mid_1[1463:1456] < top_2[1471:1464]) ? 1 : 0;
assign detect_min[181][9] = (mid_1[1463:1456] < mid_0[1455:1448]) ? 1 : 0;
assign detect_min[181][10] = (mid_1[1463:1456] < mid_0[1463:1456]) ? 1 : 0;
assign detect_min[181][11] = (mid_1[1463:1456] < mid_0[1471:1464]) ? 1 : 0;
assign detect_min[181][12] = (mid_1[1463:1456] < mid_1[1455:1448]) ? 1 : 0;
assign detect_min[181][13] = (mid_1[1463:1456] < mid_1[1471:1464]) ? 1 : 0;
assign detect_min[181][14] = (mid_1[1463:1456] < mid_2[1455:1448]) ? 1 : 0;
assign detect_min[181][15] = (mid_1[1463:1456] < mid_2[1463:1456]) ? 1 : 0;
assign detect_min[181][16] = (mid_1[1463:1456] < mid_2[1471:1464]) ? 1 : 0;
assign detect_min[181][17] = (mid_1[1463:1456] < btm_0[1455:1448]) ? 1 : 0;
assign detect_min[181][18] = (mid_1[1463:1456] < btm_0[1463:1456]) ? 1 : 0;
assign detect_min[181][19] = (mid_1[1463:1456] < btm_0[1471:1464]) ? 1 : 0;
assign detect_min[181][20] = (mid_1[1463:1456] < btm_1[1455:1448]) ? 1 : 0;
assign detect_min[181][21] = (mid_1[1463:1456] < btm_1[1463:1456]) ? 1 : 0;
assign detect_min[181][22] = (mid_1[1463:1456] < btm_1[1471:1464]) ? 1 : 0;
assign detect_min[181][23] = (mid_1[1463:1456] < btm_2[1455:1448]) ? 1 : 0;
assign detect_min[181][24] = (mid_1[1463:1456] < btm_2[1463:1456]) ? 1 : 0;
assign detect_min[181][25] = (mid_1[1463:1456] < btm_2[1471:1464]) ? 1 : 0;

assign detect_min[182][0] = (mid_1[1471:1464] < top_0[1463:1456]) ? 1 : 0;
assign detect_min[182][1] = (mid_1[1471:1464] < top_0[1471:1464]) ? 1 : 0;
assign detect_min[182][2] = (mid_1[1471:1464] < top_0[1479:1472]) ? 1 : 0;
assign detect_min[182][3] = (mid_1[1471:1464] < top_1[1463:1456]) ? 1 : 0;
assign detect_min[182][4] = (mid_1[1471:1464] < top_1[1471:1464]) ? 1 : 0;
assign detect_min[182][5] = (mid_1[1471:1464] < top_1[1479:1472]) ? 1 : 0;
assign detect_min[182][6] = (mid_1[1471:1464] < top_2[1463:1456]) ? 1 : 0;
assign detect_min[182][7] = (mid_1[1471:1464] < top_2[1471:1464]) ? 1 : 0;
assign detect_min[182][8] = (mid_1[1471:1464] < top_2[1479:1472]) ? 1 : 0;
assign detect_min[182][9] = (mid_1[1471:1464] < mid_0[1463:1456]) ? 1 : 0;
assign detect_min[182][10] = (mid_1[1471:1464] < mid_0[1471:1464]) ? 1 : 0;
assign detect_min[182][11] = (mid_1[1471:1464] < mid_0[1479:1472]) ? 1 : 0;
assign detect_min[182][12] = (mid_1[1471:1464] < mid_1[1463:1456]) ? 1 : 0;
assign detect_min[182][13] = (mid_1[1471:1464] < mid_1[1479:1472]) ? 1 : 0;
assign detect_min[182][14] = (mid_1[1471:1464] < mid_2[1463:1456]) ? 1 : 0;
assign detect_min[182][15] = (mid_1[1471:1464] < mid_2[1471:1464]) ? 1 : 0;
assign detect_min[182][16] = (mid_1[1471:1464] < mid_2[1479:1472]) ? 1 : 0;
assign detect_min[182][17] = (mid_1[1471:1464] < btm_0[1463:1456]) ? 1 : 0;
assign detect_min[182][18] = (mid_1[1471:1464] < btm_0[1471:1464]) ? 1 : 0;
assign detect_min[182][19] = (mid_1[1471:1464] < btm_0[1479:1472]) ? 1 : 0;
assign detect_min[182][20] = (mid_1[1471:1464] < btm_1[1463:1456]) ? 1 : 0;
assign detect_min[182][21] = (mid_1[1471:1464] < btm_1[1471:1464]) ? 1 : 0;
assign detect_min[182][22] = (mid_1[1471:1464] < btm_1[1479:1472]) ? 1 : 0;
assign detect_min[182][23] = (mid_1[1471:1464] < btm_2[1463:1456]) ? 1 : 0;
assign detect_min[182][24] = (mid_1[1471:1464] < btm_2[1471:1464]) ? 1 : 0;
assign detect_min[182][25] = (mid_1[1471:1464] < btm_2[1479:1472]) ? 1 : 0;

assign detect_min[183][0] = (mid_1[1479:1472] < top_0[1471:1464]) ? 1 : 0;
assign detect_min[183][1] = (mid_1[1479:1472] < top_0[1479:1472]) ? 1 : 0;
assign detect_min[183][2] = (mid_1[1479:1472] < top_0[1487:1480]) ? 1 : 0;
assign detect_min[183][3] = (mid_1[1479:1472] < top_1[1471:1464]) ? 1 : 0;
assign detect_min[183][4] = (mid_1[1479:1472] < top_1[1479:1472]) ? 1 : 0;
assign detect_min[183][5] = (mid_1[1479:1472] < top_1[1487:1480]) ? 1 : 0;
assign detect_min[183][6] = (mid_1[1479:1472] < top_2[1471:1464]) ? 1 : 0;
assign detect_min[183][7] = (mid_1[1479:1472] < top_2[1479:1472]) ? 1 : 0;
assign detect_min[183][8] = (mid_1[1479:1472] < top_2[1487:1480]) ? 1 : 0;
assign detect_min[183][9] = (mid_1[1479:1472] < mid_0[1471:1464]) ? 1 : 0;
assign detect_min[183][10] = (mid_1[1479:1472] < mid_0[1479:1472]) ? 1 : 0;
assign detect_min[183][11] = (mid_1[1479:1472] < mid_0[1487:1480]) ? 1 : 0;
assign detect_min[183][12] = (mid_1[1479:1472] < mid_1[1471:1464]) ? 1 : 0;
assign detect_min[183][13] = (mid_1[1479:1472] < mid_1[1487:1480]) ? 1 : 0;
assign detect_min[183][14] = (mid_1[1479:1472] < mid_2[1471:1464]) ? 1 : 0;
assign detect_min[183][15] = (mid_1[1479:1472] < mid_2[1479:1472]) ? 1 : 0;
assign detect_min[183][16] = (mid_1[1479:1472] < mid_2[1487:1480]) ? 1 : 0;
assign detect_min[183][17] = (mid_1[1479:1472] < btm_0[1471:1464]) ? 1 : 0;
assign detect_min[183][18] = (mid_1[1479:1472] < btm_0[1479:1472]) ? 1 : 0;
assign detect_min[183][19] = (mid_1[1479:1472] < btm_0[1487:1480]) ? 1 : 0;
assign detect_min[183][20] = (mid_1[1479:1472] < btm_1[1471:1464]) ? 1 : 0;
assign detect_min[183][21] = (mid_1[1479:1472] < btm_1[1479:1472]) ? 1 : 0;
assign detect_min[183][22] = (mid_1[1479:1472] < btm_1[1487:1480]) ? 1 : 0;
assign detect_min[183][23] = (mid_1[1479:1472] < btm_2[1471:1464]) ? 1 : 0;
assign detect_min[183][24] = (mid_1[1479:1472] < btm_2[1479:1472]) ? 1 : 0;
assign detect_min[183][25] = (mid_1[1479:1472] < btm_2[1487:1480]) ? 1 : 0;

assign detect_min[184][0] = (mid_1[1487:1480] < top_0[1479:1472]) ? 1 : 0;
assign detect_min[184][1] = (mid_1[1487:1480] < top_0[1487:1480]) ? 1 : 0;
assign detect_min[184][2] = (mid_1[1487:1480] < top_0[1495:1488]) ? 1 : 0;
assign detect_min[184][3] = (mid_1[1487:1480] < top_1[1479:1472]) ? 1 : 0;
assign detect_min[184][4] = (mid_1[1487:1480] < top_1[1487:1480]) ? 1 : 0;
assign detect_min[184][5] = (mid_1[1487:1480] < top_1[1495:1488]) ? 1 : 0;
assign detect_min[184][6] = (mid_1[1487:1480] < top_2[1479:1472]) ? 1 : 0;
assign detect_min[184][7] = (mid_1[1487:1480] < top_2[1487:1480]) ? 1 : 0;
assign detect_min[184][8] = (mid_1[1487:1480] < top_2[1495:1488]) ? 1 : 0;
assign detect_min[184][9] = (mid_1[1487:1480] < mid_0[1479:1472]) ? 1 : 0;
assign detect_min[184][10] = (mid_1[1487:1480] < mid_0[1487:1480]) ? 1 : 0;
assign detect_min[184][11] = (mid_1[1487:1480] < mid_0[1495:1488]) ? 1 : 0;
assign detect_min[184][12] = (mid_1[1487:1480] < mid_1[1479:1472]) ? 1 : 0;
assign detect_min[184][13] = (mid_1[1487:1480] < mid_1[1495:1488]) ? 1 : 0;
assign detect_min[184][14] = (mid_1[1487:1480] < mid_2[1479:1472]) ? 1 : 0;
assign detect_min[184][15] = (mid_1[1487:1480] < mid_2[1487:1480]) ? 1 : 0;
assign detect_min[184][16] = (mid_1[1487:1480] < mid_2[1495:1488]) ? 1 : 0;
assign detect_min[184][17] = (mid_1[1487:1480] < btm_0[1479:1472]) ? 1 : 0;
assign detect_min[184][18] = (mid_1[1487:1480] < btm_0[1487:1480]) ? 1 : 0;
assign detect_min[184][19] = (mid_1[1487:1480] < btm_0[1495:1488]) ? 1 : 0;
assign detect_min[184][20] = (mid_1[1487:1480] < btm_1[1479:1472]) ? 1 : 0;
assign detect_min[184][21] = (mid_1[1487:1480] < btm_1[1487:1480]) ? 1 : 0;
assign detect_min[184][22] = (mid_1[1487:1480] < btm_1[1495:1488]) ? 1 : 0;
assign detect_min[184][23] = (mid_1[1487:1480] < btm_2[1479:1472]) ? 1 : 0;
assign detect_min[184][24] = (mid_1[1487:1480] < btm_2[1487:1480]) ? 1 : 0;
assign detect_min[184][25] = (mid_1[1487:1480] < btm_2[1495:1488]) ? 1 : 0;

assign detect_min[185][0] = (mid_1[1495:1488] < top_0[1487:1480]) ? 1 : 0;
assign detect_min[185][1] = (mid_1[1495:1488] < top_0[1495:1488]) ? 1 : 0;
assign detect_min[185][2] = (mid_1[1495:1488] < top_0[1503:1496]) ? 1 : 0;
assign detect_min[185][3] = (mid_1[1495:1488] < top_1[1487:1480]) ? 1 : 0;
assign detect_min[185][4] = (mid_1[1495:1488] < top_1[1495:1488]) ? 1 : 0;
assign detect_min[185][5] = (mid_1[1495:1488] < top_1[1503:1496]) ? 1 : 0;
assign detect_min[185][6] = (mid_1[1495:1488] < top_2[1487:1480]) ? 1 : 0;
assign detect_min[185][7] = (mid_1[1495:1488] < top_2[1495:1488]) ? 1 : 0;
assign detect_min[185][8] = (mid_1[1495:1488] < top_2[1503:1496]) ? 1 : 0;
assign detect_min[185][9] = (mid_1[1495:1488] < mid_0[1487:1480]) ? 1 : 0;
assign detect_min[185][10] = (mid_1[1495:1488] < mid_0[1495:1488]) ? 1 : 0;
assign detect_min[185][11] = (mid_1[1495:1488] < mid_0[1503:1496]) ? 1 : 0;
assign detect_min[185][12] = (mid_1[1495:1488] < mid_1[1487:1480]) ? 1 : 0;
assign detect_min[185][13] = (mid_1[1495:1488] < mid_1[1503:1496]) ? 1 : 0;
assign detect_min[185][14] = (mid_1[1495:1488] < mid_2[1487:1480]) ? 1 : 0;
assign detect_min[185][15] = (mid_1[1495:1488] < mid_2[1495:1488]) ? 1 : 0;
assign detect_min[185][16] = (mid_1[1495:1488] < mid_2[1503:1496]) ? 1 : 0;
assign detect_min[185][17] = (mid_1[1495:1488] < btm_0[1487:1480]) ? 1 : 0;
assign detect_min[185][18] = (mid_1[1495:1488] < btm_0[1495:1488]) ? 1 : 0;
assign detect_min[185][19] = (mid_1[1495:1488] < btm_0[1503:1496]) ? 1 : 0;
assign detect_min[185][20] = (mid_1[1495:1488] < btm_1[1487:1480]) ? 1 : 0;
assign detect_min[185][21] = (mid_1[1495:1488] < btm_1[1495:1488]) ? 1 : 0;
assign detect_min[185][22] = (mid_1[1495:1488] < btm_1[1503:1496]) ? 1 : 0;
assign detect_min[185][23] = (mid_1[1495:1488] < btm_2[1487:1480]) ? 1 : 0;
assign detect_min[185][24] = (mid_1[1495:1488] < btm_2[1495:1488]) ? 1 : 0;
assign detect_min[185][25] = (mid_1[1495:1488] < btm_2[1503:1496]) ? 1 : 0;

assign detect_min[186][0] = (mid_1[1503:1496] < top_0[1495:1488]) ? 1 : 0;
assign detect_min[186][1] = (mid_1[1503:1496] < top_0[1503:1496]) ? 1 : 0;
assign detect_min[186][2] = (mid_1[1503:1496] < top_0[1511:1504]) ? 1 : 0;
assign detect_min[186][3] = (mid_1[1503:1496] < top_1[1495:1488]) ? 1 : 0;
assign detect_min[186][4] = (mid_1[1503:1496] < top_1[1503:1496]) ? 1 : 0;
assign detect_min[186][5] = (mid_1[1503:1496] < top_1[1511:1504]) ? 1 : 0;
assign detect_min[186][6] = (mid_1[1503:1496] < top_2[1495:1488]) ? 1 : 0;
assign detect_min[186][7] = (mid_1[1503:1496] < top_2[1503:1496]) ? 1 : 0;
assign detect_min[186][8] = (mid_1[1503:1496] < top_2[1511:1504]) ? 1 : 0;
assign detect_min[186][9] = (mid_1[1503:1496] < mid_0[1495:1488]) ? 1 : 0;
assign detect_min[186][10] = (mid_1[1503:1496] < mid_0[1503:1496]) ? 1 : 0;
assign detect_min[186][11] = (mid_1[1503:1496] < mid_0[1511:1504]) ? 1 : 0;
assign detect_min[186][12] = (mid_1[1503:1496] < mid_1[1495:1488]) ? 1 : 0;
assign detect_min[186][13] = (mid_1[1503:1496] < mid_1[1511:1504]) ? 1 : 0;
assign detect_min[186][14] = (mid_1[1503:1496] < mid_2[1495:1488]) ? 1 : 0;
assign detect_min[186][15] = (mid_1[1503:1496] < mid_2[1503:1496]) ? 1 : 0;
assign detect_min[186][16] = (mid_1[1503:1496] < mid_2[1511:1504]) ? 1 : 0;
assign detect_min[186][17] = (mid_1[1503:1496] < btm_0[1495:1488]) ? 1 : 0;
assign detect_min[186][18] = (mid_1[1503:1496] < btm_0[1503:1496]) ? 1 : 0;
assign detect_min[186][19] = (mid_1[1503:1496] < btm_0[1511:1504]) ? 1 : 0;
assign detect_min[186][20] = (mid_1[1503:1496] < btm_1[1495:1488]) ? 1 : 0;
assign detect_min[186][21] = (mid_1[1503:1496] < btm_1[1503:1496]) ? 1 : 0;
assign detect_min[186][22] = (mid_1[1503:1496] < btm_1[1511:1504]) ? 1 : 0;
assign detect_min[186][23] = (mid_1[1503:1496] < btm_2[1495:1488]) ? 1 : 0;
assign detect_min[186][24] = (mid_1[1503:1496] < btm_2[1503:1496]) ? 1 : 0;
assign detect_min[186][25] = (mid_1[1503:1496] < btm_2[1511:1504]) ? 1 : 0;

assign detect_min[187][0] = (mid_1[1511:1504] < top_0[1503:1496]) ? 1 : 0;
assign detect_min[187][1] = (mid_1[1511:1504] < top_0[1511:1504]) ? 1 : 0;
assign detect_min[187][2] = (mid_1[1511:1504] < top_0[1519:1512]) ? 1 : 0;
assign detect_min[187][3] = (mid_1[1511:1504] < top_1[1503:1496]) ? 1 : 0;
assign detect_min[187][4] = (mid_1[1511:1504] < top_1[1511:1504]) ? 1 : 0;
assign detect_min[187][5] = (mid_1[1511:1504] < top_1[1519:1512]) ? 1 : 0;
assign detect_min[187][6] = (mid_1[1511:1504] < top_2[1503:1496]) ? 1 : 0;
assign detect_min[187][7] = (mid_1[1511:1504] < top_2[1511:1504]) ? 1 : 0;
assign detect_min[187][8] = (mid_1[1511:1504] < top_2[1519:1512]) ? 1 : 0;
assign detect_min[187][9] = (mid_1[1511:1504] < mid_0[1503:1496]) ? 1 : 0;
assign detect_min[187][10] = (mid_1[1511:1504] < mid_0[1511:1504]) ? 1 : 0;
assign detect_min[187][11] = (mid_1[1511:1504] < mid_0[1519:1512]) ? 1 : 0;
assign detect_min[187][12] = (mid_1[1511:1504] < mid_1[1503:1496]) ? 1 : 0;
assign detect_min[187][13] = (mid_1[1511:1504] < mid_1[1519:1512]) ? 1 : 0;
assign detect_min[187][14] = (mid_1[1511:1504] < mid_2[1503:1496]) ? 1 : 0;
assign detect_min[187][15] = (mid_1[1511:1504] < mid_2[1511:1504]) ? 1 : 0;
assign detect_min[187][16] = (mid_1[1511:1504] < mid_2[1519:1512]) ? 1 : 0;
assign detect_min[187][17] = (mid_1[1511:1504] < btm_0[1503:1496]) ? 1 : 0;
assign detect_min[187][18] = (mid_1[1511:1504] < btm_0[1511:1504]) ? 1 : 0;
assign detect_min[187][19] = (mid_1[1511:1504] < btm_0[1519:1512]) ? 1 : 0;
assign detect_min[187][20] = (mid_1[1511:1504] < btm_1[1503:1496]) ? 1 : 0;
assign detect_min[187][21] = (mid_1[1511:1504] < btm_1[1511:1504]) ? 1 : 0;
assign detect_min[187][22] = (mid_1[1511:1504] < btm_1[1519:1512]) ? 1 : 0;
assign detect_min[187][23] = (mid_1[1511:1504] < btm_2[1503:1496]) ? 1 : 0;
assign detect_min[187][24] = (mid_1[1511:1504] < btm_2[1511:1504]) ? 1 : 0;
assign detect_min[187][25] = (mid_1[1511:1504] < btm_2[1519:1512]) ? 1 : 0;

assign detect_min[188][0] = (mid_1[1519:1512] < top_0[1511:1504]) ? 1 : 0;
assign detect_min[188][1] = (mid_1[1519:1512] < top_0[1519:1512]) ? 1 : 0;
assign detect_min[188][2] = (mid_1[1519:1512] < top_0[1527:1520]) ? 1 : 0;
assign detect_min[188][3] = (mid_1[1519:1512] < top_1[1511:1504]) ? 1 : 0;
assign detect_min[188][4] = (mid_1[1519:1512] < top_1[1519:1512]) ? 1 : 0;
assign detect_min[188][5] = (mid_1[1519:1512] < top_1[1527:1520]) ? 1 : 0;
assign detect_min[188][6] = (mid_1[1519:1512] < top_2[1511:1504]) ? 1 : 0;
assign detect_min[188][7] = (mid_1[1519:1512] < top_2[1519:1512]) ? 1 : 0;
assign detect_min[188][8] = (mid_1[1519:1512] < top_2[1527:1520]) ? 1 : 0;
assign detect_min[188][9] = (mid_1[1519:1512] < mid_0[1511:1504]) ? 1 : 0;
assign detect_min[188][10] = (mid_1[1519:1512] < mid_0[1519:1512]) ? 1 : 0;
assign detect_min[188][11] = (mid_1[1519:1512] < mid_0[1527:1520]) ? 1 : 0;
assign detect_min[188][12] = (mid_1[1519:1512] < mid_1[1511:1504]) ? 1 : 0;
assign detect_min[188][13] = (mid_1[1519:1512] < mid_1[1527:1520]) ? 1 : 0;
assign detect_min[188][14] = (mid_1[1519:1512] < mid_2[1511:1504]) ? 1 : 0;
assign detect_min[188][15] = (mid_1[1519:1512] < mid_2[1519:1512]) ? 1 : 0;
assign detect_min[188][16] = (mid_1[1519:1512] < mid_2[1527:1520]) ? 1 : 0;
assign detect_min[188][17] = (mid_1[1519:1512] < btm_0[1511:1504]) ? 1 : 0;
assign detect_min[188][18] = (mid_1[1519:1512] < btm_0[1519:1512]) ? 1 : 0;
assign detect_min[188][19] = (mid_1[1519:1512] < btm_0[1527:1520]) ? 1 : 0;
assign detect_min[188][20] = (mid_1[1519:1512] < btm_1[1511:1504]) ? 1 : 0;
assign detect_min[188][21] = (mid_1[1519:1512] < btm_1[1519:1512]) ? 1 : 0;
assign detect_min[188][22] = (mid_1[1519:1512] < btm_1[1527:1520]) ? 1 : 0;
assign detect_min[188][23] = (mid_1[1519:1512] < btm_2[1511:1504]) ? 1 : 0;
assign detect_min[188][24] = (mid_1[1519:1512] < btm_2[1519:1512]) ? 1 : 0;
assign detect_min[188][25] = (mid_1[1519:1512] < btm_2[1527:1520]) ? 1 : 0;

assign detect_min[189][0] = (mid_1[1527:1520] < top_0[1519:1512]) ? 1 : 0;
assign detect_min[189][1] = (mid_1[1527:1520] < top_0[1527:1520]) ? 1 : 0;
assign detect_min[189][2] = (mid_1[1527:1520] < top_0[1535:1528]) ? 1 : 0;
assign detect_min[189][3] = (mid_1[1527:1520] < top_1[1519:1512]) ? 1 : 0;
assign detect_min[189][4] = (mid_1[1527:1520] < top_1[1527:1520]) ? 1 : 0;
assign detect_min[189][5] = (mid_1[1527:1520] < top_1[1535:1528]) ? 1 : 0;
assign detect_min[189][6] = (mid_1[1527:1520] < top_2[1519:1512]) ? 1 : 0;
assign detect_min[189][7] = (mid_1[1527:1520] < top_2[1527:1520]) ? 1 : 0;
assign detect_min[189][8] = (mid_1[1527:1520] < top_2[1535:1528]) ? 1 : 0;
assign detect_min[189][9] = (mid_1[1527:1520] < mid_0[1519:1512]) ? 1 : 0;
assign detect_min[189][10] = (mid_1[1527:1520] < mid_0[1527:1520]) ? 1 : 0;
assign detect_min[189][11] = (mid_1[1527:1520] < mid_0[1535:1528]) ? 1 : 0;
assign detect_min[189][12] = (mid_1[1527:1520] < mid_1[1519:1512]) ? 1 : 0;
assign detect_min[189][13] = (mid_1[1527:1520] < mid_1[1535:1528]) ? 1 : 0;
assign detect_min[189][14] = (mid_1[1527:1520] < mid_2[1519:1512]) ? 1 : 0;
assign detect_min[189][15] = (mid_1[1527:1520] < mid_2[1527:1520]) ? 1 : 0;
assign detect_min[189][16] = (mid_1[1527:1520] < mid_2[1535:1528]) ? 1 : 0;
assign detect_min[189][17] = (mid_1[1527:1520] < btm_0[1519:1512]) ? 1 : 0;
assign detect_min[189][18] = (mid_1[1527:1520] < btm_0[1527:1520]) ? 1 : 0;
assign detect_min[189][19] = (mid_1[1527:1520] < btm_0[1535:1528]) ? 1 : 0;
assign detect_min[189][20] = (mid_1[1527:1520] < btm_1[1519:1512]) ? 1 : 0;
assign detect_min[189][21] = (mid_1[1527:1520] < btm_1[1527:1520]) ? 1 : 0;
assign detect_min[189][22] = (mid_1[1527:1520] < btm_1[1535:1528]) ? 1 : 0;
assign detect_min[189][23] = (mid_1[1527:1520] < btm_2[1519:1512]) ? 1 : 0;
assign detect_min[189][24] = (mid_1[1527:1520] < btm_2[1527:1520]) ? 1 : 0;
assign detect_min[189][25] = (mid_1[1527:1520] < btm_2[1535:1528]) ? 1 : 0;

assign detect_min[190][0] = (mid_1[1535:1528] < top_0[1527:1520]) ? 1 : 0;
assign detect_min[190][1] = (mid_1[1535:1528] < top_0[1535:1528]) ? 1 : 0;
assign detect_min[190][2] = (mid_1[1535:1528] < top_0[1543:1536]) ? 1 : 0;
assign detect_min[190][3] = (mid_1[1535:1528] < top_1[1527:1520]) ? 1 : 0;
assign detect_min[190][4] = (mid_1[1535:1528] < top_1[1535:1528]) ? 1 : 0;
assign detect_min[190][5] = (mid_1[1535:1528] < top_1[1543:1536]) ? 1 : 0;
assign detect_min[190][6] = (mid_1[1535:1528] < top_2[1527:1520]) ? 1 : 0;
assign detect_min[190][7] = (mid_1[1535:1528] < top_2[1535:1528]) ? 1 : 0;
assign detect_min[190][8] = (mid_1[1535:1528] < top_2[1543:1536]) ? 1 : 0;
assign detect_min[190][9] = (mid_1[1535:1528] < mid_0[1527:1520]) ? 1 : 0;
assign detect_min[190][10] = (mid_1[1535:1528] < mid_0[1535:1528]) ? 1 : 0;
assign detect_min[190][11] = (mid_1[1535:1528] < mid_0[1543:1536]) ? 1 : 0;
assign detect_min[190][12] = (mid_1[1535:1528] < mid_1[1527:1520]) ? 1 : 0;
assign detect_min[190][13] = (mid_1[1535:1528] < mid_1[1543:1536]) ? 1 : 0;
assign detect_min[190][14] = (mid_1[1535:1528] < mid_2[1527:1520]) ? 1 : 0;
assign detect_min[190][15] = (mid_1[1535:1528] < mid_2[1535:1528]) ? 1 : 0;
assign detect_min[190][16] = (mid_1[1535:1528] < mid_2[1543:1536]) ? 1 : 0;
assign detect_min[190][17] = (mid_1[1535:1528] < btm_0[1527:1520]) ? 1 : 0;
assign detect_min[190][18] = (mid_1[1535:1528] < btm_0[1535:1528]) ? 1 : 0;
assign detect_min[190][19] = (mid_1[1535:1528] < btm_0[1543:1536]) ? 1 : 0;
assign detect_min[190][20] = (mid_1[1535:1528] < btm_1[1527:1520]) ? 1 : 0;
assign detect_min[190][21] = (mid_1[1535:1528] < btm_1[1535:1528]) ? 1 : 0;
assign detect_min[190][22] = (mid_1[1535:1528] < btm_1[1543:1536]) ? 1 : 0;
assign detect_min[190][23] = (mid_1[1535:1528] < btm_2[1527:1520]) ? 1 : 0;
assign detect_min[190][24] = (mid_1[1535:1528] < btm_2[1535:1528]) ? 1 : 0;
assign detect_min[190][25] = (mid_1[1535:1528] < btm_2[1543:1536]) ? 1 : 0;

assign detect_min[191][0] = (mid_1[1543:1536] < top_0[1535:1528]) ? 1 : 0;
assign detect_min[191][1] = (mid_1[1543:1536] < top_0[1543:1536]) ? 1 : 0;
assign detect_min[191][2] = (mid_1[1543:1536] < top_0[1551:1544]) ? 1 : 0;
assign detect_min[191][3] = (mid_1[1543:1536] < top_1[1535:1528]) ? 1 : 0;
assign detect_min[191][4] = (mid_1[1543:1536] < top_1[1543:1536]) ? 1 : 0;
assign detect_min[191][5] = (mid_1[1543:1536] < top_1[1551:1544]) ? 1 : 0;
assign detect_min[191][6] = (mid_1[1543:1536] < top_2[1535:1528]) ? 1 : 0;
assign detect_min[191][7] = (mid_1[1543:1536] < top_2[1543:1536]) ? 1 : 0;
assign detect_min[191][8] = (mid_1[1543:1536] < top_2[1551:1544]) ? 1 : 0;
assign detect_min[191][9] = (mid_1[1543:1536] < mid_0[1535:1528]) ? 1 : 0;
assign detect_min[191][10] = (mid_1[1543:1536] < mid_0[1543:1536]) ? 1 : 0;
assign detect_min[191][11] = (mid_1[1543:1536] < mid_0[1551:1544]) ? 1 : 0;
assign detect_min[191][12] = (mid_1[1543:1536] < mid_1[1535:1528]) ? 1 : 0;
assign detect_min[191][13] = (mid_1[1543:1536] < mid_1[1551:1544]) ? 1 : 0;
assign detect_min[191][14] = (mid_1[1543:1536] < mid_2[1535:1528]) ? 1 : 0;
assign detect_min[191][15] = (mid_1[1543:1536] < mid_2[1543:1536]) ? 1 : 0;
assign detect_min[191][16] = (mid_1[1543:1536] < mid_2[1551:1544]) ? 1 : 0;
assign detect_min[191][17] = (mid_1[1543:1536] < btm_0[1535:1528]) ? 1 : 0;
assign detect_min[191][18] = (mid_1[1543:1536] < btm_0[1543:1536]) ? 1 : 0;
assign detect_min[191][19] = (mid_1[1543:1536] < btm_0[1551:1544]) ? 1 : 0;
assign detect_min[191][20] = (mid_1[1543:1536] < btm_1[1535:1528]) ? 1 : 0;
assign detect_min[191][21] = (mid_1[1543:1536] < btm_1[1543:1536]) ? 1 : 0;
assign detect_min[191][22] = (mid_1[1543:1536] < btm_1[1551:1544]) ? 1 : 0;
assign detect_min[191][23] = (mid_1[1543:1536] < btm_2[1535:1528]) ? 1 : 0;
assign detect_min[191][24] = (mid_1[1543:1536] < btm_2[1543:1536]) ? 1 : 0;
assign detect_min[191][25] = (mid_1[1543:1536] < btm_2[1551:1544]) ? 1 : 0;

assign detect_min[192][0] = (mid_1[1551:1544] < top_0[1543:1536]) ? 1 : 0;
assign detect_min[192][1] = (mid_1[1551:1544] < top_0[1551:1544]) ? 1 : 0;
assign detect_min[192][2] = (mid_1[1551:1544] < top_0[1559:1552]) ? 1 : 0;
assign detect_min[192][3] = (mid_1[1551:1544] < top_1[1543:1536]) ? 1 : 0;
assign detect_min[192][4] = (mid_1[1551:1544] < top_1[1551:1544]) ? 1 : 0;
assign detect_min[192][5] = (mid_1[1551:1544] < top_1[1559:1552]) ? 1 : 0;
assign detect_min[192][6] = (mid_1[1551:1544] < top_2[1543:1536]) ? 1 : 0;
assign detect_min[192][7] = (mid_1[1551:1544] < top_2[1551:1544]) ? 1 : 0;
assign detect_min[192][8] = (mid_1[1551:1544] < top_2[1559:1552]) ? 1 : 0;
assign detect_min[192][9] = (mid_1[1551:1544] < mid_0[1543:1536]) ? 1 : 0;
assign detect_min[192][10] = (mid_1[1551:1544] < mid_0[1551:1544]) ? 1 : 0;
assign detect_min[192][11] = (mid_1[1551:1544] < mid_0[1559:1552]) ? 1 : 0;
assign detect_min[192][12] = (mid_1[1551:1544] < mid_1[1543:1536]) ? 1 : 0;
assign detect_min[192][13] = (mid_1[1551:1544] < mid_1[1559:1552]) ? 1 : 0;
assign detect_min[192][14] = (mid_1[1551:1544] < mid_2[1543:1536]) ? 1 : 0;
assign detect_min[192][15] = (mid_1[1551:1544] < mid_2[1551:1544]) ? 1 : 0;
assign detect_min[192][16] = (mid_1[1551:1544] < mid_2[1559:1552]) ? 1 : 0;
assign detect_min[192][17] = (mid_1[1551:1544] < btm_0[1543:1536]) ? 1 : 0;
assign detect_min[192][18] = (mid_1[1551:1544] < btm_0[1551:1544]) ? 1 : 0;
assign detect_min[192][19] = (mid_1[1551:1544] < btm_0[1559:1552]) ? 1 : 0;
assign detect_min[192][20] = (mid_1[1551:1544] < btm_1[1543:1536]) ? 1 : 0;
assign detect_min[192][21] = (mid_1[1551:1544] < btm_1[1551:1544]) ? 1 : 0;
assign detect_min[192][22] = (mid_1[1551:1544] < btm_1[1559:1552]) ? 1 : 0;
assign detect_min[192][23] = (mid_1[1551:1544] < btm_2[1543:1536]) ? 1 : 0;
assign detect_min[192][24] = (mid_1[1551:1544] < btm_2[1551:1544]) ? 1 : 0;
assign detect_min[192][25] = (mid_1[1551:1544] < btm_2[1559:1552]) ? 1 : 0;

assign detect_min[193][0] = (mid_1[1559:1552] < top_0[1551:1544]) ? 1 : 0;
assign detect_min[193][1] = (mid_1[1559:1552] < top_0[1559:1552]) ? 1 : 0;
assign detect_min[193][2] = (mid_1[1559:1552] < top_0[1567:1560]) ? 1 : 0;
assign detect_min[193][3] = (mid_1[1559:1552] < top_1[1551:1544]) ? 1 : 0;
assign detect_min[193][4] = (mid_1[1559:1552] < top_1[1559:1552]) ? 1 : 0;
assign detect_min[193][5] = (mid_1[1559:1552] < top_1[1567:1560]) ? 1 : 0;
assign detect_min[193][6] = (mid_1[1559:1552] < top_2[1551:1544]) ? 1 : 0;
assign detect_min[193][7] = (mid_1[1559:1552] < top_2[1559:1552]) ? 1 : 0;
assign detect_min[193][8] = (mid_1[1559:1552] < top_2[1567:1560]) ? 1 : 0;
assign detect_min[193][9] = (mid_1[1559:1552] < mid_0[1551:1544]) ? 1 : 0;
assign detect_min[193][10] = (mid_1[1559:1552] < mid_0[1559:1552]) ? 1 : 0;
assign detect_min[193][11] = (mid_1[1559:1552] < mid_0[1567:1560]) ? 1 : 0;
assign detect_min[193][12] = (mid_1[1559:1552] < mid_1[1551:1544]) ? 1 : 0;
assign detect_min[193][13] = (mid_1[1559:1552] < mid_1[1567:1560]) ? 1 : 0;
assign detect_min[193][14] = (mid_1[1559:1552] < mid_2[1551:1544]) ? 1 : 0;
assign detect_min[193][15] = (mid_1[1559:1552] < mid_2[1559:1552]) ? 1 : 0;
assign detect_min[193][16] = (mid_1[1559:1552] < mid_2[1567:1560]) ? 1 : 0;
assign detect_min[193][17] = (mid_1[1559:1552] < btm_0[1551:1544]) ? 1 : 0;
assign detect_min[193][18] = (mid_1[1559:1552] < btm_0[1559:1552]) ? 1 : 0;
assign detect_min[193][19] = (mid_1[1559:1552] < btm_0[1567:1560]) ? 1 : 0;
assign detect_min[193][20] = (mid_1[1559:1552] < btm_1[1551:1544]) ? 1 : 0;
assign detect_min[193][21] = (mid_1[1559:1552] < btm_1[1559:1552]) ? 1 : 0;
assign detect_min[193][22] = (mid_1[1559:1552] < btm_1[1567:1560]) ? 1 : 0;
assign detect_min[193][23] = (mid_1[1559:1552] < btm_2[1551:1544]) ? 1 : 0;
assign detect_min[193][24] = (mid_1[1559:1552] < btm_2[1559:1552]) ? 1 : 0;
assign detect_min[193][25] = (mid_1[1559:1552] < btm_2[1567:1560]) ? 1 : 0;

assign detect_min[194][0] = (mid_1[1567:1560] < top_0[1559:1552]) ? 1 : 0;
assign detect_min[194][1] = (mid_1[1567:1560] < top_0[1567:1560]) ? 1 : 0;
assign detect_min[194][2] = (mid_1[1567:1560] < top_0[1575:1568]) ? 1 : 0;
assign detect_min[194][3] = (mid_1[1567:1560] < top_1[1559:1552]) ? 1 : 0;
assign detect_min[194][4] = (mid_1[1567:1560] < top_1[1567:1560]) ? 1 : 0;
assign detect_min[194][5] = (mid_1[1567:1560] < top_1[1575:1568]) ? 1 : 0;
assign detect_min[194][6] = (mid_1[1567:1560] < top_2[1559:1552]) ? 1 : 0;
assign detect_min[194][7] = (mid_1[1567:1560] < top_2[1567:1560]) ? 1 : 0;
assign detect_min[194][8] = (mid_1[1567:1560] < top_2[1575:1568]) ? 1 : 0;
assign detect_min[194][9] = (mid_1[1567:1560] < mid_0[1559:1552]) ? 1 : 0;
assign detect_min[194][10] = (mid_1[1567:1560] < mid_0[1567:1560]) ? 1 : 0;
assign detect_min[194][11] = (mid_1[1567:1560] < mid_0[1575:1568]) ? 1 : 0;
assign detect_min[194][12] = (mid_1[1567:1560] < mid_1[1559:1552]) ? 1 : 0;
assign detect_min[194][13] = (mid_1[1567:1560] < mid_1[1575:1568]) ? 1 : 0;
assign detect_min[194][14] = (mid_1[1567:1560] < mid_2[1559:1552]) ? 1 : 0;
assign detect_min[194][15] = (mid_1[1567:1560] < mid_2[1567:1560]) ? 1 : 0;
assign detect_min[194][16] = (mid_1[1567:1560] < mid_2[1575:1568]) ? 1 : 0;
assign detect_min[194][17] = (mid_1[1567:1560] < btm_0[1559:1552]) ? 1 : 0;
assign detect_min[194][18] = (mid_1[1567:1560] < btm_0[1567:1560]) ? 1 : 0;
assign detect_min[194][19] = (mid_1[1567:1560] < btm_0[1575:1568]) ? 1 : 0;
assign detect_min[194][20] = (mid_1[1567:1560] < btm_1[1559:1552]) ? 1 : 0;
assign detect_min[194][21] = (mid_1[1567:1560] < btm_1[1567:1560]) ? 1 : 0;
assign detect_min[194][22] = (mid_1[1567:1560] < btm_1[1575:1568]) ? 1 : 0;
assign detect_min[194][23] = (mid_1[1567:1560] < btm_2[1559:1552]) ? 1 : 0;
assign detect_min[194][24] = (mid_1[1567:1560] < btm_2[1567:1560]) ? 1 : 0;
assign detect_min[194][25] = (mid_1[1567:1560] < btm_2[1575:1568]) ? 1 : 0;

assign detect_min[195][0] = (mid_1[1575:1568] < top_0[1567:1560]) ? 1 : 0;
assign detect_min[195][1] = (mid_1[1575:1568] < top_0[1575:1568]) ? 1 : 0;
assign detect_min[195][2] = (mid_1[1575:1568] < top_0[1583:1576]) ? 1 : 0;
assign detect_min[195][3] = (mid_1[1575:1568] < top_1[1567:1560]) ? 1 : 0;
assign detect_min[195][4] = (mid_1[1575:1568] < top_1[1575:1568]) ? 1 : 0;
assign detect_min[195][5] = (mid_1[1575:1568] < top_1[1583:1576]) ? 1 : 0;
assign detect_min[195][6] = (mid_1[1575:1568] < top_2[1567:1560]) ? 1 : 0;
assign detect_min[195][7] = (mid_1[1575:1568] < top_2[1575:1568]) ? 1 : 0;
assign detect_min[195][8] = (mid_1[1575:1568] < top_2[1583:1576]) ? 1 : 0;
assign detect_min[195][9] = (mid_1[1575:1568] < mid_0[1567:1560]) ? 1 : 0;
assign detect_min[195][10] = (mid_1[1575:1568] < mid_0[1575:1568]) ? 1 : 0;
assign detect_min[195][11] = (mid_1[1575:1568] < mid_0[1583:1576]) ? 1 : 0;
assign detect_min[195][12] = (mid_1[1575:1568] < mid_1[1567:1560]) ? 1 : 0;
assign detect_min[195][13] = (mid_1[1575:1568] < mid_1[1583:1576]) ? 1 : 0;
assign detect_min[195][14] = (mid_1[1575:1568] < mid_2[1567:1560]) ? 1 : 0;
assign detect_min[195][15] = (mid_1[1575:1568] < mid_2[1575:1568]) ? 1 : 0;
assign detect_min[195][16] = (mid_1[1575:1568] < mid_2[1583:1576]) ? 1 : 0;
assign detect_min[195][17] = (mid_1[1575:1568] < btm_0[1567:1560]) ? 1 : 0;
assign detect_min[195][18] = (mid_1[1575:1568] < btm_0[1575:1568]) ? 1 : 0;
assign detect_min[195][19] = (mid_1[1575:1568] < btm_0[1583:1576]) ? 1 : 0;
assign detect_min[195][20] = (mid_1[1575:1568] < btm_1[1567:1560]) ? 1 : 0;
assign detect_min[195][21] = (mid_1[1575:1568] < btm_1[1575:1568]) ? 1 : 0;
assign detect_min[195][22] = (mid_1[1575:1568] < btm_1[1583:1576]) ? 1 : 0;
assign detect_min[195][23] = (mid_1[1575:1568] < btm_2[1567:1560]) ? 1 : 0;
assign detect_min[195][24] = (mid_1[1575:1568] < btm_2[1575:1568]) ? 1 : 0;
assign detect_min[195][25] = (mid_1[1575:1568] < btm_2[1583:1576]) ? 1 : 0;

assign detect_min[196][0] = (mid_1[1583:1576] < top_0[1575:1568]) ? 1 : 0;
assign detect_min[196][1] = (mid_1[1583:1576] < top_0[1583:1576]) ? 1 : 0;
assign detect_min[196][2] = (mid_1[1583:1576] < top_0[1591:1584]) ? 1 : 0;
assign detect_min[196][3] = (mid_1[1583:1576] < top_1[1575:1568]) ? 1 : 0;
assign detect_min[196][4] = (mid_1[1583:1576] < top_1[1583:1576]) ? 1 : 0;
assign detect_min[196][5] = (mid_1[1583:1576] < top_1[1591:1584]) ? 1 : 0;
assign detect_min[196][6] = (mid_1[1583:1576] < top_2[1575:1568]) ? 1 : 0;
assign detect_min[196][7] = (mid_1[1583:1576] < top_2[1583:1576]) ? 1 : 0;
assign detect_min[196][8] = (mid_1[1583:1576] < top_2[1591:1584]) ? 1 : 0;
assign detect_min[196][9] = (mid_1[1583:1576] < mid_0[1575:1568]) ? 1 : 0;
assign detect_min[196][10] = (mid_1[1583:1576] < mid_0[1583:1576]) ? 1 : 0;
assign detect_min[196][11] = (mid_1[1583:1576] < mid_0[1591:1584]) ? 1 : 0;
assign detect_min[196][12] = (mid_1[1583:1576] < mid_1[1575:1568]) ? 1 : 0;
assign detect_min[196][13] = (mid_1[1583:1576] < mid_1[1591:1584]) ? 1 : 0;
assign detect_min[196][14] = (mid_1[1583:1576] < mid_2[1575:1568]) ? 1 : 0;
assign detect_min[196][15] = (mid_1[1583:1576] < mid_2[1583:1576]) ? 1 : 0;
assign detect_min[196][16] = (mid_1[1583:1576] < mid_2[1591:1584]) ? 1 : 0;
assign detect_min[196][17] = (mid_1[1583:1576] < btm_0[1575:1568]) ? 1 : 0;
assign detect_min[196][18] = (mid_1[1583:1576] < btm_0[1583:1576]) ? 1 : 0;
assign detect_min[196][19] = (mid_1[1583:1576] < btm_0[1591:1584]) ? 1 : 0;
assign detect_min[196][20] = (mid_1[1583:1576] < btm_1[1575:1568]) ? 1 : 0;
assign detect_min[196][21] = (mid_1[1583:1576] < btm_1[1583:1576]) ? 1 : 0;
assign detect_min[196][22] = (mid_1[1583:1576] < btm_1[1591:1584]) ? 1 : 0;
assign detect_min[196][23] = (mid_1[1583:1576] < btm_2[1575:1568]) ? 1 : 0;
assign detect_min[196][24] = (mid_1[1583:1576] < btm_2[1583:1576]) ? 1 : 0;
assign detect_min[196][25] = (mid_1[1583:1576] < btm_2[1591:1584]) ? 1 : 0;

assign detect_min[197][0] = (mid_1[1591:1584] < top_0[1583:1576]) ? 1 : 0;
assign detect_min[197][1] = (mid_1[1591:1584] < top_0[1591:1584]) ? 1 : 0;
assign detect_min[197][2] = (mid_1[1591:1584] < top_0[1599:1592]) ? 1 : 0;
assign detect_min[197][3] = (mid_1[1591:1584] < top_1[1583:1576]) ? 1 : 0;
assign detect_min[197][4] = (mid_1[1591:1584] < top_1[1591:1584]) ? 1 : 0;
assign detect_min[197][5] = (mid_1[1591:1584] < top_1[1599:1592]) ? 1 : 0;
assign detect_min[197][6] = (mid_1[1591:1584] < top_2[1583:1576]) ? 1 : 0;
assign detect_min[197][7] = (mid_1[1591:1584] < top_2[1591:1584]) ? 1 : 0;
assign detect_min[197][8] = (mid_1[1591:1584] < top_2[1599:1592]) ? 1 : 0;
assign detect_min[197][9] = (mid_1[1591:1584] < mid_0[1583:1576]) ? 1 : 0;
assign detect_min[197][10] = (mid_1[1591:1584] < mid_0[1591:1584]) ? 1 : 0;
assign detect_min[197][11] = (mid_1[1591:1584] < mid_0[1599:1592]) ? 1 : 0;
assign detect_min[197][12] = (mid_1[1591:1584] < mid_1[1583:1576]) ? 1 : 0;
assign detect_min[197][13] = (mid_1[1591:1584] < mid_1[1599:1592]) ? 1 : 0;
assign detect_min[197][14] = (mid_1[1591:1584] < mid_2[1583:1576]) ? 1 : 0;
assign detect_min[197][15] = (mid_1[1591:1584] < mid_2[1591:1584]) ? 1 : 0;
assign detect_min[197][16] = (mid_1[1591:1584] < mid_2[1599:1592]) ? 1 : 0;
assign detect_min[197][17] = (mid_1[1591:1584] < btm_0[1583:1576]) ? 1 : 0;
assign detect_min[197][18] = (mid_1[1591:1584] < btm_0[1591:1584]) ? 1 : 0;
assign detect_min[197][19] = (mid_1[1591:1584] < btm_0[1599:1592]) ? 1 : 0;
assign detect_min[197][20] = (mid_1[1591:1584] < btm_1[1583:1576]) ? 1 : 0;
assign detect_min[197][21] = (mid_1[1591:1584] < btm_1[1591:1584]) ? 1 : 0;
assign detect_min[197][22] = (mid_1[1591:1584] < btm_1[1599:1592]) ? 1 : 0;
assign detect_min[197][23] = (mid_1[1591:1584] < btm_2[1583:1576]) ? 1 : 0;
assign detect_min[197][24] = (mid_1[1591:1584] < btm_2[1591:1584]) ? 1 : 0;
assign detect_min[197][25] = (mid_1[1591:1584] < btm_2[1599:1592]) ? 1 : 0;

assign detect_min[198][0] = (mid_1[1599:1592] < top_0[1591:1584]) ? 1 : 0;
assign detect_min[198][1] = (mid_1[1599:1592] < top_0[1599:1592]) ? 1 : 0;
assign detect_min[198][2] = (mid_1[1599:1592] < top_0[1607:1600]) ? 1 : 0;
assign detect_min[198][3] = (mid_1[1599:1592] < top_1[1591:1584]) ? 1 : 0;
assign detect_min[198][4] = (mid_1[1599:1592] < top_1[1599:1592]) ? 1 : 0;
assign detect_min[198][5] = (mid_1[1599:1592] < top_1[1607:1600]) ? 1 : 0;
assign detect_min[198][6] = (mid_1[1599:1592] < top_2[1591:1584]) ? 1 : 0;
assign detect_min[198][7] = (mid_1[1599:1592] < top_2[1599:1592]) ? 1 : 0;
assign detect_min[198][8] = (mid_1[1599:1592] < top_2[1607:1600]) ? 1 : 0;
assign detect_min[198][9] = (mid_1[1599:1592] < mid_0[1591:1584]) ? 1 : 0;
assign detect_min[198][10] = (mid_1[1599:1592] < mid_0[1599:1592]) ? 1 : 0;
assign detect_min[198][11] = (mid_1[1599:1592] < mid_0[1607:1600]) ? 1 : 0;
assign detect_min[198][12] = (mid_1[1599:1592] < mid_1[1591:1584]) ? 1 : 0;
assign detect_min[198][13] = (mid_1[1599:1592] < mid_1[1607:1600]) ? 1 : 0;
assign detect_min[198][14] = (mid_1[1599:1592] < mid_2[1591:1584]) ? 1 : 0;
assign detect_min[198][15] = (mid_1[1599:1592] < mid_2[1599:1592]) ? 1 : 0;
assign detect_min[198][16] = (mid_1[1599:1592] < mid_2[1607:1600]) ? 1 : 0;
assign detect_min[198][17] = (mid_1[1599:1592] < btm_0[1591:1584]) ? 1 : 0;
assign detect_min[198][18] = (mid_1[1599:1592] < btm_0[1599:1592]) ? 1 : 0;
assign detect_min[198][19] = (mid_1[1599:1592] < btm_0[1607:1600]) ? 1 : 0;
assign detect_min[198][20] = (mid_1[1599:1592] < btm_1[1591:1584]) ? 1 : 0;
assign detect_min[198][21] = (mid_1[1599:1592] < btm_1[1599:1592]) ? 1 : 0;
assign detect_min[198][22] = (mid_1[1599:1592] < btm_1[1607:1600]) ? 1 : 0;
assign detect_min[198][23] = (mid_1[1599:1592] < btm_2[1591:1584]) ? 1 : 0;
assign detect_min[198][24] = (mid_1[1599:1592] < btm_2[1599:1592]) ? 1 : 0;
assign detect_min[198][25] = (mid_1[1599:1592] < btm_2[1607:1600]) ? 1 : 0;

assign detect_min[199][0] = (mid_1[1607:1600] < top_0[1599:1592]) ? 1 : 0;
assign detect_min[199][1] = (mid_1[1607:1600] < top_0[1607:1600]) ? 1 : 0;
assign detect_min[199][2] = (mid_1[1607:1600] < top_0[1615:1608]) ? 1 : 0;
assign detect_min[199][3] = (mid_1[1607:1600] < top_1[1599:1592]) ? 1 : 0;
assign detect_min[199][4] = (mid_1[1607:1600] < top_1[1607:1600]) ? 1 : 0;
assign detect_min[199][5] = (mid_1[1607:1600] < top_1[1615:1608]) ? 1 : 0;
assign detect_min[199][6] = (mid_1[1607:1600] < top_2[1599:1592]) ? 1 : 0;
assign detect_min[199][7] = (mid_1[1607:1600] < top_2[1607:1600]) ? 1 : 0;
assign detect_min[199][8] = (mid_1[1607:1600] < top_2[1615:1608]) ? 1 : 0;
assign detect_min[199][9] = (mid_1[1607:1600] < mid_0[1599:1592]) ? 1 : 0;
assign detect_min[199][10] = (mid_1[1607:1600] < mid_0[1607:1600]) ? 1 : 0;
assign detect_min[199][11] = (mid_1[1607:1600] < mid_0[1615:1608]) ? 1 : 0;
assign detect_min[199][12] = (mid_1[1607:1600] < mid_1[1599:1592]) ? 1 : 0;
assign detect_min[199][13] = (mid_1[1607:1600] < mid_1[1615:1608]) ? 1 : 0;
assign detect_min[199][14] = (mid_1[1607:1600] < mid_2[1599:1592]) ? 1 : 0;
assign detect_min[199][15] = (mid_1[1607:1600] < mid_2[1607:1600]) ? 1 : 0;
assign detect_min[199][16] = (mid_1[1607:1600] < mid_2[1615:1608]) ? 1 : 0;
assign detect_min[199][17] = (mid_1[1607:1600] < btm_0[1599:1592]) ? 1 : 0;
assign detect_min[199][18] = (mid_1[1607:1600] < btm_0[1607:1600]) ? 1 : 0;
assign detect_min[199][19] = (mid_1[1607:1600] < btm_0[1615:1608]) ? 1 : 0;
assign detect_min[199][20] = (mid_1[1607:1600] < btm_1[1599:1592]) ? 1 : 0;
assign detect_min[199][21] = (mid_1[1607:1600] < btm_1[1607:1600]) ? 1 : 0;
assign detect_min[199][22] = (mid_1[1607:1600] < btm_1[1615:1608]) ? 1 : 0;
assign detect_min[199][23] = (mid_1[1607:1600] < btm_2[1599:1592]) ? 1 : 0;
assign detect_min[199][24] = (mid_1[1607:1600] < btm_2[1607:1600]) ? 1 : 0;
assign detect_min[199][25] = (mid_1[1607:1600] < btm_2[1615:1608]) ? 1 : 0;

assign detect_min[200][0] = (mid_1[1615:1608] < top_0[1607:1600]) ? 1 : 0;
assign detect_min[200][1] = (mid_1[1615:1608] < top_0[1615:1608]) ? 1 : 0;
assign detect_min[200][2] = (mid_1[1615:1608] < top_0[1623:1616]) ? 1 : 0;
assign detect_min[200][3] = (mid_1[1615:1608] < top_1[1607:1600]) ? 1 : 0;
assign detect_min[200][4] = (mid_1[1615:1608] < top_1[1615:1608]) ? 1 : 0;
assign detect_min[200][5] = (mid_1[1615:1608] < top_1[1623:1616]) ? 1 : 0;
assign detect_min[200][6] = (mid_1[1615:1608] < top_2[1607:1600]) ? 1 : 0;
assign detect_min[200][7] = (mid_1[1615:1608] < top_2[1615:1608]) ? 1 : 0;
assign detect_min[200][8] = (mid_1[1615:1608] < top_2[1623:1616]) ? 1 : 0;
assign detect_min[200][9] = (mid_1[1615:1608] < mid_0[1607:1600]) ? 1 : 0;
assign detect_min[200][10] = (mid_1[1615:1608] < mid_0[1615:1608]) ? 1 : 0;
assign detect_min[200][11] = (mid_1[1615:1608] < mid_0[1623:1616]) ? 1 : 0;
assign detect_min[200][12] = (mid_1[1615:1608] < mid_1[1607:1600]) ? 1 : 0;
assign detect_min[200][13] = (mid_1[1615:1608] < mid_1[1623:1616]) ? 1 : 0;
assign detect_min[200][14] = (mid_1[1615:1608] < mid_2[1607:1600]) ? 1 : 0;
assign detect_min[200][15] = (mid_1[1615:1608] < mid_2[1615:1608]) ? 1 : 0;
assign detect_min[200][16] = (mid_1[1615:1608] < mid_2[1623:1616]) ? 1 : 0;
assign detect_min[200][17] = (mid_1[1615:1608] < btm_0[1607:1600]) ? 1 : 0;
assign detect_min[200][18] = (mid_1[1615:1608] < btm_0[1615:1608]) ? 1 : 0;
assign detect_min[200][19] = (mid_1[1615:1608] < btm_0[1623:1616]) ? 1 : 0;
assign detect_min[200][20] = (mid_1[1615:1608] < btm_1[1607:1600]) ? 1 : 0;
assign detect_min[200][21] = (mid_1[1615:1608] < btm_1[1615:1608]) ? 1 : 0;
assign detect_min[200][22] = (mid_1[1615:1608] < btm_1[1623:1616]) ? 1 : 0;
assign detect_min[200][23] = (mid_1[1615:1608] < btm_2[1607:1600]) ? 1 : 0;
assign detect_min[200][24] = (mid_1[1615:1608] < btm_2[1615:1608]) ? 1 : 0;
assign detect_min[200][25] = (mid_1[1615:1608] < btm_2[1623:1616]) ? 1 : 0;

assign detect_min[201][0] = (mid_1[1623:1616] < top_0[1615:1608]) ? 1 : 0;
assign detect_min[201][1] = (mid_1[1623:1616] < top_0[1623:1616]) ? 1 : 0;
assign detect_min[201][2] = (mid_1[1623:1616] < top_0[1631:1624]) ? 1 : 0;
assign detect_min[201][3] = (mid_1[1623:1616] < top_1[1615:1608]) ? 1 : 0;
assign detect_min[201][4] = (mid_1[1623:1616] < top_1[1623:1616]) ? 1 : 0;
assign detect_min[201][5] = (mid_1[1623:1616] < top_1[1631:1624]) ? 1 : 0;
assign detect_min[201][6] = (mid_1[1623:1616] < top_2[1615:1608]) ? 1 : 0;
assign detect_min[201][7] = (mid_1[1623:1616] < top_2[1623:1616]) ? 1 : 0;
assign detect_min[201][8] = (mid_1[1623:1616] < top_2[1631:1624]) ? 1 : 0;
assign detect_min[201][9] = (mid_1[1623:1616] < mid_0[1615:1608]) ? 1 : 0;
assign detect_min[201][10] = (mid_1[1623:1616] < mid_0[1623:1616]) ? 1 : 0;
assign detect_min[201][11] = (mid_1[1623:1616] < mid_0[1631:1624]) ? 1 : 0;
assign detect_min[201][12] = (mid_1[1623:1616] < mid_1[1615:1608]) ? 1 : 0;
assign detect_min[201][13] = (mid_1[1623:1616] < mid_1[1631:1624]) ? 1 : 0;
assign detect_min[201][14] = (mid_1[1623:1616] < mid_2[1615:1608]) ? 1 : 0;
assign detect_min[201][15] = (mid_1[1623:1616] < mid_2[1623:1616]) ? 1 : 0;
assign detect_min[201][16] = (mid_1[1623:1616] < mid_2[1631:1624]) ? 1 : 0;
assign detect_min[201][17] = (mid_1[1623:1616] < btm_0[1615:1608]) ? 1 : 0;
assign detect_min[201][18] = (mid_1[1623:1616] < btm_0[1623:1616]) ? 1 : 0;
assign detect_min[201][19] = (mid_1[1623:1616] < btm_0[1631:1624]) ? 1 : 0;
assign detect_min[201][20] = (mid_1[1623:1616] < btm_1[1615:1608]) ? 1 : 0;
assign detect_min[201][21] = (mid_1[1623:1616] < btm_1[1623:1616]) ? 1 : 0;
assign detect_min[201][22] = (mid_1[1623:1616] < btm_1[1631:1624]) ? 1 : 0;
assign detect_min[201][23] = (mid_1[1623:1616] < btm_2[1615:1608]) ? 1 : 0;
assign detect_min[201][24] = (mid_1[1623:1616] < btm_2[1623:1616]) ? 1 : 0;
assign detect_min[201][25] = (mid_1[1623:1616] < btm_2[1631:1624]) ? 1 : 0;

assign detect_min[202][0] = (mid_1[1631:1624] < top_0[1623:1616]) ? 1 : 0;
assign detect_min[202][1] = (mid_1[1631:1624] < top_0[1631:1624]) ? 1 : 0;
assign detect_min[202][2] = (mid_1[1631:1624] < top_0[1639:1632]) ? 1 : 0;
assign detect_min[202][3] = (mid_1[1631:1624] < top_1[1623:1616]) ? 1 : 0;
assign detect_min[202][4] = (mid_1[1631:1624] < top_1[1631:1624]) ? 1 : 0;
assign detect_min[202][5] = (mid_1[1631:1624] < top_1[1639:1632]) ? 1 : 0;
assign detect_min[202][6] = (mid_1[1631:1624] < top_2[1623:1616]) ? 1 : 0;
assign detect_min[202][7] = (mid_1[1631:1624] < top_2[1631:1624]) ? 1 : 0;
assign detect_min[202][8] = (mid_1[1631:1624] < top_2[1639:1632]) ? 1 : 0;
assign detect_min[202][9] = (mid_1[1631:1624] < mid_0[1623:1616]) ? 1 : 0;
assign detect_min[202][10] = (mid_1[1631:1624] < mid_0[1631:1624]) ? 1 : 0;
assign detect_min[202][11] = (mid_1[1631:1624] < mid_0[1639:1632]) ? 1 : 0;
assign detect_min[202][12] = (mid_1[1631:1624] < mid_1[1623:1616]) ? 1 : 0;
assign detect_min[202][13] = (mid_1[1631:1624] < mid_1[1639:1632]) ? 1 : 0;
assign detect_min[202][14] = (mid_1[1631:1624] < mid_2[1623:1616]) ? 1 : 0;
assign detect_min[202][15] = (mid_1[1631:1624] < mid_2[1631:1624]) ? 1 : 0;
assign detect_min[202][16] = (mid_1[1631:1624] < mid_2[1639:1632]) ? 1 : 0;
assign detect_min[202][17] = (mid_1[1631:1624] < btm_0[1623:1616]) ? 1 : 0;
assign detect_min[202][18] = (mid_1[1631:1624] < btm_0[1631:1624]) ? 1 : 0;
assign detect_min[202][19] = (mid_1[1631:1624] < btm_0[1639:1632]) ? 1 : 0;
assign detect_min[202][20] = (mid_1[1631:1624] < btm_1[1623:1616]) ? 1 : 0;
assign detect_min[202][21] = (mid_1[1631:1624] < btm_1[1631:1624]) ? 1 : 0;
assign detect_min[202][22] = (mid_1[1631:1624] < btm_1[1639:1632]) ? 1 : 0;
assign detect_min[202][23] = (mid_1[1631:1624] < btm_2[1623:1616]) ? 1 : 0;
assign detect_min[202][24] = (mid_1[1631:1624] < btm_2[1631:1624]) ? 1 : 0;
assign detect_min[202][25] = (mid_1[1631:1624] < btm_2[1639:1632]) ? 1 : 0;

assign detect_min[203][0] = (mid_1[1639:1632] < top_0[1631:1624]) ? 1 : 0;
assign detect_min[203][1] = (mid_1[1639:1632] < top_0[1639:1632]) ? 1 : 0;
assign detect_min[203][2] = (mid_1[1639:1632] < top_0[1647:1640]) ? 1 : 0;
assign detect_min[203][3] = (mid_1[1639:1632] < top_1[1631:1624]) ? 1 : 0;
assign detect_min[203][4] = (mid_1[1639:1632] < top_1[1639:1632]) ? 1 : 0;
assign detect_min[203][5] = (mid_1[1639:1632] < top_1[1647:1640]) ? 1 : 0;
assign detect_min[203][6] = (mid_1[1639:1632] < top_2[1631:1624]) ? 1 : 0;
assign detect_min[203][7] = (mid_1[1639:1632] < top_2[1639:1632]) ? 1 : 0;
assign detect_min[203][8] = (mid_1[1639:1632] < top_2[1647:1640]) ? 1 : 0;
assign detect_min[203][9] = (mid_1[1639:1632] < mid_0[1631:1624]) ? 1 : 0;
assign detect_min[203][10] = (mid_1[1639:1632] < mid_0[1639:1632]) ? 1 : 0;
assign detect_min[203][11] = (mid_1[1639:1632] < mid_0[1647:1640]) ? 1 : 0;
assign detect_min[203][12] = (mid_1[1639:1632] < mid_1[1631:1624]) ? 1 : 0;
assign detect_min[203][13] = (mid_1[1639:1632] < mid_1[1647:1640]) ? 1 : 0;
assign detect_min[203][14] = (mid_1[1639:1632] < mid_2[1631:1624]) ? 1 : 0;
assign detect_min[203][15] = (mid_1[1639:1632] < mid_2[1639:1632]) ? 1 : 0;
assign detect_min[203][16] = (mid_1[1639:1632] < mid_2[1647:1640]) ? 1 : 0;
assign detect_min[203][17] = (mid_1[1639:1632] < btm_0[1631:1624]) ? 1 : 0;
assign detect_min[203][18] = (mid_1[1639:1632] < btm_0[1639:1632]) ? 1 : 0;
assign detect_min[203][19] = (mid_1[1639:1632] < btm_0[1647:1640]) ? 1 : 0;
assign detect_min[203][20] = (mid_1[1639:1632] < btm_1[1631:1624]) ? 1 : 0;
assign detect_min[203][21] = (mid_1[1639:1632] < btm_1[1639:1632]) ? 1 : 0;
assign detect_min[203][22] = (mid_1[1639:1632] < btm_1[1647:1640]) ? 1 : 0;
assign detect_min[203][23] = (mid_1[1639:1632] < btm_2[1631:1624]) ? 1 : 0;
assign detect_min[203][24] = (mid_1[1639:1632] < btm_2[1639:1632]) ? 1 : 0;
assign detect_min[203][25] = (mid_1[1639:1632] < btm_2[1647:1640]) ? 1 : 0;

assign detect_min[204][0] = (mid_1[1647:1640] < top_0[1639:1632]) ? 1 : 0;
assign detect_min[204][1] = (mid_1[1647:1640] < top_0[1647:1640]) ? 1 : 0;
assign detect_min[204][2] = (mid_1[1647:1640] < top_0[1655:1648]) ? 1 : 0;
assign detect_min[204][3] = (mid_1[1647:1640] < top_1[1639:1632]) ? 1 : 0;
assign detect_min[204][4] = (mid_1[1647:1640] < top_1[1647:1640]) ? 1 : 0;
assign detect_min[204][5] = (mid_1[1647:1640] < top_1[1655:1648]) ? 1 : 0;
assign detect_min[204][6] = (mid_1[1647:1640] < top_2[1639:1632]) ? 1 : 0;
assign detect_min[204][7] = (mid_1[1647:1640] < top_2[1647:1640]) ? 1 : 0;
assign detect_min[204][8] = (mid_1[1647:1640] < top_2[1655:1648]) ? 1 : 0;
assign detect_min[204][9] = (mid_1[1647:1640] < mid_0[1639:1632]) ? 1 : 0;
assign detect_min[204][10] = (mid_1[1647:1640] < mid_0[1647:1640]) ? 1 : 0;
assign detect_min[204][11] = (mid_1[1647:1640] < mid_0[1655:1648]) ? 1 : 0;
assign detect_min[204][12] = (mid_1[1647:1640] < mid_1[1639:1632]) ? 1 : 0;
assign detect_min[204][13] = (mid_1[1647:1640] < mid_1[1655:1648]) ? 1 : 0;
assign detect_min[204][14] = (mid_1[1647:1640] < mid_2[1639:1632]) ? 1 : 0;
assign detect_min[204][15] = (mid_1[1647:1640] < mid_2[1647:1640]) ? 1 : 0;
assign detect_min[204][16] = (mid_1[1647:1640] < mid_2[1655:1648]) ? 1 : 0;
assign detect_min[204][17] = (mid_1[1647:1640] < btm_0[1639:1632]) ? 1 : 0;
assign detect_min[204][18] = (mid_1[1647:1640] < btm_0[1647:1640]) ? 1 : 0;
assign detect_min[204][19] = (mid_1[1647:1640] < btm_0[1655:1648]) ? 1 : 0;
assign detect_min[204][20] = (mid_1[1647:1640] < btm_1[1639:1632]) ? 1 : 0;
assign detect_min[204][21] = (mid_1[1647:1640] < btm_1[1647:1640]) ? 1 : 0;
assign detect_min[204][22] = (mid_1[1647:1640] < btm_1[1655:1648]) ? 1 : 0;
assign detect_min[204][23] = (mid_1[1647:1640] < btm_2[1639:1632]) ? 1 : 0;
assign detect_min[204][24] = (mid_1[1647:1640] < btm_2[1647:1640]) ? 1 : 0;
assign detect_min[204][25] = (mid_1[1647:1640] < btm_2[1655:1648]) ? 1 : 0;

assign detect_min[205][0] = (mid_1[1655:1648] < top_0[1647:1640]) ? 1 : 0;
assign detect_min[205][1] = (mid_1[1655:1648] < top_0[1655:1648]) ? 1 : 0;
assign detect_min[205][2] = (mid_1[1655:1648] < top_0[1663:1656]) ? 1 : 0;
assign detect_min[205][3] = (mid_1[1655:1648] < top_1[1647:1640]) ? 1 : 0;
assign detect_min[205][4] = (mid_1[1655:1648] < top_1[1655:1648]) ? 1 : 0;
assign detect_min[205][5] = (mid_1[1655:1648] < top_1[1663:1656]) ? 1 : 0;
assign detect_min[205][6] = (mid_1[1655:1648] < top_2[1647:1640]) ? 1 : 0;
assign detect_min[205][7] = (mid_1[1655:1648] < top_2[1655:1648]) ? 1 : 0;
assign detect_min[205][8] = (mid_1[1655:1648] < top_2[1663:1656]) ? 1 : 0;
assign detect_min[205][9] = (mid_1[1655:1648] < mid_0[1647:1640]) ? 1 : 0;
assign detect_min[205][10] = (mid_1[1655:1648] < mid_0[1655:1648]) ? 1 : 0;
assign detect_min[205][11] = (mid_1[1655:1648] < mid_0[1663:1656]) ? 1 : 0;
assign detect_min[205][12] = (mid_1[1655:1648] < mid_1[1647:1640]) ? 1 : 0;
assign detect_min[205][13] = (mid_1[1655:1648] < mid_1[1663:1656]) ? 1 : 0;
assign detect_min[205][14] = (mid_1[1655:1648] < mid_2[1647:1640]) ? 1 : 0;
assign detect_min[205][15] = (mid_1[1655:1648] < mid_2[1655:1648]) ? 1 : 0;
assign detect_min[205][16] = (mid_1[1655:1648] < mid_2[1663:1656]) ? 1 : 0;
assign detect_min[205][17] = (mid_1[1655:1648] < btm_0[1647:1640]) ? 1 : 0;
assign detect_min[205][18] = (mid_1[1655:1648] < btm_0[1655:1648]) ? 1 : 0;
assign detect_min[205][19] = (mid_1[1655:1648] < btm_0[1663:1656]) ? 1 : 0;
assign detect_min[205][20] = (mid_1[1655:1648] < btm_1[1647:1640]) ? 1 : 0;
assign detect_min[205][21] = (mid_1[1655:1648] < btm_1[1655:1648]) ? 1 : 0;
assign detect_min[205][22] = (mid_1[1655:1648] < btm_1[1663:1656]) ? 1 : 0;
assign detect_min[205][23] = (mid_1[1655:1648] < btm_2[1647:1640]) ? 1 : 0;
assign detect_min[205][24] = (mid_1[1655:1648] < btm_2[1655:1648]) ? 1 : 0;
assign detect_min[205][25] = (mid_1[1655:1648] < btm_2[1663:1656]) ? 1 : 0;

assign detect_min[206][0] = (mid_1[1663:1656] < top_0[1655:1648]) ? 1 : 0;
assign detect_min[206][1] = (mid_1[1663:1656] < top_0[1663:1656]) ? 1 : 0;
assign detect_min[206][2] = (mid_1[1663:1656] < top_0[1671:1664]) ? 1 : 0;
assign detect_min[206][3] = (mid_1[1663:1656] < top_1[1655:1648]) ? 1 : 0;
assign detect_min[206][4] = (mid_1[1663:1656] < top_1[1663:1656]) ? 1 : 0;
assign detect_min[206][5] = (mid_1[1663:1656] < top_1[1671:1664]) ? 1 : 0;
assign detect_min[206][6] = (mid_1[1663:1656] < top_2[1655:1648]) ? 1 : 0;
assign detect_min[206][7] = (mid_1[1663:1656] < top_2[1663:1656]) ? 1 : 0;
assign detect_min[206][8] = (mid_1[1663:1656] < top_2[1671:1664]) ? 1 : 0;
assign detect_min[206][9] = (mid_1[1663:1656] < mid_0[1655:1648]) ? 1 : 0;
assign detect_min[206][10] = (mid_1[1663:1656] < mid_0[1663:1656]) ? 1 : 0;
assign detect_min[206][11] = (mid_1[1663:1656] < mid_0[1671:1664]) ? 1 : 0;
assign detect_min[206][12] = (mid_1[1663:1656] < mid_1[1655:1648]) ? 1 : 0;
assign detect_min[206][13] = (mid_1[1663:1656] < mid_1[1671:1664]) ? 1 : 0;
assign detect_min[206][14] = (mid_1[1663:1656] < mid_2[1655:1648]) ? 1 : 0;
assign detect_min[206][15] = (mid_1[1663:1656] < mid_2[1663:1656]) ? 1 : 0;
assign detect_min[206][16] = (mid_1[1663:1656] < mid_2[1671:1664]) ? 1 : 0;
assign detect_min[206][17] = (mid_1[1663:1656] < btm_0[1655:1648]) ? 1 : 0;
assign detect_min[206][18] = (mid_1[1663:1656] < btm_0[1663:1656]) ? 1 : 0;
assign detect_min[206][19] = (mid_1[1663:1656] < btm_0[1671:1664]) ? 1 : 0;
assign detect_min[206][20] = (mid_1[1663:1656] < btm_1[1655:1648]) ? 1 : 0;
assign detect_min[206][21] = (mid_1[1663:1656] < btm_1[1663:1656]) ? 1 : 0;
assign detect_min[206][22] = (mid_1[1663:1656] < btm_1[1671:1664]) ? 1 : 0;
assign detect_min[206][23] = (mid_1[1663:1656] < btm_2[1655:1648]) ? 1 : 0;
assign detect_min[206][24] = (mid_1[1663:1656] < btm_2[1663:1656]) ? 1 : 0;
assign detect_min[206][25] = (mid_1[1663:1656] < btm_2[1671:1664]) ? 1 : 0;

assign detect_min[207][0] = (mid_1[1671:1664] < top_0[1663:1656]) ? 1 : 0;
assign detect_min[207][1] = (mid_1[1671:1664] < top_0[1671:1664]) ? 1 : 0;
assign detect_min[207][2] = (mid_1[1671:1664] < top_0[1679:1672]) ? 1 : 0;
assign detect_min[207][3] = (mid_1[1671:1664] < top_1[1663:1656]) ? 1 : 0;
assign detect_min[207][4] = (mid_1[1671:1664] < top_1[1671:1664]) ? 1 : 0;
assign detect_min[207][5] = (mid_1[1671:1664] < top_1[1679:1672]) ? 1 : 0;
assign detect_min[207][6] = (mid_1[1671:1664] < top_2[1663:1656]) ? 1 : 0;
assign detect_min[207][7] = (mid_1[1671:1664] < top_2[1671:1664]) ? 1 : 0;
assign detect_min[207][8] = (mid_1[1671:1664] < top_2[1679:1672]) ? 1 : 0;
assign detect_min[207][9] = (mid_1[1671:1664] < mid_0[1663:1656]) ? 1 : 0;
assign detect_min[207][10] = (mid_1[1671:1664] < mid_0[1671:1664]) ? 1 : 0;
assign detect_min[207][11] = (mid_1[1671:1664] < mid_0[1679:1672]) ? 1 : 0;
assign detect_min[207][12] = (mid_1[1671:1664] < mid_1[1663:1656]) ? 1 : 0;
assign detect_min[207][13] = (mid_1[1671:1664] < mid_1[1679:1672]) ? 1 : 0;
assign detect_min[207][14] = (mid_1[1671:1664] < mid_2[1663:1656]) ? 1 : 0;
assign detect_min[207][15] = (mid_1[1671:1664] < mid_2[1671:1664]) ? 1 : 0;
assign detect_min[207][16] = (mid_1[1671:1664] < mid_2[1679:1672]) ? 1 : 0;
assign detect_min[207][17] = (mid_1[1671:1664] < btm_0[1663:1656]) ? 1 : 0;
assign detect_min[207][18] = (mid_1[1671:1664] < btm_0[1671:1664]) ? 1 : 0;
assign detect_min[207][19] = (mid_1[1671:1664] < btm_0[1679:1672]) ? 1 : 0;
assign detect_min[207][20] = (mid_1[1671:1664] < btm_1[1663:1656]) ? 1 : 0;
assign detect_min[207][21] = (mid_1[1671:1664] < btm_1[1671:1664]) ? 1 : 0;
assign detect_min[207][22] = (mid_1[1671:1664] < btm_1[1679:1672]) ? 1 : 0;
assign detect_min[207][23] = (mid_1[1671:1664] < btm_2[1663:1656]) ? 1 : 0;
assign detect_min[207][24] = (mid_1[1671:1664] < btm_2[1671:1664]) ? 1 : 0;
assign detect_min[207][25] = (mid_1[1671:1664] < btm_2[1679:1672]) ? 1 : 0;

assign detect_min[208][0] = (mid_1[1679:1672] < top_0[1671:1664]) ? 1 : 0;
assign detect_min[208][1] = (mid_1[1679:1672] < top_0[1679:1672]) ? 1 : 0;
assign detect_min[208][2] = (mid_1[1679:1672] < top_0[1687:1680]) ? 1 : 0;
assign detect_min[208][3] = (mid_1[1679:1672] < top_1[1671:1664]) ? 1 : 0;
assign detect_min[208][4] = (mid_1[1679:1672] < top_1[1679:1672]) ? 1 : 0;
assign detect_min[208][5] = (mid_1[1679:1672] < top_1[1687:1680]) ? 1 : 0;
assign detect_min[208][6] = (mid_1[1679:1672] < top_2[1671:1664]) ? 1 : 0;
assign detect_min[208][7] = (mid_1[1679:1672] < top_2[1679:1672]) ? 1 : 0;
assign detect_min[208][8] = (mid_1[1679:1672] < top_2[1687:1680]) ? 1 : 0;
assign detect_min[208][9] = (mid_1[1679:1672] < mid_0[1671:1664]) ? 1 : 0;
assign detect_min[208][10] = (mid_1[1679:1672] < mid_0[1679:1672]) ? 1 : 0;
assign detect_min[208][11] = (mid_1[1679:1672] < mid_0[1687:1680]) ? 1 : 0;
assign detect_min[208][12] = (mid_1[1679:1672] < mid_1[1671:1664]) ? 1 : 0;
assign detect_min[208][13] = (mid_1[1679:1672] < mid_1[1687:1680]) ? 1 : 0;
assign detect_min[208][14] = (mid_1[1679:1672] < mid_2[1671:1664]) ? 1 : 0;
assign detect_min[208][15] = (mid_1[1679:1672] < mid_2[1679:1672]) ? 1 : 0;
assign detect_min[208][16] = (mid_1[1679:1672] < mid_2[1687:1680]) ? 1 : 0;
assign detect_min[208][17] = (mid_1[1679:1672] < btm_0[1671:1664]) ? 1 : 0;
assign detect_min[208][18] = (mid_1[1679:1672] < btm_0[1679:1672]) ? 1 : 0;
assign detect_min[208][19] = (mid_1[1679:1672] < btm_0[1687:1680]) ? 1 : 0;
assign detect_min[208][20] = (mid_1[1679:1672] < btm_1[1671:1664]) ? 1 : 0;
assign detect_min[208][21] = (mid_1[1679:1672] < btm_1[1679:1672]) ? 1 : 0;
assign detect_min[208][22] = (mid_1[1679:1672] < btm_1[1687:1680]) ? 1 : 0;
assign detect_min[208][23] = (mid_1[1679:1672] < btm_2[1671:1664]) ? 1 : 0;
assign detect_min[208][24] = (mid_1[1679:1672] < btm_2[1679:1672]) ? 1 : 0;
assign detect_min[208][25] = (mid_1[1679:1672] < btm_2[1687:1680]) ? 1 : 0;

assign detect_min[209][0] = (mid_1[1687:1680] < top_0[1679:1672]) ? 1 : 0;
assign detect_min[209][1] = (mid_1[1687:1680] < top_0[1687:1680]) ? 1 : 0;
assign detect_min[209][2] = (mid_1[1687:1680] < top_0[1695:1688]) ? 1 : 0;
assign detect_min[209][3] = (mid_1[1687:1680] < top_1[1679:1672]) ? 1 : 0;
assign detect_min[209][4] = (mid_1[1687:1680] < top_1[1687:1680]) ? 1 : 0;
assign detect_min[209][5] = (mid_1[1687:1680] < top_1[1695:1688]) ? 1 : 0;
assign detect_min[209][6] = (mid_1[1687:1680] < top_2[1679:1672]) ? 1 : 0;
assign detect_min[209][7] = (mid_1[1687:1680] < top_2[1687:1680]) ? 1 : 0;
assign detect_min[209][8] = (mid_1[1687:1680] < top_2[1695:1688]) ? 1 : 0;
assign detect_min[209][9] = (mid_1[1687:1680] < mid_0[1679:1672]) ? 1 : 0;
assign detect_min[209][10] = (mid_1[1687:1680] < mid_0[1687:1680]) ? 1 : 0;
assign detect_min[209][11] = (mid_1[1687:1680] < mid_0[1695:1688]) ? 1 : 0;
assign detect_min[209][12] = (mid_1[1687:1680] < mid_1[1679:1672]) ? 1 : 0;
assign detect_min[209][13] = (mid_1[1687:1680] < mid_1[1695:1688]) ? 1 : 0;
assign detect_min[209][14] = (mid_1[1687:1680] < mid_2[1679:1672]) ? 1 : 0;
assign detect_min[209][15] = (mid_1[1687:1680] < mid_2[1687:1680]) ? 1 : 0;
assign detect_min[209][16] = (mid_1[1687:1680] < mid_2[1695:1688]) ? 1 : 0;
assign detect_min[209][17] = (mid_1[1687:1680] < btm_0[1679:1672]) ? 1 : 0;
assign detect_min[209][18] = (mid_1[1687:1680] < btm_0[1687:1680]) ? 1 : 0;
assign detect_min[209][19] = (mid_1[1687:1680] < btm_0[1695:1688]) ? 1 : 0;
assign detect_min[209][20] = (mid_1[1687:1680] < btm_1[1679:1672]) ? 1 : 0;
assign detect_min[209][21] = (mid_1[1687:1680] < btm_1[1687:1680]) ? 1 : 0;
assign detect_min[209][22] = (mid_1[1687:1680] < btm_1[1695:1688]) ? 1 : 0;
assign detect_min[209][23] = (mid_1[1687:1680] < btm_2[1679:1672]) ? 1 : 0;
assign detect_min[209][24] = (mid_1[1687:1680] < btm_2[1687:1680]) ? 1 : 0;
assign detect_min[209][25] = (mid_1[1687:1680] < btm_2[1695:1688]) ? 1 : 0;

assign detect_min[210][0] = (mid_1[1695:1688] < top_0[1687:1680]) ? 1 : 0;
assign detect_min[210][1] = (mid_1[1695:1688] < top_0[1695:1688]) ? 1 : 0;
assign detect_min[210][2] = (mid_1[1695:1688] < top_0[1703:1696]) ? 1 : 0;
assign detect_min[210][3] = (mid_1[1695:1688] < top_1[1687:1680]) ? 1 : 0;
assign detect_min[210][4] = (mid_1[1695:1688] < top_1[1695:1688]) ? 1 : 0;
assign detect_min[210][5] = (mid_1[1695:1688] < top_1[1703:1696]) ? 1 : 0;
assign detect_min[210][6] = (mid_1[1695:1688] < top_2[1687:1680]) ? 1 : 0;
assign detect_min[210][7] = (mid_1[1695:1688] < top_2[1695:1688]) ? 1 : 0;
assign detect_min[210][8] = (mid_1[1695:1688] < top_2[1703:1696]) ? 1 : 0;
assign detect_min[210][9] = (mid_1[1695:1688] < mid_0[1687:1680]) ? 1 : 0;
assign detect_min[210][10] = (mid_1[1695:1688] < mid_0[1695:1688]) ? 1 : 0;
assign detect_min[210][11] = (mid_1[1695:1688] < mid_0[1703:1696]) ? 1 : 0;
assign detect_min[210][12] = (mid_1[1695:1688] < mid_1[1687:1680]) ? 1 : 0;
assign detect_min[210][13] = (mid_1[1695:1688] < mid_1[1703:1696]) ? 1 : 0;
assign detect_min[210][14] = (mid_1[1695:1688] < mid_2[1687:1680]) ? 1 : 0;
assign detect_min[210][15] = (mid_1[1695:1688] < mid_2[1695:1688]) ? 1 : 0;
assign detect_min[210][16] = (mid_1[1695:1688] < mid_2[1703:1696]) ? 1 : 0;
assign detect_min[210][17] = (mid_1[1695:1688] < btm_0[1687:1680]) ? 1 : 0;
assign detect_min[210][18] = (mid_1[1695:1688] < btm_0[1695:1688]) ? 1 : 0;
assign detect_min[210][19] = (mid_1[1695:1688] < btm_0[1703:1696]) ? 1 : 0;
assign detect_min[210][20] = (mid_1[1695:1688] < btm_1[1687:1680]) ? 1 : 0;
assign detect_min[210][21] = (mid_1[1695:1688] < btm_1[1695:1688]) ? 1 : 0;
assign detect_min[210][22] = (mid_1[1695:1688] < btm_1[1703:1696]) ? 1 : 0;
assign detect_min[210][23] = (mid_1[1695:1688] < btm_2[1687:1680]) ? 1 : 0;
assign detect_min[210][24] = (mid_1[1695:1688] < btm_2[1695:1688]) ? 1 : 0;
assign detect_min[210][25] = (mid_1[1695:1688] < btm_2[1703:1696]) ? 1 : 0;

assign detect_min[211][0] = (mid_1[1703:1696] < top_0[1695:1688]) ? 1 : 0;
assign detect_min[211][1] = (mid_1[1703:1696] < top_0[1703:1696]) ? 1 : 0;
assign detect_min[211][2] = (mid_1[1703:1696] < top_0[1711:1704]) ? 1 : 0;
assign detect_min[211][3] = (mid_1[1703:1696] < top_1[1695:1688]) ? 1 : 0;
assign detect_min[211][4] = (mid_1[1703:1696] < top_1[1703:1696]) ? 1 : 0;
assign detect_min[211][5] = (mid_1[1703:1696] < top_1[1711:1704]) ? 1 : 0;
assign detect_min[211][6] = (mid_1[1703:1696] < top_2[1695:1688]) ? 1 : 0;
assign detect_min[211][7] = (mid_1[1703:1696] < top_2[1703:1696]) ? 1 : 0;
assign detect_min[211][8] = (mid_1[1703:1696] < top_2[1711:1704]) ? 1 : 0;
assign detect_min[211][9] = (mid_1[1703:1696] < mid_0[1695:1688]) ? 1 : 0;
assign detect_min[211][10] = (mid_1[1703:1696] < mid_0[1703:1696]) ? 1 : 0;
assign detect_min[211][11] = (mid_1[1703:1696] < mid_0[1711:1704]) ? 1 : 0;
assign detect_min[211][12] = (mid_1[1703:1696] < mid_1[1695:1688]) ? 1 : 0;
assign detect_min[211][13] = (mid_1[1703:1696] < mid_1[1711:1704]) ? 1 : 0;
assign detect_min[211][14] = (mid_1[1703:1696] < mid_2[1695:1688]) ? 1 : 0;
assign detect_min[211][15] = (mid_1[1703:1696] < mid_2[1703:1696]) ? 1 : 0;
assign detect_min[211][16] = (mid_1[1703:1696] < mid_2[1711:1704]) ? 1 : 0;
assign detect_min[211][17] = (mid_1[1703:1696] < btm_0[1695:1688]) ? 1 : 0;
assign detect_min[211][18] = (mid_1[1703:1696] < btm_0[1703:1696]) ? 1 : 0;
assign detect_min[211][19] = (mid_1[1703:1696] < btm_0[1711:1704]) ? 1 : 0;
assign detect_min[211][20] = (mid_1[1703:1696] < btm_1[1695:1688]) ? 1 : 0;
assign detect_min[211][21] = (mid_1[1703:1696] < btm_1[1703:1696]) ? 1 : 0;
assign detect_min[211][22] = (mid_1[1703:1696] < btm_1[1711:1704]) ? 1 : 0;
assign detect_min[211][23] = (mid_1[1703:1696] < btm_2[1695:1688]) ? 1 : 0;
assign detect_min[211][24] = (mid_1[1703:1696] < btm_2[1703:1696]) ? 1 : 0;
assign detect_min[211][25] = (mid_1[1703:1696] < btm_2[1711:1704]) ? 1 : 0;

assign detect_min[212][0] = (mid_1[1711:1704] < top_0[1703:1696]) ? 1 : 0;
assign detect_min[212][1] = (mid_1[1711:1704] < top_0[1711:1704]) ? 1 : 0;
assign detect_min[212][2] = (mid_1[1711:1704] < top_0[1719:1712]) ? 1 : 0;
assign detect_min[212][3] = (mid_1[1711:1704] < top_1[1703:1696]) ? 1 : 0;
assign detect_min[212][4] = (mid_1[1711:1704] < top_1[1711:1704]) ? 1 : 0;
assign detect_min[212][5] = (mid_1[1711:1704] < top_1[1719:1712]) ? 1 : 0;
assign detect_min[212][6] = (mid_1[1711:1704] < top_2[1703:1696]) ? 1 : 0;
assign detect_min[212][7] = (mid_1[1711:1704] < top_2[1711:1704]) ? 1 : 0;
assign detect_min[212][8] = (mid_1[1711:1704] < top_2[1719:1712]) ? 1 : 0;
assign detect_min[212][9] = (mid_1[1711:1704] < mid_0[1703:1696]) ? 1 : 0;
assign detect_min[212][10] = (mid_1[1711:1704] < mid_0[1711:1704]) ? 1 : 0;
assign detect_min[212][11] = (mid_1[1711:1704] < mid_0[1719:1712]) ? 1 : 0;
assign detect_min[212][12] = (mid_1[1711:1704] < mid_1[1703:1696]) ? 1 : 0;
assign detect_min[212][13] = (mid_1[1711:1704] < mid_1[1719:1712]) ? 1 : 0;
assign detect_min[212][14] = (mid_1[1711:1704] < mid_2[1703:1696]) ? 1 : 0;
assign detect_min[212][15] = (mid_1[1711:1704] < mid_2[1711:1704]) ? 1 : 0;
assign detect_min[212][16] = (mid_1[1711:1704] < mid_2[1719:1712]) ? 1 : 0;
assign detect_min[212][17] = (mid_1[1711:1704] < btm_0[1703:1696]) ? 1 : 0;
assign detect_min[212][18] = (mid_1[1711:1704] < btm_0[1711:1704]) ? 1 : 0;
assign detect_min[212][19] = (mid_1[1711:1704] < btm_0[1719:1712]) ? 1 : 0;
assign detect_min[212][20] = (mid_1[1711:1704] < btm_1[1703:1696]) ? 1 : 0;
assign detect_min[212][21] = (mid_1[1711:1704] < btm_1[1711:1704]) ? 1 : 0;
assign detect_min[212][22] = (mid_1[1711:1704] < btm_1[1719:1712]) ? 1 : 0;
assign detect_min[212][23] = (mid_1[1711:1704] < btm_2[1703:1696]) ? 1 : 0;
assign detect_min[212][24] = (mid_1[1711:1704] < btm_2[1711:1704]) ? 1 : 0;
assign detect_min[212][25] = (mid_1[1711:1704] < btm_2[1719:1712]) ? 1 : 0;

assign detect_min[213][0] = (mid_1[1719:1712] < top_0[1711:1704]) ? 1 : 0;
assign detect_min[213][1] = (mid_1[1719:1712] < top_0[1719:1712]) ? 1 : 0;
assign detect_min[213][2] = (mid_1[1719:1712] < top_0[1727:1720]) ? 1 : 0;
assign detect_min[213][3] = (mid_1[1719:1712] < top_1[1711:1704]) ? 1 : 0;
assign detect_min[213][4] = (mid_1[1719:1712] < top_1[1719:1712]) ? 1 : 0;
assign detect_min[213][5] = (mid_1[1719:1712] < top_1[1727:1720]) ? 1 : 0;
assign detect_min[213][6] = (mid_1[1719:1712] < top_2[1711:1704]) ? 1 : 0;
assign detect_min[213][7] = (mid_1[1719:1712] < top_2[1719:1712]) ? 1 : 0;
assign detect_min[213][8] = (mid_1[1719:1712] < top_2[1727:1720]) ? 1 : 0;
assign detect_min[213][9] = (mid_1[1719:1712] < mid_0[1711:1704]) ? 1 : 0;
assign detect_min[213][10] = (mid_1[1719:1712] < mid_0[1719:1712]) ? 1 : 0;
assign detect_min[213][11] = (mid_1[1719:1712] < mid_0[1727:1720]) ? 1 : 0;
assign detect_min[213][12] = (mid_1[1719:1712] < mid_1[1711:1704]) ? 1 : 0;
assign detect_min[213][13] = (mid_1[1719:1712] < mid_1[1727:1720]) ? 1 : 0;
assign detect_min[213][14] = (mid_1[1719:1712] < mid_2[1711:1704]) ? 1 : 0;
assign detect_min[213][15] = (mid_1[1719:1712] < mid_2[1719:1712]) ? 1 : 0;
assign detect_min[213][16] = (mid_1[1719:1712] < mid_2[1727:1720]) ? 1 : 0;
assign detect_min[213][17] = (mid_1[1719:1712] < btm_0[1711:1704]) ? 1 : 0;
assign detect_min[213][18] = (mid_1[1719:1712] < btm_0[1719:1712]) ? 1 : 0;
assign detect_min[213][19] = (mid_1[1719:1712] < btm_0[1727:1720]) ? 1 : 0;
assign detect_min[213][20] = (mid_1[1719:1712] < btm_1[1711:1704]) ? 1 : 0;
assign detect_min[213][21] = (mid_1[1719:1712] < btm_1[1719:1712]) ? 1 : 0;
assign detect_min[213][22] = (mid_1[1719:1712] < btm_1[1727:1720]) ? 1 : 0;
assign detect_min[213][23] = (mid_1[1719:1712] < btm_2[1711:1704]) ? 1 : 0;
assign detect_min[213][24] = (mid_1[1719:1712] < btm_2[1719:1712]) ? 1 : 0;
assign detect_min[213][25] = (mid_1[1719:1712] < btm_2[1727:1720]) ? 1 : 0;

assign detect_min[214][0] = (mid_1[1727:1720] < top_0[1719:1712]) ? 1 : 0;
assign detect_min[214][1] = (mid_1[1727:1720] < top_0[1727:1720]) ? 1 : 0;
assign detect_min[214][2] = (mid_1[1727:1720] < top_0[1735:1728]) ? 1 : 0;
assign detect_min[214][3] = (mid_1[1727:1720] < top_1[1719:1712]) ? 1 : 0;
assign detect_min[214][4] = (mid_1[1727:1720] < top_1[1727:1720]) ? 1 : 0;
assign detect_min[214][5] = (mid_1[1727:1720] < top_1[1735:1728]) ? 1 : 0;
assign detect_min[214][6] = (mid_1[1727:1720] < top_2[1719:1712]) ? 1 : 0;
assign detect_min[214][7] = (mid_1[1727:1720] < top_2[1727:1720]) ? 1 : 0;
assign detect_min[214][8] = (mid_1[1727:1720] < top_2[1735:1728]) ? 1 : 0;
assign detect_min[214][9] = (mid_1[1727:1720] < mid_0[1719:1712]) ? 1 : 0;
assign detect_min[214][10] = (mid_1[1727:1720] < mid_0[1727:1720]) ? 1 : 0;
assign detect_min[214][11] = (mid_1[1727:1720] < mid_0[1735:1728]) ? 1 : 0;
assign detect_min[214][12] = (mid_1[1727:1720] < mid_1[1719:1712]) ? 1 : 0;
assign detect_min[214][13] = (mid_1[1727:1720] < mid_1[1735:1728]) ? 1 : 0;
assign detect_min[214][14] = (mid_1[1727:1720] < mid_2[1719:1712]) ? 1 : 0;
assign detect_min[214][15] = (mid_1[1727:1720] < mid_2[1727:1720]) ? 1 : 0;
assign detect_min[214][16] = (mid_1[1727:1720] < mid_2[1735:1728]) ? 1 : 0;
assign detect_min[214][17] = (mid_1[1727:1720] < btm_0[1719:1712]) ? 1 : 0;
assign detect_min[214][18] = (mid_1[1727:1720] < btm_0[1727:1720]) ? 1 : 0;
assign detect_min[214][19] = (mid_1[1727:1720] < btm_0[1735:1728]) ? 1 : 0;
assign detect_min[214][20] = (mid_1[1727:1720] < btm_1[1719:1712]) ? 1 : 0;
assign detect_min[214][21] = (mid_1[1727:1720] < btm_1[1727:1720]) ? 1 : 0;
assign detect_min[214][22] = (mid_1[1727:1720] < btm_1[1735:1728]) ? 1 : 0;
assign detect_min[214][23] = (mid_1[1727:1720] < btm_2[1719:1712]) ? 1 : 0;
assign detect_min[214][24] = (mid_1[1727:1720] < btm_2[1727:1720]) ? 1 : 0;
assign detect_min[214][25] = (mid_1[1727:1720] < btm_2[1735:1728]) ? 1 : 0;

assign detect_min[215][0] = (mid_1[1735:1728] < top_0[1727:1720]) ? 1 : 0;
assign detect_min[215][1] = (mid_1[1735:1728] < top_0[1735:1728]) ? 1 : 0;
assign detect_min[215][2] = (mid_1[1735:1728] < top_0[1743:1736]) ? 1 : 0;
assign detect_min[215][3] = (mid_1[1735:1728] < top_1[1727:1720]) ? 1 : 0;
assign detect_min[215][4] = (mid_1[1735:1728] < top_1[1735:1728]) ? 1 : 0;
assign detect_min[215][5] = (mid_1[1735:1728] < top_1[1743:1736]) ? 1 : 0;
assign detect_min[215][6] = (mid_1[1735:1728] < top_2[1727:1720]) ? 1 : 0;
assign detect_min[215][7] = (mid_1[1735:1728] < top_2[1735:1728]) ? 1 : 0;
assign detect_min[215][8] = (mid_1[1735:1728] < top_2[1743:1736]) ? 1 : 0;
assign detect_min[215][9] = (mid_1[1735:1728] < mid_0[1727:1720]) ? 1 : 0;
assign detect_min[215][10] = (mid_1[1735:1728] < mid_0[1735:1728]) ? 1 : 0;
assign detect_min[215][11] = (mid_1[1735:1728] < mid_0[1743:1736]) ? 1 : 0;
assign detect_min[215][12] = (mid_1[1735:1728] < mid_1[1727:1720]) ? 1 : 0;
assign detect_min[215][13] = (mid_1[1735:1728] < mid_1[1743:1736]) ? 1 : 0;
assign detect_min[215][14] = (mid_1[1735:1728] < mid_2[1727:1720]) ? 1 : 0;
assign detect_min[215][15] = (mid_1[1735:1728] < mid_2[1735:1728]) ? 1 : 0;
assign detect_min[215][16] = (mid_1[1735:1728] < mid_2[1743:1736]) ? 1 : 0;
assign detect_min[215][17] = (mid_1[1735:1728] < btm_0[1727:1720]) ? 1 : 0;
assign detect_min[215][18] = (mid_1[1735:1728] < btm_0[1735:1728]) ? 1 : 0;
assign detect_min[215][19] = (mid_1[1735:1728] < btm_0[1743:1736]) ? 1 : 0;
assign detect_min[215][20] = (mid_1[1735:1728] < btm_1[1727:1720]) ? 1 : 0;
assign detect_min[215][21] = (mid_1[1735:1728] < btm_1[1735:1728]) ? 1 : 0;
assign detect_min[215][22] = (mid_1[1735:1728] < btm_1[1743:1736]) ? 1 : 0;
assign detect_min[215][23] = (mid_1[1735:1728] < btm_2[1727:1720]) ? 1 : 0;
assign detect_min[215][24] = (mid_1[1735:1728] < btm_2[1735:1728]) ? 1 : 0;
assign detect_min[215][25] = (mid_1[1735:1728] < btm_2[1743:1736]) ? 1 : 0;

assign detect_min[216][0] = (mid_1[1743:1736] < top_0[1735:1728]) ? 1 : 0;
assign detect_min[216][1] = (mid_1[1743:1736] < top_0[1743:1736]) ? 1 : 0;
assign detect_min[216][2] = (mid_1[1743:1736] < top_0[1751:1744]) ? 1 : 0;
assign detect_min[216][3] = (mid_1[1743:1736] < top_1[1735:1728]) ? 1 : 0;
assign detect_min[216][4] = (mid_1[1743:1736] < top_1[1743:1736]) ? 1 : 0;
assign detect_min[216][5] = (mid_1[1743:1736] < top_1[1751:1744]) ? 1 : 0;
assign detect_min[216][6] = (mid_1[1743:1736] < top_2[1735:1728]) ? 1 : 0;
assign detect_min[216][7] = (mid_1[1743:1736] < top_2[1743:1736]) ? 1 : 0;
assign detect_min[216][8] = (mid_1[1743:1736] < top_2[1751:1744]) ? 1 : 0;
assign detect_min[216][9] = (mid_1[1743:1736] < mid_0[1735:1728]) ? 1 : 0;
assign detect_min[216][10] = (mid_1[1743:1736] < mid_0[1743:1736]) ? 1 : 0;
assign detect_min[216][11] = (mid_1[1743:1736] < mid_0[1751:1744]) ? 1 : 0;
assign detect_min[216][12] = (mid_1[1743:1736] < mid_1[1735:1728]) ? 1 : 0;
assign detect_min[216][13] = (mid_1[1743:1736] < mid_1[1751:1744]) ? 1 : 0;
assign detect_min[216][14] = (mid_1[1743:1736] < mid_2[1735:1728]) ? 1 : 0;
assign detect_min[216][15] = (mid_1[1743:1736] < mid_2[1743:1736]) ? 1 : 0;
assign detect_min[216][16] = (mid_1[1743:1736] < mid_2[1751:1744]) ? 1 : 0;
assign detect_min[216][17] = (mid_1[1743:1736] < btm_0[1735:1728]) ? 1 : 0;
assign detect_min[216][18] = (mid_1[1743:1736] < btm_0[1743:1736]) ? 1 : 0;
assign detect_min[216][19] = (mid_1[1743:1736] < btm_0[1751:1744]) ? 1 : 0;
assign detect_min[216][20] = (mid_1[1743:1736] < btm_1[1735:1728]) ? 1 : 0;
assign detect_min[216][21] = (mid_1[1743:1736] < btm_1[1743:1736]) ? 1 : 0;
assign detect_min[216][22] = (mid_1[1743:1736] < btm_1[1751:1744]) ? 1 : 0;
assign detect_min[216][23] = (mid_1[1743:1736] < btm_2[1735:1728]) ? 1 : 0;
assign detect_min[216][24] = (mid_1[1743:1736] < btm_2[1743:1736]) ? 1 : 0;
assign detect_min[216][25] = (mid_1[1743:1736] < btm_2[1751:1744]) ? 1 : 0;

assign detect_min[217][0] = (mid_1[1751:1744] < top_0[1743:1736]) ? 1 : 0;
assign detect_min[217][1] = (mid_1[1751:1744] < top_0[1751:1744]) ? 1 : 0;
assign detect_min[217][2] = (mid_1[1751:1744] < top_0[1759:1752]) ? 1 : 0;
assign detect_min[217][3] = (mid_1[1751:1744] < top_1[1743:1736]) ? 1 : 0;
assign detect_min[217][4] = (mid_1[1751:1744] < top_1[1751:1744]) ? 1 : 0;
assign detect_min[217][5] = (mid_1[1751:1744] < top_1[1759:1752]) ? 1 : 0;
assign detect_min[217][6] = (mid_1[1751:1744] < top_2[1743:1736]) ? 1 : 0;
assign detect_min[217][7] = (mid_1[1751:1744] < top_2[1751:1744]) ? 1 : 0;
assign detect_min[217][8] = (mid_1[1751:1744] < top_2[1759:1752]) ? 1 : 0;
assign detect_min[217][9] = (mid_1[1751:1744] < mid_0[1743:1736]) ? 1 : 0;
assign detect_min[217][10] = (mid_1[1751:1744] < mid_0[1751:1744]) ? 1 : 0;
assign detect_min[217][11] = (mid_1[1751:1744] < mid_0[1759:1752]) ? 1 : 0;
assign detect_min[217][12] = (mid_1[1751:1744] < mid_1[1743:1736]) ? 1 : 0;
assign detect_min[217][13] = (mid_1[1751:1744] < mid_1[1759:1752]) ? 1 : 0;
assign detect_min[217][14] = (mid_1[1751:1744] < mid_2[1743:1736]) ? 1 : 0;
assign detect_min[217][15] = (mid_1[1751:1744] < mid_2[1751:1744]) ? 1 : 0;
assign detect_min[217][16] = (mid_1[1751:1744] < mid_2[1759:1752]) ? 1 : 0;
assign detect_min[217][17] = (mid_1[1751:1744] < btm_0[1743:1736]) ? 1 : 0;
assign detect_min[217][18] = (mid_1[1751:1744] < btm_0[1751:1744]) ? 1 : 0;
assign detect_min[217][19] = (mid_1[1751:1744] < btm_0[1759:1752]) ? 1 : 0;
assign detect_min[217][20] = (mid_1[1751:1744] < btm_1[1743:1736]) ? 1 : 0;
assign detect_min[217][21] = (mid_1[1751:1744] < btm_1[1751:1744]) ? 1 : 0;
assign detect_min[217][22] = (mid_1[1751:1744] < btm_1[1759:1752]) ? 1 : 0;
assign detect_min[217][23] = (mid_1[1751:1744] < btm_2[1743:1736]) ? 1 : 0;
assign detect_min[217][24] = (mid_1[1751:1744] < btm_2[1751:1744]) ? 1 : 0;
assign detect_min[217][25] = (mid_1[1751:1744] < btm_2[1759:1752]) ? 1 : 0;

assign detect_min[218][0] = (mid_1[1759:1752] < top_0[1751:1744]) ? 1 : 0;
assign detect_min[218][1] = (mid_1[1759:1752] < top_0[1759:1752]) ? 1 : 0;
assign detect_min[218][2] = (mid_1[1759:1752] < top_0[1767:1760]) ? 1 : 0;
assign detect_min[218][3] = (mid_1[1759:1752] < top_1[1751:1744]) ? 1 : 0;
assign detect_min[218][4] = (mid_1[1759:1752] < top_1[1759:1752]) ? 1 : 0;
assign detect_min[218][5] = (mid_1[1759:1752] < top_1[1767:1760]) ? 1 : 0;
assign detect_min[218][6] = (mid_1[1759:1752] < top_2[1751:1744]) ? 1 : 0;
assign detect_min[218][7] = (mid_1[1759:1752] < top_2[1759:1752]) ? 1 : 0;
assign detect_min[218][8] = (mid_1[1759:1752] < top_2[1767:1760]) ? 1 : 0;
assign detect_min[218][9] = (mid_1[1759:1752] < mid_0[1751:1744]) ? 1 : 0;
assign detect_min[218][10] = (mid_1[1759:1752] < mid_0[1759:1752]) ? 1 : 0;
assign detect_min[218][11] = (mid_1[1759:1752] < mid_0[1767:1760]) ? 1 : 0;
assign detect_min[218][12] = (mid_1[1759:1752] < mid_1[1751:1744]) ? 1 : 0;
assign detect_min[218][13] = (mid_1[1759:1752] < mid_1[1767:1760]) ? 1 : 0;
assign detect_min[218][14] = (mid_1[1759:1752] < mid_2[1751:1744]) ? 1 : 0;
assign detect_min[218][15] = (mid_1[1759:1752] < mid_2[1759:1752]) ? 1 : 0;
assign detect_min[218][16] = (mid_1[1759:1752] < mid_2[1767:1760]) ? 1 : 0;
assign detect_min[218][17] = (mid_1[1759:1752] < btm_0[1751:1744]) ? 1 : 0;
assign detect_min[218][18] = (mid_1[1759:1752] < btm_0[1759:1752]) ? 1 : 0;
assign detect_min[218][19] = (mid_1[1759:1752] < btm_0[1767:1760]) ? 1 : 0;
assign detect_min[218][20] = (mid_1[1759:1752] < btm_1[1751:1744]) ? 1 : 0;
assign detect_min[218][21] = (mid_1[1759:1752] < btm_1[1759:1752]) ? 1 : 0;
assign detect_min[218][22] = (mid_1[1759:1752] < btm_1[1767:1760]) ? 1 : 0;
assign detect_min[218][23] = (mid_1[1759:1752] < btm_2[1751:1744]) ? 1 : 0;
assign detect_min[218][24] = (mid_1[1759:1752] < btm_2[1759:1752]) ? 1 : 0;
assign detect_min[218][25] = (mid_1[1759:1752] < btm_2[1767:1760]) ? 1 : 0;

assign detect_min[219][0] = (mid_1[1767:1760] < top_0[1759:1752]) ? 1 : 0;
assign detect_min[219][1] = (mid_1[1767:1760] < top_0[1767:1760]) ? 1 : 0;
assign detect_min[219][2] = (mid_1[1767:1760] < top_0[1775:1768]) ? 1 : 0;
assign detect_min[219][3] = (mid_1[1767:1760] < top_1[1759:1752]) ? 1 : 0;
assign detect_min[219][4] = (mid_1[1767:1760] < top_1[1767:1760]) ? 1 : 0;
assign detect_min[219][5] = (mid_1[1767:1760] < top_1[1775:1768]) ? 1 : 0;
assign detect_min[219][6] = (mid_1[1767:1760] < top_2[1759:1752]) ? 1 : 0;
assign detect_min[219][7] = (mid_1[1767:1760] < top_2[1767:1760]) ? 1 : 0;
assign detect_min[219][8] = (mid_1[1767:1760] < top_2[1775:1768]) ? 1 : 0;
assign detect_min[219][9] = (mid_1[1767:1760] < mid_0[1759:1752]) ? 1 : 0;
assign detect_min[219][10] = (mid_1[1767:1760] < mid_0[1767:1760]) ? 1 : 0;
assign detect_min[219][11] = (mid_1[1767:1760] < mid_0[1775:1768]) ? 1 : 0;
assign detect_min[219][12] = (mid_1[1767:1760] < mid_1[1759:1752]) ? 1 : 0;
assign detect_min[219][13] = (mid_1[1767:1760] < mid_1[1775:1768]) ? 1 : 0;
assign detect_min[219][14] = (mid_1[1767:1760] < mid_2[1759:1752]) ? 1 : 0;
assign detect_min[219][15] = (mid_1[1767:1760] < mid_2[1767:1760]) ? 1 : 0;
assign detect_min[219][16] = (mid_1[1767:1760] < mid_2[1775:1768]) ? 1 : 0;
assign detect_min[219][17] = (mid_1[1767:1760] < btm_0[1759:1752]) ? 1 : 0;
assign detect_min[219][18] = (mid_1[1767:1760] < btm_0[1767:1760]) ? 1 : 0;
assign detect_min[219][19] = (mid_1[1767:1760] < btm_0[1775:1768]) ? 1 : 0;
assign detect_min[219][20] = (mid_1[1767:1760] < btm_1[1759:1752]) ? 1 : 0;
assign detect_min[219][21] = (mid_1[1767:1760] < btm_1[1767:1760]) ? 1 : 0;
assign detect_min[219][22] = (mid_1[1767:1760] < btm_1[1775:1768]) ? 1 : 0;
assign detect_min[219][23] = (mid_1[1767:1760] < btm_2[1759:1752]) ? 1 : 0;
assign detect_min[219][24] = (mid_1[1767:1760] < btm_2[1767:1760]) ? 1 : 0;
assign detect_min[219][25] = (mid_1[1767:1760] < btm_2[1775:1768]) ? 1 : 0;

assign detect_min[220][0] = (mid_1[1775:1768] < top_0[1767:1760]) ? 1 : 0;
assign detect_min[220][1] = (mid_1[1775:1768] < top_0[1775:1768]) ? 1 : 0;
assign detect_min[220][2] = (mid_1[1775:1768] < top_0[1783:1776]) ? 1 : 0;
assign detect_min[220][3] = (mid_1[1775:1768] < top_1[1767:1760]) ? 1 : 0;
assign detect_min[220][4] = (mid_1[1775:1768] < top_1[1775:1768]) ? 1 : 0;
assign detect_min[220][5] = (mid_1[1775:1768] < top_1[1783:1776]) ? 1 : 0;
assign detect_min[220][6] = (mid_1[1775:1768] < top_2[1767:1760]) ? 1 : 0;
assign detect_min[220][7] = (mid_1[1775:1768] < top_2[1775:1768]) ? 1 : 0;
assign detect_min[220][8] = (mid_1[1775:1768] < top_2[1783:1776]) ? 1 : 0;
assign detect_min[220][9] = (mid_1[1775:1768] < mid_0[1767:1760]) ? 1 : 0;
assign detect_min[220][10] = (mid_1[1775:1768] < mid_0[1775:1768]) ? 1 : 0;
assign detect_min[220][11] = (mid_1[1775:1768] < mid_0[1783:1776]) ? 1 : 0;
assign detect_min[220][12] = (mid_1[1775:1768] < mid_1[1767:1760]) ? 1 : 0;
assign detect_min[220][13] = (mid_1[1775:1768] < mid_1[1783:1776]) ? 1 : 0;
assign detect_min[220][14] = (mid_1[1775:1768] < mid_2[1767:1760]) ? 1 : 0;
assign detect_min[220][15] = (mid_1[1775:1768] < mid_2[1775:1768]) ? 1 : 0;
assign detect_min[220][16] = (mid_1[1775:1768] < mid_2[1783:1776]) ? 1 : 0;
assign detect_min[220][17] = (mid_1[1775:1768] < btm_0[1767:1760]) ? 1 : 0;
assign detect_min[220][18] = (mid_1[1775:1768] < btm_0[1775:1768]) ? 1 : 0;
assign detect_min[220][19] = (mid_1[1775:1768] < btm_0[1783:1776]) ? 1 : 0;
assign detect_min[220][20] = (mid_1[1775:1768] < btm_1[1767:1760]) ? 1 : 0;
assign detect_min[220][21] = (mid_1[1775:1768] < btm_1[1775:1768]) ? 1 : 0;
assign detect_min[220][22] = (mid_1[1775:1768] < btm_1[1783:1776]) ? 1 : 0;
assign detect_min[220][23] = (mid_1[1775:1768] < btm_2[1767:1760]) ? 1 : 0;
assign detect_min[220][24] = (mid_1[1775:1768] < btm_2[1775:1768]) ? 1 : 0;
assign detect_min[220][25] = (mid_1[1775:1768] < btm_2[1783:1776]) ? 1 : 0;

assign detect_min[221][0] = (mid_1[1783:1776] < top_0[1775:1768]) ? 1 : 0;
assign detect_min[221][1] = (mid_1[1783:1776] < top_0[1783:1776]) ? 1 : 0;
assign detect_min[221][2] = (mid_1[1783:1776] < top_0[1791:1784]) ? 1 : 0;
assign detect_min[221][3] = (mid_1[1783:1776] < top_1[1775:1768]) ? 1 : 0;
assign detect_min[221][4] = (mid_1[1783:1776] < top_1[1783:1776]) ? 1 : 0;
assign detect_min[221][5] = (mid_1[1783:1776] < top_1[1791:1784]) ? 1 : 0;
assign detect_min[221][6] = (mid_1[1783:1776] < top_2[1775:1768]) ? 1 : 0;
assign detect_min[221][7] = (mid_1[1783:1776] < top_2[1783:1776]) ? 1 : 0;
assign detect_min[221][8] = (mid_1[1783:1776] < top_2[1791:1784]) ? 1 : 0;
assign detect_min[221][9] = (mid_1[1783:1776] < mid_0[1775:1768]) ? 1 : 0;
assign detect_min[221][10] = (mid_1[1783:1776] < mid_0[1783:1776]) ? 1 : 0;
assign detect_min[221][11] = (mid_1[1783:1776] < mid_0[1791:1784]) ? 1 : 0;
assign detect_min[221][12] = (mid_1[1783:1776] < mid_1[1775:1768]) ? 1 : 0;
assign detect_min[221][13] = (mid_1[1783:1776] < mid_1[1791:1784]) ? 1 : 0;
assign detect_min[221][14] = (mid_1[1783:1776] < mid_2[1775:1768]) ? 1 : 0;
assign detect_min[221][15] = (mid_1[1783:1776] < mid_2[1783:1776]) ? 1 : 0;
assign detect_min[221][16] = (mid_1[1783:1776] < mid_2[1791:1784]) ? 1 : 0;
assign detect_min[221][17] = (mid_1[1783:1776] < btm_0[1775:1768]) ? 1 : 0;
assign detect_min[221][18] = (mid_1[1783:1776] < btm_0[1783:1776]) ? 1 : 0;
assign detect_min[221][19] = (mid_1[1783:1776] < btm_0[1791:1784]) ? 1 : 0;
assign detect_min[221][20] = (mid_1[1783:1776] < btm_1[1775:1768]) ? 1 : 0;
assign detect_min[221][21] = (mid_1[1783:1776] < btm_1[1783:1776]) ? 1 : 0;
assign detect_min[221][22] = (mid_1[1783:1776] < btm_1[1791:1784]) ? 1 : 0;
assign detect_min[221][23] = (mid_1[1783:1776] < btm_2[1775:1768]) ? 1 : 0;
assign detect_min[221][24] = (mid_1[1783:1776] < btm_2[1783:1776]) ? 1 : 0;
assign detect_min[221][25] = (mid_1[1783:1776] < btm_2[1791:1784]) ? 1 : 0;

assign detect_min[222][0] = (mid_1[1791:1784] < top_0[1783:1776]) ? 1 : 0;
assign detect_min[222][1] = (mid_1[1791:1784] < top_0[1791:1784]) ? 1 : 0;
assign detect_min[222][2] = (mid_1[1791:1784] < top_0[1799:1792]) ? 1 : 0;
assign detect_min[222][3] = (mid_1[1791:1784] < top_1[1783:1776]) ? 1 : 0;
assign detect_min[222][4] = (mid_1[1791:1784] < top_1[1791:1784]) ? 1 : 0;
assign detect_min[222][5] = (mid_1[1791:1784] < top_1[1799:1792]) ? 1 : 0;
assign detect_min[222][6] = (mid_1[1791:1784] < top_2[1783:1776]) ? 1 : 0;
assign detect_min[222][7] = (mid_1[1791:1784] < top_2[1791:1784]) ? 1 : 0;
assign detect_min[222][8] = (mid_1[1791:1784] < top_2[1799:1792]) ? 1 : 0;
assign detect_min[222][9] = (mid_1[1791:1784] < mid_0[1783:1776]) ? 1 : 0;
assign detect_min[222][10] = (mid_1[1791:1784] < mid_0[1791:1784]) ? 1 : 0;
assign detect_min[222][11] = (mid_1[1791:1784] < mid_0[1799:1792]) ? 1 : 0;
assign detect_min[222][12] = (mid_1[1791:1784] < mid_1[1783:1776]) ? 1 : 0;
assign detect_min[222][13] = (mid_1[1791:1784] < mid_1[1799:1792]) ? 1 : 0;
assign detect_min[222][14] = (mid_1[1791:1784] < mid_2[1783:1776]) ? 1 : 0;
assign detect_min[222][15] = (mid_1[1791:1784] < mid_2[1791:1784]) ? 1 : 0;
assign detect_min[222][16] = (mid_1[1791:1784] < mid_2[1799:1792]) ? 1 : 0;
assign detect_min[222][17] = (mid_1[1791:1784] < btm_0[1783:1776]) ? 1 : 0;
assign detect_min[222][18] = (mid_1[1791:1784] < btm_0[1791:1784]) ? 1 : 0;
assign detect_min[222][19] = (mid_1[1791:1784] < btm_0[1799:1792]) ? 1 : 0;
assign detect_min[222][20] = (mid_1[1791:1784] < btm_1[1783:1776]) ? 1 : 0;
assign detect_min[222][21] = (mid_1[1791:1784] < btm_1[1791:1784]) ? 1 : 0;
assign detect_min[222][22] = (mid_1[1791:1784] < btm_1[1799:1792]) ? 1 : 0;
assign detect_min[222][23] = (mid_1[1791:1784] < btm_2[1783:1776]) ? 1 : 0;
assign detect_min[222][24] = (mid_1[1791:1784] < btm_2[1791:1784]) ? 1 : 0;
assign detect_min[222][25] = (mid_1[1791:1784] < btm_2[1799:1792]) ? 1 : 0;

assign detect_min[223][0] = (mid_1[1799:1792] < top_0[1791:1784]) ? 1 : 0;
assign detect_min[223][1] = (mid_1[1799:1792] < top_0[1799:1792]) ? 1 : 0;
assign detect_min[223][2] = (mid_1[1799:1792] < top_0[1807:1800]) ? 1 : 0;
assign detect_min[223][3] = (mid_1[1799:1792] < top_1[1791:1784]) ? 1 : 0;
assign detect_min[223][4] = (mid_1[1799:1792] < top_1[1799:1792]) ? 1 : 0;
assign detect_min[223][5] = (mid_1[1799:1792] < top_1[1807:1800]) ? 1 : 0;
assign detect_min[223][6] = (mid_1[1799:1792] < top_2[1791:1784]) ? 1 : 0;
assign detect_min[223][7] = (mid_1[1799:1792] < top_2[1799:1792]) ? 1 : 0;
assign detect_min[223][8] = (mid_1[1799:1792] < top_2[1807:1800]) ? 1 : 0;
assign detect_min[223][9] = (mid_1[1799:1792] < mid_0[1791:1784]) ? 1 : 0;
assign detect_min[223][10] = (mid_1[1799:1792] < mid_0[1799:1792]) ? 1 : 0;
assign detect_min[223][11] = (mid_1[1799:1792] < mid_0[1807:1800]) ? 1 : 0;
assign detect_min[223][12] = (mid_1[1799:1792] < mid_1[1791:1784]) ? 1 : 0;
assign detect_min[223][13] = (mid_1[1799:1792] < mid_1[1807:1800]) ? 1 : 0;
assign detect_min[223][14] = (mid_1[1799:1792] < mid_2[1791:1784]) ? 1 : 0;
assign detect_min[223][15] = (mid_1[1799:1792] < mid_2[1799:1792]) ? 1 : 0;
assign detect_min[223][16] = (mid_1[1799:1792] < mid_2[1807:1800]) ? 1 : 0;
assign detect_min[223][17] = (mid_1[1799:1792] < btm_0[1791:1784]) ? 1 : 0;
assign detect_min[223][18] = (mid_1[1799:1792] < btm_0[1799:1792]) ? 1 : 0;
assign detect_min[223][19] = (mid_1[1799:1792] < btm_0[1807:1800]) ? 1 : 0;
assign detect_min[223][20] = (mid_1[1799:1792] < btm_1[1791:1784]) ? 1 : 0;
assign detect_min[223][21] = (mid_1[1799:1792] < btm_1[1799:1792]) ? 1 : 0;
assign detect_min[223][22] = (mid_1[1799:1792] < btm_1[1807:1800]) ? 1 : 0;
assign detect_min[223][23] = (mid_1[1799:1792] < btm_2[1791:1784]) ? 1 : 0;
assign detect_min[223][24] = (mid_1[1799:1792] < btm_2[1799:1792]) ? 1 : 0;
assign detect_min[223][25] = (mid_1[1799:1792] < btm_2[1807:1800]) ? 1 : 0;

assign detect_min[224][0] = (mid_1[1807:1800] < top_0[1799:1792]) ? 1 : 0;
assign detect_min[224][1] = (mid_1[1807:1800] < top_0[1807:1800]) ? 1 : 0;
assign detect_min[224][2] = (mid_1[1807:1800] < top_0[1815:1808]) ? 1 : 0;
assign detect_min[224][3] = (mid_1[1807:1800] < top_1[1799:1792]) ? 1 : 0;
assign detect_min[224][4] = (mid_1[1807:1800] < top_1[1807:1800]) ? 1 : 0;
assign detect_min[224][5] = (mid_1[1807:1800] < top_1[1815:1808]) ? 1 : 0;
assign detect_min[224][6] = (mid_1[1807:1800] < top_2[1799:1792]) ? 1 : 0;
assign detect_min[224][7] = (mid_1[1807:1800] < top_2[1807:1800]) ? 1 : 0;
assign detect_min[224][8] = (mid_1[1807:1800] < top_2[1815:1808]) ? 1 : 0;
assign detect_min[224][9] = (mid_1[1807:1800] < mid_0[1799:1792]) ? 1 : 0;
assign detect_min[224][10] = (mid_1[1807:1800] < mid_0[1807:1800]) ? 1 : 0;
assign detect_min[224][11] = (mid_1[1807:1800] < mid_0[1815:1808]) ? 1 : 0;
assign detect_min[224][12] = (mid_1[1807:1800] < mid_1[1799:1792]) ? 1 : 0;
assign detect_min[224][13] = (mid_1[1807:1800] < mid_1[1815:1808]) ? 1 : 0;
assign detect_min[224][14] = (mid_1[1807:1800] < mid_2[1799:1792]) ? 1 : 0;
assign detect_min[224][15] = (mid_1[1807:1800] < mid_2[1807:1800]) ? 1 : 0;
assign detect_min[224][16] = (mid_1[1807:1800] < mid_2[1815:1808]) ? 1 : 0;
assign detect_min[224][17] = (mid_1[1807:1800] < btm_0[1799:1792]) ? 1 : 0;
assign detect_min[224][18] = (mid_1[1807:1800] < btm_0[1807:1800]) ? 1 : 0;
assign detect_min[224][19] = (mid_1[1807:1800] < btm_0[1815:1808]) ? 1 : 0;
assign detect_min[224][20] = (mid_1[1807:1800] < btm_1[1799:1792]) ? 1 : 0;
assign detect_min[224][21] = (mid_1[1807:1800] < btm_1[1807:1800]) ? 1 : 0;
assign detect_min[224][22] = (mid_1[1807:1800] < btm_1[1815:1808]) ? 1 : 0;
assign detect_min[224][23] = (mid_1[1807:1800] < btm_2[1799:1792]) ? 1 : 0;
assign detect_min[224][24] = (mid_1[1807:1800] < btm_2[1807:1800]) ? 1 : 0;
assign detect_min[224][25] = (mid_1[1807:1800] < btm_2[1815:1808]) ? 1 : 0;

assign detect_min[225][0] = (mid_1[1815:1808] < top_0[1807:1800]) ? 1 : 0;
assign detect_min[225][1] = (mid_1[1815:1808] < top_0[1815:1808]) ? 1 : 0;
assign detect_min[225][2] = (mid_1[1815:1808] < top_0[1823:1816]) ? 1 : 0;
assign detect_min[225][3] = (mid_1[1815:1808] < top_1[1807:1800]) ? 1 : 0;
assign detect_min[225][4] = (mid_1[1815:1808] < top_1[1815:1808]) ? 1 : 0;
assign detect_min[225][5] = (mid_1[1815:1808] < top_1[1823:1816]) ? 1 : 0;
assign detect_min[225][6] = (mid_1[1815:1808] < top_2[1807:1800]) ? 1 : 0;
assign detect_min[225][7] = (mid_1[1815:1808] < top_2[1815:1808]) ? 1 : 0;
assign detect_min[225][8] = (mid_1[1815:1808] < top_2[1823:1816]) ? 1 : 0;
assign detect_min[225][9] = (mid_1[1815:1808] < mid_0[1807:1800]) ? 1 : 0;
assign detect_min[225][10] = (mid_1[1815:1808] < mid_0[1815:1808]) ? 1 : 0;
assign detect_min[225][11] = (mid_1[1815:1808] < mid_0[1823:1816]) ? 1 : 0;
assign detect_min[225][12] = (mid_1[1815:1808] < mid_1[1807:1800]) ? 1 : 0;
assign detect_min[225][13] = (mid_1[1815:1808] < mid_1[1823:1816]) ? 1 : 0;
assign detect_min[225][14] = (mid_1[1815:1808] < mid_2[1807:1800]) ? 1 : 0;
assign detect_min[225][15] = (mid_1[1815:1808] < mid_2[1815:1808]) ? 1 : 0;
assign detect_min[225][16] = (mid_1[1815:1808] < mid_2[1823:1816]) ? 1 : 0;
assign detect_min[225][17] = (mid_1[1815:1808] < btm_0[1807:1800]) ? 1 : 0;
assign detect_min[225][18] = (mid_1[1815:1808] < btm_0[1815:1808]) ? 1 : 0;
assign detect_min[225][19] = (mid_1[1815:1808] < btm_0[1823:1816]) ? 1 : 0;
assign detect_min[225][20] = (mid_1[1815:1808] < btm_1[1807:1800]) ? 1 : 0;
assign detect_min[225][21] = (mid_1[1815:1808] < btm_1[1815:1808]) ? 1 : 0;
assign detect_min[225][22] = (mid_1[1815:1808] < btm_1[1823:1816]) ? 1 : 0;
assign detect_min[225][23] = (mid_1[1815:1808] < btm_2[1807:1800]) ? 1 : 0;
assign detect_min[225][24] = (mid_1[1815:1808] < btm_2[1815:1808]) ? 1 : 0;
assign detect_min[225][25] = (mid_1[1815:1808] < btm_2[1823:1816]) ? 1 : 0;

assign detect_min[226][0] = (mid_1[1823:1816] < top_0[1815:1808]) ? 1 : 0;
assign detect_min[226][1] = (mid_1[1823:1816] < top_0[1823:1816]) ? 1 : 0;
assign detect_min[226][2] = (mid_1[1823:1816] < top_0[1831:1824]) ? 1 : 0;
assign detect_min[226][3] = (mid_1[1823:1816] < top_1[1815:1808]) ? 1 : 0;
assign detect_min[226][4] = (mid_1[1823:1816] < top_1[1823:1816]) ? 1 : 0;
assign detect_min[226][5] = (mid_1[1823:1816] < top_1[1831:1824]) ? 1 : 0;
assign detect_min[226][6] = (mid_1[1823:1816] < top_2[1815:1808]) ? 1 : 0;
assign detect_min[226][7] = (mid_1[1823:1816] < top_2[1823:1816]) ? 1 : 0;
assign detect_min[226][8] = (mid_1[1823:1816] < top_2[1831:1824]) ? 1 : 0;
assign detect_min[226][9] = (mid_1[1823:1816] < mid_0[1815:1808]) ? 1 : 0;
assign detect_min[226][10] = (mid_1[1823:1816] < mid_0[1823:1816]) ? 1 : 0;
assign detect_min[226][11] = (mid_1[1823:1816] < mid_0[1831:1824]) ? 1 : 0;
assign detect_min[226][12] = (mid_1[1823:1816] < mid_1[1815:1808]) ? 1 : 0;
assign detect_min[226][13] = (mid_1[1823:1816] < mid_1[1831:1824]) ? 1 : 0;
assign detect_min[226][14] = (mid_1[1823:1816] < mid_2[1815:1808]) ? 1 : 0;
assign detect_min[226][15] = (mid_1[1823:1816] < mid_2[1823:1816]) ? 1 : 0;
assign detect_min[226][16] = (mid_1[1823:1816] < mid_2[1831:1824]) ? 1 : 0;
assign detect_min[226][17] = (mid_1[1823:1816] < btm_0[1815:1808]) ? 1 : 0;
assign detect_min[226][18] = (mid_1[1823:1816] < btm_0[1823:1816]) ? 1 : 0;
assign detect_min[226][19] = (mid_1[1823:1816] < btm_0[1831:1824]) ? 1 : 0;
assign detect_min[226][20] = (mid_1[1823:1816] < btm_1[1815:1808]) ? 1 : 0;
assign detect_min[226][21] = (mid_1[1823:1816] < btm_1[1823:1816]) ? 1 : 0;
assign detect_min[226][22] = (mid_1[1823:1816] < btm_1[1831:1824]) ? 1 : 0;
assign detect_min[226][23] = (mid_1[1823:1816] < btm_2[1815:1808]) ? 1 : 0;
assign detect_min[226][24] = (mid_1[1823:1816] < btm_2[1823:1816]) ? 1 : 0;
assign detect_min[226][25] = (mid_1[1823:1816] < btm_2[1831:1824]) ? 1 : 0;

assign detect_min[227][0] = (mid_1[1831:1824] < top_0[1823:1816]) ? 1 : 0;
assign detect_min[227][1] = (mid_1[1831:1824] < top_0[1831:1824]) ? 1 : 0;
assign detect_min[227][2] = (mid_1[1831:1824] < top_0[1839:1832]) ? 1 : 0;
assign detect_min[227][3] = (mid_1[1831:1824] < top_1[1823:1816]) ? 1 : 0;
assign detect_min[227][4] = (mid_1[1831:1824] < top_1[1831:1824]) ? 1 : 0;
assign detect_min[227][5] = (mid_1[1831:1824] < top_1[1839:1832]) ? 1 : 0;
assign detect_min[227][6] = (mid_1[1831:1824] < top_2[1823:1816]) ? 1 : 0;
assign detect_min[227][7] = (mid_1[1831:1824] < top_2[1831:1824]) ? 1 : 0;
assign detect_min[227][8] = (mid_1[1831:1824] < top_2[1839:1832]) ? 1 : 0;
assign detect_min[227][9] = (mid_1[1831:1824] < mid_0[1823:1816]) ? 1 : 0;
assign detect_min[227][10] = (mid_1[1831:1824] < mid_0[1831:1824]) ? 1 : 0;
assign detect_min[227][11] = (mid_1[1831:1824] < mid_0[1839:1832]) ? 1 : 0;
assign detect_min[227][12] = (mid_1[1831:1824] < mid_1[1823:1816]) ? 1 : 0;
assign detect_min[227][13] = (mid_1[1831:1824] < mid_1[1839:1832]) ? 1 : 0;
assign detect_min[227][14] = (mid_1[1831:1824] < mid_2[1823:1816]) ? 1 : 0;
assign detect_min[227][15] = (mid_1[1831:1824] < mid_2[1831:1824]) ? 1 : 0;
assign detect_min[227][16] = (mid_1[1831:1824] < mid_2[1839:1832]) ? 1 : 0;
assign detect_min[227][17] = (mid_1[1831:1824] < btm_0[1823:1816]) ? 1 : 0;
assign detect_min[227][18] = (mid_1[1831:1824] < btm_0[1831:1824]) ? 1 : 0;
assign detect_min[227][19] = (mid_1[1831:1824] < btm_0[1839:1832]) ? 1 : 0;
assign detect_min[227][20] = (mid_1[1831:1824] < btm_1[1823:1816]) ? 1 : 0;
assign detect_min[227][21] = (mid_1[1831:1824] < btm_1[1831:1824]) ? 1 : 0;
assign detect_min[227][22] = (mid_1[1831:1824] < btm_1[1839:1832]) ? 1 : 0;
assign detect_min[227][23] = (mid_1[1831:1824] < btm_2[1823:1816]) ? 1 : 0;
assign detect_min[227][24] = (mid_1[1831:1824] < btm_2[1831:1824]) ? 1 : 0;
assign detect_min[227][25] = (mid_1[1831:1824] < btm_2[1839:1832]) ? 1 : 0;

assign detect_min[228][0] = (mid_1[1839:1832] < top_0[1831:1824]) ? 1 : 0;
assign detect_min[228][1] = (mid_1[1839:1832] < top_0[1839:1832]) ? 1 : 0;
assign detect_min[228][2] = (mid_1[1839:1832] < top_0[1847:1840]) ? 1 : 0;
assign detect_min[228][3] = (mid_1[1839:1832] < top_1[1831:1824]) ? 1 : 0;
assign detect_min[228][4] = (mid_1[1839:1832] < top_1[1839:1832]) ? 1 : 0;
assign detect_min[228][5] = (mid_1[1839:1832] < top_1[1847:1840]) ? 1 : 0;
assign detect_min[228][6] = (mid_1[1839:1832] < top_2[1831:1824]) ? 1 : 0;
assign detect_min[228][7] = (mid_1[1839:1832] < top_2[1839:1832]) ? 1 : 0;
assign detect_min[228][8] = (mid_1[1839:1832] < top_2[1847:1840]) ? 1 : 0;
assign detect_min[228][9] = (mid_1[1839:1832] < mid_0[1831:1824]) ? 1 : 0;
assign detect_min[228][10] = (mid_1[1839:1832] < mid_0[1839:1832]) ? 1 : 0;
assign detect_min[228][11] = (mid_1[1839:1832] < mid_0[1847:1840]) ? 1 : 0;
assign detect_min[228][12] = (mid_1[1839:1832] < mid_1[1831:1824]) ? 1 : 0;
assign detect_min[228][13] = (mid_1[1839:1832] < mid_1[1847:1840]) ? 1 : 0;
assign detect_min[228][14] = (mid_1[1839:1832] < mid_2[1831:1824]) ? 1 : 0;
assign detect_min[228][15] = (mid_1[1839:1832] < mid_2[1839:1832]) ? 1 : 0;
assign detect_min[228][16] = (mid_1[1839:1832] < mid_2[1847:1840]) ? 1 : 0;
assign detect_min[228][17] = (mid_1[1839:1832] < btm_0[1831:1824]) ? 1 : 0;
assign detect_min[228][18] = (mid_1[1839:1832] < btm_0[1839:1832]) ? 1 : 0;
assign detect_min[228][19] = (mid_1[1839:1832] < btm_0[1847:1840]) ? 1 : 0;
assign detect_min[228][20] = (mid_1[1839:1832] < btm_1[1831:1824]) ? 1 : 0;
assign detect_min[228][21] = (mid_1[1839:1832] < btm_1[1839:1832]) ? 1 : 0;
assign detect_min[228][22] = (mid_1[1839:1832] < btm_1[1847:1840]) ? 1 : 0;
assign detect_min[228][23] = (mid_1[1839:1832] < btm_2[1831:1824]) ? 1 : 0;
assign detect_min[228][24] = (mid_1[1839:1832] < btm_2[1839:1832]) ? 1 : 0;
assign detect_min[228][25] = (mid_1[1839:1832] < btm_2[1847:1840]) ? 1 : 0;

assign detect_min[229][0] = (mid_1[1847:1840] < top_0[1839:1832]) ? 1 : 0;
assign detect_min[229][1] = (mid_1[1847:1840] < top_0[1847:1840]) ? 1 : 0;
assign detect_min[229][2] = (mid_1[1847:1840] < top_0[1855:1848]) ? 1 : 0;
assign detect_min[229][3] = (mid_1[1847:1840] < top_1[1839:1832]) ? 1 : 0;
assign detect_min[229][4] = (mid_1[1847:1840] < top_1[1847:1840]) ? 1 : 0;
assign detect_min[229][5] = (mid_1[1847:1840] < top_1[1855:1848]) ? 1 : 0;
assign detect_min[229][6] = (mid_1[1847:1840] < top_2[1839:1832]) ? 1 : 0;
assign detect_min[229][7] = (mid_1[1847:1840] < top_2[1847:1840]) ? 1 : 0;
assign detect_min[229][8] = (mid_1[1847:1840] < top_2[1855:1848]) ? 1 : 0;
assign detect_min[229][9] = (mid_1[1847:1840] < mid_0[1839:1832]) ? 1 : 0;
assign detect_min[229][10] = (mid_1[1847:1840] < mid_0[1847:1840]) ? 1 : 0;
assign detect_min[229][11] = (mid_1[1847:1840] < mid_0[1855:1848]) ? 1 : 0;
assign detect_min[229][12] = (mid_1[1847:1840] < mid_1[1839:1832]) ? 1 : 0;
assign detect_min[229][13] = (mid_1[1847:1840] < mid_1[1855:1848]) ? 1 : 0;
assign detect_min[229][14] = (mid_1[1847:1840] < mid_2[1839:1832]) ? 1 : 0;
assign detect_min[229][15] = (mid_1[1847:1840] < mid_2[1847:1840]) ? 1 : 0;
assign detect_min[229][16] = (mid_1[1847:1840] < mid_2[1855:1848]) ? 1 : 0;
assign detect_min[229][17] = (mid_1[1847:1840] < btm_0[1839:1832]) ? 1 : 0;
assign detect_min[229][18] = (mid_1[1847:1840] < btm_0[1847:1840]) ? 1 : 0;
assign detect_min[229][19] = (mid_1[1847:1840] < btm_0[1855:1848]) ? 1 : 0;
assign detect_min[229][20] = (mid_1[1847:1840] < btm_1[1839:1832]) ? 1 : 0;
assign detect_min[229][21] = (mid_1[1847:1840] < btm_1[1847:1840]) ? 1 : 0;
assign detect_min[229][22] = (mid_1[1847:1840] < btm_1[1855:1848]) ? 1 : 0;
assign detect_min[229][23] = (mid_1[1847:1840] < btm_2[1839:1832]) ? 1 : 0;
assign detect_min[229][24] = (mid_1[1847:1840] < btm_2[1847:1840]) ? 1 : 0;
assign detect_min[229][25] = (mid_1[1847:1840] < btm_2[1855:1848]) ? 1 : 0;

assign detect_min[230][0] = (mid_1[1855:1848] < top_0[1847:1840]) ? 1 : 0;
assign detect_min[230][1] = (mid_1[1855:1848] < top_0[1855:1848]) ? 1 : 0;
assign detect_min[230][2] = (mid_1[1855:1848] < top_0[1863:1856]) ? 1 : 0;
assign detect_min[230][3] = (mid_1[1855:1848] < top_1[1847:1840]) ? 1 : 0;
assign detect_min[230][4] = (mid_1[1855:1848] < top_1[1855:1848]) ? 1 : 0;
assign detect_min[230][5] = (mid_1[1855:1848] < top_1[1863:1856]) ? 1 : 0;
assign detect_min[230][6] = (mid_1[1855:1848] < top_2[1847:1840]) ? 1 : 0;
assign detect_min[230][7] = (mid_1[1855:1848] < top_2[1855:1848]) ? 1 : 0;
assign detect_min[230][8] = (mid_1[1855:1848] < top_2[1863:1856]) ? 1 : 0;
assign detect_min[230][9] = (mid_1[1855:1848] < mid_0[1847:1840]) ? 1 : 0;
assign detect_min[230][10] = (mid_1[1855:1848] < mid_0[1855:1848]) ? 1 : 0;
assign detect_min[230][11] = (mid_1[1855:1848] < mid_0[1863:1856]) ? 1 : 0;
assign detect_min[230][12] = (mid_1[1855:1848] < mid_1[1847:1840]) ? 1 : 0;
assign detect_min[230][13] = (mid_1[1855:1848] < mid_1[1863:1856]) ? 1 : 0;
assign detect_min[230][14] = (mid_1[1855:1848] < mid_2[1847:1840]) ? 1 : 0;
assign detect_min[230][15] = (mid_1[1855:1848] < mid_2[1855:1848]) ? 1 : 0;
assign detect_min[230][16] = (mid_1[1855:1848] < mid_2[1863:1856]) ? 1 : 0;
assign detect_min[230][17] = (mid_1[1855:1848] < btm_0[1847:1840]) ? 1 : 0;
assign detect_min[230][18] = (mid_1[1855:1848] < btm_0[1855:1848]) ? 1 : 0;
assign detect_min[230][19] = (mid_1[1855:1848] < btm_0[1863:1856]) ? 1 : 0;
assign detect_min[230][20] = (mid_1[1855:1848] < btm_1[1847:1840]) ? 1 : 0;
assign detect_min[230][21] = (mid_1[1855:1848] < btm_1[1855:1848]) ? 1 : 0;
assign detect_min[230][22] = (mid_1[1855:1848] < btm_1[1863:1856]) ? 1 : 0;
assign detect_min[230][23] = (mid_1[1855:1848] < btm_2[1847:1840]) ? 1 : 0;
assign detect_min[230][24] = (mid_1[1855:1848] < btm_2[1855:1848]) ? 1 : 0;
assign detect_min[230][25] = (mid_1[1855:1848] < btm_2[1863:1856]) ? 1 : 0;

assign detect_min[231][0] = (mid_1[1863:1856] < top_0[1855:1848]) ? 1 : 0;
assign detect_min[231][1] = (mid_1[1863:1856] < top_0[1863:1856]) ? 1 : 0;
assign detect_min[231][2] = (mid_1[1863:1856] < top_0[1871:1864]) ? 1 : 0;
assign detect_min[231][3] = (mid_1[1863:1856] < top_1[1855:1848]) ? 1 : 0;
assign detect_min[231][4] = (mid_1[1863:1856] < top_1[1863:1856]) ? 1 : 0;
assign detect_min[231][5] = (mid_1[1863:1856] < top_1[1871:1864]) ? 1 : 0;
assign detect_min[231][6] = (mid_1[1863:1856] < top_2[1855:1848]) ? 1 : 0;
assign detect_min[231][7] = (mid_1[1863:1856] < top_2[1863:1856]) ? 1 : 0;
assign detect_min[231][8] = (mid_1[1863:1856] < top_2[1871:1864]) ? 1 : 0;
assign detect_min[231][9] = (mid_1[1863:1856] < mid_0[1855:1848]) ? 1 : 0;
assign detect_min[231][10] = (mid_1[1863:1856] < mid_0[1863:1856]) ? 1 : 0;
assign detect_min[231][11] = (mid_1[1863:1856] < mid_0[1871:1864]) ? 1 : 0;
assign detect_min[231][12] = (mid_1[1863:1856] < mid_1[1855:1848]) ? 1 : 0;
assign detect_min[231][13] = (mid_1[1863:1856] < mid_1[1871:1864]) ? 1 : 0;
assign detect_min[231][14] = (mid_1[1863:1856] < mid_2[1855:1848]) ? 1 : 0;
assign detect_min[231][15] = (mid_1[1863:1856] < mid_2[1863:1856]) ? 1 : 0;
assign detect_min[231][16] = (mid_1[1863:1856] < mid_2[1871:1864]) ? 1 : 0;
assign detect_min[231][17] = (mid_1[1863:1856] < btm_0[1855:1848]) ? 1 : 0;
assign detect_min[231][18] = (mid_1[1863:1856] < btm_0[1863:1856]) ? 1 : 0;
assign detect_min[231][19] = (mid_1[1863:1856] < btm_0[1871:1864]) ? 1 : 0;
assign detect_min[231][20] = (mid_1[1863:1856] < btm_1[1855:1848]) ? 1 : 0;
assign detect_min[231][21] = (mid_1[1863:1856] < btm_1[1863:1856]) ? 1 : 0;
assign detect_min[231][22] = (mid_1[1863:1856] < btm_1[1871:1864]) ? 1 : 0;
assign detect_min[231][23] = (mid_1[1863:1856] < btm_2[1855:1848]) ? 1 : 0;
assign detect_min[231][24] = (mid_1[1863:1856] < btm_2[1863:1856]) ? 1 : 0;
assign detect_min[231][25] = (mid_1[1863:1856] < btm_2[1871:1864]) ? 1 : 0;

assign detect_min[232][0] = (mid_1[1871:1864] < top_0[1863:1856]) ? 1 : 0;
assign detect_min[232][1] = (mid_1[1871:1864] < top_0[1871:1864]) ? 1 : 0;
assign detect_min[232][2] = (mid_1[1871:1864] < top_0[1879:1872]) ? 1 : 0;
assign detect_min[232][3] = (mid_1[1871:1864] < top_1[1863:1856]) ? 1 : 0;
assign detect_min[232][4] = (mid_1[1871:1864] < top_1[1871:1864]) ? 1 : 0;
assign detect_min[232][5] = (mid_1[1871:1864] < top_1[1879:1872]) ? 1 : 0;
assign detect_min[232][6] = (mid_1[1871:1864] < top_2[1863:1856]) ? 1 : 0;
assign detect_min[232][7] = (mid_1[1871:1864] < top_2[1871:1864]) ? 1 : 0;
assign detect_min[232][8] = (mid_1[1871:1864] < top_2[1879:1872]) ? 1 : 0;
assign detect_min[232][9] = (mid_1[1871:1864] < mid_0[1863:1856]) ? 1 : 0;
assign detect_min[232][10] = (mid_1[1871:1864] < mid_0[1871:1864]) ? 1 : 0;
assign detect_min[232][11] = (mid_1[1871:1864] < mid_0[1879:1872]) ? 1 : 0;
assign detect_min[232][12] = (mid_1[1871:1864] < mid_1[1863:1856]) ? 1 : 0;
assign detect_min[232][13] = (mid_1[1871:1864] < mid_1[1879:1872]) ? 1 : 0;
assign detect_min[232][14] = (mid_1[1871:1864] < mid_2[1863:1856]) ? 1 : 0;
assign detect_min[232][15] = (mid_1[1871:1864] < mid_2[1871:1864]) ? 1 : 0;
assign detect_min[232][16] = (mid_1[1871:1864] < mid_2[1879:1872]) ? 1 : 0;
assign detect_min[232][17] = (mid_1[1871:1864] < btm_0[1863:1856]) ? 1 : 0;
assign detect_min[232][18] = (mid_1[1871:1864] < btm_0[1871:1864]) ? 1 : 0;
assign detect_min[232][19] = (mid_1[1871:1864] < btm_0[1879:1872]) ? 1 : 0;
assign detect_min[232][20] = (mid_1[1871:1864] < btm_1[1863:1856]) ? 1 : 0;
assign detect_min[232][21] = (mid_1[1871:1864] < btm_1[1871:1864]) ? 1 : 0;
assign detect_min[232][22] = (mid_1[1871:1864] < btm_1[1879:1872]) ? 1 : 0;
assign detect_min[232][23] = (mid_1[1871:1864] < btm_2[1863:1856]) ? 1 : 0;
assign detect_min[232][24] = (mid_1[1871:1864] < btm_2[1871:1864]) ? 1 : 0;
assign detect_min[232][25] = (mid_1[1871:1864] < btm_2[1879:1872]) ? 1 : 0;

assign detect_min[233][0] = (mid_1[1879:1872] < top_0[1871:1864]) ? 1 : 0;
assign detect_min[233][1] = (mid_1[1879:1872] < top_0[1879:1872]) ? 1 : 0;
assign detect_min[233][2] = (mid_1[1879:1872] < top_0[1887:1880]) ? 1 : 0;
assign detect_min[233][3] = (mid_1[1879:1872] < top_1[1871:1864]) ? 1 : 0;
assign detect_min[233][4] = (mid_1[1879:1872] < top_1[1879:1872]) ? 1 : 0;
assign detect_min[233][5] = (mid_1[1879:1872] < top_1[1887:1880]) ? 1 : 0;
assign detect_min[233][6] = (mid_1[1879:1872] < top_2[1871:1864]) ? 1 : 0;
assign detect_min[233][7] = (mid_1[1879:1872] < top_2[1879:1872]) ? 1 : 0;
assign detect_min[233][8] = (mid_1[1879:1872] < top_2[1887:1880]) ? 1 : 0;
assign detect_min[233][9] = (mid_1[1879:1872] < mid_0[1871:1864]) ? 1 : 0;
assign detect_min[233][10] = (mid_1[1879:1872] < mid_0[1879:1872]) ? 1 : 0;
assign detect_min[233][11] = (mid_1[1879:1872] < mid_0[1887:1880]) ? 1 : 0;
assign detect_min[233][12] = (mid_1[1879:1872] < mid_1[1871:1864]) ? 1 : 0;
assign detect_min[233][13] = (mid_1[1879:1872] < mid_1[1887:1880]) ? 1 : 0;
assign detect_min[233][14] = (mid_1[1879:1872] < mid_2[1871:1864]) ? 1 : 0;
assign detect_min[233][15] = (mid_1[1879:1872] < mid_2[1879:1872]) ? 1 : 0;
assign detect_min[233][16] = (mid_1[1879:1872] < mid_2[1887:1880]) ? 1 : 0;
assign detect_min[233][17] = (mid_1[1879:1872] < btm_0[1871:1864]) ? 1 : 0;
assign detect_min[233][18] = (mid_1[1879:1872] < btm_0[1879:1872]) ? 1 : 0;
assign detect_min[233][19] = (mid_1[1879:1872] < btm_0[1887:1880]) ? 1 : 0;
assign detect_min[233][20] = (mid_1[1879:1872] < btm_1[1871:1864]) ? 1 : 0;
assign detect_min[233][21] = (mid_1[1879:1872] < btm_1[1879:1872]) ? 1 : 0;
assign detect_min[233][22] = (mid_1[1879:1872] < btm_1[1887:1880]) ? 1 : 0;
assign detect_min[233][23] = (mid_1[1879:1872] < btm_2[1871:1864]) ? 1 : 0;
assign detect_min[233][24] = (mid_1[1879:1872] < btm_2[1879:1872]) ? 1 : 0;
assign detect_min[233][25] = (mid_1[1879:1872] < btm_2[1887:1880]) ? 1 : 0;

assign detect_min[234][0] = (mid_1[1887:1880] < top_0[1879:1872]) ? 1 : 0;
assign detect_min[234][1] = (mid_1[1887:1880] < top_0[1887:1880]) ? 1 : 0;
assign detect_min[234][2] = (mid_1[1887:1880] < top_0[1895:1888]) ? 1 : 0;
assign detect_min[234][3] = (mid_1[1887:1880] < top_1[1879:1872]) ? 1 : 0;
assign detect_min[234][4] = (mid_1[1887:1880] < top_1[1887:1880]) ? 1 : 0;
assign detect_min[234][5] = (mid_1[1887:1880] < top_1[1895:1888]) ? 1 : 0;
assign detect_min[234][6] = (mid_1[1887:1880] < top_2[1879:1872]) ? 1 : 0;
assign detect_min[234][7] = (mid_1[1887:1880] < top_2[1887:1880]) ? 1 : 0;
assign detect_min[234][8] = (mid_1[1887:1880] < top_2[1895:1888]) ? 1 : 0;
assign detect_min[234][9] = (mid_1[1887:1880] < mid_0[1879:1872]) ? 1 : 0;
assign detect_min[234][10] = (mid_1[1887:1880] < mid_0[1887:1880]) ? 1 : 0;
assign detect_min[234][11] = (mid_1[1887:1880] < mid_0[1895:1888]) ? 1 : 0;
assign detect_min[234][12] = (mid_1[1887:1880] < mid_1[1879:1872]) ? 1 : 0;
assign detect_min[234][13] = (mid_1[1887:1880] < mid_1[1895:1888]) ? 1 : 0;
assign detect_min[234][14] = (mid_1[1887:1880] < mid_2[1879:1872]) ? 1 : 0;
assign detect_min[234][15] = (mid_1[1887:1880] < mid_2[1887:1880]) ? 1 : 0;
assign detect_min[234][16] = (mid_1[1887:1880] < mid_2[1895:1888]) ? 1 : 0;
assign detect_min[234][17] = (mid_1[1887:1880] < btm_0[1879:1872]) ? 1 : 0;
assign detect_min[234][18] = (mid_1[1887:1880] < btm_0[1887:1880]) ? 1 : 0;
assign detect_min[234][19] = (mid_1[1887:1880] < btm_0[1895:1888]) ? 1 : 0;
assign detect_min[234][20] = (mid_1[1887:1880] < btm_1[1879:1872]) ? 1 : 0;
assign detect_min[234][21] = (mid_1[1887:1880] < btm_1[1887:1880]) ? 1 : 0;
assign detect_min[234][22] = (mid_1[1887:1880] < btm_1[1895:1888]) ? 1 : 0;
assign detect_min[234][23] = (mid_1[1887:1880] < btm_2[1879:1872]) ? 1 : 0;
assign detect_min[234][24] = (mid_1[1887:1880] < btm_2[1887:1880]) ? 1 : 0;
assign detect_min[234][25] = (mid_1[1887:1880] < btm_2[1895:1888]) ? 1 : 0;

assign detect_min[235][0] = (mid_1[1895:1888] < top_0[1887:1880]) ? 1 : 0;
assign detect_min[235][1] = (mid_1[1895:1888] < top_0[1895:1888]) ? 1 : 0;
assign detect_min[235][2] = (mid_1[1895:1888] < top_0[1903:1896]) ? 1 : 0;
assign detect_min[235][3] = (mid_1[1895:1888] < top_1[1887:1880]) ? 1 : 0;
assign detect_min[235][4] = (mid_1[1895:1888] < top_1[1895:1888]) ? 1 : 0;
assign detect_min[235][5] = (mid_1[1895:1888] < top_1[1903:1896]) ? 1 : 0;
assign detect_min[235][6] = (mid_1[1895:1888] < top_2[1887:1880]) ? 1 : 0;
assign detect_min[235][7] = (mid_1[1895:1888] < top_2[1895:1888]) ? 1 : 0;
assign detect_min[235][8] = (mid_1[1895:1888] < top_2[1903:1896]) ? 1 : 0;
assign detect_min[235][9] = (mid_1[1895:1888] < mid_0[1887:1880]) ? 1 : 0;
assign detect_min[235][10] = (mid_1[1895:1888] < mid_0[1895:1888]) ? 1 : 0;
assign detect_min[235][11] = (mid_1[1895:1888] < mid_0[1903:1896]) ? 1 : 0;
assign detect_min[235][12] = (mid_1[1895:1888] < mid_1[1887:1880]) ? 1 : 0;
assign detect_min[235][13] = (mid_1[1895:1888] < mid_1[1903:1896]) ? 1 : 0;
assign detect_min[235][14] = (mid_1[1895:1888] < mid_2[1887:1880]) ? 1 : 0;
assign detect_min[235][15] = (mid_1[1895:1888] < mid_2[1895:1888]) ? 1 : 0;
assign detect_min[235][16] = (mid_1[1895:1888] < mid_2[1903:1896]) ? 1 : 0;
assign detect_min[235][17] = (mid_1[1895:1888] < btm_0[1887:1880]) ? 1 : 0;
assign detect_min[235][18] = (mid_1[1895:1888] < btm_0[1895:1888]) ? 1 : 0;
assign detect_min[235][19] = (mid_1[1895:1888] < btm_0[1903:1896]) ? 1 : 0;
assign detect_min[235][20] = (mid_1[1895:1888] < btm_1[1887:1880]) ? 1 : 0;
assign detect_min[235][21] = (mid_1[1895:1888] < btm_1[1895:1888]) ? 1 : 0;
assign detect_min[235][22] = (mid_1[1895:1888] < btm_1[1903:1896]) ? 1 : 0;
assign detect_min[235][23] = (mid_1[1895:1888] < btm_2[1887:1880]) ? 1 : 0;
assign detect_min[235][24] = (mid_1[1895:1888] < btm_2[1895:1888]) ? 1 : 0;
assign detect_min[235][25] = (mid_1[1895:1888] < btm_2[1903:1896]) ? 1 : 0;

assign detect_min[236][0] = (mid_1[1903:1896] < top_0[1895:1888]) ? 1 : 0;
assign detect_min[236][1] = (mid_1[1903:1896] < top_0[1903:1896]) ? 1 : 0;
assign detect_min[236][2] = (mid_1[1903:1896] < top_0[1911:1904]) ? 1 : 0;
assign detect_min[236][3] = (mid_1[1903:1896] < top_1[1895:1888]) ? 1 : 0;
assign detect_min[236][4] = (mid_1[1903:1896] < top_1[1903:1896]) ? 1 : 0;
assign detect_min[236][5] = (mid_1[1903:1896] < top_1[1911:1904]) ? 1 : 0;
assign detect_min[236][6] = (mid_1[1903:1896] < top_2[1895:1888]) ? 1 : 0;
assign detect_min[236][7] = (mid_1[1903:1896] < top_2[1903:1896]) ? 1 : 0;
assign detect_min[236][8] = (mid_1[1903:1896] < top_2[1911:1904]) ? 1 : 0;
assign detect_min[236][9] = (mid_1[1903:1896] < mid_0[1895:1888]) ? 1 : 0;
assign detect_min[236][10] = (mid_1[1903:1896] < mid_0[1903:1896]) ? 1 : 0;
assign detect_min[236][11] = (mid_1[1903:1896] < mid_0[1911:1904]) ? 1 : 0;
assign detect_min[236][12] = (mid_1[1903:1896] < mid_1[1895:1888]) ? 1 : 0;
assign detect_min[236][13] = (mid_1[1903:1896] < mid_1[1911:1904]) ? 1 : 0;
assign detect_min[236][14] = (mid_1[1903:1896] < mid_2[1895:1888]) ? 1 : 0;
assign detect_min[236][15] = (mid_1[1903:1896] < mid_2[1903:1896]) ? 1 : 0;
assign detect_min[236][16] = (mid_1[1903:1896] < mid_2[1911:1904]) ? 1 : 0;
assign detect_min[236][17] = (mid_1[1903:1896] < btm_0[1895:1888]) ? 1 : 0;
assign detect_min[236][18] = (mid_1[1903:1896] < btm_0[1903:1896]) ? 1 : 0;
assign detect_min[236][19] = (mid_1[1903:1896] < btm_0[1911:1904]) ? 1 : 0;
assign detect_min[236][20] = (mid_1[1903:1896] < btm_1[1895:1888]) ? 1 : 0;
assign detect_min[236][21] = (mid_1[1903:1896] < btm_1[1903:1896]) ? 1 : 0;
assign detect_min[236][22] = (mid_1[1903:1896] < btm_1[1911:1904]) ? 1 : 0;
assign detect_min[236][23] = (mid_1[1903:1896] < btm_2[1895:1888]) ? 1 : 0;
assign detect_min[236][24] = (mid_1[1903:1896] < btm_2[1903:1896]) ? 1 : 0;
assign detect_min[236][25] = (mid_1[1903:1896] < btm_2[1911:1904]) ? 1 : 0;

assign detect_min[237][0] = (mid_1[1911:1904] < top_0[1903:1896]) ? 1 : 0;
assign detect_min[237][1] = (mid_1[1911:1904] < top_0[1911:1904]) ? 1 : 0;
assign detect_min[237][2] = (mid_1[1911:1904] < top_0[1919:1912]) ? 1 : 0;
assign detect_min[237][3] = (mid_1[1911:1904] < top_1[1903:1896]) ? 1 : 0;
assign detect_min[237][4] = (mid_1[1911:1904] < top_1[1911:1904]) ? 1 : 0;
assign detect_min[237][5] = (mid_1[1911:1904] < top_1[1919:1912]) ? 1 : 0;
assign detect_min[237][6] = (mid_1[1911:1904] < top_2[1903:1896]) ? 1 : 0;
assign detect_min[237][7] = (mid_1[1911:1904] < top_2[1911:1904]) ? 1 : 0;
assign detect_min[237][8] = (mid_1[1911:1904] < top_2[1919:1912]) ? 1 : 0;
assign detect_min[237][9] = (mid_1[1911:1904] < mid_0[1903:1896]) ? 1 : 0;
assign detect_min[237][10] = (mid_1[1911:1904] < mid_0[1911:1904]) ? 1 : 0;
assign detect_min[237][11] = (mid_1[1911:1904] < mid_0[1919:1912]) ? 1 : 0;
assign detect_min[237][12] = (mid_1[1911:1904] < mid_1[1903:1896]) ? 1 : 0;
assign detect_min[237][13] = (mid_1[1911:1904] < mid_1[1919:1912]) ? 1 : 0;
assign detect_min[237][14] = (mid_1[1911:1904] < mid_2[1903:1896]) ? 1 : 0;
assign detect_min[237][15] = (mid_1[1911:1904] < mid_2[1911:1904]) ? 1 : 0;
assign detect_min[237][16] = (mid_1[1911:1904] < mid_2[1919:1912]) ? 1 : 0;
assign detect_min[237][17] = (mid_1[1911:1904] < btm_0[1903:1896]) ? 1 : 0;
assign detect_min[237][18] = (mid_1[1911:1904] < btm_0[1911:1904]) ? 1 : 0;
assign detect_min[237][19] = (mid_1[1911:1904] < btm_0[1919:1912]) ? 1 : 0;
assign detect_min[237][20] = (mid_1[1911:1904] < btm_1[1903:1896]) ? 1 : 0;
assign detect_min[237][21] = (mid_1[1911:1904] < btm_1[1911:1904]) ? 1 : 0;
assign detect_min[237][22] = (mid_1[1911:1904] < btm_1[1919:1912]) ? 1 : 0;
assign detect_min[237][23] = (mid_1[1911:1904] < btm_2[1903:1896]) ? 1 : 0;
assign detect_min[237][24] = (mid_1[1911:1904] < btm_2[1911:1904]) ? 1 : 0;
assign detect_min[237][25] = (mid_1[1911:1904] < btm_2[1919:1912]) ? 1 : 0;

assign detect_min[238][0] = (mid_1[1919:1912] < top_0[1911:1904]) ? 1 : 0;
assign detect_min[238][1] = (mid_1[1919:1912] < top_0[1919:1912]) ? 1 : 0;
assign detect_min[238][2] = (mid_1[1919:1912] < top_0[1927:1920]) ? 1 : 0;
assign detect_min[238][3] = (mid_1[1919:1912] < top_1[1911:1904]) ? 1 : 0;
assign detect_min[238][4] = (mid_1[1919:1912] < top_1[1919:1912]) ? 1 : 0;
assign detect_min[238][5] = (mid_1[1919:1912] < top_1[1927:1920]) ? 1 : 0;
assign detect_min[238][6] = (mid_1[1919:1912] < top_2[1911:1904]) ? 1 : 0;
assign detect_min[238][7] = (mid_1[1919:1912] < top_2[1919:1912]) ? 1 : 0;
assign detect_min[238][8] = (mid_1[1919:1912] < top_2[1927:1920]) ? 1 : 0;
assign detect_min[238][9] = (mid_1[1919:1912] < mid_0[1911:1904]) ? 1 : 0;
assign detect_min[238][10] = (mid_1[1919:1912] < mid_0[1919:1912]) ? 1 : 0;
assign detect_min[238][11] = (mid_1[1919:1912] < mid_0[1927:1920]) ? 1 : 0;
assign detect_min[238][12] = (mid_1[1919:1912] < mid_1[1911:1904]) ? 1 : 0;
assign detect_min[238][13] = (mid_1[1919:1912] < mid_1[1927:1920]) ? 1 : 0;
assign detect_min[238][14] = (mid_1[1919:1912] < mid_2[1911:1904]) ? 1 : 0;
assign detect_min[238][15] = (mid_1[1919:1912] < mid_2[1919:1912]) ? 1 : 0;
assign detect_min[238][16] = (mid_1[1919:1912] < mid_2[1927:1920]) ? 1 : 0;
assign detect_min[238][17] = (mid_1[1919:1912] < btm_0[1911:1904]) ? 1 : 0;
assign detect_min[238][18] = (mid_1[1919:1912] < btm_0[1919:1912]) ? 1 : 0;
assign detect_min[238][19] = (mid_1[1919:1912] < btm_0[1927:1920]) ? 1 : 0;
assign detect_min[238][20] = (mid_1[1919:1912] < btm_1[1911:1904]) ? 1 : 0;
assign detect_min[238][21] = (mid_1[1919:1912] < btm_1[1919:1912]) ? 1 : 0;
assign detect_min[238][22] = (mid_1[1919:1912] < btm_1[1927:1920]) ? 1 : 0;
assign detect_min[238][23] = (mid_1[1919:1912] < btm_2[1911:1904]) ? 1 : 0;
assign detect_min[238][24] = (mid_1[1919:1912] < btm_2[1919:1912]) ? 1 : 0;
assign detect_min[238][25] = (mid_1[1919:1912] < btm_2[1927:1920]) ? 1 : 0;

assign detect_min[239][0] = (mid_1[1927:1920] < top_0[1919:1912]) ? 1 : 0;
assign detect_min[239][1] = (mid_1[1927:1920] < top_0[1927:1920]) ? 1 : 0;
assign detect_min[239][2] = (mid_1[1927:1920] < top_0[1935:1928]) ? 1 : 0;
assign detect_min[239][3] = (mid_1[1927:1920] < top_1[1919:1912]) ? 1 : 0;
assign detect_min[239][4] = (mid_1[1927:1920] < top_1[1927:1920]) ? 1 : 0;
assign detect_min[239][5] = (mid_1[1927:1920] < top_1[1935:1928]) ? 1 : 0;
assign detect_min[239][6] = (mid_1[1927:1920] < top_2[1919:1912]) ? 1 : 0;
assign detect_min[239][7] = (mid_1[1927:1920] < top_2[1927:1920]) ? 1 : 0;
assign detect_min[239][8] = (mid_1[1927:1920] < top_2[1935:1928]) ? 1 : 0;
assign detect_min[239][9] = (mid_1[1927:1920] < mid_0[1919:1912]) ? 1 : 0;
assign detect_min[239][10] = (mid_1[1927:1920] < mid_0[1927:1920]) ? 1 : 0;
assign detect_min[239][11] = (mid_1[1927:1920] < mid_0[1935:1928]) ? 1 : 0;
assign detect_min[239][12] = (mid_1[1927:1920] < mid_1[1919:1912]) ? 1 : 0;
assign detect_min[239][13] = (mid_1[1927:1920] < mid_1[1935:1928]) ? 1 : 0;
assign detect_min[239][14] = (mid_1[1927:1920] < mid_2[1919:1912]) ? 1 : 0;
assign detect_min[239][15] = (mid_1[1927:1920] < mid_2[1927:1920]) ? 1 : 0;
assign detect_min[239][16] = (mid_1[1927:1920] < mid_2[1935:1928]) ? 1 : 0;
assign detect_min[239][17] = (mid_1[1927:1920] < btm_0[1919:1912]) ? 1 : 0;
assign detect_min[239][18] = (mid_1[1927:1920] < btm_0[1927:1920]) ? 1 : 0;
assign detect_min[239][19] = (mid_1[1927:1920] < btm_0[1935:1928]) ? 1 : 0;
assign detect_min[239][20] = (mid_1[1927:1920] < btm_1[1919:1912]) ? 1 : 0;
assign detect_min[239][21] = (mid_1[1927:1920] < btm_1[1927:1920]) ? 1 : 0;
assign detect_min[239][22] = (mid_1[1927:1920] < btm_1[1935:1928]) ? 1 : 0;
assign detect_min[239][23] = (mid_1[1927:1920] < btm_2[1919:1912]) ? 1 : 0;
assign detect_min[239][24] = (mid_1[1927:1920] < btm_2[1927:1920]) ? 1 : 0;
assign detect_min[239][25] = (mid_1[1927:1920] < btm_2[1935:1928]) ? 1 : 0;

assign detect_min[240][0] = (mid_1[1935:1928] < top_0[1927:1920]) ? 1 : 0;
assign detect_min[240][1] = (mid_1[1935:1928] < top_0[1935:1928]) ? 1 : 0;
assign detect_min[240][2] = (mid_1[1935:1928] < top_0[1943:1936]) ? 1 : 0;
assign detect_min[240][3] = (mid_1[1935:1928] < top_1[1927:1920]) ? 1 : 0;
assign detect_min[240][4] = (mid_1[1935:1928] < top_1[1935:1928]) ? 1 : 0;
assign detect_min[240][5] = (mid_1[1935:1928] < top_1[1943:1936]) ? 1 : 0;
assign detect_min[240][6] = (mid_1[1935:1928] < top_2[1927:1920]) ? 1 : 0;
assign detect_min[240][7] = (mid_1[1935:1928] < top_2[1935:1928]) ? 1 : 0;
assign detect_min[240][8] = (mid_1[1935:1928] < top_2[1943:1936]) ? 1 : 0;
assign detect_min[240][9] = (mid_1[1935:1928] < mid_0[1927:1920]) ? 1 : 0;
assign detect_min[240][10] = (mid_1[1935:1928] < mid_0[1935:1928]) ? 1 : 0;
assign detect_min[240][11] = (mid_1[1935:1928] < mid_0[1943:1936]) ? 1 : 0;
assign detect_min[240][12] = (mid_1[1935:1928] < mid_1[1927:1920]) ? 1 : 0;
assign detect_min[240][13] = (mid_1[1935:1928] < mid_1[1943:1936]) ? 1 : 0;
assign detect_min[240][14] = (mid_1[1935:1928] < mid_2[1927:1920]) ? 1 : 0;
assign detect_min[240][15] = (mid_1[1935:1928] < mid_2[1935:1928]) ? 1 : 0;
assign detect_min[240][16] = (mid_1[1935:1928] < mid_2[1943:1936]) ? 1 : 0;
assign detect_min[240][17] = (mid_1[1935:1928] < btm_0[1927:1920]) ? 1 : 0;
assign detect_min[240][18] = (mid_1[1935:1928] < btm_0[1935:1928]) ? 1 : 0;
assign detect_min[240][19] = (mid_1[1935:1928] < btm_0[1943:1936]) ? 1 : 0;
assign detect_min[240][20] = (mid_1[1935:1928] < btm_1[1927:1920]) ? 1 : 0;
assign detect_min[240][21] = (mid_1[1935:1928] < btm_1[1935:1928]) ? 1 : 0;
assign detect_min[240][22] = (mid_1[1935:1928] < btm_1[1943:1936]) ? 1 : 0;
assign detect_min[240][23] = (mid_1[1935:1928] < btm_2[1927:1920]) ? 1 : 0;
assign detect_min[240][24] = (mid_1[1935:1928] < btm_2[1935:1928]) ? 1 : 0;
assign detect_min[240][25] = (mid_1[1935:1928] < btm_2[1943:1936]) ? 1 : 0;

assign detect_min[241][0] = (mid_1[1943:1936] < top_0[1935:1928]) ? 1 : 0;
assign detect_min[241][1] = (mid_1[1943:1936] < top_0[1943:1936]) ? 1 : 0;
assign detect_min[241][2] = (mid_1[1943:1936] < top_0[1951:1944]) ? 1 : 0;
assign detect_min[241][3] = (mid_1[1943:1936] < top_1[1935:1928]) ? 1 : 0;
assign detect_min[241][4] = (mid_1[1943:1936] < top_1[1943:1936]) ? 1 : 0;
assign detect_min[241][5] = (mid_1[1943:1936] < top_1[1951:1944]) ? 1 : 0;
assign detect_min[241][6] = (mid_1[1943:1936] < top_2[1935:1928]) ? 1 : 0;
assign detect_min[241][7] = (mid_1[1943:1936] < top_2[1943:1936]) ? 1 : 0;
assign detect_min[241][8] = (mid_1[1943:1936] < top_2[1951:1944]) ? 1 : 0;
assign detect_min[241][9] = (mid_1[1943:1936] < mid_0[1935:1928]) ? 1 : 0;
assign detect_min[241][10] = (mid_1[1943:1936] < mid_0[1943:1936]) ? 1 : 0;
assign detect_min[241][11] = (mid_1[1943:1936] < mid_0[1951:1944]) ? 1 : 0;
assign detect_min[241][12] = (mid_1[1943:1936] < mid_1[1935:1928]) ? 1 : 0;
assign detect_min[241][13] = (mid_1[1943:1936] < mid_1[1951:1944]) ? 1 : 0;
assign detect_min[241][14] = (mid_1[1943:1936] < mid_2[1935:1928]) ? 1 : 0;
assign detect_min[241][15] = (mid_1[1943:1936] < mid_2[1943:1936]) ? 1 : 0;
assign detect_min[241][16] = (mid_1[1943:1936] < mid_2[1951:1944]) ? 1 : 0;
assign detect_min[241][17] = (mid_1[1943:1936] < btm_0[1935:1928]) ? 1 : 0;
assign detect_min[241][18] = (mid_1[1943:1936] < btm_0[1943:1936]) ? 1 : 0;
assign detect_min[241][19] = (mid_1[1943:1936] < btm_0[1951:1944]) ? 1 : 0;
assign detect_min[241][20] = (mid_1[1943:1936] < btm_1[1935:1928]) ? 1 : 0;
assign detect_min[241][21] = (mid_1[1943:1936] < btm_1[1943:1936]) ? 1 : 0;
assign detect_min[241][22] = (mid_1[1943:1936] < btm_1[1951:1944]) ? 1 : 0;
assign detect_min[241][23] = (mid_1[1943:1936] < btm_2[1935:1928]) ? 1 : 0;
assign detect_min[241][24] = (mid_1[1943:1936] < btm_2[1943:1936]) ? 1 : 0;
assign detect_min[241][25] = (mid_1[1943:1936] < btm_2[1951:1944]) ? 1 : 0;

assign detect_min[242][0] = (mid_1[1951:1944] < top_0[1943:1936]) ? 1 : 0;
assign detect_min[242][1] = (mid_1[1951:1944] < top_0[1951:1944]) ? 1 : 0;
assign detect_min[242][2] = (mid_1[1951:1944] < top_0[1959:1952]) ? 1 : 0;
assign detect_min[242][3] = (mid_1[1951:1944] < top_1[1943:1936]) ? 1 : 0;
assign detect_min[242][4] = (mid_1[1951:1944] < top_1[1951:1944]) ? 1 : 0;
assign detect_min[242][5] = (mid_1[1951:1944] < top_1[1959:1952]) ? 1 : 0;
assign detect_min[242][6] = (mid_1[1951:1944] < top_2[1943:1936]) ? 1 : 0;
assign detect_min[242][7] = (mid_1[1951:1944] < top_2[1951:1944]) ? 1 : 0;
assign detect_min[242][8] = (mid_1[1951:1944] < top_2[1959:1952]) ? 1 : 0;
assign detect_min[242][9] = (mid_1[1951:1944] < mid_0[1943:1936]) ? 1 : 0;
assign detect_min[242][10] = (mid_1[1951:1944] < mid_0[1951:1944]) ? 1 : 0;
assign detect_min[242][11] = (mid_1[1951:1944] < mid_0[1959:1952]) ? 1 : 0;
assign detect_min[242][12] = (mid_1[1951:1944] < mid_1[1943:1936]) ? 1 : 0;
assign detect_min[242][13] = (mid_1[1951:1944] < mid_1[1959:1952]) ? 1 : 0;
assign detect_min[242][14] = (mid_1[1951:1944] < mid_2[1943:1936]) ? 1 : 0;
assign detect_min[242][15] = (mid_1[1951:1944] < mid_2[1951:1944]) ? 1 : 0;
assign detect_min[242][16] = (mid_1[1951:1944] < mid_2[1959:1952]) ? 1 : 0;
assign detect_min[242][17] = (mid_1[1951:1944] < btm_0[1943:1936]) ? 1 : 0;
assign detect_min[242][18] = (mid_1[1951:1944] < btm_0[1951:1944]) ? 1 : 0;
assign detect_min[242][19] = (mid_1[1951:1944] < btm_0[1959:1952]) ? 1 : 0;
assign detect_min[242][20] = (mid_1[1951:1944] < btm_1[1943:1936]) ? 1 : 0;
assign detect_min[242][21] = (mid_1[1951:1944] < btm_1[1951:1944]) ? 1 : 0;
assign detect_min[242][22] = (mid_1[1951:1944] < btm_1[1959:1952]) ? 1 : 0;
assign detect_min[242][23] = (mid_1[1951:1944] < btm_2[1943:1936]) ? 1 : 0;
assign detect_min[242][24] = (mid_1[1951:1944] < btm_2[1951:1944]) ? 1 : 0;
assign detect_min[242][25] = (mid_1[1951:1944] < btm_2[1959:1952]) ? 1 : 0;

assign detect_min[243][0] = (mid_1[1959:1952] < top_0[1951:1944]) ? 1 : 0;
assign detect_min[243][1] = (mid_1[1959:1952] < top_0[1959:1952]) ? 1 : 0;
assign detect_min[243][2] = (mid_1[1959:1952] < top_0[1967:1960]) ? 1 : 0;
assign detect_min[243][3] = (mid_1[1959:1952] < top_1[1951:1944]) ? 1 : 0;
assign detect_min[243][4] = (mid_1[1959:1952] < top_1[1959:1952]) ? 1 : 0;
assign detect_min[243][5] = (mid_1[1959:1952] < top_1[1967:1960]) ? 1 : 0;
assign detect_min[243][6] = (mid_1[1959:1952] < top_2[1951:1944]) ? 1 : 0;
assign detect_min[243][7] = (mid_1[1959:1952] < top_2[1959:1952]) ? 1 : 0;
assign detect_min[243][8] = (mid_1[1959:1952] < top_2[1967:1960]) ? 1 : 0;
assign detect_min[243][9] = (mid_1[1959:1952] < mid_0[1951:1944]) ? 1 : 0;
assign detect_min[243][10] = (mid_1[1959:1952] < mid_0[1959:1952]) ? 1 : 0;
assign detect_min[243][11] = (mid_1[1959:1952] < mid_0[1967:1960]) ? 1 : 0;
assign detect_min[243][12] = (mid_1[1959:1952] < mid_1[1951:1944]) ? 1 : 0;
assign detect_min[243][13] = (mid_1[1959:1952] < mid_1[1967:1960]) ? 1 : 0;
assign detect_min[243][14] = (mid_1[1959:1952] < mid_2[1951:1944]) ? 1 : 0;
assign detect_min[243][15] = (mid_1[1959:1952] < mid_2[1959:1952]) ? 1 : 0;
assign detect_min[243][16] = (mid_1[1959:1952] < mid_2[1967:1960]) ? 1 : 0;
assign detect_min[243][17] = (mid_1[1959:1952] < btm_0[1951:1944]) ? 1 : 0;
assign detect_min[243][18] = (mid_1[1959:1952] < btm_0[1959:1952]) ? 1 : 0;
assign detect_min[243][19] = (mid_1[1959:1952] < btm_0[1967:1960]) ? 1 : 0;
assign detect_min[243][20] = (mid_1[1959:1952] < btm_1[1951:1944]) ? 1 : 0;
assign detect_min[243][21] = (mid_1[1959:1952] < btm_1[1959:1952]) ? 1 : 0;
assign detect_min[243][22] = (mid_1[1959:1952] < btm_1[1967:1960]) ? 1 : 0;
assign detect_min[243][23] = (mid_1[1959:1952] < btm_2[1951:1944]) ? 1 : 0;
assign detect_min[243][24] = (mid_1[1959:1952] < btm_2[1959:1952]) ? 1 : 0;
assign detect_min[243][25] = (mid_1[1959:1952] < btm_2[1967:1960]) ? 1 : 0;

assign detect_min[244][0] = (mid_1[1967:1960] < top_0[1959:1952]) ? 1 : 0;
assign detect_min[244][1] = (mid_1[1967:1960] < top_0[1967:1960]) ? 1 : 0;
assign detect_min[244][2] = (mid_1[1967:1960] < top_0[1975:1968]) ? 1 : 0;
assign detect_min[244][3] = (mid_1[1967:1960] < top_1[1959:1952]) ? 1 : 0;
assign detect_min[244][4] = (mid_1[1967:1960] < top_1[1967:1960]) ? 1 : 0;
assign detect_min[244][5] = (mid_1[1967:1960] < top_1[1975:1968]) ? 1 : 0;
assign detect_min[244][6] = (mid_1[1967:1960] < top_2[1959:1952]) ? 1 : 0;
assign detect_min[244][7] = (mid_1[1967:1960] < top_2[1967:1960]) ? 1 : 0;
assign detect_min[244][8] = (mid_1[1967:1960] < top_2[1975:1968]) ? 1 : 0;
assign detect_min[244][9] = (mid_1[1967:1960] < mid_0[1959:1952]) ? 1 : 0;
assign detect_min[244][10] = (mid_1[1967:1960] < mid_0[1967:1960]) ? 1 : 0;
assign detect_min[244][11] = (mid_1[1967:1960] < mid_0[1975:1968]) ? 1 : 0;
assign detect_min[244][12] = (mid_1[1967:1960] < mid_1[1959:1952]) ? 1 : 0;
assign detect_min[244][13] = (mid_1[1967:1960] < mid_1[1975:1968]) ? 1 : 0;
assign detect_min[244][14] = (mid_1[1967:1960] < mid_2[1959:1952]) ? 1 : 0;
assign detect_min[244][15] = (mid_1[1967:1960] < mid_2[1967:1960]) ? 1 : 0;
assign detect_min[244][16] = (mid_1[1967:1960] < mid_2[1975:1968]) ? 1 : 0;
assign detect_min[244][17] = (mid_1[1967:1960] < btm_0[1959:1952]) ? 1 : 0;
assign detect_min[244][18] = (mid_1[1967:1960] < btm_0[1967:1960]) ? 1 : 0;
assign detect_min[244][19] = (mid_1[1967:1960] < btm_0[1975:1968]) ? 1 : 0;
assign detect_min[244][20] = (mid_1[1967:1960] < btm_1[1959:1952]) ? 1 : 0;
assign detect_min[244][21] = (mid_1[1967:1960] < btm_1[1967:1960]) ? 1 : 0;
assign detect_min[244][22] = (mid_1[1967:1960] < btm_1[1975:1968]) ? 1 : 0;
assign detect_min[244][23] = (mid_1[1967:1960] < btm_2[1959:1952]) ? 1 : 0;
assign detect_min[244][24] = (mid_1[1967:1960] < btm_2[1967:1960]) ? 1 : 0;
assign detect_min[244][25] = (mid_1[1967:1960] < btm_2[1975:1968]) ? 1 : 0;

assign detect_min[245][0] = (mid_1[1975:1968] < top_0[1967:1960]) ? 1 : 0;
assign detect_min[245][1] = (mid_1[1975:1968] < top_0[1975:1968]) ? 1 : 0;
assign detect_min[245][2] = (mid_1[1975:1968] < top_0[1983:1976]) ? 1 : 0;
assign detect_min[245][3] = (mid_1[1975:1968] < top_1[1967:1960]) ? 1 : 0;
assign detect_min[245][4] = (mid_1[1975:1968] < top_1[1975:1968]) ? 1 : 0;
assign detect_min[245][5] = (mid_1[1975:1968] < top_1[1983:1976]) ? 1 : 0;
assign detect_min[245][6] = (mid_1[1975:1968] < top_2[1967:1960]) ? 1 : 0;
assign detect_min[245][7] = (mid_1[1975:1968] < top_2[1975:1968]) ? 1 : 0;
assign detect_min[245][8] = (mid_1[1975:1968] < top_2[1983:1976]) ? 1 : 0;
assign detect_min[245][9] = (mid_1[1975:1968] < mid_0[1967:1960]) ? 1 : 0;
assign detect_min[245][10] = (mid_1[1975:1968] < mid_0[1975:1968]) ? 1 : 0;
assign detect_min[245][11] = (mid_1[1975:1968] < mid_0[1983:1976]) ? 1 : 0;
assign detect_min[245][12] = (mid_1[1975:1968] < mid_1[1967:1960]) ? 1 : 0;
assign detect_min[245][13] = (mid_1[1975:1968] < mid_1[1983:1976]) ? 1 : 0;
assign detect_min[245][14] = (mid_1[1975:1968] < mid_2[1967:1960]) ? 1 : 0;
assign detect_min[245][15] = (mid_1[1975:1968] < mid_2[1975:1968]) ? 1 : 0;
assign detect_min[245][16] = (mid_1[1975:1968] < mid_2[1983:1976]) ? 1 : 0;
assign detect_min[245][17] = (mid_1[1975:1968] < btm_0[1967:1960]) ? 1 : 0;
assign detect_min[245][18] = (mid_1[1975:1968] < btm_0[1975:1968]) ? 1 : 0;
assign detect_min[245][19] = (mid_1[1975:1968] < btm_0[1983:1976]) ? 1 : 0;
assign detect_min[245][20] = (mid_1[1975:1968] < btm_1[1967:1960]) ? 1 : 0;
assign detect_min[245][21] = (mid_1[1975:1968] < btm_1[1975:1968]) ? 1 : 0;
assign detect_min[245][22] = (mid_1[1975:1968] < btm_1[1983:1976]) ? 1 : 0;
assign detect_min[245][23] = (mid_1[1975:1968] < btm_2[1967:1960]) ? 1 : 0;
assign detect_min[245][24] = (mid_1[1975:1968] < btm_2[1975:1968]) ? 1 : 0;
assign detect_min[245][25] = (mid_1[1975:1968] < btm_2[1983:1976]) ? 1 : 0;

assign detect_min[246][0] = (mid_1[1983:1976] < top_0[1975:1968]) ? 1 : 0;
assign detect_min[246][1] = (mid_1[1983:1976] < top_0[1983:1976]) ? 1 : 0;
assign detect_min[246][2] = (mid_1[1983:1976] < top_0[1991:1984]) ? 1 : 0;
assign detect_min[246][3] = (mid_1[1983:1976] < top_1[1975:1968]) ? 1 : 0;
assign detect_min[246][4] = (mid_1[1983:1976] < top_1[1983:1976]) ? 1 : 0;
assign detect_min[246][5] = (mid_1[1983:1976] < top_1[1991:1984]) ? 1 : 0;
assign detect_min[246][6] = (mid_1[1983:1976] < top_2[1975:1968]) ? 1 : 0;
assign detect_min[246][7] = (mid_1[1983:1976] < top_2[1983:1976]) ? 1 : 0;
assign detect_min[246][8] = (mid_1[1983:1976] < top_2[1991:1984]) ? 1 : 0;
assign detect_min[246][9] = (mid_1[1983:1976] < mid_0[1975:1968]) ? 1 : 0;
assign detect_min[246][10] = (mid_1[1983:1976] < mid_0[1983:1976]) ? 1 : 0;
assign detect_min[246][11] = (mid_1[1983:1976] < mid_0[1991:1984]) ? 1 : 0;
assign detect_min[246][12] = (mid_1[1983:1976] < mid_1[1975:1968]) ? 1 : 0;
assign detect_min[246][13] = (mid_1[1983:1976] < mid_1[1991:1984]) ? 1 : 0;
assign detect_min[246][14] = (mid_1[1983:1976] < mid_2[1975:1968]) ? 1 : 0;
assign detect_min[246][15] = (mid_1[1983:1976] < mid_2[1983:1976]) ? 1 : 0;
assign detect_min[246][16] = (mid_1[1983:1976] < mid_2[1991:1984]) ? 1 : 0;
assign detect_min[246][17] = (mid_1[1983:1976] < btm_0[1975:1968]) ? 1 : 0;
assign detect_min[246][18] = (mid_1[1983:1976] < btm_0[1983:1976]) ? 1 : 0;
assign detect_min[246][19] = (mid_1[1983:1976] < btm_0[1991:1984]) ? 1 : 0;
assign detect_min[246][20] = (mid_1[1983:1976] < btm_1[1975:1968]) ? 1 : 0;
assign detect_min[246][21] = (mid_1[1983:1976] < btm_1[1983:1976]) ? 1 : 0;
assign detect_min[246][22] = (mid_1[1983:1976] < btm_1[1991:1984]) ? 1 : 0;
assign detect_min[246][23] = (mid_1[1983:1976] < btm_2[1975:1968]) ? 1 : 0;
assign detect_min[246][24] = (mid_1[1983:1976] < btm_2[1983:1976]) ? 1 : 0;
assign detect_min[246][25] = (mid_1[1983:1976] < btm_2[1991:1984]) ? 1 : 0;

assign detect_min[247][0] = (mid_1[1991:1984] < top_0[1983:1976]) ? 1 : 0;
assign detect_min[247][1] = (mid_1[1991:1984] < top_0[1991:1984]) ? 1 : 0;
assign detect_min[247][2] = (mid_1[1991:1984] < top_0[1999:1992]) ? 1 : 0;
assign detect_min[247][3] = (mid_1[1991:1984] < top_1[1983:1976]) ? 1 : 0;
assign detect_min[247][4] = (mid_1[1991:1984] < top_1[1991:1984]) ? 1 : 0;
assign detect_min[247][5] = (mid_1[1991:1984] < top_1[1999:1992]) ? 1 : 0;
assign detect_min[247][6] = (mid_1[1991:1984] < top_2[1983:1976]) ? 1 : 0;
assign detect_min[247][7] = (mid_1[1991:1984] < top_2[1991:1984]) ? 1 : 0;
assign detect_min[247][8] = (mid_1[1991:1984] < top_2[1999:1992]) ? 1 : 0;
assign detect_min[247][9] = (mid_1[1991:1984] < mid_0[1983:1976]) ? 1 : 0;
assign detect_min[247][10] = (mid_1[1991:1984] < mid_0[1991:1984]) ? 1 : 0;
assign detect_min[247][11] = (mid_1[1991:1984] < mid_0[1999:1992]) ? 1 : 0;
assign detect_min[247][12] = (mid_1[1991:1984] < mid_1[1983:1976]) ? 1 : 0;
assign detect_min[247][13] = (mid_1[1991:1984] < mid_1[1999:1992]) ? 1 : 0;
assign detect_min[247][14] = (mid_1[1991:1984] < mid_2[1983:1976]) ? 1 : 0;
assign detect_min[247][15] = (mid_1[1991:1984] < mid_2[1991:1984]) ? 1 : 0;
assign detect_min[247][16] = (mid_1[1991:1984] < mid_2[1999:1992]) ? 1 : 0;
assign detect_min[247][17] = (mid_1[1991:1984] < btm_0[1983:1976]) ? 1 : 0;
assign detect_min[247][18] = (mid_1[1991:1984] < btm_0[1991:1984]) ? 1 : 0;
assign detect_min[247][19] = (mid_1[1991:1984] < btm_0[1999:1992]) ? 1 : 0;
assign detect_min[247][20] = (mid_1[1991:1984] < btm_1[1983:1976]) ? 1 : 0;
assign detect_min[247][21] = (mid_1[1991:1984] < btm_1[1991:1984]) ? 1 : 0;
assign detect_min[247][22] = (mid_1[1991:1984] < btm_1[1999:1992]) ? 1 : 0;
assign detect_min[247][23] = (mid_1[1991:1984] < btm_2[1983:1976]) ? 1 : 0;
assign detect_min[247][24] = (mid_1[1991:1984] < btm_2[1991:1984]) ? 1 : 0;
assign detect_min[247][25] = (mid_1[1991:1984] < btm_2[1999:1992]) ? 1 : 0;

assign detect_min[248][0] = (mid_1[1999:1992] < top_0[1991:1984]) ? 1 : 0;
assign detect_min[248][1] = (mid_1[1999:1992] < top_0[1999:1992]) ? 1 : 0;
assign detect_min[248][2] = (mid_1[1999:1992] < top_0[2007:2000]) ? 1 : 0;
assign detect_min[248][3] = (mid_1[1999:1992] < top_1[1991:1984]) ? 1 : 0;
assign detect_min[248][4] = (mid_1[1999:1992] < top_1[1999:1992]) ? 1 : 0;
assign detect_min[248][5] = (mid_1[1999:1992] < top_1[2007:2000]) ? 1 : 0;
assign detect_min[248][6] = (mid_1[1999:1992] < top_2[1991:1984]) ? 1 : 0;
assign detect_min[248][7] = (mid_1[1999:1992] < top_2[1999:1992]) ? 1 : 0;
assign detect_min[248][8] = (mid_1[1999:1992] < top_2[2007:2000]) ? 1 : 0;
assign detect_min[248][9] = (mid_1[1999:1992] < mid_0[1991:1984]) ? 1 : 0;
assign detect_min[248][10] = (mid_1[1999:1992] < mid_0[1999:1992]) ? 1 : 0;
assign detect_min[248][11] = (mid_1[1999:1992] < mid_0[2007:2000]) ? 1 : 0;
assign detect_min[248][12] = (mid_1[1999:1992] < mid_1[1991:1984]) ? 1 : 0;
assign detect_min[248][13] = (mid_1[1999:1992] < mid_1[2007:2000]) ? 1 : 0;
assign detect_min[248][14] = (mid_1[1999:1992] < mid_2[1991:1984]) ? 1 : 0;
assign detect_min[248][15] = (mid_1[1999:1992] < mid_2[1999:1992]) ? 1 : 0;
assign detect_min[248][16] = (mid_1[1999:1992] < mid_2[2007:2000]) ? 1 : 0;
assign detect_min[248][17] = (mid_1[1999:1992] < btm_0[1991:1984]) ? 1 : 0;
assign detect_min[248][18] = (mid_1[1999:1992] < btm_0[1999:1992]) ? 1 : 0;
assign detect_min[248][19] = (mid_1[1999:1992] < btm_0[2007:2000]) ? 1 : 0;
assign detect_min[248][20] = (mid_1[1999:1992] < btm_1[1991:1984]) ? 1 : 0;
assign detect_min[248][21] = (mid_1[1999:1992] < btm_1[1999:1992]) ? 1 : 0;
assign detect_min[248][22] = (mid_1[1999:1992] < btm_1[2007:2000]) ? 1 : 0;
assign detect_min[248][23] = (mid_1[1999:1992] < btm_2[1991:1984]) ? 1 : 0;
assign detect_min[248][24] = (mid_1[1999:1992] < btm_2[1999:1992]) ? 1 : 0;
assign detect_min[248][25] = (mid_1[1999:1992] < btm_2[2007:2000]) ? 1 : 0;

assign detect_min[249][0] = (mid_1[2007:2000] < top_0[1999:1992]) ? 1 : 0;
assign detect_min[249][1] = (mid_1[2007:2000] < top_0[2007:2000]) ? 1 : 0;
assign detect_min[249][2] = (mid_1[2007:2000] < top_0[2015:2008]) ? 1 : 0;
assign detect_min[249][3] = (mid_1[2007:2000] < top_1[1999:1992]) ? 1 : 0;
assign detect_min[249][4] = (mid_1[2007:2000] < top_1[2007:2000]) ? 1 : 0;
assign detect_min[249][5] = (mid_1[2007:2000] < top_1[2015:2008]) ? 1 : 0;
assign detect_min[249][6] = (mid_1[2007:2000] < top_2[1999:1992]) ? 1 : 0;
assign detect_min[249][7] = (mid_1[2007:2000] < top_2[2007:2000]) ? 1 : 0;
assign detect_min[249][8] = (mid_1[2007:2000] < top_2[2015:2008]) ? 1 : 0;
assign detect_min[249][9] = (mid_1[2007:2000] < mid_0[1999:1992]) ? 1 : 0;
assign detect_min[249][10] = (mid_1[2007:2000] < mid_0[2007:2000]) ? 1 : 0;
assign detect_min[249][11] = (mid_1[2007:2000] < mid_0[2015:2008]) ? 1 : 0;
assign detect_min[249][12] = (mid_1[2007:2000] < mid_1[1999:1992]) ? 1 : 0;
assign detect_min[249][13] = (mid_1[2007:2000] < mid_1[2015:2008]) ? 1 : 0;
assign detect_min[249][14] = (mid_1[2007:2000] < mid_2[1999:1992]) ? 1 : 0;
assign detect_min[249][15] = (mid_1[2007:2000] < mid_2[2007:2000]) ? 1 : 0;
assign detect_min[249][16] = (mid_1[2007:2000] < mid_2[2015:2008]) ? 1 : 0;
assign detect_min[249][17] = (mid_1[2007:2000] < btm_0[1999:1992]) ? 1 : 0;
assign detect_min[249][18] = (mid_1[2007:2000] < btm_0[2007:2000]) ? 1 : 0;
assign detect_min[249][19] = (mid_1[2007:2000] < btm_0[2015:2008]) ? 1 : 0;
assign detect_min[249][20] = (mid_1[2007:2000] < btm_1[1999:1992]) ? 1 : 0;
assign detect_min[249][21] = (mid_1[2007:2000] < btm_1[2007:2000]) ? 1 : 0;
assign detect_min[249][22] = (mid_1[2007:2000] < btm_1[2015:2008]) ? 1 : 0;
assign detect_min[249][23] = (mid_1[2007:2000] < btm_2[1999:1992]) ? 1 : 0;
assign detect_min[249][24] = (mid_1[2007:2000] < btm_2[2007:2000]) ? 1 : 0;
assign detect_min[249][25] = (mid_1[2007:2000] < btm_2[2015:2008]) ? 1 : 0;

assign detect_min[250][0] = (mid_1[2015:2008] < top_0[2007:2000]) ? 1 : 0;
assign detect_min[250][1] = (mid_1[2015:2008] < top_0[2015:2008]) ? 1 : 0;
assign detect_min[250][2] = (mid_1[2015:2008] < top_0[2023:2016]) ? 1 : 0;
assign detect_min[250][3] = (mid_1[2015:2008] < top_1[2007:2000]) ? 1 : 0;
assign detect_min[250][4] = (mid_1[2015:2008] < top_1[2015:2008]) ? 1 : 0;
assign detect_min[250][5] = (mid_1[2015:2008] < top_1[2023:2016]) ? 1 : 0;
assign detect_min[250][6] = (mid_1[2015:2008] < top_2[2007:2000]) ? 1 : 0;
assign detect_min[250][7] = (mid_1[2015:2008] < top_2[2015:2008]) ? 1 : 0;
assign detect_min[250][8] = (mid_1[2015:2008] < top_2[2023:2016]) ? 1 : 0;
assign detect_min[250][9] = (mid_1[2015:2008] < mid_0[2007:2000]) ? 1 : 0;
assign detect_min[250][10] = (mid_1[2015:2008] < mid_0[2015:2008]) ? 1 : 0;
assign detect_min[250][11] = (mid_1[2015:2008] < mid_0[2023:2016]) ? 1 : 0;
assign detect_min[250][12] = (mid_1[2015:2008] < mid_1[2007:2000]) ? 1 : 0;
assign detect_min[250][13] = (mid_1[2015:2008] < mid_1[2023:2016]) ? 1 : 0;
assign detect_min[250][14] = (mid_1[2015:2008] < mid_2[2007:2000]) ? 1 : 0;
assign detect_min[250][15] = (mid_1[2015:2008] < mid_2[2015:2008]) ? 1 : 0;
assign detect_min[250][16] = (mid_1[2015:2008] < mid_2[2023:2016]) ? 1 : 0;
assign detect_min[250][17] = (mid_1[2015:2008] < btm_0[2007:2000]) ? 1 : 0;
assign detect_min[250][18] = (mid_1[2015:2008] < btm_0[2015:2008]) ? 1 : 0;
assign detect_min[250][19] = (mid_1[2015:2008] < btm_0[2023:2016]) ? 1 : 0;
assign detect_min[250][20] = (mid_1[2015:2008] < btm_1[2007:2000]) ? 1 : 0;
assign detect_min[250][21] = (mid_1[2015:2008] < btm_1[2015:2008]) ? 1 : 0;
assign detect_min[250][22] = (mid_1[2015:2008] < btm_1[2023:2016]) ? 1 : 0;
assign detect_min[250][23] = (mid_1[2015:2008] < btm_2[2007:2000]) ? 1 : 0;
assign detect_min[250][24] = (mid_1[2015:2008] < btm_2[2015:2008]) ? 1 : 0;
assign detect_min[250][25] = (mid_1[2015:2008] < btm_2[2023:2016]) ? 1 : 0;

assign detect_min[251][0] = (mid_1[2023:2016] < top_0[2015:2008]) ? 1 : 0;
assign detect_min[251][1] = (mid_1[2023:2016] < top_0[2023:2016]) ? 1 : 0;
assign detect_min[251][2] = (mid_1[2023:2016] < top_0[2031:2024]) ? 1 : 0;
assign detect_min[251][3] = (mid_1[2023:2016] < top_1[2015:2008]) ? 1 : 0;
assign detect_min[251][4] = (mid_1[2023:2016] < top_1[2023:2016]) ? 1 : 0;
assign detect_min[251][5] = (mid_1[2023:2016] < top_1[2031:2024]) ? 1 : 0;
assign detect_min[251][6] = (mid_1[2023:2016] < top_2[2015:2008]) ? 1 : 0;
assign detect_min[251][7] = (mid_1[2023:2016] < top_2[2023:2016]) ? 1 : 0;
assign detect_min[251][8] = (mid_1[2023:2016] < top_2[2031:2024]) ? 1 : 0;
assign detect_min[251][9] = (mid_1[2023:2016] < mid_0[2015:2008]) ? 1 : 0;
assign detect_min[251][10] = (mid_1[2023:2016] < mid_0[2023:2016]) ? 1 : 0;
assign detect_min[251][11] = (mid_1[2023:2016] < mid_0[2031:2024]) ? 1 : 0;
assign detect_min[251][12] = (mid_1[2023:2016] < mid_1[2015:2008]) ? 1 : 0;
assign detect_min[251][13] = (mid_1[2023:2016] < mid_1[2031:2024]) ? 1 : 0;
assign detect_min[251][14] = (mid_1[2023:2016] < mid_2[2015:2008]) ? 1 : 0;
assign detect_min[251][15] = (mid_1[2023:2016] < mid_2[2023:2016]) ? 1 : 0;
assign detect_min[251][16] = (mid_1[2023:2016] < mid_2[2031:2024]) ? 1 : 0;
assign detect_min[251][17] = (mid_1[2023:2016] < btm_0[2015:2008]) ? 1 : 0;
assign detect_min[251][18] = (mid_1[2023:2016] < btm_0[2023:2016]) ? 1 : 0;
assign detect_min[251][19] = (mid_1[2023:2016] < btm_0[2031:2024]) ? 1 : 0;
assign detect_min[251][20] = (mid_1[2023:2016] < btm_1[2015:2008]) ? 1 : 0;
assign detect_min[251][21] = (mid_1[2023:2016] < btm_1[2023:2016]) ? 1 : 0;
assign detect_min[251][22] = (mid_1[2023:2016] < btm_1[2031:2024]) ? 1 : 0;
assign detect_min[251][23] = (mid_1[2023:2016] < btm_2[2015:2008]) ? 1 : 0;
assign detect_min[251][24] = (mid_1[2023:2016] < btm_2[2023:2016]) ? 1 : 0;
assign detect_min[251][25] = (mid_1[2023:2016] < btm_2[2031:2024]) ? 1 : 0;

assign detect_min[252][0] = (mid_1[2031:2024] < top_0[2023:2016]) ? 1 : 0;
assign detect_min[252][1] = (mid_1[2031:2024] < top_0[2031:2024]) ? 1 : 0;
assign detect_min[252][2] = (mid_1[2031:2024] < top_0[2039:2032]) ? 1 : 0;
assign detect_min[252][3] = (mid_1[2031:2024] < top_1[2023:2016]) ? 1 : 0;
assign detect_min[252][4] = (mid_1[2031:2024] < top_1[2031:2024]) ? 1 : 0;
assign detect_min[252][5] = (mid_1[2031:2024] < top_1[2039:2032]) ? 1 : 0;
assign detect_min[252][6] = (mid_1[2031:2024] < top_2[2023:2016]) ? 1 : 0;
assign detect_min[252][7] = (mid_1[2031:2024] < top_2[2031:2024]) ? 1 : 0;
assign detect_min[252][8] = (mid_1[2031:2024] < top_2[2039:2032]) ? 1 : 0;
assign detect_min[252][9] = (mid_1[2031:2024] < mid_0[2023:2016]) ? 1 : 0;
assign detect_min[252][10] = (mid_1[2031:2024] < mid_0[2031:2024]) ? 1 : 0;
assign detect_min[252][11] = (mid_1[2031:2024] < mid_0[2039:2032]) ? 1 : 0;
assign detect_min[252][12] = (mid_1[2031:2024] < mid_1[2023:2016]) ? 1 : 0;
assign detect_min[252][13] = (mid_1[2031:2024] < mid_1[2039:2032]) ? 1 : 0;
assign detect_min[252][14] = (mid_1[2031:2024] < mid_2[2023:2016]) ? 1 : 0;
assign detect_min[252][15] = (mid_1[2031:2024] < mid_2[2031:2024]) ? 1 : 0;
assign detect_min[252][16] = (mid_1[2031:2024] < mid_2[2039:2032]) ? 1 : 0;
assign detect_min[252][17] = (mid_1[2031:2024] < btm_0[2023:2016]) ? 1 : 0;
assign detect_min[252][18] = (mid_1[2031:2024] < btm_0[2031:2024]) ? 1 : 0;
assign detect_min[252][19] = (mid_1[2031:2024] < btm_0[2039:2032]) ? 1 : 0;
assign detect_min[252][20] = (mid_1[2031:2024] < btm_1[2023:2016]) ? 1 : 0;
assign detect_min[252][21] = (mid_1[2031:2024] < btm_1[2031:2024]) ? 1 : 0;
assign detect_min[252][22] = (mid_1[2031:2024] < btm_1[2039:2032]) ? 1 : 0;
assign detect_min[252][23] = (mid_1[2031:2024] < btm_2[2023:2016]) ? 1 : 0;
assign detect_min[252][24] = (mid_1[2031:2024] < btm_2[2031:2024]) ? 1 : 0;
assign detect_min[252][25] = (mid_1[2031:2024] < btm_2[2039:2032]) ? 1 : 0;

assign detect_min[253][0] = (mid_1[2039:2032] < top_0[2031:2024]) ? 1 : 0;
assign detect_min[253][1] = (mid_1[2039:2032] < top_0[2039:2032]) ? 1 : 0;
assign detect_min[253][2] = (mid_1[2039:2032] < top_0[2047:2040]) ? 1 : 0;
assign detect_min[253][3] = (mid_1[2039:2032] < top_1[2031:2024]) ? 1 : 0;
assign detect_min[253][4] = (mid_1[2039:2032] < top_1[2039:2032]) ? 1 : 0;
assign detect_min[253][5] = (mid_1[2039:2032] < top_1[2047:2040]) ? 1 : 0;
assign detect_min[253][6] = (mid_1[2039:2032] < top_2[2031:2024]) ? 1 : 0;
assign detect_min[253][7] = (mid_1[2039:2032] < top_2[2039:2032]) ? 1 : 0;
assign detect_min[253][8] = (mid_1[2039:2032] < top_2[2047:2040]) ? 1 : 0;
assign detect_min[253][9] = (mid_1[2039:2032] < mid_0[2031:2024]) ? 1 : 0;
assign detect_min[253][10] = (mid_1[2039:2032] < mid_0[2039:2032]) ? 1 : 0;
assign detect_min[253][11] = (mid_1[2039:2032] < mid_0[2047:2040]) ? 1 : 0;
assign detect_min[253][12] = (mid_1[2039:2032] < mid_1[2031:2024]) ? 1 : 0;
assign detect_min[253][13] = (mid_1[2039:2032] < mid_1[2047:2040]) ? 1 : 0;
assign detect_min[253][14] = (mid_1[2039:2032] < mid_2[2031:2024]) ? 1 : 0;
assign detect_min[253][15] = (mid_1[2039:2032] < mid_2[2039:2032]) ? 1 : 0;
assign detect_min[253][16] = (mid_1[2039:2032] < mid_2[2047:2040]) ? 1 : 0;
assign detect_min[253][17] = (mid_1[2039:2032] < btm_0[2031:2024]) ? 1 : 0;
assign detect_min[253][18] = (mid_1[2039:2032] < btm_0[2039:2032]) ? 1 : 0;
assign detect_min[253][19] = (mid_1[2039:2032] < btm_0[2047:2040]) ? 1 : 0;
assign detect_min[253][20] = (mid_1[2039:2032] < btm_1[2031:2024]) ? 1 : 0;
assign detect_min[253][21] = (mid_1[2039:2032] < btm_1[2039:2032]) ? 1 : 0;
assign detect_min[253][22] = (mid_1[2039:2032] < btm_1[2047:2040]) ? 1 : 0;
assign detect_min[253][23] = (mid_1[2039:2032] < btm_2[2031:2024]) ? 1 : 0;
assign detect_min[253][24] = (mid_1[2039:2032] < btm_2[2039:2032]) ? 1 : 0;
assign detect_min[253][25] = (mid_1[2039:2032] < btm_2[2047:2040]) ? 1 : 0;

assign detect_min[254][0] = (mid_1[2047:2040] < top_0[2039:2032]) ? 1 : 0;
assign detect_min[254][1] = (mid_1[2047:2040] < top_0[2047:2040]) ? 1 : 0;
assign detect_min[254][2] = (mid_1[2047:2040] < top_0[2055:2048]) ? 1 : 0;
assign detect_min[254][3] = (mid_1[2047:2040] < top_1[2039:2032]) ? 1 : 0;
assign detect_min[254][4] = (mid_1[2047:2040] < top_1[2047:2040]) ? 1 : 0;
assign detect_min[254][5] = (mid_1[2047:2040] < top_1[2055:2048]) ? 1 : 0;
assign detect_min[254][6] = (mid_1[2047:2040] < top_2[2039:2032]) ? 1 : 0;
assign detect_min[254][7] = (mid_1[2047:2040] < top_2[2047:2040]) ? 1 : 0;
assign detect_min[254][8] = (mid_1[2047:2040] < top_2[2055:2048]) ? 1 : 0;
assign detect_min[254][9] = (mid_1[2047:2040] < mid_0[2039:2032]) ? 1 : 0;
assign detect_min[254][10] = (mid_1[2047:2040] < mid_0[2047:2040]) ? 1 : 0;
assign detect_min[254][11] = (mid_1[2047:2040] < mid_0[2055:2048]) ? 1 : 0;
assign detect_min[254][12] = (mid_1[2047:2040] < mid_1[2039:2032]) ? 1 : 0;
assign detect_min[254][13] = (mid_1[2047:2040] < mid_1[2055:2048]) ? 1 : 0;
assign detect_min[254][14] = (mid_1[2047:2040] < mid_2[2039:2032]) ? 1 : 0;
assign detect_min[254][15] = (mid_1[2047:2040] < mid_2[2047:2040]) ? 1 : 0;
assign detect_min[254][16] = (mid_1[2047:2040] < mid_2[2055:2048]) ? 1 : 0;
assign detect_min[254][17] = (mid_1[2047:2040] < btm_0[2039:2032]) ? 1 : 0;
assign detect_min[254][18] = (mid_1[2047:2040] < btm_0[2047:2040]) ? 1 : 0;
assign detect_min[254][19] = (mid_1[2047:2040] < btm_0[2055:2048]) ? 1 : 0;
assign detect_min[254][20] = (mid_1[2047:2040] < btm_1[2039:2032]) ? 1 : 0;
assign detect_min[254][21] = (mid_1[2047:2040] < btm_1[2047:2040]) ? 1 : 0;
assign detect_min[254][22] = (mid_1[2047:2040] < btm_1[2055:2048]) ? 1 : 0;
assign detect_min[254][23] = (mid_1[2047:2040] < btm_2[2039:2032]) ? 1 : 0;
assign detect_min[254][24] = (mid_1[2047:2040] < btm_2[2047:2040]) ? 1 : 0;
assign detect_min[254][25] = (mid_1[2047:2040] < btm_2[2055:2048]) ? 1 : 0;

assign detect_min[255][0] = (mid_1[2055:2048] < top_0[2047:2040]) ? 1 : 0;
assign detect_min[255][1] = (mid_1[2055:2048] < top_0[2055:2048]) ? 1 : 0;
assign detect_min[255][2] = (mid_1[2055:2048] < top_0[2063:2056]) ? 1 : 0;
assign detect_min[255][3] = (mid_1[2055:2048] < top_1[2047:2040]) ? 1 : 0;
assign detect_min[255][4] = (mid_1[2055:2048] < top_1[2055:2048]) ? 1 : 0;
assign detect_min[255][5] = (mid_1[2055:2048] < top_1[2063:2056]) ? 1 : 0;
assign detect_min[255][6] = (mid_1[2055:2048] < top_2[2047:2040]) ? 1 : 0;
assign detect_min[255][7] = (mid_1[2055:2048] < top_2[2055:2048]) ? 1 : 0;
assign detect_min[255][8] = (mid_1[2055:2048] < top_2[2063:2056]) ? 1 : 0;
assign detect_min[255][9] = (mid_1[2055:2048] < mid_0[2047:2040]) ? 1 : 0;
assign detect_min[255][10] = (mid_1[2055:2048] < mid_0[2055:2048]) ? 1 : 0;
assign detect_min[255][11] = (mid_1[2055:2048] < mid_0[2063:2056]) ? 1 : 0;
assign detect_min[255][12] = (mid_1[2055:2048] < mid_1[2047:2040]) ? 1 : 0;
assign detect_min[255][13] = (mid_1[2055:2048] < mid_1[2063:2056]) ? 1 : 0;
assign detect_min[255][14] = (mid_1[2055:2048] < mid_2[2047:2040]) ? 1 : 0;
assign detect_min[255][15] = (mid_1[2055:2048] < mid_2[2055:2048]) ? 1 : 0;
assign detect_min[255][16] = (mid_1[2055:2048] < mid_2[2063:2056]) ? 1 : 0;
assign detect_min[255][17] = (mid_1[2055:2048] < btm_0[2047:2040]) ? 1 : 0;
assign detect_min[255][18] = (mid_1[2055:2048] < btm_0[2055:2048]) ? 1 : 0;
assign detect_min[255][19] = (mid_1[2055:2048] < btm_0[2063:2056]) ? 1 : 0;
assign detect_min[255][20] = (mid_1[2055:2048] < btm_1[2047:2040]) ? 1 : 0;
assign detect_min[255][21] = (mid_1[2055:2048] < btm_1[2055:2048]) ? 1 : 0;
assign detect_min[255][22] = (mid_1[2055:2048] < btm_1[2063:2056]) ? 1 : 0;
assign detect_min[255][23] = (mid_1[2055:2048] < btm_2[2047:2040]) ? 1 : 0;
assign detect_min[255][24] = (mid_1[2055:2048] < btm_2[2055:2048]) ? 1 : 0;
assign detect_min[255][25] = (mid_1[2055:2048] < btm_2[2063:2056]) ? 1 : 0;

assign detect_min[256][0] = (mid_1[2063:2056] < top_0[2055:2048]) ? 1 : 0;
assign detect_min[256][1] = (mid_1[2063:2056] < top_0[2063:2056]) ? 1 : 0;
assign detect_min[256][2] = (mid_1[2063:2056] < top_0[2071:2064]) ? 1 : 0;
assign detect_min[256][3] = (mid_1[2063:2056] < top_1[2055:2048]) ? 1 : 0;
assign detect_min[256][4] = (mid_1[2063:2056] < top_1[2063:2056]) ? 1 : 0;
assign detect_min[256][5] = (mid_1[2063:2056] < top_1[2071:2064]) ? 1 : 0;
assign detect_min[256][6] = (mid_1[2063:2056] < top_2[2055:2048]) ? 1 : 0;
assign detect_min[256][7] = (mid_1[2063:2056] < top_2[2063:2056]) ? 1 : 0;
assign detect_min[256][8] = (mid_1[2063:2056] < top_2[2071:2064]) ? 1 : 0;
assign detect_min[256][9] = (mid_1[2063:2056] < mid_0[2055:2048]) ? 1 : 0;
assign detect_min[256][10] = (mid_1[2063:2056] < mid_0[2063:2056]) ? 1 : 0;
assign detect_min[256][11] = (mid_1[2063:2056] < mid_0[2071:2064]) ? 1 : 0;
assign detect_min[256][12] = (mid_1[2063:2056] < mid_1[2055:2048]) ? 1 : 0;
assign detect_min[256][13] = (mid_1[2063:2056] < mid_1[2071:2064]) ? 1 : 0;
assign detect_min[256][14] = (mid_1[2063:2056] < mid_2[2055:2048]) ? 1 : 0;
assign detect_min[256][15] = (mid_1[2063:2056] < mid_2[2063:2056]) ? 1 : 0;
assign detect_min[256][16] = (mid_1[2063:2056] < mid_2[2071:2064]) ? 1 : 0;
assign detect_min[256][17] = (mid_1[2063:2056] < btm_0[2055:2048]) ? 1 : 0;
assign detect_min[256][18] = (mid_1[2063:2056] < btm_0[2063:2056]) ? 1 : 0;
assign detect_min[256][19] = (mid_1[2063:2056] < btm_0[2071:2064]) ? 1 : 0;
assign detect_min[256][20] = (mid_1[2063:2056] < btm_1[2055:2048]) ? 1 : 0;
assign detect_min[256][21] = (mid_1[2063:2056] < btm_1[2063:2056]) ? 1 : 0;
assign detect_min[256][22] = (mid_1[2063:2056] < btm_1[2071:2064]) ? 1 : 0;
assign detect_min[256][23] = (mid_1[2063:2056] < btm_2[2055:2048]) ? 1 : 0;
assign detect_min[256][24] = (mid_1[2063:2056] < btm_2[2063:2056]) ? 1 : 0;
assign detect_min[256][25] = (mid_1[2063:2056] < btm_2[2071:2064]) ? 1 : 0;

assign detect_min[257][0] = (mid_1[2071:2064] < top_0[2063:2056]) ? 1 : 0;
assign detect_min[257][1] = (mid_1[2071:2064] < top_0[2071:2064]) ? 1 : 0;
assign detect_min[257][2] = (mid_1[2071:2064] < top_0[2079:2072]) ? 1 : 0;
assign detect_min[257][3] = (mid_1[2071:2064] < top_1[2063:2056]) ? 1 : 0;
assign detect_min[257][4] = (mid_1[2071:2064] < top_1[2071:2064]) ? 1 : 0;
assign detect_min[257][5] = (mid_1[2071:2064] < top_1[2079:2072]) ? 1 : 0;
assign detect_min[257][6] = (mid_1[2071:2064] < top_2[2063:2056]) ? 1 : 0;
assign detect_min[257][7] = (mid_1[2071:2064] < top_2[2071:2064]) ? 1 : 0;
assign detect_min[257][8] = (mid_1[2071:2064] < top_2[2079:2072]) ? 1 : 0;
assign detect_min[257][9] = (mid_1[2071:2064] < mid_0[2063:2056]) ? 1 : 0;
assign detect_min[257][10] = (mid_1[2071:2064] < mid_0[2071:2064]) ? 1 : 0;
assign detect_min[257][11] = (mid_1[2071:2064] < mid_0[2079:2072]) ? 1 : 0;
assign detect_min[257][12] = (mid_1[2071:2064] < mid_1[2063:2056]) ? 1 : 0;
assign detect_min[257][13] = (mid_1[2071:2064] < mid_1[2079:2072]) ? 1 : 0;
assign detect_min[257][14] = (mid_1[2071:2064] < mid_2[2063:2056]) ? 1 : 0;
assign detect_min[257][15] = (mid_1[2071:2064] < mid_2[2071:2064]) ? 1 : 0;
assign detect_min[257][16] = (mid_1[2071:2064] < mid_2[2079:2072]) ? 1 : 0;
assign detect_min[257][17] = (mid_1[2071:2064] < btm_0[2063:2056]) ? 1 : 0;
assign detect_min[257][18] = (mid_1[2071:2064] < btm_0[2071:2064]) ? 1 : 0;
assign detect_min[257][19] = (mid_1[2071:2064] < btm_0[2079:2072]) ? 1 : 0;
assign detect_min[257][20] = (mid_1[2071:2064] < btm_1[2063:2056]) ? 1 : 0;
assign detect_min[257][21] = (mid_1[2071:2064] < btm_1[2071:2064]) ? 1 : 0;
assign detect_min[257][22] = (mid_1[2071:2064] < btm_1[2079:2072]) ? 1 : 0;
assign detect_min[257][23] = (mid_1[2071:2064] < btm_2[2063:2056]) ? 1 : 0;
assign detect_min[257][24] = (mid_1[2071:2064] < btm_2[2071:2064]) ? 1 : 0;
assign detect_min[257][25] = (mid_1[2071:2064] < btm_2[2079:2072]) ? 1 : 0;

assign detect_min[258][0] = (mid_1[2079:2072] < top_0[2071:2064]) ? 1 : 0;
assign detect_min[258][1] = (mid_1[2079:2072] < top_0[2079:2072]) ? 1 : 0;
assign detect_min[258][2] = (mid_1[2079:2072] < top_0[2087:2080]) ? 1 : 0;
assign detect_min[258][3] = (mid_1[2079:2072] < top_1[2071:2064]) ? 1 : 0;
assign detect_min[258][4] = (mid_1[2079:2072] < top_1[2079:2072]) ? 1 : 0;
assign detect_min[258][5] = (mid_1[2079:2072] < top_1[2087:2080]) ? 1 : 0;
assign detect_min[258][6] = (mid_1[2079:2072] < top_2[2071:2064]) ? 1 : 0;
assign detect_min[258][7] = (mid_1[2079:2072] < top_2[2079:2072]) ? 1 : 0;
assign detect_min[258][8] = (mid_1[2079:2072] < top_2[2087:2080]) ? 1 : 0;
assign detect_min[258][9] = (mid_1[2079:2072] < mid_0[2071:2064]) ? 1 : 0;
assign detect_min[258][10] = (mid_1[2079:2072] < mid_0[2079:2072]) ? 1 : 0;
assign detect_min[258][11] = (mid_1[2079:2072] < mid_0[2087:2080]) ? 1 : 0;
assign detect_min[258][12] = (mid_1[2079:2072] < mid_1[2071:2064]) ? 1 : 0;
assign detect_min[258][13] = (mid_1[2079:2072] < mid_1[2087:2080]) ? 1 : 0;
assign detect_min[258][14] = (mid_1[2079:2072] < mid_2[2071:2064]) ? 1 : 0;
assign detect_min[258][15] = (mid_1[2079:2072] < mid_2[2079:2072]) ? 1 : 0;
assign detect_min[258][16] = (mid_1[2079:2072] < mid_2[2087:2080]) ? 1 : 0;
assign detect_min[258][17] = (mid_1[2079:2072] < btm_0[2071:2064]) ? 1 : 0;
assign detect_min[258][18] = (mid_1[2079:2072] < btm_0[2079:2072]) ? 1 : 0;
assign detect_min[258][19] = (mid_1[2079:2072] < btm_0[2087:2080]) ? 1 : 0;
assign detect_min[258][20] = (mid_1[2079:2072] < btm_1[2071:2064]) ? 1 : 0;
assign detect_min[258][21] = (mid_1[2079:2072] < btm_1[2079:2072]) ? 1 : 0;
assign detect_min[258][22] = (mid_1[2079:2072] < btm_1[2087:2080]) ? 1 : 0;
assign detect_min[258][23] = (mid_1[2079:2072] < btm_2[2071:2064]) ? 1 : 0;
assign detect_min[258][24] = (mid_1[2079:2072] < btm_2[2079:2072]) ? 1 : 0;
assign detect_min[258][25] = (mid_1[2079:2072] < btm_2[2087:2080]) ? 1 : 0;

assign detect_min[259][0] = (mid_1[2087:2080] < top_0[2079:2072]) ? 1 : 0;
assign detect_min[259][1] = (mid_1[2087:2080] < top_0[2087:2080]) ? 1 : 0;
assign detect_min[259][2] = (mid_1[2087:2080] < top_0[2095:2088]) ? 1 : 0;
assign detect_min[259][3] = (mid_1[2087:2080] < top_1[2079:2072]) ? 1 : 0;
assign detect_min[259][4] = (mid_1[2087:2080] < top_1[2087:2080]) ? 1 : 0;
assign detect_min[259][5] = (mid_1[2087:2080] < top_1[2095:2088]) ? 1 : 0;
assign detect_min[259][6] = (mid_1[2087:2080] < top_2[2079:2072]) ? 1 : 0;
assign detect_min[259][7] = (mid_1[2087:2080] < top_2[2087:2080]) ? 1 : 0;
assign detect_min[259][8] = (mid_1[2087:2080] < top_2[2095:2088]) ? 1 : 0;
assign detect_min[259][9] = (mid_1[2087:2080] < mid_0[2079:2072]) ? 1 : 0;
assign detect_min[259][10] = (mid_1[2087:2080] < mid_0[2087:2080]) ? 1 : 0;
assign detect_min[259][11] = (mid_1[2087:2080] < mid_0[2095:2088]) ? 1 : 0;
assign detect_min[259][12] = (mid_1[2087:2080] < mid_1[2079:2072]) ? 1 : 0;
assign detect_min[259][13] = (mid_1[2087:2080] < mid_1[2095:2088]) ? 1 : 0;
assign detect_min[259][14] = (mid_1[2087:2080] < mid_2[2079:2072]) ? 1 : 0;
assign detect_min[259][15] = (mid_1[2087:2080] < mid_2[2087:2080]) ? 1 : 0;
assign detect_min[259][16] = (mid_1[2087:2080] < mid_2[2095:2088]) ? 1 : 0;
assign detect_min[259][17] = (mid_1[2087:2080] < btm_0[2079:2072]) ? 1 : 0;
assign detect_min[259][18] = (mid_1[2087:2080] < btm_0[2087:2080]) ? 1 : 0;
assign detect_min[259][19] = (mid_1[2087:2080] < btm_0[2095:2088]) ? 1 : 0;
assign detect_min[259][20] = (mid_1[2087:2080] < btm_1[2079:2072]) ? 1 : 0;
assign detect_min[259][21] = (mid_1[2087:2080] < btm_1[2087:2080]) ? 1 : 0;
assign detect_min[259][22] = (mid_1[2087:2080] < btm_1[2095:2088]) ? 1 : 0;
assign detect_min[259][23] = (mid_1[2087:2080] < btm_2[2079:2072]) ? 1 : 0;
assign detect_min[259][24] = (mid_1[2087:2080] < btm_2[2087:2080]) ? 1 : 0;
assign detect_min[259][25] = (mid_1[2087:2080] < btm_2[2095:2088]) ? 1 : 0;

assign detect_min[260][0] = (mid_1[2095:2088] < top_0[2087:2080]) ? 1 : 0;
assign detect_min[260][1] = (mid_1[2095:2088] < top_0[2095:2088]) ? 1 : 0;
assign detect_min[260][2] = (mid_1[2095:2088] < top_0[2103:2096]) ? 1 : 0;
assign detect_min[260][3] = (mid_1[2095:2088] < top_1[2087:2080]) ? 1 : 0;
assign detect_min[260][4] = (mid_1[2095:2088] < top_1[2095:2088]) ? 1 : 0;
assign detect_min[260][5] = (mid_1[2095:2088] < top_1[2103:2096]) ? 1 : 0;
assign detect_min[260][6] = (mid_1[2095:2088] < top_2[2087:2080]) ? 1 : 0;
assign detect_min[260][7] = (mid_1[2095:2088] < top_2[2095:2088]) ? 1 : 0;
assign detect_min[260][8] = (mid_1[2095:2088] < top_2[2103:2096]) ? 1 : 0;
assign detect_min[260][9] = (mid_1[2095:2088] < mid_0[2087:2080]) ? 1 : 0;
assign detect_min[260][10] = (mid_1[2095:2088] < mid_0[2095:2088]) ? 1 : 0;
assign detect_min[260][11] = (mid_1[2095:2088] < mid_0[2103:2096]) ? 1 : 0;
assign detect_min[260][12] = (mid_1[2095:2088] < mid_1[2087:2080]) ? 1 : 0;
assign detect_min[260][13] = (mid_1[2095:2088] < mid_1[2103:2096]) ? 1 : 0;
assign detect_min[260][14] = (mid_1[2095:2088] < mid_2[2087:2080]) ? 1 : 0;
assign detect_min[260][15] = (mid_1[2095:2088] < mid_2[2095:2088]) ? 1 : 0;
assign detect_min[260][16] = (mid_1[2095:2088] < mid_2[2103:2096]) ? 1 : 0;
assign detect_min[260][17] = (mid_1[2095:2088] < btm_0[2087:2080]) ? 1 : 0;
assign detect_min[260][18] = (mid_1[2095:2088] < btm_0[2095:2088]) ? 1 : 0;
assign detect_min[260][19] = (mid_1[2095:2088] < btm_0[2103:2096]) ? 1 : 0;
assign detect_min[260][20] = (mid_1[2095:2088] < btm_1[2087:2080]) ? 1 : 0;
assign detect_min[260][21] = (mid_1[2095:2088] < btm_1[2095:2088]) ? 1 : 0;
assign detect_min[260][22] = (mid_1[2095:2088] < btm_1[2103:2096]) ? 1 : 0;
assign detect_min[260][23] = (mid_1[2095:2088] < btm_2[2087:2080]) ? 1 : 0;
assign detect_min[260][24] = (mid_1[2095:2088] < btm_2[2095:2088]) ? 1 : 0;
assign detect_min[260][25] = (mid_1[2095:2088] < btm_2[2103:2096]) ? 1 : 0;

assign detect_min[261][0] = (mid_1[2103:2096] < top_0[2095:2088]) ? 1 : 0;
assign detect_min[261][1] = (mid_1[2103:2096] < top_0[2103:2096]) ? 1 : 0;
assign detect_min[261][2] = (mid_1[2103:2096] < top_0[2111:2104]) ? 1 : 0;
assign detect_min[261][3] = (mid_1[2103:2096] < top_1[2095:2088]) ? 1 : 0;
assign detect_min[261][4] = (mid_1[2103:2096] < top_1[2103:2096]) ? 1 : 0;
assign detect_min[261][5] = (mid_1[2103:2096] < top_1[2111:2104]) ? 1 : 0;
assign detect_min[261][6] = (mid_1[2103:2096] < top_2[2095:2088]) ? 1 : 0;
assign detect_min[261][7] = (mid_1[2103:2096] < top_2[2103:2096]) ? 1 : 0;
assign detect_min[261][8] = (mid_1[2103:2096] < top_2[2111:2104]) ? 1 : 0;
assign detect_min[261][9] = (mid_1[2103:2096] < mid_0[2095:2088]) ? 1 : 0;
assign detect_min[261][10] = (mid_1[2103:2096] < mid_0[2103:2096]) ? 1 : 0;
assign detect_min[261][11] = (mid_1[2103:2096] < mid_0[2111:2104]) ? 1 : 0;
assign detect_min[261][12] = (mid_1[2103:2096] < mid_1[2095:2088]) ? 1 : 0;
assign detect_min[261][13] = (mid_1[2103:2096] < mid_1[2111:2104]) ? 1 : 0;
assign detect_min[261][14] = (mid_1[2103:2096] < mid_2[2095:2088]) ? 1 : 0;
assign detect_min[261][15] = (mid_1[2103:2096] < mid_2[2103:2096]) ? 1 : 0;
assign detect_min[261][16] = (mid_1[2103:2096] < mid_2[2111:2104]) ? 1 : 0;
assign detect_min[261][17] = (mid_1[2103:2096] < btm_0[2095:2088]) ? 1 : 0;
assign detect_min[261][18] = (mid_1[2103:2096] < btm_0[2103:2096]) ? 1 : 0;
assign detect_min[261][19] = (mid_1[2103:2096] < btm_0[2111:2104]) ? 1 : 0;
assign detect_min[261][20] = (mid_1[2103:2096] < btm_1[2095:2088]) ? 1 : 0;
assign detect_min[261][21] = (mid_1[2103:2096] < btm_1[2103:2096]) ? 1 : 0;
assign detect_min[261][22] = (mid_1[2103:2096] < btm_1[2111:2104]) ? 1 : 0;
assign detect_min[261][23] = (mid_1[2103:2096] < btm_2[2095:2088]) ? 1 : 0;
assign detect_min[261][24] = (mid_1[2103:2096] < btm_2[2103:2096]) ? 1 : 0;
assign detect_min[261][25] = (mid_1[2103:2096] < btm_2[2111:2104]) ? 1 : 0;

assign detect_min[262][0] = (mid_1[2111:2104] < top_0[2103:2096]) ? 1 : 0;
assign detect_min[262][1] = (mid_1[2111:2104] < top_0[2111:2104]) ? 1 : 0;
assign detect_min[262][2] = (mid_1[2111:2104] < top_0[2119:2112]) ? 1 : 0;
assign detect_min[262][3] = (mid_1[2111:2104] < top_1[2103:2096]) ? 1 : 0;
assign detect_min[262][4] = (mid_1[2111:2104] < top_1[2111:2104]) ? 1 : 0;
assign detect_min[262][5] = (mid_1[2111:2104] < top_1[2119:2112]) ? 1 : 0;
assign detect_min[262][6] = (mid_1[2111:2104] < top_2[2103:2096]) ? 1 : 0;
assign detect_min[262][7] = (mid_1[2111:2104] < top_2[2111:2104]) ? 1 : 0;
assign detect_min[262][8] = (mid_1[2111:2104] < top_2[2119:2112]) ? 1 : 0;
assign detect_min[262][9] = (mid_1[2111:2104] < mid_0[2103:2096]) ? 1 : 0;
assign detect_min[262][10] = (mid_1[2111:2104] < mid_0[2111:2104]) ? 1 : 0;
assign detect_min[262][11] = (mid_1[2111:2104] < mid_0[2119:2112]) ? 1 : 0;
assign detect_min[262][12] = (mid_1[2111:2104] < mid_1[2103:2096]) ? 1 : 0;
assign detect_min[262][13] = (mid_1[2111:2104] < mid_1[2119:2112]) ? 1 : 0;
assign detect_min[262][14] = (mid_1[2111:2104] < mid_2[2103:2096]) ? 1 : 0;
assign detect_min[262][15] = (mid_1[2111:2104] < mid_2[2111:2104]) ? 1 : 0;
assign detect_min[262][16] = (mid_1[2111:2104] < mid_2[2119:2112]) ? 1 : 0;
assign detect_min[262][17] = (mid_1[2111:2104] < btm_0[2103:2096]) ? 1 : 0;
assign detect_min[262][18] = (mid_1[2111:2104] < btm_0[2111:2104]) ? 1 : 0;
assign detect_min[262][19] = (mid_1[2111:2104] < btm_0[2119:2112]) ? 1 : 0;
assign detect_min[262][20] = (mid_1[2111:2104] < btm_1[2103:2096]) ? 1 : 0;
assign detect_min[262][21] = (mid_1[2111:2104] < btm_1[2111:2104]) ? 1 : 0;
assign detect_min[262][22] = (mid_1[2111:2104] < btm_1[2119:2112]) ? 1 : 0;
assign detect_min[262][23] = (mid_1[2111:2104] < btm_2[2103:2096]) ? 1 : 0;
assign detect_min[262][24] = (mid_1[2111:2104] < btm_2[2111:2104]) ? 1 : 0;
assign detect_min[262][25] = (mid_1[2111:2104] < btm_2[2119:2112]) ? 1 : 0;

assign detect_min[263][0] = (mid_1[2119:2112] < top_0[2111:2104]) ? 1 : 0;
assign detect_min[263][1] = (mid_1[2119:2112] < top_0[2119:2112]) ? 1 : 0;
assign detect_min[263][2] = (mid_1[2119:2112] < top_0[2127:2120]) ? 1 : 0;
assign detect_min[263][3] = (mid_1[2119:2112] < top_1[2111:2104]) ? 1 : 0;
assign detect_min[263][4] = (mid_1[2119:2112] < top_1[2119:2112]) ? 1 : 0;
assign detect_min[263][5] = (mid_1[2119:2112] < top_1[2127:2120]) ? 1 : 0;
assign detect_min[263][6] = (mid_1[2119:2112] < top_2[2111:2104]) ? 1 : 0;
assign detect_min[263][7] = (mid_1[2119:2112] < top_2[2119:2112]) ? 1 : 0;
assign detect_min[263][8] = (mid_1[2119:2112] < top_2[2127:2120]) ? 1 : 0;
assign detect_min[263][9] = (mid_1[2119:2112] < mid_0[2111:2104]) ? 1 : 0;
assign detect_min[263][10] = (mid_1[2119:2112] < mid_0[2119:2112]) ? 1 : 0;
assign detect_min[263][11] = (mid_1[2119:2112] < mid_0[2127:2120]) ? 1 : 0;
assign detect_min[263][12] = (mid_1[2119:2112] < mid_1[2111:2104]) ? 1 : 0;
assign detect_min[263][13] = (mid_1[2119:2112] < mid_1[2127:2120]) ? 1 : 0;
assign detect_min[263][14] = (mid_1[2119:2112] < mid_2[2111:2104]) ? 1 : 0;
assign detect_min[263][15] = (mid_1[2119:2112] < mid_2[2119:2112]) ? 1 : 0;
assign detect_min[263][16] = (mid_1[2119:2112] < mid_2[2127:2120]) ? 1 : 0;
assign detect_min[263][17] = (mid_1[2119:2112] < btm_0[2111:2104]) ? 1 : 0;
assign detect_min[263][18] = (mid_1[2119:2112] < btm_0[2119:2112]) ? 1 : 0;
assign detect_min[263][19] = (mid_1[2119:2112] < btm_0[2127:2120]) ? 1 : 0;
assign detect_min[263][20] = (mid_1[2119:2112] < btm_1[2111:2104]) ? 1 : 0;
assign detect_min[263][21] = (mid_1[2119:2112] < btm_1[2119:2112]) ? 1 : 0;
assign detect_min[263][22] = (mid_1[2119:2112] < btm_1[2127:2120]) ? 1 : 0;
assign detect_min[263][23] = (mid_1[2119:2112] < btm_2[2111:2104]) ? 1 : 0;
assign detect_min[263][24] = (mid_1[2119:2112] < btm_2[2119:2112]) ? 1 : 0;
assign detect_min[263][25] = (mid_1[2119:2112] < btm_2[2127:2120]) ? 1 : 0;

assign detect_min[264][0] = (mid_1[2127:2120] < top_0[2119:2112]) ? 1 : 0;
assign detect_min[264][1] = (mid_1[2127:2120] < top_0[2127:2120]) ? 1 : 0;
assign detect_min[264][2] = (mid_1[2127:2120] < top_0[2135:2128]) ? 1 : 0;
assign detect_min[264][3] = (mid_1[2127:2120] < top_1[2119:2112]) ? 1 : 0;
assign detect_min[264][4] = (mid_1[2127:2120] < top_1[2127:2120]) ? 1 : 0;
assign detect_min[264][5] = (mid_1[2127:2120] < top_1[2135:2128]) ? 1 : 0;
assign detect_min[264][6] = (mid_1[2127:2120] < top_2[2119:2112]) ? 1 : 0;
assign detect_min[264][7] = (mid_1[2127:2120] < top_2[2127:2120]) ? 1 : 0;
assign detect_min[264][8] = (mid_1[2127:2120] < top_2[2135:2128]) ? 1 : 0;
assign detect_min[264][9] = (mid_1[2127:2120] < mid_0[2119:2112]) ? 1 : 0;
assign detect_min[264][10] = (mid_1[2127:2120] < mid_0[2127:2120]) ? 1 : 0;
assign detect_min[264][11] = (mid_1[2127:2120] < mid_0[2135:2128]) ? 1 : 0;
assign detect_min[264][12] = (mid_1[2127:2120] < mid_1[2119:2112]) ? 1 : 0;
assign detect_min[264][13] = (mid_1[2127:2120] < mid_1[2135:2128]) ? 1 : 0;
assign detect_min[264][14] = (mid_1[2127:2120] < mid_2[2119:2112]) ? 1 : 0;
assign detect_min[264][15] = (mid_1[2127:2120] < mid_2[2127:2120]) ? 1 : 0;
assign detect_min[264][16] = (mid_1[2127:2120] < mid_2[2135:2128]) ? 1 : 0;
assign detect_min[264][17] = (mid_1[2127:2120] < btm_0[2119:2112]) ? 1 : 0;
assign detect_min[264][18] = (mid_1[2127:2120] < btm_0[2127:2120]) ? 1 : 0;
assign detect_min[264][19] = (mid_1[2127:2120] < btm_0[2135:2128]) ? 1 : 0;
assign detect_min[264][20] = (mid_1[2127:2120] < btm_1[2119:2112]) ? 1 : 0;
assign detect_min[264][21] = (mid_1[2127:2120] < btm_1[2127:2120]) ? 1 : 0;
assign detect_min[264][22] = (mid_1[2127:2120] < btm_1[2135:2128]) ? 1 : 0;
assign detect_min[264][23] = (mid_1[2127:2120] < btm_2[2119:2112]) ? 1 : 0;
assign detect_min[264][24] = (mid_1[2127:2120] < btm_2[2127:2120]) ? 1 : 0;
assign detect_min[264][25] = (mid_1[2127:2120] < btm_2[2135:2128]) ? 1 : 0;

assign detect_min[265][0] = (mid_1[2135:2128] < top_0[2127:2120]) ? 1 : 0;
assign detect_min[265][1] = (mid_1[2135:2128] < top_0[2135:2128]) ? 1 : 0;
assign detect_min[265][2] = (mid_1[2135:2128] < top_0[2143:2136]) ? 1 : 0;
assign detect_min[265][3] = (mid_1[2135:2128] < top_1[2127:2120]) ? 1 : 0;
assign detect_min[265][4] = (mid_1[2135:2128] < top_1[2135:2128]) ? 1 : 0;
assign detect_min[265][5] = (mid_1[2135:2128] < top_1[2143:2136]) ? 1 : 0;
assign detect_min[265][6] = (mid_1[2135:2128] < top_2[2127:2120]) ? 1 : 0;
assign detect_min[265][7] = (mid_1[2135:2128] < top_2[2135:2128]) ? 1 : 0;
assign detect_min[265][8] = (mid_1[2135:2128] < top_2[2143:2136]) ? 1 : 0;
assign detect_min[265][9] = (mid_1[2135:2128] < mid_0[2127:2120]) ? 1 : 0;
assign detect_min[265][10] = (mid_1[2135:2128] < mid_0[2135:2128]) ? 1 : 0;
assign detect_min[265][11] = (mid_1[2135:2128] < mid_0[2143:2136]) ? 1 : 0;
assign detect_min[265][12] = (mid_1[2135:2128] < mid_1[2127:2120]) ? 1 : 0;
assign detect_min[265][13] = (mid_1[2135:2128] < mid_1[2143:2136]) ? 1 : 0;
assign detect_min[265][14] = (mid_1[2135:2128] < mid_2[2127:2120]) ? 1 : 0;
assign detect_min[265][15] = (mid_1[2135:2128] < mid_2[2135:2128]) ? 1 : 0;
assign detect_min[265][16] = (mid_1[2135:2128] < mid_2[2143:2136]) ? 1 : 0;
assign detect_min[265][17] = (mid_1[2135:2128] < btm_0[2127:2120]) ? 1 : 0;
assign detect_min[265][18] = (mid_1[2135:2128] < btm_0[2135:2128]) ? 1 : 0;
assign detect_min[265][19] = (mid_1[2135:2128] < btm_0[2143:2136]) ? 1 : 0;
assign detect_min[265][20] = (mid_1[2135:2128] < btm_1[2127:2120]) ? 1 : 0;
assign detect_min[265][21] = (mid_1[2135:2128] < btm_1[2135:2128]) ? 1 : 0;
assign detect_min[265][22] = (mid_1[2135:2128] < btm_1[2143:2136]) ? 1 : 0;
assign detect_min[265][23] = (mid_1[2135:2128] < btm_2[2127:2120]) ? 1 : 0;
assign detect_min[265][24] = (mid_1[2135:2128] < btm_2[2135:2128]) ? 1 : 0;
assign detect_min[265][25] = (mid_1[2135:2128] < btm_2[2143:2136]) ? 1 : 0;

assign detect_min[266][0] = (mid_1[2143:2136] < top_0[2135:2128]) ? 1 : 0;
assign detect_min[266][1] = (mid_1[2143:2136] < top_0[2143:2136]) ? 1 : 0;
assign detect_min[266][2] = (mid_1[2143:2136] < top_0[2151:2144]) ? 1 : 0;
assign detect_min[266][3] = (mid_1[2143:2136] < top_1[2135:2128]) ? 1 : 0;
assign detect_min[266][4] = (mid_1[2143:2136] < top_1[2143:2136]) ? 1 : 0;
assign detect_min[266][5] = (mid_1[2143:2136] < top_1[2151:2144]) ? 1 : 0;
assign detect_min[266][6] = (mid_1[2143:2136] < top_2[2135:2128]) ? 1 : 0;
assign detect_min[266][7] = (mid_1[2143:2136] < top_2[2143:2136]) ? 1 : 0;
assign detect_min[266][8] = (mid_1[2143:2136] < top_2[2151:2144]) ? 1 : 0;
assign detect_min[266][9] = (mid_1[2143:2136] < mid_0[2135:2128]) ? 1 : 0;
assign detect_min[266][10] = (mid_1[2143:2136] < mid_0[2143:2136]) ? 1 : 0;
assign detect_min[266][11] = (mid_1[2143:2136] < mid_0[2151:2144]) ? 1 : 0;
assign detect_min[266][12] = (mid_1[2143:2136] < mid_1[2135:2128]) ? 1 : 0;
assign detect_min[266][13] = (mid_1[2143:2136] < mid_1[2151:2144]) ? 1 : 0;
assign detect_min[266][14] = (mid_1[2143:2136] < mid_2[2135:2128]) ? 1 : 0;
assign detect_min[266][15] = (mid_1[2143:2136] < mid_2[2143:2136]) ? 1 : 0;
assign detect_min[266][16] = (mid_1[2143:2136] < mid_2[2151:2144]) ? 1 : 0;
assign detect_min[266][17] = (mid_1[2143:2136] < btm_0[2135:2128]) ? 1 : 0;
assign detect_min[266][18] = (mid_1[2143:2136] < btm_0[2143:2136]) ? 1 : 0;
assign detect_min[266][19] = (mid_1[2143:2136] < btm_0[2151:2144]) ? 1 : 0;
assign detect_min[266][20] = (mid_1[2143:2136] < btm_1[2135:2128]) ? 1 : 0;
assign detect_min[266][21] = (mid_1[2143:2136] < btm_1[2143:2136]) ? 1 : 0;
assign detect_min[266][22] = (mid_1[2143:2136] < btm_1[2151:2144]) ? 1 : 0;
assign detect_min[266][23] = (mid_1[2143:2136] < btm_2[2135:2128]) ? 1 : 0;
assign detect_min[266][24] = (mid_1[2143:2136] < btm_2[2143:2136]) ? 1 : 0;
assign detect_min[266][25] = (mid_1[2143:2136] < btm_2[2151:2144]) ? 1 : 0;

assign detect_min[267][0] = (mid_1[2151:2144] < top_0[2143:2136]) ? 1 : 0;
assign detect_min[267][1] = (mid_1[2151:2144] < top_0[2151:2144]) ? 1 : 0;
assign detect_min[267][2] = (mid_1[2151:2144] < top_0[2159:2152]) ? 1 : 0;
assign detect_min[267][3] = (mid_1[2151:2144] < top_1[2143:2136]) ? 1 : 0;
assign detect_min[267][4] = (mid_1[2151:2144] < top_1[2151:2144]) ? 1 : 0;
assign detect_min[267][5] = (mid_1[2151:2144] < top_1[2159:2152]) ? 1 : 0;
assign detect_min[267][6] = (mid_1[2151:2144] < top_2[2143:2136]) ? 1 : 0;
assign detect_min[267][7] = (mid_1[2151:2144] < top_2[2151:2144]) ? 1 : 0;
assign detect_min[267][8] = (mid_1[2151:2144] < top_2[2159:2152]) ? 1 : 0;
assign detect_min[267][9] = (mid_1[2151:2144] < mid_0[2143:2136]) ? 1 : 0;
assign detect_min[267][10] = (mid_1[2151:2144] < mid_0[2151:2144]) ? 1 : 0;
assign detect_min[267][11] = (mid_1[2151:2144] < mid_0[2159:2152]) ? 1 : 0;
assign detect_min[267][12] = (mid_1[2151:2144] < mid_1[2143:2136]) ? 1 : 0;
assign detect_min[267][13] = (mid_1[2151:2144] < mid_1[2159:2152]) ? 1 : 0;
assign detect_min[267][14] = (mid_1[2151:2144] < mid_2[2143:2136]) ? 1 : 0;
assign detect_min[267][15] = (mid_1[2151:2144] < mid_2[2151:2144]) ? 1 : 0;
assign detect_min[267][16] = (mid_1[2151:2144] < mid_2[2159:2152]) ? 1 : 0;
assign detect_min[267][17] = (mid_1[2151:2144] < btm_0[2143:2136]) ? 1 : 0;
assign detect_min[267][18] = (mid_1[2151:2144] < btm_0[2151:2144]) ? 1 : 0;
assign detect_min[267][19] = (mid_1[2151:2144] < btm_0[2159:2152]) ? 1 : 0;
assign detect_min[267][20] = (mid_1[2151:2144] < btm_1[2143:2136]) ? 1 : 0;
assign detect_min[267][21] = (mid_1[2151:2144] < btm_1[2151:2144]) ? 1 : 0;
assign detect_min[267][22] = (mid_1[2151:2144] < btm_1[2159:2152]) ? 1 : 0;
assign detect_min[267][23] = (mid_1[2151:2144] < btm_2[2143:2136]) ? 1 : 0;
assign detect_min[267][24] = (mid_1[2151:2144] < btm_2[2151:2144]) ? 1 : 0;
assign detect_min[267][25] = (mid_1[2151:2144] < btm_2[2159:2152]) ? 1 : 0;

assign detect_min[268][0] = (mid_1[2159:2152] < top_0[2151:2144]) ? 1 : 0;
assign detect_min[268][1] = (mid_1[2159:2152] < top_0[2159:2152]) ? 1 : 0;
assign detect_min[268][2] = (mid_1[2159:2152] < top_0[2167:2160]) ? 1 : 0;
assign detect_min[268][3] = (mid_1[2159:2152] < top_1[2151:2144]) ? 1 : 0;
assign detect_min[268][4] = (mid_1[2159:2152] < top_1[2159:2152]) ? 1 : 0;
assign detect_min[268][5] = (mid_1[2159:2152] < top_1[2167:2160]) ? 1 : 0;
assign detect_min[268][6] = (mid_1[2159:2152] < top_2[2151:2144]) ? 1 : 0;
assign detect_min[268][7] = (mid_1[2159:2152] < top_2[2159:2152]) ? 1 : 0;
assign detect_min[268][8] = (mid_1[2159:2152] < top_2[2167:2160]) ? 1 : 0;
assign detect_min[268][9] = (mid_1[2159:2152] < mid_0[2151:2144]) ? 1 : 0;
assign detect_min[268][10] = (mid_1[2159:2152] < mid_0[2159:2152]) ? 1 : 0;
assign detect_min[268][11] = (mid_1[2159:2152] < mid_0[2167:2160]) ? 1 : 0;
assign detect_min[268][12] = (mid_1[2159:2152] < mid_1[2151:2144]) ? 1 : 0;
assign detect_min[268][13] = (mid_1[2159:2152] < mid_1[2167:2160]) ? 1 : 0;
assign detect_min[268][14] = (mid_1[2159:2152] < mid_2[2151:2144]) ? 1 : 0;
assign detect_min[268][15] = (mid_1[2159:2152] < mid_2[2159:2152]) ? 1 : 0;
assign detect_min[268][16] = (mid_1[2159:2152] < mid_2[2167:2160]) ? 1 : 0;
assign detect_min[268][17] = (mid_1[2159:2152] < btm_0[2151:2144]) ? 1 : 0;
assign detect_min[268][18] = (mid_1[2159:2152] < btm_0[2159:2152]) ? 1 : 0;
assign detect_min[268][19] = (mid_1[2159:2152] < btm_0[2167:2160]) ? 1 : 0;
assign detect_min[268][20] = (mid_1[2159:2152] < btm_1[2151:2144]) ? 1 : 0;
assign detect_min[268][21] = (mid_1[2159:2152] < btm_1[2159:2152]) ? 1 : 0;
assign detect_min[268][22] = (mid_1[2159:2152] < btm_1[2167:2160]) ? 1 : 0;
assign detect_min[268][23] = (mid_1[2159:2152] < btm_2[2151:2144]) ? 1 : 0;
assign detect_min[268][24] = (mid_1[2159:2152] < btm_2[2159:2152]) ? 1 : 0;
assign detect_min[268][25] = (mid_1[2159:2152] < btm_2[2167:2160]) ? 1 : 0;

assign detect_min[269][0] = (mid_1[2167:2160] < top_0[2159:2152]) ? 1 : 0;
assign detect_min[269][1] = (mid_1[2167:2160] < top_0[2167:2160]) ? 1 : 0;
assign detect_min[269][2] = (mid_1[2167:2160] < top_0[2175:2168]) ? 1 : 0;
assign detect_min[269][3] = (mid_1[2167:2160] < top_1[2159:2152]) ? 1 : 0;
assign detect_min[269][4] = (mid_1[2167:2160] < top_1[2167:2160]) ? 1 : 0;
assign detect_min[269][5] = (mid_1[2167:2160] < top_1[2175:2168]) ? 1 : 0;
assign detect_min[269][6] = (mid_1[2167:2160] < top_2[2159:2152]) ? 1 : 0;
assign detect_min[269][7] = (mid_1[2167:2160] < top_2[2167:2160]) ? 1 : 0;
assign detect_min[269][8] = (mid_1[2167:2160] < top_2[2175:2168]) ? 1 : 0;
assign detect_min[269][9] = (mid_1[2167:2160] < mid_0[2159:2152]) ? 1 : 0;
assign detect_min[269][10] = (mid_1[2167:2160] < mid_0[2167:2160]) ? 1 : 0;
assign detect_min[269][11] = (mid_1[2167:2160] < mid_0[2175:2168]) ? 1 : 0;
assign detect_min[269][12] = (mid_1[2167:2160] < mid_1[2159:2152]) ? 1 : 0;
assign detect_min[269][13] = (mid_1[2167:2160] < mid_1[2175:2168]) ? 1 : 0;
assign detect_min[269][14] = (mid_1[2167:2160] < mid_2[2159:2152]) ? 1 : 0;
assign detect_min[269][15] = (mid_1[2167:2160] < mid_2[2167:2160]) ? 1 : 0;
assign detect_min[269][16] = (mid_1[2167:2160] < mid_2[2175:2168]) ? 1 : 0;
assign detect_min[269][17] = (mid_1[2167:2160] < btm_0[2159:2152]) ? 1 : 0;
assign detect_min[269][18] = (mid_1[2167:2160] < btm_0[2167:2160]) ? 1 : 0;
assign detect_min[269][19] = (mid_1[2167:2160] < btm_0[2175:2168]) ? 1 : 0;
assign detect_min[269][20] = (mid_1[2167:2160] < btm_1[2159:2152]) ? 1 : 0;
assign detect_min[269][21] = (mid_1[2167:2160] < btm_1[2167:2160]) ? 1 : 0;
assign detect_min[269][22] = (mid_1[2167:2160] < btm_1[2175:2168]) ? 1 : 0;
assign detect_min[269][23] = (mid_1[2167:2160] < btm_2[2159:2152]) ? 1 : 0;
assign detect_min[269][24] = (mid_1[2167:2160] < btm_2[2167:2160]) ? 1 : 0;
assign detect_min[269][25] = (mid_1[2167:2160] < btm_2[2175:2168]) ? 1 : 0;

assign detect_min[270][0] = (mid_1[2175:2168] < top_0[2167:2160]) ? 1 : 0;
assign detect_min[270][1] = (mid_1[2175:2168] < top_0[2175:2168]) ? 1 : 0;
assign detect_min[270][2] = (mid_1[2175:2168] < top_0[2183:2176]) ? 1 : 0;
assign detect_min[270][3] = (mid_1[2175:2168] < top_1[2167:2160]) ? 1 : 0;
assign detect_min[270][4] = (mid_1[2175:2168] < top_1[2175:2168]) ? 1 : 0;
assign detect_min[270][5] = (mid_1[2175:2168] < top_1[2183:2176]) ? 1 : 0;
assign detect_min[270][6] = (mid_1[2175:2168] < top_2[2167:2160]) ? 1 : 0;
assign detect_min[270][7] = (mid_1[2175:2168] < top_2[2175:2168]) ? 1 : 0;
assign detect_min[270][8] = (mid_1[2175:2168] < top_2[2183:2176]) ? 1 : 0;
assign detect_min[270][9] = (mid_1[2175:2168] < mid_0[2167:2160]) ? 1 : 0;
assign detect_min[270][10] = (mid_1[2175:2168] < mid_0[2175:2168]) ? 1 : 0;
assign detect_min[270][11] = (mid_1[2175:2168] < mid_0[2183:2176]) ? 1 : 0;
assign detect_min[270][12] = (mid_1[2175:2168] < mid_1[2167:2160]) ? 1 : 0;
assign detect_min[270][13] = (mid_1[2175:2168] < mid_1[2183:2176]) ? 1 : 0;
assign detect_min[270][14] = (mid_1[2175:2168] < mid_2[2167:2160]) ? 1 : 0;
assign detect_min[270][15] = (mid_1[2175:2168] < mid_2[2175:2168]) ? 1 : 0;
assign detect_min[270][16] = (mid_1[2175:2168] < mid_2[2183:2176]) ? 1 : 0;
assign detect_min[270][17] = (mid_1[2175:2168] < btm_0[2167:2160]) ? 1 : 0;
assign detect_min[270][18] = (mid_1[2175:2168] < btm_0[2175:2168]) ? 1 : 0;
assign detect_min[270][19] = (mid_1[2175:2168] < btm_0[2183:2176]) ? 1 : 0;
assign detect_min[270][20] = (mid_1[2175:2168] < btm_1[2167:2160]) ? 1 : 0;
assign detect_min[270][21] = (mid_1[2175:2168] < btm_1[2175:2168]) ? 1 : 0;
assign detect_min[270][22] = (mid_1[2175:2168] < btm_1[2183:2176]) ? 1 : 0;
assign detect_min[270][23] = (mid_1[2175:2168] < btm_2[2167:2160]) ? 1 : 0;
assign detect_min[270][24] = (mid_1[2175:2168] < btm_2[2175:2168]) ? 1 : 0;
assign detect_min[270][25] = (mid_1[2175:2168] < btm_2[2183:2176]) ? 1 : 0;

assign detect_min[271][0] = (mid_1[2183:2176] < top_0[2175:2168]) ? 1 : 0;
assign detect_min[271][1] = (mid_1[2183:2176] < top_0[2183:2176]) ? 1 : 0;
assign detect_min[271][2] = (mid_1[2183:2176] < top_0[2191:2184]) ? 1 : 0;
assign detect_min[271][3] = (mid_1[2183:2176] < top_1[2175:2168]) ? 1 : 0;
assign detect_min[271][4] = (mid_1[2183:2176] < top_1[2183:2176]) ? 1 : 0;
assign detect_min[271][5] = (mid_1[2183:2176] < top_1[2191:2184]) ? 1 : 0;
assign detect_min[271][6] = (mid_1[2183:2176] < top_2[2175:2168]) ? 1 : 0;
assign detect_min[271][7] = (mid_1[2183:2176] < top_2[2183:2176]) ? 1 : 0;
assign detect_min[271][8] = (mid_1[2183:2176] < top_2[2191:2184]) ? 1 : 0;
assign detect_min[271][9] = (mid_1[2183:2176] < mid_0[2175:2168]) ? 1 : 0;
assign detect_min[271][10] = (mid_1[2183:2176] < mid_0[2183:2176]) ? 1 : 0;
assign detect_min[271][11] = (mid_1[2183:2176] < mid_0[2191:2184]) ? 1 : 0;
assign detect_min[271][12] = (mid_1[2183:2176] < mid_1[2175:2168]) ? 1 : 0;
assign detect_min[271][13] = (mid_1[2183:2176] < mid_1[2191:2184]) ? 1 : 0;
assign detect_min[271][14] = (mid_1[2183:2176] < mid_2[2175:2168]) ? 1 : 0;
assign detect_min[271][15] = (mid_1[2183:2176] < mid_2[2183:2176]) ? 1 : 0;
assign detect_min[271][16] = (mid_1[2183:2176] < mid_2[2191:2184]) ? 1 : 0;
assign detect_min[271][17] = (mid_1[2183:2176] < btm_0[2175:2168]) ? 1 : 0;
assign detect_min[271][18] = (mid_1[2183:2176] < btm_0[2183:2176]) ? 1 : 0;
assign detect_min[271][19] = (mid_1[2183:2176] < btm_0[2191:2184]) ? 1 : 0;
assign detect_min[271][20] = (mid_1[2183:2176] < btm_1[2175:2168]) ? 1 : 0;
assign detect_min[271][21] = (mid_1[2183:2176] < btm_1[2183:2176]) ? 1 : 0;
assign detect_min[271][22] = (mid_1[2183:2176] < btm_1[2191:2184]) ? 1 : 0;
assign detect_min[271][23] = (mid_1[2183:2176] < btm_2[2175:2168]) ? 1 : 0;
assign detect_min[271][24] = (mid_1[2183:2176] < btm_2[2183:2176]) ? 1 : 0;
assign detect_min[271][25] = (mid_1[2183:2176] < btm_2[2191:2184]) ? 1 : 0;

assign detect_min[272][0] = (mid_1[2191:2184] < top_0[2183:2176]) ? 1 : 0;
assign detect_min[272][1] = (mid_1[2191:2184] < top_0[2191:2184]) ? 1 : 0;
assign detect_min[272][2] = (mid_1[2191:2184] < top_0[2199:2192]) ? 1 : 0;
assign detect_min[272][3] = (mid_1[2191:2184] < top_1[2183:2176]) ? 1 : 0;
assign detect_min[272][4] = (mid_1[2191:2184] < top_1[2191:2184]) ? 1 : 0;
assign detect_min[272][5] = (mid_1[2191:2184] < top_1[2199:2192]) ? 1 : 0;
assign detect_min[272][6] = (mid_1[2191:2184] < top_2[2183:2176]) ? 1 : 0;
assign detect_min[272][7] = (mid_1[2191:2184] < top_2[2191:2184]) ? 1 : 0;
assign detect_min[272][8] = (mid_1[2191:2184] < top_2[2199:2192]) ? 1 : 0;
assign detect_min[272][9] = (mid_1[2191:2184] < mid_0[2183:2176]) ? 1 : 0;
assign detect_min[272][10] = (mid_1[2191:2184] < mid_0[2191:2184]) ? 1 : 0;
assign detect_min[272][11] = (mid_1[2191:2184] < mid_0[2199:2192]) ? 1 : 0;
assign detect_min[272][12] = (mid_1[2191:2184] < mid_1[2183:2176]) ? 1 : 0;
assign detect_min[272][13] = (mid_1[2191:2184] < mid_1[2199:2192]) ? 1 : 0;
assign detect_min[272][14] = (mid_1[2191:2184] < mid_2[2183:2176]) ? 1 : 0;
assign detect_min[272][15] = (mid_1[2191:2184] < mid_2[2191:2184]) ? 1 : 0;
assign detect_min[272][16] = (mid_1[2191:2184] < mid_2[2199:2192]) ? 1 : 0;
assign detect_min[272][17] = (mid_1[2191:2184] < btm_0[2183:2176]) ? 1 : 0;
assign detect_min[272][18] = (mid_1[2191:2184] < btm_0[2191:2184]) ? 1 : 0;
assign detect_min[272][19] = (mid_1[2191:2184] < btm_0[2199:2192]) ? 1 : 0;
assign detect_min[272][20] = (mid_1[2191:2184] < btm_1[2183:2176]) ? 1 : 0;
assign detect_min[272][21] = (mid_1[2191:2184] < btm_1[2191:2184]) ? 1 : 0;
assign detect_min[272][22] = (mid_1[2191:2184] < btm_1[2199:2192]) ? 1 : 0;
assign detect_min[272][23] = (mid_1[2191:2184] < btm_2[2183:2176]) ? 1 : 0;
assign detect_min[272][24] = (mid_1[2191:2184] < btm_2[2191:2184]) ? 1 : 0;
assign detect_min[272][25] = (mid_1[2191:2184] < btm_2[2199:2192]) ? 1 : 0;

assign detect_min[273][0] = (mid_1[2199:2192] < top_0[2191:2184]) ? 1 : 0;
assign detect_min[273][1] = (mid_1[2199:2192] < top_0[2199:2192]) ? 1 : 0;
assign detect_min[273][2] = (mid_1[2199:2192] < top_0[2207:2200]) ? 1 : 0;
assign detect_min[273][3] = (mid_1[2199:2192] < top_1[2191:2184]) ? 1 : 0;
assign detect_min[273][4] = (mid_1[2199:2192] < top_1[2199:2192]) ? 1 : 0;
assign detect_min[273][5] = (mid_1[2199:2192] < top_1[2207:2200]) ? 1 : 0;
assign detect_min[273][6] = (mid_1[2199:2192] < top_2[2191:2184]) ? 1 : 0;
assign detect_min[273][7] = (mid_1[2199:2192] < top_2[2199:2192]) ? 1 : 0;
assign detect_min[273][8] = (mid_1[2199:2192] < top_2[2207:2200]) ? 1 : 0;
assign detect_min[273][9] = (mid_1[2199:2192] < mid_0[2191:2184]) ? 1 : 0;
assign detect_min[273][10] = (mid_1[2199:2192] < mid_0[2199:2192]) ? 1 : 0;
assign detect_min[273][11] = (mid_1[2199:2192] < mid_0[2207:2200]) ? 1 : 0;
assign detect_min[273][12] = (mid_1[2199:2192] < mid_1[2191:2184]) ? 1 : 0;
assign detect_min[273][13] = (mid_1[2199:2192] < mid_1[2207:2200]) ? 1 : 0;
assign detect_min[273][14] = (mid_1[2199:2192] < mid_2[2191:2184]) ? 1 : 0;
assign detect_min[273][15] = (mid_1[2199:2192] < mid_2[2199:2192]) ? 1 : 0;
assign detect_min[273][16] = (mid_1[2199:2192] < mid_2[2207:2200]) ? 1 : 0;
assign detect_min[273][17] = (mid_1[2199:2192] < btm_0[2191:2184]) ? 1 : 0;
assign detect_min[273][18] = (mid_1[2199:2192] < btm_0[2199:2192]) ? 1 : 0;
assign detect_min[273][19] = (mid_1[2199:2192] < btm_0[2207:2200]) ? 1 : 0;
assign detect_min[273][20] = (mid_1[2199:2192] < btm_1[2191:2184]) ? 1 : 0;
assign detect_min[273][21] = (mid_1[2199:2192] < btm_1[2199:2192]) ? 1 : 0;
assign detect_min[273][22] = (mid_1[2199:2192] < btm_1[2207:2200]) ? 1 : 0;
assign detect_min[273][23] = (mid_1[2199:2192] < btm_2[2191:2184]) ? 1 : 0;
assign detect_min[273][24] = (mid_1[2199:2192] < btm_2[2199:2192]) ? 1 : 0;
assign detect_min[273][25] = (mid_1[2199:2192] < btm_2[2207:2200]) ? 1 : 0;

assign detect_min[274][0] = (mid_1[2207:2200] < top_0[2199:2192]) ? 1 : 0;
assign detect_min[274][1] = (mid_1[2207:2200] < top_0[2207:2200]) ? 1 : 0;
assign detect_min[274][2] = (mid_1[2207:2200] < top_0[2215:2208]) ? 1 : 0;
assign detect_min[274][3] = (mid_1[2207:2200] < top_1[2199:2192]) ? 1 : 0;
assign detect_min[274][4] = (mid_1[2207:2200] < top_1[2207:2200]) ? 1 : 0;
assign detect_min[274][5] = (mid_1[2207:2200] < top_1[2215:2208]) ? 1 : 0;
assign detect_min[274][6] = (mid_1[2207:2200] < top_2[2199:2192]) ? 1 : 0;
assign detect_min[274][7] = (mid_1[2207:2200] < top_2[2207:2200]) ? 1 : 0;
assign detect_min[274][8] = (mid_1[2207:2200] < top_2[2215:2208]) ? 1 : 0;
assign detect_min[274][9] = (mid_1[2207:2200] < mid_0[2199:2192]) ? 1 : 0;
assign detect_min[274][10] = (mid_1[2207:2200] < mid_0[2207:2200]) ? 1 : 0;
assign detect_min[274][11] = (mid_1[2207:2200] < mid_0[2215:2208]) ? 1 : 0;
assign detect_min[274][12] = (mid_1[2207:2200] < mid_1[2199:2192]) ? 1 : 0;
assign detect_min[274][13] = (mid_1[2207:2200] < mid_1[2215:2208]) ? 1 : 0;
assign detect_min[274][14] = (mid_1[2207:2200] < mid_2[2199:2192]) ? 1 : 0;
assign detect_min[274][15] = (mid_1[2207:2200] < mid_2[2207:2200]) ? 1 : 0;
assign detect_min[274][16] = (mid_1[2207:2200] < mid_2[2215:2208]) ? 1 : 0;
assign detect_min[274][17] = (mid_1[2207:2200] < btm_0[2199:2192]) ? 1 : 0;
assign detect_min[274][18] = (mid_1[2207:2200] < btm_0[2207:2200]) ? 1 : 0;
assign detect_min[274][19] = (mid_1[2207:2200] < btm_0[2215:2208]) ? 1 : 0;
assign detect_min[274][20] = (mid_1[2207:2200] < btm_1[2199:2192]) ? 1 : 0;
assign detect_min[274][21] = (mid_1[2207:2200] < btm_1[2207:2200]) ? 1 : 0;
assign detect_min[274][22] = (mid_1[2207:2200] < btm_1[2215:2208]) ? 1 : 0;
assign detect_min[274][23] = (mid_1[2207:2200] < btm_2[2199:2192]) ? 1 : 0;
assign detect_min[274][24] = (mid_1[2207:2200] < btm_2[2207:2200]) ? 1 : 0;
assign detect_min[274][25] = (mid_1[2207:2200] < btm_2[2215:2208]) ? 1 : 0;

assign detect_min[275][0] = (mid_1[2215:2208] < top_0[2207:2200]) ? 1 : 0;
assign detect_min[275][1] = (mid_1[2215:2208] < top_0[2215:2208]) ? 1 : 0;
assign detect_min[275][2] = (mid_1[2215:2208] < top_0[2223:2216]) ? 1 : 0;
assign detect_min[275][3] = (mid_1[2215:2208] < top_1[2207:2200]) ? 1 : 0;
assign detect_min[275][4] = (mid_1[2215:2208] < top_1[2215:2208]) ? 1 : 0;
assign detect_min[275][5] = (mid_1[2215:2208] < top_1[2223:2216]) ? 1 : 0;
assign detect_min[275][6] = (mid_1[2215:2208] < top_2[2207:2200]) ? 1 : 0;
assign detect_min[275][7] = (mid_1[2215:2208] < top_2[2215:2208]) ? 1 : 0;
assign detect_min[275][8] = (mid_1[2215:2208] < top_2[2223:2216]) ? 1 : 0;
assign detect_min[275][9] = (mid_1[2215:2208] < mid_0[2207:2200]) ? 1 : 0;
assign detect_min[275][10] = (mid_1[2215:2208] < mid_0[2215:2208]) ? 1 : 0;
assign detect_min[275][11] = (mid_1[2215:2208] < mid_0[2223:2216]) ? 1 : 0;
assign detect_min[275][12] = (mid_1[2215:2208] < mid_1[2207:2200]) ? 1 : 0;
assign detect_min[275][13] = (mid_1[2215:2208] < mid_1[2223:2216]) ? 1 : 0;
assign detect_min[275][14] = (mid_1[2215:2208] < mid_2[2207:2200]) ? 1 : 0;
assign detect_min[275][15] = (mid_1[2215:2208] < mid_2[2215:2208]) ? 1 : 0;
assign detect_min[275][16] = (mid_1[2215:2208] < mid_2[2223:2216]) ? 1 : 0;
assign detect_min[275][17] = (mid_1[2215:2208] < btm_0[2207:2200]) ? 1 : 0;
assign detect_min[275][18] = (mid_1[2215:2208] < btm_0[2215:2208]) ? 1 : 0;
assign detect_min[275][19] = (mid_1[2215:2208] < btm_0[2223:2216]) ? 1 : 0;
assign detect_min[275][20] = (mid_1[2215:2208] < btm_1[2207:2200]) ? 1 : 0;
assign detect_min[275][21] = (mid_1[2215:2208] < btm_1[2215:2208]) ? 1 : 0;
assign detect_min[275][22] = (mid_1[2215:2208] < btm_1[2223:2216]) ? 1 : 0;
assign detect_min[275][23] = (mid_1[2215:2208] < btm_2[2207:2200]) ? 1 : 0;
assign detect_min[275][24] = (mid_1[2215:2208] < btm_2[2215:2208]) ? 1 : 0;
assign detect_min[275][25] = (mid_1[2215:2208] < btm_2[2223:2216]) ? 1 : 0;

assign detect_min[276][0] = (mid_1[2223:2216] < top_0[2215:2208]) ? 1 : 0;
assign detect_min[276][1] = (mid_1[2223:2216] < top_0[2223:2216]) ? 1 : 0;
assign detect_min[276][2] = (mid_1[2223:2216] < top_0[2231:2224]) ? 1 : 0;
assign detect_min[276][3] = (mid_1[2223:2216] < top_1[2215:2208]) ? 1 : 0;
assign detect_min[276][4] = (mid_1[2223:2216] < top_1[2223:2216]) ? 1 : 0;
assign detect_min[276][5] = (mid_1[2223:2216] < top_1[2231:2224]) ? 1 : 0;
assign detect_min[276][6] = (mid_1[2223:2216] < top_2[2215:2208]) ? 1 : 0;
assign detect_min[276][7] = (mid_1[2223:2216] < top_2[2223:2216]) ? 1 : 0;
assign detect_min[276][8] = (mid_1[2223:2216] < top_2[2231:2224]) ? 1 : 0;
assign detect_min[276][9] = (mid_1[2223:2216] < mid_0[2215:2208]) ? 1 : 0;
assign detect_min[276][10] = (mid_1[2223:2216] < mid_0[2223:2216]) ? 1 : 0;
assign detect_min[276][11] = (mid_1[2223:2216] < mid_0[2231:2224]) ? 1 : 0;
assign detect_min[276][12] = (mid_1[2223:2216] < mid_1[2215:2208]) ? 1 : 0;
assign detect_min[276][13] = (mid_1[2223:2216] < mid_1[2231:2224]) ? 1 : 0;
assign detect_min[276][14] = (mid_1[2223:2216] < mid_2[2215:2208]) ? 1 : 0;
assign detect_min[276][15] = (mid_1[2223:2216] < mid_2[2223:2216]) ? 1 : 0;
assign detect_min[276][16] = (mid_1[2223:2216] < mid_2[2231:2224]) ? 1 : 0;
assign detect_min[276][17] = (mid_1[2223:2216] < btm_0[2215:2208]) ? 1 : 0;
assign detect_min[276][18] = (mid_1[2223:2216] < btm_0[2223:2216]) ? 1 : 0;
assign detect_min[276][19] = (mid_1[2223:2216] < btm_0[2231:2224]) ? 1 : 0;
assign detect_min[276][20] = (mid_1[2223:2216] < btm_1[2215:2208]) ? 1 : 0;
assign detect_min[276][21] = (mid_1[2223:2216] < btm_1[2223:2216]) ? 1 : 0;
assign detect_min[276][22] = (mid_1[2223:2216] < btm_1[2231:2224]) ? 1 : 0;
assign detect_min[276][23] = (mid_1[2223:2216] < btm_2[2215:2208]) ? 1 : 0;
assign detect_min[276][24] = (mid_1[2223:2216] < btm_2[2223:2216]) ? 1 : 0;
assign detect_min[276][25] = (mid_1[2223:2216] < btm_2[2231:2224]) ? 1 : 0;

assign detect_min[277][0] = (mid_1[2231:2224] < top_0[2223:2216]) ? 1 : 0;
assign detect_min[277][1] = (mid_1[2231:2224] < top_0[2231:2224]) ? 1 : 0;
assign detect_min[277][2] = (mid_1[2231:2224] < top_0[2239:2232]) ? 1 : 0;
assign detect_min[277][3] = (mid_1[2231:2224] < top_1[2223:2216]) ? 1 : 0;
assign detect_min[277][4] = (mid_1[2231:2224] < top_1[2231:2224]) ? 1 : 0;
assign detect_min[277][5] = (mid_1[2231:2224] < top_1[2239:2232]) ? 1 : 0;
assign detect_min[277][6] = (mid_1[2231:2224] < top_2[2223:2216]) ? 1 : 0;
assign detect_min[277][7] = (mid_1[2231:2224] < top_2[2231:2224]) ? 1 : 0;
assign detect_min[277][8] = (mid_1[2231:2224] < top_2[2239:2232]) ? 1 : 0;
assign detect_min[277][9] = (mid_1[2231:2224] < mid_0[2223:2216]) ? 1 : 0;
assign detect_min[277][10] = (mid_1[2231:2224] < mid_0[2231:2224]) ? 1 : 0;
assign detect_min[277][11] = (mid_1[2231:2224] < mid_0[2239:2232]) ? 1 : 0;
assign detect_min[277][12] = (mid_1[2231:2224] < mid_1[2223:2216]) ? 1 : 0;
assign detect_min[277][13] = (mid_1[2231:2224] < mid_1[2239:2232]) ? 1 : 0;
assign detect_min[277][14] = (mid_1[2231:2224] < mid_2[2223:2216]) ? 1 : 0;
assign detect_min[277][15] = (mid_1[2231:2224] < mid_2[2231:2224]) ? 1 : 0;
assign detect_min[277][16] = (mid_1[2231:2224] < mid_2[2239:2232]) ? 1 : 0;
assign detect_min[277][17] = (mid_1[2231:2224] < btm_0[2223:2216]) ? 1 : 0;
assign detect_min[277][18] = (mid_1[2231:2224] < btm_0[2231:2224]) ? 1 : 0;
assign detect_min[277][19] = (mid_1[2231:2224] < btm_0[2239:2232]) ? 1 : 0;
assign detect_min[277][20] = (mid_1[2231:2224] < btm_1[2223:2216]) ? 1 : 0;
assign detect_min[277][21] = (mid_1[2231:2224] < btm_1[2231:2224]) ? 1 : 0;
assign detect_min[277][22] = (mid_1[2231:2224] < btm_1[2239:2232]) ? 1 : 0;
assign detect_min[277][23] = (mid_1[2231:2224] < btm_2[2223:2216]) ? 1 : 0;
assign detect_min[277][24] = (mid_1[2231:2224] < btm_2[2231:2224]) ? 1 : 0;
assign detect_min[277][25] = (mid_1[2231:2224] < btm_2[2239:2232]) ? 1 : 0;

assign detect_min[278][0] = (mid_1[2239:2232] < top_0[2231:2224]) ? 1 : 0;
assign detect_min[278][1] = (mid_1[2239:2232] < top_0[2239:2232]) ? 1 : 0;
assign detect_min[278][2] = (mid_1[2239:2232] < top_0[2247:2240]) ? 1 : 0;
assign detect_min[278][3] = (mid_1[2239:2232] < top_1[2231:2224]) ? 1 : 0;
assign detect_min[278][4] = (mid_1[2239:2232] < top_1[2239:2232]) ? 1 : 0;
assign detect_min[278][5] = (mid_1[2239:2232] < top_1[2247:2240]) ? 1 : 0;
assign detect_min[278][6] = (mid_1[2239:2232] < top_2[2231:2224]) ? 1 : 0;
assign detect_min[278][7] = (mid_1[2239:2232] < top_2[2239:2232]) ? 1 : 0;
assign detect_min[278][8] = (mid_1[2239:2232] < top_2[2247:2240]) ? 1 : 0;
assign detect_min[278][9] = (mid_1[2239:2232] < mid_0[2231:2224]) ? 1 : 0;
assign detect_min[278][10] = (mid_1[2239:2232] < mid_0[2239:2232]) ? 1 : 0;
assign detect_min[278][11] = (mid_1[2239:2232] < mid_0[2247:2240]) ? 1 : 0;
assign detect_min[278][12] = (mid_1[2239:2232] < mid_1[2231:2224]) ? 1 : 0;
assign detect_min[278][13] = (mid_1[2239:2232] < mid_1[2247:2240]) ? 1 : 0;
assign detect_min[278][14] = (mid_1[2239:2232] < mid_2[2231:2224]) ? 1 : 0;
assign detect_min[278][15] = (mid_1[2239:2232] < mid_2[2239:2232]) ? 1 : 0;
assign detect_min[278][16] = (mid_1[2239:2232] < mid_2[2247:2240]) ? 1 : 0;
assign detect_min[278][17] = (mid_1[2239:2232] < btm_0[2231:2224]) ? 1 : 0;
assign detect_min[278][18] = (mid_1[2239:2232] < btm_0[2239:2232]) ? 1 : 0;
assign detect_min[278][19] = (mid_1[2239:2232] < btm_0[2247:2240]) ? 1 : 0;
assign detect_min[278][20] = (mid_1[2239:2232] < btm_1[2231:2224]) ? 1 : 0;
assign detect_min[278][21] = (mid_1[2239:2232] < btm_1[2239:2232]) ? 1 : 0;
assign detect_min[278][22] = (mid_1[2239:2232] < btm_1[2247:2240]) ? 1 : 0;
assign detect_min[278][23] = (mid_1[2239:2232] < btm_2[2231:2224]) ? 1 : 0;
assign detect_min[278][24] = (mid_1[2239:2232] < btm_2[2239:2232]) ? 1 : 0;
assign detect_min[278][25] = (mid_1[2239:2232] < btm_2[2247:2240]) ? 1 : 0;

assign detect_min[279][0] = (mid_1[2247:2240] < top_0[2239:2232]) ? 1 : 0;
assign detect_min[279][1] = (mid_1[2247:2240] < top_0[2247:2240]) ? 1 : 0;
assign detect_min[279][2] = (mid_1[2247:2240] < top_0[2255:2248]) ? 1 : 0;
assign detect_min[279][3] = (mid_1[2247:2240] < top_1[2239:2232]) ? 1 : 0;
assign detect_min[279][4] = (mid_1[2247:2240] < top_1[2247:2240]) ? 1 : 0;
assign detect_min[279][5] = (mid_1[2247:2240] < top_1[2255:2248]) ? 1 : 0;
assign detect_min[279][6] = (mid_1[2247:2240] < top_2[2239:2232]) ? 1 : 0;
assign detect_min[279][7] = (mid_1[2247:2240] < top_2[2247:2240]) ? 1 : 0;
assign detect_min[279][8] = (mid_1[2247:2240] < top_2[2255:2248]) ? 1 : 0;
assign detect_min[279][9] = (mid_1[2247:2240] < mid_0[2239:2232]) ? 1 : 0;
assign detect_min[279][10] = (mid_1[2247:2240] < mid_0[2247:2240]) ? 1 : 0;
assign detect_min[279][11] = (mid_1[2247:2240] < mid_0[2255:2248]) ? 1 : 0;
assign detect_min[279][12] = (mid_1[2247:2240] < mid_1[2239:2232]) ? 1 : 0;
assign detect_min[279][13] = (mid_1[2247:2240] < mid_1[2255:2248]) ? 1 : 0;
assign detect_min[279][14] = (mid_1[2247:2240] < mid_2[2239:2232]) ? 1 : 0;
assign detect_min[279][15] = (mid_1[2247:2240] < mid_2[2247:2240]) ? 1 : 0;
assign detect_min[279][16] = (mid_1[2247:2240] < mid_2[2255:2248]) ? 1 : 0;
assign detect_min[279][17] = (mid_1[2247:2240] < btm_0[2239:2232]) ? 1 : 0;
assign detect_min[279][18] = (mid_1[2247:2240] < btm_0[2247:2240]) ? 1 : 0;
assign detect_min[279][19] = (mid_1[2247:2240] < btm_0[2255:2248]) ? 1 : 0;
assign detect_min[279][20] = (mid_1[2247:2240] < btm_1[2239:2232]) ? 1 : 0;
assign detect_min[279][21] = (mid_1[2247:2240] < btm_1[2247:2240]) ? 1 : 0;
assign detect_min[279][22] = (mid_1[2247:2240] < btm_1[2255:2248]) ? 1 : 0;
assign detect_min[279][23] = (mid_1[2247:2240] < btm_2[2239:2232]) ? 1 : 0;
assign detect_min[279][24] = (mid_1[2247:2240] < btm_2[2247:2240]) ? 1 : 0;
assign detect_min[279][25] = (mid_1[2247:2240] < btm_2[2255:2248]) ? 1 : 0;

assign detect_min[280][0] = (mid_1[2255:2248] < top_0[2247:2240]) ? 1 : 0;
assign detect_min[280][1] = (mid_1[2255:2248] < top_0[2255:2248]) ? 1 : 0;
assign detect_min[280][2] = (mid_1[2255:2248] < top_0[2263:2256]) ? 1 : 0;
assign detect_min[280][3] = (mid_1[2255:2248] < top_1[2247:2240]) ? 1 : 0;
assign detect_min[280][4] = (mid_1[2255:2248] < top_1[2255:2248]) ? 1 : 0;
assign detect_min[280][5] = (mid_1[2255:2248] < top_1[2263:2256]) ? 1 : 0;
assign detect_min[280][6] = (mid_1[2255:2248] < top_2[2247:2240]) ? 1 : 0;
assign detect_min[280][7] = (mid_1[2255:2248] < top_2[2255:2248]) ? 1 : 0;
assign detect_min[280][8] = (mid_1[2255:2248] < top_2[2263:2256]) ? 1 : 0;
assign detect_min[280][9] = (mid_1[2255:2248] < mid_0[2247:2240]) ? 1 : 0;
assign detect_min[280][10] = (mid_1[2255:2248] < mid_0[2255:2248]) ? 1 : 0;
assign detect_min[280][11] = (mid_1[2255:2248] < mid_0[2263:2256]) ? 1 : 0;
assign detect_min[280][12] = (mid_1[2255:2248] < mid_1[2247:2240]) ? 1 : 0;
assign detect_min[280][13] = (mid_1[2255:2248] < mid_1[2263:2256]) ? 1 : 0;
assign detect_min[280][14] = (mid_1[2255:2248] < mid_2[2247:2240]) ? 1 : 0;
assign detect_min[280][15] = (mid_1[2255:2248] < mid_2[2255:2248]) ? 1 : 0;
assign detect_min[280][16] = (mid_1[2255:2248] < mid_2[2263:2256]) ? 1 : 0;
assign detect_min[280][17] = (mid_1[2255:2248] < btm_0[2247:2240]) ? 1 : 0;
assign detect_min[280][18] = (mid_1[2255:2248] < btm_0[2255:2248]) ? 1 : 0;
assign detect_min[280][19] = (mid_1[2255:2248] < btm_0[2263:2256]) ? 1 : 0;
assign detect_min[280][20] = (mid_1[2255:2248] < btm_1[2247:2240]) ? 1 : 0;
assign detect_min[280][21] = (mid_1[2255:2248] < btm_1[2255:2248]) ? 1 : 0;
assign detect_min[280][22] = (mid_1[2255:2248] < btm_1[2263:2256]) ? 1 : 0;
assign detect_min[280][23] = (mid_1[2255:2248] < btm_2[2247:2240]) ? 1 : 0;
assign detect_min[280][24] = (mid_1[2255:2248] < btm_2[2255:2248]) ? 1 : 0;
assign detect_min[280][25] = (mid_1[2255:2248] < btm_2[2263:2256]) ? 1 : 0;

assign detect_min[281][0] = (mid_1[2263:2256] < top_0[2255:2248]) ? 1 : 0;
assign detect_min[281][1] = (mid_1[2263:2256] < top_0[2263:2256]) ? 1 : 0;
assign detect_min[281][2] = (mid_1[2263:2256] < top_0[2271:2264]) ? 1 : 0;
assign detect_min[281][3] = (mid_1[2263:2256] < top_1[2255:2248]) ? 1 : 0;
assign detect_min[281][4] = (mid_1[2263:2256] < top_1[2263:2256]) ? 1 : 0;
assign detect_min[281][5] = (mid_1[2263:2256] < top_1[2271:2264]) ? 1 : 0;
assign detect_min[281][6] = (mid_1[2263:2256] < top_2[2255:2248]) ? 1 : 0;
assign detect_min[281][7] = (mid_1[2263:2256] < top_2[2263:2256]) ? 1 : 0;
assign detect_min[281][8] = (mid_1[2263:2256] < top_2[2271:2264]) ? 1 : 0;
assign detect_min[281][9] = (mid_1[2263:2256] < mid_0[2255:2248]) ? 1 : 0;
assign detect_min[281][10] = (mid_1[2263:2256] < mid_0[2263:2256]) ? 1 : 0;
assign detect_min[281][11] = (mid_1[2263:2256] < mid_0[2271:2264]) ? 1 : 0;
assign detect_min[281][12] = (mid_1[2263:2256] < mid_1[2255:2248]) ? 1 : 0;
assign detect_min[281][13] = (mid_1[2263:2256] < mid_1[2271:2264]) ? 1 : 0;
assign detect_min[281][14] = (mid_1[2263:2256] < mid_2[2255:2248]) ? 1 : 0;
assign detect_min[281][15] = (mid_1[2263:2256] < mid_2[2263:2256]) ? 1 : 0;
assign detect_min[281][16] = (mid_1[2263:2256] < mid_2[2271:2264]) ? 1 : 0;
assign detect_min[281][17] = (mid_1[2263:2256] < btm_0[2255:2248]) ? 1 : 0;
assign detect_min[281][18] = (mid_1[2263:2256] < btm_0[2263:2256]) ? 1 : 0;
assign detect_min[281][19] = (mid_1[2263:2256] < btm_0[2271:2264]) ? 1 : 0;
assign detect_min[281][20] = (mid_1[2263:2256] < btm_1[2255:2248]) ? 1 : 0;
assign detect_min[281][21] = (mid_1[2263:2256] < btm_1[2263:2256]) ? 1 : 0;
assign detect_min[281][22] = (mid_1[2263:2256] < btm_1[2271:2264]) ? 1 : 0;
assign detect_min[281][23] = (mid_1[2263:2256] < btm_2[2255:2248]) ? 1 : 0;
assign detect_min[281][24] = (mid_1[2263:2256] < btm_2[2263:2256]) ? 1 : 0;
assign detect_min[281][25] = (mid_1[2263:2256] < btm_2[2271:2264]) ? 1 : 0;

assign detect_min[282][0] = (mid_1[2271:2264] < top_0[2263:2256]) ? 1 : 0;
assign detect_min[282][1] = (mid_1[2271:2264] < top_0[2271:2264]) ? 1 : 0;
assign detect_min[282][2] = (mid_1[2271:2264] < top_0[2279:2272]) ? 1 : 0;
assign detect_min[282][3] = (mid_1[2271:2264] < top_1[2263:2256]) ? 1 : 0;
assign detect_min[282][4] = (mid_1[2271:2264] < top_1[2271:2264]) ? 1 : 0;
assign detect_min[282][5] = (mid_1[2271:2264] < top_1[2279:2272]) ? 1 : 0;
assign detect_min[282][6] = (mid_1[2271:2264] < top_2[2263:2256]) ? 1 : 0;
assign detect_min[282][7] = (mid_1[2271:2264] < top_2[2271:2264]) ? 1 : 0;
assign detect_min[282][8] = (mid_1[2271:2264] < top_2[2279:2272]) ? 1 : 0;
assign detect_min[282][9] = (mid_1[2271:2264] < mid_0[2263:2256]) ? 1 : 0;
assign detect_min[282][10] = (mid_1[2271:2264] < mid_0[2271:2264]) ? 1 : 0;
assign detect_min[282][11] = (mid_1[2271:2264] < mid_0[2279:2272]) ? 1 : 0;
assign detect_min[282][12] = (mid_1[2271:2264] < mid_1[2263:2256]) ? 1 : 0;
assign detect_min[282][13] = (mid_1[2271:2264] < mid_1[2279:2272]) ? 1 : 0;
assign detect_min[282][14] = (mid_1[2271:2264] < mid_2[2263:2256]) ? 1 : 0;
assign detect_min[282][15] = (mid_1[2271:2264] < mid_2[2271:2264]) ? 1 : 0;
assign detect_min[282][16] = (mid_1[2271:2264] < mid_2[2279:2272]) ? 1 : 0;
assign detect_min[282][17] = (mid_1[2271:2264] < btm_0[2263:2256]) ? 1 : 0;
assign detect_min[282][18] = (mid_1[2271:2264] < btm_0[2271:2264]) ? 1 : 0;
assign detect_min[282][19] = (mid_1[2271:2264] < btm_0[2279:2272]) ? 1 : 0;
assign detect_min[282][20] = (mid_1[2271:2264] < btm_1[2263:2256]) ? 1 : 0;
assign detect_min[282][21] = (mid_1[2271:2264] < btm_1[2271:2264]) ? 1 : 0;
assign detect_min[282][22] = (mid_1[2271:2264] < btm_1[2279:2272]) ? 1 : 0;
assign detect_min[282][23] = (mid_1[2271:2264] < btm_2[2263:2256]) ? 1 : 0;
assign detect_min[282][24] = (mid_1[2271:2264] < btm_2[2271:2264]) ? 1 : 0;
assign detect_min[282][25] = (mid_1[2271:2264] < btm_2[2279:2272]) ? 1 : 0;

assign detect_min[283][0] = (mid_1[2279:2272] < top_0[2271:2264]) ? 1 : 0;
assign detect_min[283][1] = (mid_1[2279:2272] < top_0[2279:2272]) ? 1 : 0;
assign detect_min[283][2] = (mid_1[2279:2272] < top_0[2287:2280]) ? 1 : 0;
assign detect_min[283][3] = (mid_1[2279:2272] < top_1[2271:2264]) ? 1 : 0;
assign detect_min[283][4] = (mid_1[2279:2272] < top_1[2279:2272]) ? 1 : 0;
assign detect_min[283][5] = (mid_1[2279:2272] < top_1[2287:2280]) ? 1 : 0;
assign detect_min[283][6] = (mid_1[2279:2272] < top_2[2271:2264]) ? 1 : 0;
assign detect_min[283][7] = (mid_1[2279:2272] < top_2[2279:2272]) ? 1 : 0;
assign detect_min[283][8] = (mid_1[2279:2272] < top_2[2287:2280]) ? 1 : 0;
assign detect_min[283][9] = (mid_1[2279:2272] < mid_0[2271:2264]) ? 1 : 0;
assign detect_min[283][10] = (mid_1[2279:2272] < mid_0[2279:2272]) ? 1 : 0;
assign detect_min[283][11] = (mid_1[2279:2272] < mid_0[2287:2280]) ? 1 : 0;
assign detect_min[283][12] = (mid_1[2279:2272] < mid_1[2271:2264]) ? 1 : 0;
assign detect_min[283][13] = (mid_1[2279:2272] < mid_1[2287:2280]) ? 1 : 0;
assign detect_min[283][14] = (mid_1[2279:2272] < mid_2[2271:2264]) ? 1 : 0;
assign detect_min[283][15] = (mid_1[2279:2272] < mid_2[2279:2272]) ? 1 : 0;
assign detect_min[283][16] = (mid_1[2279:2272] < mid_2[2287:2280]) ? 1 : 0;
assign detect_min[283][17] = (mid_1[2279:2272] < btm_0[2271:2264]) ? 1 : 0;
assign detect_min[283][18] = (mid_1[2279:2272] < btm_0[2279:2272]) ? 1 : 0;
assign detect_min[283][19] = (mid_1[2279:2272] < btm_0[2287:2280]) ? 1 : 0;
assign detect_min[283][20] = (mid_1[2279:2272] < btm_1[2271:2264]) ? 1 : 0;
assign detect_min[283][21] = (mid_1[2279:2272] < btm_1[2279:2272]) ? 1 : 0;
assign detect_min[283][22] = (mid_1[2279:2272] < btm_1[2287:2280]) ? 1 : 0;
assign detect_min[283][23] = (mid_1[2279:2272] < btm_2[2271:2264]) ? 1 : 0;
assign detect_min[283][24] = (mid_1[2279:2272] < btm_2[2279:2272]) ? 1 : 0;
assign detect_min[283][25] = (mid_1[2279:2272] < btm_2[2287:2280]) ? 1 : 0;

assign detect_min[284][0] = (mid_1[2287:2280] < top_0[2279:2272]) ? 1 : 0;
assign detect_min[284][1] = (mid_1[2287:2280] < top_0[2287:2280]) ? 1 : 0;
assign detect_min[284][2] = (mid_1[2287:2280] < top_0[2295:2288]) ? 1 : 0;
assign detect_min[284][3] = (mid_1[2287:2280] < top_1[2279:2272]) ? 1 : 0;
assign detect_min[284][4] = (mid_1[2287:2280] < top_1[2287:2280]) ? 1 : 0;
assign detect_min[284][5] = (mid_1[2287:2280] < top_1[2295:2288]) ? 1 : 0;
assign detect_min[284][6] = (mid_1[2287:2280] < top_2[2279:2272]) ? 1 : 0;
assign detect_min[284][7] = (mid_1[2287:2280] < top_2[2287:2280]) ? 1 : 0;
assign detect_min[284][8] = (mid_1[2287:2280] < top_2[2295:2288]) ? 1 : 0;
assign detect_min[284][9] = (mid_1[2287:2280] < mid_0[2279:2272]) ? 1 : 0;
assign detect_min[284][10] = (mid_1[2287:2280] < mid_0[2287:2280]) ? 1 : 0;
assign detect_min[284][11] = (mid_1[2287:2280] < mid_0[2295:2288]) ? 1 : 0;
assign detect_min[284][12] = (mid_1[2287:2280] < mid_1[2279:2272]) ? 1 : 0;
assign detect_min[284][13] = (mid_1[2287:2280] < mid_1[2295:2288]) ? 1 : 0;
assign detect_min[284][14] = (mid_1[2287:2280] < mid_2[2279:2272]) ? 1 : 0;
assign detect_min[284][15] = (mid_1[2287:2280] < mid_2[2287:2280]) ? 1 : 0;
assign detect_min[284][16] = (mid_1[2287:2280] < mid_2[2295:2288]) ? 1 : 0;
assign detect_min[284][17] = (mid_1[2287:2280] < btm_0[2279:2272]) ? 1 : 0;
assign detect_min[284][18] = (mid_1[2287:2280] < btm_0[2287:2280]) ? 1 : 0;
assign detect_min[284][19] = (mid_1[2287:2280] < btm_0[2295:2288]) ? 1 : 0;
assign detect_min[284][20] = (mid_1[2287:2280] < btm_1[2279:2272]) ? 1 : 0;
assign detect_min[284][21] = (mid_1[2287:2280] < btm_1[2287:2280]) ? 1 : 0;
assign detect_min[284][22] = (mid_1[2287:2280] < btm_1[2295:2288]) ? 1 : 0;
assign detect_min[284][23] = (mid_1[2287:2280] < btm_2[2279:2272]) ? 1 : 0;
assign detect_min[284][24] = (mid_1[2287:2280] < btm_2[2287:2280]) ? 1 : 0;
assign detect_min[284][25] = (mid_1[2287:2280] < btm_2[2295:2288]) ? 1 : 0;

assign detect_min[285][0] = (mid_1[2295:2288] < top_0[2287:2280]) ? 1 : 0;
assign detect_min[285][1] = (mid_1[2295:2288] < top_0[2295:2288]) ? 1 : 0;
assign detect_min[285][2] = (mid_1[2295:2288] < top_0[2303:2296]) ? 1 : 0;
assign detect_min[285][3] = (mid_1[2295:2288] < top_1[2287:2280]) ? 1 : 0;
assign detect_min[285][4] = (mid_1[2295:2288] < top_1[2295:2288]) ? 1 : 0;
assign detect_min[285][5] = (mid_1[2295:2288] < top_1[2303:2296]) ? 1 : 0;
assign detect_min[285][6] = (mid_1[2295:2288] < top_2[2287:2280]) ? 1 : 0;
assign detect_min[285][7] = (mid_1[2295:2288] < top_2[2295:2288]) ? 1 : 0;
assign detect_min[285][8] = (mid_1[2295:2288] < top_2[2303:2296]) ? 1 : 0;
assign detect_min[285][9] = (mid_1[2295:2288] < mid_0[2287:2280]) ? 1 : 0;
assign detect_min[285][10] = (mid_1[2295:2288] < mid_0[2295:2288]) ? 1 : 0;
assign detect_min[285][11] = (mid_1[2295:2288] < mid_0[2303:2296]) ? 1 : 0;
assign detect_min[285][12] = (mid_1[2295:2288] < mid_1[2287:2280]) ? 1 : 0;
assign detect_min[285][13] = (mid_1[2295:2288] < mid_1[2303:2296]) ? 1 : 0;
assign detect_min[285][14] = (mid_1[2295:2288] < mid_2[2287:2280]) ? 1 : 0;
assign detect_min[285][15] = (mid_1[2295:2288] < mid_2[2295:2288]) ? 1 : 0;
assign detect_min[285][16] = (mid_1[2295:2288] < mid_2[2303:2296]) ? 1 : 0;
assign detect_min[285][17] = (mid_1[2295:2288] < btm_0[2287:2280]) ? 1 : 0;
assign detect_min[285][18] = (mid_1[2295:2288] < btm_0[2295:2288]) ? 1 : 0;
assign detect_min[285][19] = (mid_1[2295:2288] < btm_0[2303:2296]) ? 1 : 0;
assign detect_min[285][20] = (mid_1[2295:2288] < btm_1[2287:2280]) ? 1 : 0;
assign detect_min[285][21] = (mid_1[2295:2288] < btm_1[2295:2288]) ? 1 : 0;
assign detect_min[285][22] = (mid_1[2295:2288] < btm_1[2303:2296]) ? 1 : 0;
assign detect_min[285][23] = (mid_1[2295:2288] < btm_2[2287:2280]) ? 1 : 0;
assign detect_min[285][24] = (mid_1[2295:2288] < btm_2[2295:2288]) ? 1 : 0;
assign detect_min[285][25] = (mid_1[2295:2288] < btm_2[2303:2296]) ? 1 : 0;

assign detect_min[286][0] = (mid_1[2303:2296] < top_0[2295:2288]) ? 1 : 0;
assign detect_min[286][1] = (mid_1[2303:2296] < top_0[2303:2296]) ? 1 : 0;
assign detect_min[286][2] = (mid_1[2303:2296] < top_0[2311:2304]) ? 1 : 0;
assign detect_min[286][3] = (mid_1[2303:2296] < top_1[2295:2288]) ? 1 : 0;
assign detect_min[286][4] = (mid_1[2303:2296] < top_1[2303:2296]) ? 1 : 0;
assign detect_min[286][5] = (mid_1[2303:2296] < top_1[2311:2304]) ? 1 : 0;
assign detect_min[286][6] = (mid_1[2303:2296] < top_2[2295:2288]) ? 1 : 0;
assign detect_min[286][7] = (mid_1[2303:2296] < top_2[2303:2296]) ? 1 : 0;
assign detect_min[286][8] = (mid_1[2303:2296] < top_2[2311:2304]) ? 1 : 0;
assign detect_min[286][9] = (mid_1[2303:2296] < mid_0[2295:2288]) ? 1 : 0;
assign detect_min[286][10] = (mid_1[2303:2296] < mid_0[2303:2296]) ? 1 : 0;
assign detect_min[286][11] = (mid_1[2303:2296] < mid_0[2311:2304]) ? 1 : 0;
assign detect_min[286][12] = (mid_1[2303:2296] < mid_1[2295:2288]) ? 1 : 0;
assign detect_min[286][13] = (mid_1[2303:2296] < mid_1[2311:2304]) ? 1 : 0;
assign detect_min[286][14] = (mid_1[2303:2296] < mid_2[2295:2288]) ? 1 : 0;
assign detect_min[286][15] = (mid_1[2303:2296] < mid_2[2303:2296]) ? 1 : 0;
assign detect_min[286][16] = (mid_1[2303:2296] < mid_2[2311:2304]) ? 1 : 0;
assign detect_min[286][17] = (mid_1[2303:2296] < btm_0[2295:2288]) ? 1 : 0;
assign detect_min[286][18] = (mid_1[2303:2296] < btm_0[2303:2296]) ? 1 : 0;
assign detect_min[286][19] = (mid_1[2303:2296] < btm_0[2311:2304]) ? 1 : 0;
assign detect_min[286][20] = (mid_1[2303:2296] < btm_1[2295:2288]) ? 1 : 0;
assign detect_min[286][21] = (mid_1[2303:2296] < btm_1[2303:2296]) ? 1 : 0;
assign detect_min[286][22] = (mid_1[2303:2296] < btm_1[2311:2304]) ? 1 : 0;
assign detect_min[286][23] = (mid_1[2303:2296] < btm_2[2295:2288]) ? 1 : 0;
assign detect_min[286][24] = (mid_1[2303:2296] < btm_2[2303:2296]) ? 1 : 0;
assign detect_min[286][25] = (mid_1[2303:2296] < btm_2[2311:2304]) ? 1 : 0;

assign detect_min[287][0] = (mid_1[2311:2304] < top_0[2303:2296]) ? 1 : 0;
assign detect_min[287][1] = (mid_1[2311:2304] < top_0[2311:2304]) ? 1 : 0;
assign detect_min[287][2] = (mid_1[2311:2304] < top_0[2319:2312]) ? 1 : 0;
assign detect_min[287][3] = (mid_1[2311:2304] < top_1[2303:2296]) ? 1 : 0;
assign detect_min[287][4] = (mid_1[2311:2304] < top_1[2311:2304]) ? 1 : 0;
assign detect_min[287][5] = (mid_1[2311:2304] < top_1[2319:2312]) ? 1 : 0;
assign detect_min[287][6] = (mid_1[2311:2304] < top_2[2303:2296]) ? 1 : 0;
assign detect_min[287][7] = (mid_1[2311:2304] < top_2[2311:2304]) ? 1 : 0;
assign detect_min[287][8] = (mid_1[2311:2304] < top_2[2319:2312]) ? 1 : 0;
assign detect_min[287][9] = (mid_1[2311:2304] < mid_0[2303:2296]) ? 1 : 0;
assign detect_min[287][10] = (mid_1[2311:2304] < mid_0[2311:2304]) ? 1 : 0;
assign detect_min[287][11] = (mid_1[2311:2304] < mid_0[2319:2312]) ? 1 : 0;
assign detect_min[287][12] = (mid_1[2311:2304] < mid_1[2303:2296]) ? 1 : 0;
assign detect_min[287][13] = (mid_1[2311:2304] < mid_1[2319:2312]) ? 1 : 0;
assign detect_min[287][14] = (mid_1[2311:2304] < mid_2[2303:2296]) ? 1 : 0;
assign detect_min[287][15] = (mid_1[2311:2304] < mid_2[2311:2304]) ? 1 : 0;
assign detect_min[287][16] = (mid_1[2311:2304] < mid_2[2319:2312]) ? 1 : 0;
assign detect_min[287][17] = (mid_1[2311:2304] < btm_0[2303:2296]) ? 1 : 0;
assign detect_min[287][18] = (mid_1[2311:2304] < btm_0[2311:2304]) ? 1 : 0;
assign detect_min[287][19] = (mid_1[2311:2304] < btm_0[2319:2312]) ? 1 : 0;
assign detect_min[287][20] = (mid_1[2311:2304] < btm_1[2303:2296]) ? 1 : 0;
assign detect_min[287][21] = (mid_1[2311:2304] < btm_1[2311:2304]) ? 1 : 0;
assign detect_min[287][22] = (mid_1[2311:2304] < btm_1[2319:2312]) ? 1 : 0;
assign detect_min[287][23] = (mid_1[2311:2304] < btm_2[2303:2296]) ? 1 : 0;
assign detect_min[287][24] = (mid_1[2311:2304] < btm_2[2311:2304]) ? 1 : 0;
assign detect_min[287][25] = (mid_1[2311:2304] < btm_2[2319:2312]) ? 1 : 0;

assign detect_min[288][0] = (mid_1[2319:2312] < top_0[2311:2304]) ? 1 : 0;
assign detect_min[288][1] = (mid_1[2319:2312] < top_0[2319:2312]) ? 1 : 0;
assign detect_min[288][2] = (mid_1[2319:2312] < top_0[2327:2320]) ? 1 : 0;
assign detect_min[288][3] = (mid_1[2319:2312] < top_1[2311:2304]) ? 1 : 0;
assign detect_min[288][4] = (mid_1[2319:2312] < top_1[2319:2312]) ? 1 : 0;
assign detect_min[288][5] = (mid_1[2319:2312] < top_1[2327:2320]) ? 1 : 0;
assign detect_min[288][6] = (mid_1[2319:2312] < top_2[2311:2304]) ? 1 : 0;
assign detect_min[288][7] = (mid_1[2319:2312] < top_2[2319:2312]) ? 1 : 0;
assign detect_min[288][8] = (mid_1[2319:2312] < top_2[2327:2320]) ? 1 : 0;
assign detect_min[288][9] = (mid_1[2319:2312] < mid_0[2311:2304]) ? 1 : 0;
assign detect_min[288][10] = (mid_1[2319:2312] < mid_0[2319:2312]) ? 1 : 0;
assign detect_min[288][11] = (mid_1[2319:2312] < mid_0[2327:2320]) ? 1 : 0;
assign detect_min[288][12] = (mid_1[2319:2312] < mid_1[2311:2304]) ? 1 : 0;
assign detect_min[288][13] = (mid_1[2319:2312] < mid_1[2327:2320]) ? 1 : 0;
assign detect_min[288][14] = (mid_1[2319:2312] < mid_2[2311:2304]) ? 1 : 0;
assign detect_min[288][15] = (mid_1[2319:2312] < mid_2[2319:2312]) ? 1 : 0;
assign detect_min[288][16] = (mid_1[2319:2312] < mid_2[2327:2320]) ? 1 : 0;
assign detect_min[288][17] = (mid_1[2319:2312] < btm_0[2311:2304]) ? 1 : 0;
assign detect_min[288][18] = (mid_1[2319:2312] < btm_0[2319:2312]) ? 1 : 0;
assign detect_min[288][19] = (mid_1[2319:2312] < btm_0[2327:2320]) ? 1 : 0;
assign detect_min[288][20] = (mid_1[2319:2312] < btm_1[2311:2304]) ? 1 : 0;
assign detect_min[288][21] = (mid_1[2319:2312] < btm_1[2319:2312]) ? 1 : 0;
assign detect_min[288][22] = (mid_1[2319:2312] < btm_1[2327:2320]) ? 1 : 0;
assign detect_min[288][23] = (mid_1[2319:2312] < btm_2[2311:2304]) ? 1 : 0;
assign detect_min[288][24] = (mid_1[2319:2312] < btm_2[2319:2312]) ? 1 : 0;
assign detect_min[288][25] = (mid_1[2319:2312] < btm_2[2327:2320]) ? 1 : 0;

assign detect_min[289][0] = (mid_1[2327:2320] < top_0[2319:2312]) ? 1 : 0;
assign detect_min[289][1] = (mid_1[2327:2320] < top_0[2327:2320]) ? 1 : 0;
assign detect_min[289][2] = (mid_1[2327:2320] < top_0[2335:2328]) ? 1 : 0;
assign detect_min[289][3] = (mid_1[2327:2320] < top_1[2319:2312]) ? 1 : 0;
assign detect_min[289][4] = (mid_1[2327:2320] < top_1[2327:2320]) ? 1 : 0;
assign detect_min[289][5] = (mid_1[2327:2320] < top_1[2335:2328]) ? 1 : 0;
assign detect_min[289][6] = (mid_1[2327:2320] < top_2[2319:2312]) ? 1 : 0;
assign detect_min[289][7] = (mid_1[2327:2320] < top_2[2327:2320]) ? 1 : 0;
assign detect_min[289][8] = (mid_1[2327:2320] < top_2[2335:2328]) ? 1 : 0;
assign detect_min[289][9] = (mid_1[2327:2320] < mid_0[2319:2312]) ? 1 : 0;
assign detect_min[289][10] = (mid_1[2327:2320] < mid_0[2327:2320]) ? 1 : 0;
assign detect_min[289][11] = (mid_1[2327:2320] < mid_0[2335:2328]) ? 1 : 0;
assign detect_min[289][12] = (mid_1[2327:2320] < mid_1[2319:2312]) ? 1 : 0;
assign detect_min[289][13] = (mid_1[2327:2320] < mid_1[2335:2328]) ? 1 : 0;
assign detect_min[289][14] = (mid_1[2327:2320] < mid_2[2319:2312]) ? 1 : 0;
assign detect_min[289][15] = (mid_1[2327:2320] < mid_2[2327:2320]) ? 1 : 0;
assign detect_min[289][16] = (mid_1[2327:2320] < mid_2[2335:2328]) ? 1 : 0;
assign detect_min[289][17] = (mid_1[2327:2320] < btm_0[2319:2312]) ? 1 : 0;
assign detect_min[289][18] = (mid_1[2327:2320] < btm_0[2327:2320]) ? 1 : 0;
assign detect_min[289][19] = (mid_1[2327:2320] < btm_0[2335:2328]) ? 1 : 0;
assign detect_min[289][20] = (mid_1[2327:2320] < btm_1[2319:2312]) ? 1 : 0;
assign detect_min[289][21] = (mid_1[2327:2320] < btm_1[2327:2320]) ? 1 : 0;
assign detect_min[289][22] = (mid_1[2327:2320] < btm_1[2335:2328]) ? 1 : 0;
assign detect_min[289][23] = (mid_1[2327:2320] < btm_2[2319:2312]) ? 1 : 0;
assign detect_min[289][24] = (mid_1[2327:2320] < btm_2[2327:2320]) ? 1 : 0;
assign detect_min[289][25] = (mid_1[2327:2320] < btm_2[2335:2328]) ? 1 : 0;

assign detect_min[290][0] = (mid_1[2335:2328] < top_0[2327:2320]) ? 1 : 0;
assign detect_min[290][1] = (mid_1[2335:2328] < top_0[2335:2328]) ? 1 : 0;
assign detect_min[290][2] = (mid_1[2335:2328] < top_0[2343:2336]) ? 1 : 0;
assign detect_min[290][3] = (mid_1[2335:2328] < top_1[2327:2320]) ? 1 : 0;
assign detect_min[290][4] = (mid_1[2335:2328] < top_1[2335:2328]) ? 1 : 0;
assign detect_min[290][5] = (mid_1[2335:2328] < top_1[2343:2336]) ? 1 : 0;
assign detect_min[290][6] = (mid_1[2335:2328] < top_2[2327:2320]) ? 1 : 0;
assign detect_min[290][7] = (mid_1[2335:2328] < top_2[2335:2328]) ? 1 : 0;
assign detect_min[290][8] = (mid_1[2335:2328] < top_2[2343:2336]) ? 1 : 0;
assign detect_min[290][9] = (mid_1[2335:2328] < mid_0[2327:2320]) ? 1 : 0;
assign detect_min[290][10] = (mid_1[2335:2328] < mid_0[2335:2328]) ? 1 : 0;
assign detect_min[290][11] = (mid_1[2335:2328] < mid_0[2343:2336]) ? 1 : 0;
assign detect_min[290][12] = (mid_1[2335:2328] < mid_1[2327:2320]) ? 1 : 0;
assign detect_min[290][13] = (mid_1[2335:2328] < mid_1[2343:2336]) ? 1 : 0;
assign detect_min[290][14] = (mid_1[2335:2328] < mid_2[2327:2320]) ? 1 : 0;
assign detect_min[290][15] = (mid_1[2335:2328] < mid_2[2335:2328]) ? 1 : 0;
assign detect_min[290][16] = (mid_1[2335:2328] < mid_2[2343:2336]) ? 1 : 0;
assign detect_min[290][17] = (mid_1[2335:2328] < btm_0[2327:2320]) ? 1 : 0;
assign detect_min[290][18] = (mid_1[2335:2328] < btm_0[2335:2328]) ? 1 : 0;
assign detect_min[290][19] = (mid_1[2335:2328] < btm_0[2343:2336]) ? 1 : 0;
assign detect_min[290][20] = (mid_1[2335:2328] < btm_1[2327:2320]) ? 1 : 0;
assign detect_min[290][21] = (mid_1[2335:2328] < btm_1[2335:2328]) ? 1 : 0;
assign detect_min[290][22] = (mid_1[2335:2328] < btm_1[2343:2336]) ? 1 : 0;
assign detect_min[290][23] = (mid_1[2335:2328] < btm_2[2327:2320]) ? 1 : 0;
assign detect_min[290][24] = (mid_1[2335:2328] < btm_2[2335:2328]) ? 1 : 0;
assign detect_min[290][25] = (mid_1[2335:2328] < btm_2[2343:2336]) ? 1 : 0;

assign detect_min[291][0] = (mid_1[2343:2336] < top_0[2335:2328]) ? 1 : 0;
assign detect_min[291][1] = (mid_1[2343:2336] < top_0[2343:2336]) ? 1 : 0;
assign detect_min[291][2] = (mid_1[2343:2336] < top_0[2351:2344]) ? 1 : 0;
assign detect_min[291][3] = (mid_1[2343:2336] < top_1[2335:2328]) ? 1 : 0;
assign detect_min[291][4] = (mid_1[2343:2336] < top_1[2343:2336]) ? 1 : 0;
assign detect_min[291][5] = (mid_1[2343:2336] < top_1[2351:2344]) ? 1 : 0;
assign detect_min[291][6] = (mid_1[2343:2336] < top_2[2335:2328]) ? 1 : 0;
assign detect_min[291][7] = (mid_1[2343:2336] < top_2[2343:2336]) ? 1 : 0;
assign detect_min[291][8] = (mid_1[2343:2336] < top_2[2351:2344]) ? 1 : 0;
assign detect_min[291][9] = (mid_1[2343:2336] < mid_0[2335:2328]) ? 1 : 0;
assign detect_min[291][10] = (mid_1[2343:2336] < mid_0[2343:2336]) ? 1 : 0;
assign detect_min[291][11] = (mid_1[2343:2336] < mid_0[2351:2344]) ? 1 : 0;
assign detect_min[291][12] = (mid_1[2343:2336] < mid_1[2335:2328]) ? 1 : 0;
assign detect_min[291][13] = (mid_1[2343:2336] < mid_1[2351:2344]) ? 1 : 0;
assign detect_min[291][14] = (mid_1[2343:2336] < mid_2[2335:2328]) ? 1 : 0;
assign detect_min[291][15] = (mid_1[2343:2336] < mid_2[2343:2336]) ? 1 : 0;
assign detect_min[291][16] = (mid_1[2343:2336] < mid_2[2351:2344]) ? 1 : 0;
assign detect_min[291][17] = (mid_1[2343:2336] < btm_0[2335:2328]) ? 1 : 0;
assign detect_min[291][18] = (mid_1[2343:2336] < btm_0[2343:2336]) ? 1 : 0;
assign detect_min[291][19] = (mid_1[2343:2336] < btm_0[2351:2344]) ? 1 : 0;
assign detect_min[291][20] = (mid_1[2343:2336] < btm_1[2335:2328]) ? 1 : 0;
assign detect_min[291][21] = (mid_1[2343:2336] < btm_1[2343:2336]) ? 1 : 0;
assign detect_min[291][22] = (mid_1[2343:2336] < btm_1[2351:2344]) ? 1 : 0;
assign detect_min[291][23] = (mid_1[2343:2336] < btm_2[2335:2328]) ? 1 : 0;
assign detect_min[291][24] = (mid_1[2343:2336] < btm_2[2343:2336]) ? 1 : 0;
assign detect_min[291][25] = (mid_1[2343:2336] < btm_2[2351:2344]) ? 1 : 0;

assign detect_min[292][0] = (mid_1[2351:2344] < top_0[2343:2336]) ? 1 : 0;
assign detect_min[292][1] = (mid_1[2351:2344] < top_0[2351:2344]) ? 1 : 0;
assign detect_min[292][2] = (mid_1[2351:2344] < top_0[2359:2352]) ? 1 : 0;
assign detect_min[292][3] = (mid_1[2351:2344] < top_1[2343:2336]) ? 1 : 0;
assign detect_min[292][4] = (mid_1[2351:2344] < top_1[2351:2344]) ? 1 : 0;
assign detect_min[292][5] = (mid_1[2351:2344] < top_1[2359:2352]) ? 1 : 0;
assign detect_min[292][6] = (mid_1[2351:2344] < top_2[2343:2336]) ? 1 : 0;
assign detect_min[292][7] = (mid_1[2351:2344] < top_2[2351:2344]) ? 1 : 0;
assign detect_min[292][8] = (mid_1[2351:2344] < top_2[2359:2352]) ? 1 : 0;
assign detect_min[292][9] = (mid_1[2351:2344] < mid_0[2343:2336]) ? 1 : 0;
assign detect_min[292][10] = (mid_1[2351:2344] < mid_0[2351:2344]) ? 1 : 0;
assign detect_min[292][11] = (mid_1[2351:2344] < mid_0[2359:2352]) ? 1 : 0;
assign detect_min[292][12] = (mid_1[2351:2344] < mid_1[2343:2336]) ? 1 : 0;
assign detect_min[292][13] = (mid_1[2351:2344] < mid_1[2359:2352]) ? 1 : 0;
assign detect_min[292][14] = (mid_1[2351:2344] < mid_2[2343:2336]) ? 1 : 0;
assign detect_min[292][15] = (mid_1[2351:2344] < mid_2[2351:2344]) ? 1 : 0;
assign detect_min[292][16] = (mid_1[2351:2344] < mid_2[2359:2352]) ? 1 : 0;
assign detect_min[292][17] = (mid_1[2351:2344] < btm_0[2343:2336]) ? 1 : 0;
assign detect_min[292][18] = (mid_1[2351:2344] < btm_0[2351:2344]) ? 1 : 0;
assign detect_min[292][19] = (mid_1[2351:2344] < btm_0[2359:2352]) ? 1 : 0;
assign detect_min[292][20] = (mid_1[2351:2344] < btm_1[2343:2336]) ? 1 : 0;
assign detect_min[292][21] = (mid_1[2351:2344] < btm_1[2351:2344]) ? 1 : 0;
assign detect_min[292][22] = (mid_1[2351:2344] < btm_1[2359:2352]) ? 1 : 0;
assign detect_min[292][23] = (mid_1[2351:2344] < btm_2[2343:2336]) ? 1 : 0;
assign detect_min[292][24] = (mid_1[2351:2344] < btm_2[2351:2344]) ? 1 : 0;
assign detect_min[292][25] = (mid_1[2351:2344] < btm_2[2359:2352]) ? 1 : 0;

assign detect_min[293][0] = (mid_1[2359:2352] < top_0[2351:2344]) ? 1 : 0;
assign detect_min[293][1] = (mid_1[2359:2352] < top_0[2359:2352]) ? 1 : 0;
assign detect_min[293][2] = (mid_1[2359:2352] < top_0[2367:2360]) ? 1 : 0;
assign detect_min[293][3] = (mid_1[2359:2352] < top_1[2351:2344]) ? 1 : 0;
assign detect_min[293][4] = (mid_1[2359:2352] < top_1[2359:2352]) ? 1 : 0;
assign detect_min[293][5] = (mid_1[2359:2352] < top_1[2367:2360]) ? 1 : 0;
assign detect_min[293][6] = (mid_1[2359:2352] < top_2[2351:2344]) ? 1 : 0;
assign detect_min[293][7] = (mid_1[2359:2352] < top_2[2359:2352]) ? 1 : 0;
assign detect_min[293][8] = (mid_1[2359:2352] < top_2[2367:2360]) ? 1 : 0;
assign detect_min[293][9] = (mid_1[2359:2352] < mid_0[2351:2344]) ? 1 : 0;
assign detect_min[293][10] = (mid_1[2359:2352] < mid_0[2359:2352]) ? 1 : 0;
assign detect_min[293][11] = (mid_1[2359:2352] < mid_0[2367:2360]) ? 1 : 0;
assign detect_min[293][12] = (mid_1[2359:2352] < mid_1[2351:2344]) ? 1 : 0;
assign detect_min[293][13] = (mid_1[2359:2352] < mid_1[2367:2360]) ? 1 : 0;
assign detect_min[293][14] = (mid_1[2359:2352] < mid_2[2351:2344]) ? 1 : 0;
assign detect_min[293][15] = (mid_1[2359:2352] < mid_2[2359:2352]) ? 1 : 0;
assign detect_min[293][16] = (mid_1[2359:2352] < mid_2[2367:2360]) ? 1 : 0;
assign detect_min[293][17] = (mid_1[2359:2352] < btm_0[2351:2344]) ? 1 : 0;
assign detect_min[293][18] = (mid_1[2359:2352] < btm_0[2359:2352]) ? 1 : 0;
assign detect_min[293][19] = (mid_1[2359:2352] < btm_0[2367:2360]) ? 1 : 0;
assign detect_min[293][20] = (mid_1[2359:2352] < btm_1[2351:2344]) ? 1 : 0;
assign detect_min[293][21] = (mid_1[2359:2352] < btm_1[2359:2352]) ? 1 : 0;
assign detect_min[293][22] = (mid_1[2359:2352] < btm_1[2367:2360]) ? 1 : 0;
assign detect_min[293][23] = (mid_1[2359:2352] < btm_2[2351:2344]) ? 1 : 0;
assign detect_min[293][24] = (mid_1[2359:2352] < btm_2[2359:2352]) ? 1 : 0;
assign detect_min[293][25] = (mid_1[2359:2352] < btm_2[2367:2360]) ? 1 : 0;

assign detect_min[294][0] = (mid_1[2367:2360] < top_0[2359:2352]) ? 1 : 0;
assign detect_min[294][1] = (mid_1[2367:2360] < top_0[2367:2360]) ? 1 : 0;
assign detect_min[294][2] = (mid_1[2367:2360] < top_0[2375:2368]) ? 1 : 0;
assign detect_min[294][3] = (mid_1[2367:2360] < top_1[2359:2352]) ? 1 : 0;
assign detect_min[294][4] = (mid_1[2367:2360] < top_1[2367:2360]) ? 1 : 0;
assign detect_min[294][5] = (mid_1[2367:2360] < top_1[2375:2368]) ? 1 : 0;
assign detect_min[294][6] = (mid_1[2367:2360] < top_2[2359:2352]) ? 1 : 0;
assign detect_min[294][7] = (mid_1[2367:2360] < top_2[2367:2360]) ? 1 : 0;
assign detect_min[294][8] = (mid_1[2367:2360] < top_2[2375:2368]) ? 1 : 0;
assign detect_min[294][9] = (mid_1[2367:2360] < mid_0[2359:2352]) ? 1 : 0;
assign detect_min[294][10] = (mid_1[2367:2360] < mid_0[2367:2360]) ? 1 : 0;
assign detect_min[294][11] = (mid_1[2367:2360] < mid_0[2375:2368]) ? 1 : 0;
assign detect_min[294][12] = (mid_1[2367:2360] < mid_1[2359:2352]) ? 1 : 0;
assign detect_min[294][13] = (mid_1[2367:2360] < mid_1[2375:2368]) ? 1 : 0;
assign detect_min[294][14] = (mid_1[2367:2360] < mid_2[2359:2352]) ? 1 : 0;
assign detect_min[294][15] = (mid_1[2367:2360] < mid_2[2367:2360]) ? 1 : 0;
assign detect_min[294][16] = (mid_1[2367:2360] < mid_2[2375:2368]) ? 1 : 0;
assign detect_min[294][17] = (mid_1[2367:2360] < btm_0[2359:2352]) ? 1 : 0;
assign detect_min[294][18] = (mid_1[2367:2360] < btm_0[2367:2360]) ? 1 : 0;
assign detect_min[294][19] = (mid_1[2367:2360] < btm_0[2375:2368]) ? 1 : 0;
assign detect_min[294][20] = (mid_1[2367:2360] < btm_1[2359:2352]) ? 1 : 0;
assign detect_min[294][21] = (mid_1[2367:2360] < btm_1[2367:2360]) ? 1 : 0;
assign detect_min[294][22] = (mid_1[2367:2360] < btm_1[2375:2368]) ? 1 : 0;
assign detect_min[294][23] = (mid_1[2367:2360] < btm_2[2359:2352]) ? 1 : 0;
assign detect_min[294][24] = (mid_1[2367:2360] < btm_2[2367:2360]) ? 1 : 0;
assign detect_min[294][25] = (mid_1[2367:2360] < btm_2[2375:2368]) ? 1 : 0;

assign detect_min[295][0] = (mid_1[2375:2368] < top_0[2367:2360]) ? 1 : 0;
assign detect_min[295][1] = (mid_1[2375:2368] < top_0[2375:2368]) ? 1 : 0;
assign detect_min[295][2] = (mid_1[2375:2368] < top_0[2383:2376]) ? 1 : 0;
assign detect_min[295][3] = (mid_1[2375:2368] < top_1[2367:2360]) ? 1 : 0;
assign detect_min[295][4] = (mid_1[2375:2368] < top_1[2375:2368]) ? 1 : 0;
assign detect_min[295][5] = (mid_1[2375:2368] < top_1[2383:2376]) ? 1 : 0;
assign detect_min[295][6] = (mid_1[2375:2368] < top_2[2367:2360]) ? 1 : 0;
assign detect_min[295][7] = (mid_1[2375:2368] < top_2[2375:2368]) ? 1 : 0;
assign detect_min[295][8] = (mid_1[2375:2368] < top_2[2383:2376]) ? 1 : 0;
assign detect_min[295][9] = (mid_1[2375:2368] < mid_0[2367:2360]) ? 1 : 0;
assign detect_min[295][10] = (mid_1[2375:2368] < mid_0[2375:2368]) ? 1 : 0;
assign detect_min[295][11] = (mid_1[2375:2368] < mid_0[2383:2376]) ? 1 : 0;
assign detect_min[295][12] = (mid_1[2375:2368] < mid_1[2367:2360]) ? 1 : 0;
assign detect_min[295][13] = (mid_1[2375:2368] < mid_1[2383:2376]) ? 1 : 0;
assign detect_min[295][14] = (mid_1[2375:2368] < mid_2[2367:2360]) ? 1 : 0;
assign detect_min[295][15] = (mid_1[2375:2368] < mid_2[2375:2368]) ? 1 : 0;
assign detect_min[295][16] = (mid_1[2375:2368] < mid_2[2383:2376]) ? 1 : 0;
assign detect_min[295][17] = (mid_1[2375:2368] < btm_0[2367:2360]) ? 1 : 0;
assign detect_min[295][18] = (mid_1[2375:2368] < btm_0[2375:2368]) ? 1 : 0;
assign detect_min[295][19] = (mid_1[2375:2368] < btm_0[2383:2376]) ? 1 : 0;
assign detect_min[295][20] = (mid_1[2375:2368] < btm_1[2367:2360]) ? 1 : 0;
assign detect_min[295][21] = (mid_1[2375:2368] < btm_1[2375:2368]) ? 1 : 0;
assign detect_min[295][22] = (mid_1[2375:2368] < btm_1[2383:2376]) ? 1 : 0;
assign detect_min[295][23] = (mid_1[2375:2368] < btm_2[2367:2360]) ? 1 : 0;
assign detect_min[295][24] = (mid_1[2375:2368] < btm_2[2375:2368]) ? 1 : 0;
assign detect_min[295][25] = (mid_1[2375:2368] < btm_2[2383:2376]) ? 1 : 0;

assign detect_min[296][0] = (mid_1[2383:2376] < top_0[2375:2368]) ? 1 : 0;
assign detect_min[296][1] = (mid_1[2383:2376] < top_0[2383:2376]) ? 1 : 0;
assign detect_min[296][2] = (mid_1[2383:2376] < top_0[2391:2384]) ? 1 : 0;
assign detect_min[296][3] = (mid_1[2383:2376] < top_1[2375:2368]) ? 1 : 0;
assign detect_min[296][4] = (mid_1[2383:2376] < top_1[2383:2376]) ? 1 : 0;
assign detect_min[296][5] = (mid_1[2383:2376] < top_1[2391:2384]) ? 1 : 0;
assign detect_min[296][6] = (mid_1[2383:2376] < top_2[2375:2368]) ? 1 : 0;
assign detect_min[296][7] = (mid_1[2383:2376] < top_2[2383:2376]) ? 1 : 0;
assign detect_min[296][8] = (mid_1[2383:2376] < top_2[2391:2384]) ? 1 : 0;
assign detect_min[296][9] = (mid_1[2383:2376] < mid_0[2375:2368]) ? 1 : 0;
assign detect_min[296][10] = (mid_1[2383:2376] < mid_0[2383:2376]) ? 1 : 0;
assign detect_min[296][11] = (mid_1[2383:2376] < mid_0[2391:2384]) ? 1 : 0;
assign detect_min[296][12] = (mid_1[2383:2376] < mid_1[2375:2368]) ? 1 : 0;
assign detect_min[296][13] = (mid_1[2383:2376] < mid_1[2391:2384]) ? 1 : 0;
assign detect_min[296][14] = (mid_1[2383:2376] < mid_2[2375:2368]) ? 1 : 0;
assign detect_min[296][15] = (mid_1[2383:2376] < mid_2[2383:2376]) ? 1 : 0;
assign detect_min[296][16] = (mid_1[2383:2376] < mid_2[2391:2384]) ? 1 : 0;
assign detect_min[296][17] = (mid_1[2383:2376] < btm_0[2375:2368]) ? 1 : 0;
assign detect_min[296][18] = (mid_1[2383:2376] < btm_0[2383:2376]) ? 1 : 0;
assign detect_min[296][19] = (mid_1[2383:2376] < btm_0[2391:2384]) ? 1 : 0;
assign detect_min[296][20] = (mid_1[2383:2376] < btm_1[2375:2368]) ? 1 : 0;
assign detect_min[296][21] = (mid_1[2383:2376] < btm_1[2383:2376]) ? 1 : 0;
assign detect_min[296][22] = (mid_1[2383:2376] < btm_1[2391:2384]) ? 1 : 0;
assign detect_min[296][23] = (mid_1[2383:2376] < btm_2[2375:2368]) ? 1 : 0;
assign detect_min[296][24] = (mid_1[2383:2376] < btm_2[2383:2376]) ? 1 : 0;
assign detect_min[296][25] = (mid_1[2383:2376] < btm_2[2391:2384]) ? 1 : 0;

assign detect_min[297][0] = (mid_1[2391:2384] < top_0[2383:2376]) ? 1 : 0;
assign detect_min[297][1] = (mid_1[2391:2384] < top_0[2391:2384]) ? 1 : 0;
assign detect_min[297][2] = (mid_1[2391:2384] < top_0[2399:2392]) ? 1 : 0;
assign detect_min[297][3] = (mid_1[2391:2384] < top_1[2383:2376]) ? 1 : 0;
assign detect_min[297][4] = (mid_1[2391:2384] < top_1[2391:2384]) ? 1 : 0;
assign detect_min[297][5] = (mid_1[2391:2384] < top_1[2399:2392]) ? 1 : 0;
assign detect_min[297][6] = (mid_1[2391:2384] < top_2[2383:2376]) ? 1 : 0;
assign detect_min[297][7] = (mid_1[2391:2384] < top_2[2391:2384]) ? 1 : 0;
assign detect_min[297][8] = (mid_1[2391:2384] < top_2[2399:2392]) ? 1 : 0;
assign detect_min[297][9] = (mid_1[2391:2384] < mid_0[2383:2376]) ? 1 : 0;
assign detect_min[297][10] = (mid_1[2391:2384] < mid_0[2391:2384]) ? 1 : 0;
assign detect_min[297][11] = (mid_1[2391:2384] < mid_0[2399:2392]) ? 1 : 0;
assign detect_min[297][12] = (mid_1[2391:2384] < mid_1[2383:2376]) ? 1 : 0;
assign detect_min[297][13] = (mid_1[2391:2384] < mid_1[2399:2392]) ? 1 : 0;
assign detect_min[297][14] = (mid_1[2391:2384] < mid_2[2383:2376]) ? 1 : 0;
assign detect_min[297][15] = (mid_1[2391:2384] < mid_2[2391:2384]) ? 1 : 0;
assign detect_min[297][16] = (mid_1[2391:2384] < mid_2[2399:2392]) ? 1 : 0;
assign detect_min[297][17] = (mid_1[2391:2384] < btm_0[2383:2376]) ? 1 : 0;
assign detect_min[297][18] = (mid_1[2391:2384] < btm_0[2391:2384]) ? 1 : 0;
assign detect_min[297][19] = (mid_1[2391:2384] < btm_0[2399:2392]) ? 1 : 0;
assign detect_min[297][20] = (mid_1[2391:2384] < btm_1[2383:2376]) ? 1 : 0;
assign detect_min[297][21] = (mid_1[2391:2384] < btm_1[2391:2384]) ? 1 : 0;
assign detect_min[297][22] = (mid_1[2391:2384] < btm_1[2399:2392]) ? 1 : 0;
assign detect_min[297][23] = (mid_1[2391:2384] < btm_2[2383:2376]) ? 1 : 0;
assign detect_min[297][24] = (mid_1[2391:2384] < btm_2[2391:2384]) ? 1 : 0;
assign detect_min[297][25] = (mid_1[2391:2384] < btm_2[2399:2392]) ? 1 : 0;

assign detect_min[298][0] = (mid_1[2399:2392] < top_0[2391:2384]) ? 1 : 0;
assign detect_min[298][1] = (mid_1[2399:2392] < top_0[2399:2392]) ? 1 : 0;
assign detect_min[298][2] = (mid_1[2399:2392] < top_0[2407:2400]) ? 1 : 0;
assign detect_min[298][3] = (mid_1[2399:2392] < top_1[2391:2384]) ? 1 : 0;
assign detect_min[298][4] = (mid_1[2399:2392] < top_1[2399:2392]) ? 1 : 0;
assign detect_min[298][5] = (mid_1[2399:2392] < top_1[2407:2400]) ? 1 : 0;
assign detect_min[298][6] = (mid_1[2399:2392] < top_2[2391:2384]) ? 1 : 0;
assign detect_min[298][7] = (mid_1[2399:2392] < top_2[2399:2392]) ? 1 : 0;
assign detect_min[298][8] = (mid_1[2399:2392] < top_2[2407:2400]) ? 1 : 0;
assign detect_min[298][9] = (mid_1[2399:2392] < mid_0[2391:2384]) ? 1 : 0;
assign detect_min[298][10] = (mid_1[2399:2392] < mid_0[2399:2392]) ? 1 : 0;
assign detect_min[298][11] = (mid_1[2399:2392] < mid_0[2407:2400]) ? 1 : 0;
assign detect_min[298][12] = (mid_1[2399:2392] < mid_1[2391:2384]) ? 1 : 0;
assign detect_min[298][13] = (mid_1[2399:2392] < mid_1[2407:2400]) ? 1 : 0;
assign detect_min[298][14] = (mid_1[2399:2392] < mid_2[2391:2384]) ? 1 : 0;
assign detect_min[298][15] = (mid_1[2399:2392] < mid_2[2399:2392]) ? 1 : 0;
assign detect_min[298][16] = (mid_1[2399:2392] < mid_2[2407:2400]) ? 1 : 0;
assign detect_min[298][17] = (mid_1[2399:2392] < btm_0[2391:2384]) ? 1 : 0;
assign detect_min[298][18] = (mid_1[2399:2392] < btm_0[2399:2392]) ? 1 : 0;
assign detect_min[298][19] = (mid_1[2399:2392] < btm_0[2407:2400]) ? 1 : 0;
assign detect_min[298][20] = (mid_1[2399:2392] < btm_1[2391:2384]) ? 1 : 0;
assign detect_min[298][21] = (mid_1[2399:2392] < btm_1[2399:2392]) ? 1 : 0;
assign detect_min[298][22] = (mid_1[2399:2392] < btm_1[2407:2400]) ? 1 : 0;
assign detect_min[298][23] = (mid_1[2399:2392] < btm_2[2391:2384]) ? 1 : 0;
assign detect_min[298][24] = (mid_1[2399:2392] < btm_2[2399:2392]) ? 1 : 0;
assign detect_min[298][25] = (mid_1[2399:2392] < btm_2[2407:2400]) ? 1 : 0;

assign detect_min[299][0] = (mid_1[2407:2400] < top_0[2399:2392]) ? 1 : 0;
assign detect_min[299][1] = (mid_1[2407:2400] < top_0[2407:2400]) ? 1 : 0;
assign detect_min[299][2] = (mid_1[2407:2400] < top_0[2415:2408]) ? 1 : 0;
assign detect_min[299][3] = (mid_1[2407:2400] < top_1[2399:2392]) ? 1 : 0;
assign detect_min[299][4] = (mid_1[2407:2400] < top_1[2407:2400]) ? 1 : 0;
assign detect_min[299][5] = (mid_1[2407:2400] < top_1[2415:2408]) ? 1 : 0;
assign detect_min[299][6] = (mid_1[2407:2400] < top_2[2399:2392]) ? 1 : 0;
assign detect_min[299][7] = (mid_1[2407:2400] < top_2[2407:2400]) ? 1 : 0;
assign detect_min[299][8] = (mid_1[2407:2400] < top_2[2415:2408]) ? 1 : 0;
assign detect_min[299][9] = (mid_1[2407:2400] < mid_0[2399:2392]) ? 1 : 0;
assign detect_min[299][10] = (mid_1[2407:2400] < mid_0[2407:2400]) ? 1 : 0;
assign detect_min[299][11] = (mid_1[2407:2400] < mid_0[2415:2408]) ? 1 : 0;
assign detect_min[299][12] = (mid_1[2407:2400] < mid_1[2399:2392]) ? 1 : 0;
assign detect_min[299][13] = (mid_1[2407:2400] < mid_1[2415:2408]) ? 1 : 0;
assign detect_min[299][14] = (mid_1[2407:2400] < mid_2[2399:2392]) ? 1 : 0;
assign detect_min[299][15] = (mid_1[2407:2400] < mid_2[2407:2400]) ? 1 : 0;
assign detect_min[299][16] = (mid_1[2407:2400] < mid_2[2415:2408]) ? 1 : 0;
assign detect_min[299][17] = (mid_1[2407:2400] < btm_0[2399:2392]) ? 1 : 0;
assign detect_min[299][18] = (mid_1[2407:2400] < btm_0[2407:2400]) ? 1 : 0;
assign detect_min[299][19] = (mid_1[2407:2400] < btm_0[2415:2408]) ? 1 : 0;
assign detect_min[299][20] = (mid_1[2407:2400] < btm_1[2399:2392]) ? 1 : 0;
assign detect_min[299][21] = (mid_1[2407:2400] < btm_1[2407:2400]) ? 1 : 0;
assign detect_min[299][22] = (mid_1[2407:2400] < btm_1[2415:2408]) ? 1 : 0;
assign detect_min[299][23] = (mid_1[2407:2400] < btm_2[2399:2392]) ? 1 : 0;
assign detect_min[299][24] = (mid_1[2407:2400] < btm_2[2407:2400]) ? 1 : 0;
assign detect_min[299][25] = (mid_1[2407:2400] < btm_2[2415:2408]) ? 1 : 0;

assign detect_min[300][0] = (mid_1[2415:2408] < top_0[2407:2400]) ? 1 : 0;
assign detect_min[300][1] = (mid_1[2415:2408] < top_0[2415:2408]) ? 1 : 0;
assign detect_min[300][2] = (mid_1[2415:2408] < top_0[2423:2416]) ? 1 : 0;
assign detect_min[300][3] = (mid_1[2415:2408] < top_1[2407:2400]) ? 1 : 0;
assign detect_min[300][4] = (mid_1[2415:2408] < top_1[2415:2408]) ? 1 : 0;
assign detect_min[300][5] = (mid_1[2415:2408] < top_1[2423:2416]) ? 1 : 0;
assign detect_min[300][6] = (mid_1[2415:2408] < top_2[2407:2400]) ? 1 : 0;
assign detect_min[300][7] = (mid_1[2415:2408] < top_2[2415:2408]) ? 1 : 0;
assign detect_min[300][8] = (mid_1[2415:2408] < top_2[2423:2416]) ? 1 : 0;
assign detect_min[300][9] = (mid_1[2415:2408] < mid_0[2407:2400]) ? 1 : 0;
assign detect_min[300][10] = (mid_1[2415:2408] < mid_0[2415:2408]) ? 1 : 0;
assign detect_min[300][11] = (mid_1[2415:2408] < mid_0[2423:2416]) ? 1 : 0;
assign detect_min[300][12] = (mid_1[2415:2408] < mid_1[2407:2400]) ? 1 : 0;
assign detect_min[300][13] = (mid_1[2415:2408] < mid_1[2423:2416]) ? 1 : 0;
assign detect_min[300][14] = (mid_1[2415:2408] < mid_2[2407:2400]) ? 1 : 0;
assign detect_min[300][15] = (mid_1[2415:2408] < mid_2[2415:2408]) ? 1 : 0;
assign detect_min[300][16] = (mid_1[2415:2408] < mid_2[2423:2416]) ? 1 : 0;
assign detect_min[300][17] = (mid_1[2415:2408] < btm_0[2407:2400]) ? 1 : 0;
assign detect_min[300][18] = (mid_1[2415:2408] < btm_0[2415:2408]) ? 1 : 0;
assign detect_min[300][19] = (mid_1[2415:2408] < btm_0[2423:2416]) ? 1 : 0;
assign detect_min[300][20] = (mid_1[2415:2408] < btm_1[2407:2400]) ? 1 : 0;
assign detect_min[300][21] = (mid_1[2415:2408] < btm_1[2415:2408]) ? 1 : 0;
assign detect_min[300][22] = (mid_1[2415:2408] < btm_1[2423:2416]) ? 1 : 0;
assign detect_min[300][23] = (mid_1[2415:2408] < btm_2[2407:2400]) ? 1 : 0;
assign detect_min[300][24] = (mid_1[2415:2408] < btm_2[2415:2408]) ? 1 : 0;
assign detect_min[300][25] = (mid_1[2415:2408] < btm_2[2423:2416]) ? 1 : 0;

assign detect_min[301][0] = (mid_1[2423:2416] < top_0[2415:2408]) ? 1 : 0;
assign detect_min[301][1] = (mid_1[2423:2416] < top_0[2423:2416]) ? 1 : 0;
assign detect_min[301][2] = (mid_1[2423:2416] < top_0[2431:2424]) ? 1 : 0;
assign detect_min[301][3] = (mid_1[2423:2416] < top_1[2415:2408]) ? 1 : 0;
assign detect_min[301][4] = (mid_1[2423:2416] < top_1[2423:2416]) ? 1 : 0;
assign detect_min[301][5] = (mid_1[2423:2416] < top_1[2431:2424]) ? 1 : 0;
assign detect_min[301][6] = (mid_1[2423:2416] < top_2[2415:2408]) ? 1 : 0;
assign detect_min[301][7] = (mid_1[2423:2416] < top_2[2423:2416]) ? 1 : 0;
assign detect_min[301][8] = (mid_1[2423:2416] < top_2[2431:2424]) ? 1 : 0;
assign detect_min[301][9] = (mid_1[2423:2416] < mid_0[2415:2408]) ? 1 : 0;
assign detect_min[301][10] = (mid_1[2423:2416] < mid_0[2423:2416]) ? 1 : 0;
assign detect_min[301][11] = (mid_1[2423:2416] < mid_0[2431:2424]) ? 1 : 0;
assign detect_min[301][12] = (mid_1[2423:2416] < mid_1[2415:2408]) ? 1 : 0;
assign detect_min[301][13] = (mid_1[2423:2416] < mid_1[2431:2424]) ? 1 : 0;
assign detect_min[301][14] = (mid_1[2423:2416] < mid_2[2415:2408]) ? 1 : 0;
assign detect_min[301][15] = (mid_1[2423:2416] < mid_2[2423:2416]) ? 1 : 0;
assign detect_min[301][16] = (mid_1[2423:2416] < mid_2[2431:2424]) ? 1 : 0;
assign detect_min[301][17] = (mid_1[2423:2416] < btm_0[2415:2408]) ? 1 : 0;
assign detect_min[301][18] = (mid_1[2423:2416] < btm_0[2423:2416]) ? 1 : 0;
assign detect_min[301][19] = (mid_1[2423:2416] < btm_0[2431:2424]) ? 1 : 0;
assign detect_min[301][20] = (mid_1[2423:2416] < btm_1[2415:2408]) ? 1 : 0;
assign detect_min[301][21] = (mid_1[2423:2416] < btm_1[2423:2416]) ? 1 : 0;
assign detect_min[301][22] = (mid_1[2423:2416] < btm_1[2431:2424]) ? 1 : 0;
assign detect_min[301][23] = (mid_1[2423:2416] < btm_2[2415:2408]) ? 1 : 0;
assign detect_min[301][24] = (mid_1[2423:2416] < btm_2[2423:2416]) ? 1 : 0;
assign detect_min[301][25] = (mid_1[2423:2416] < btm_2[2431:2424]) ? 1 : 0;

assign detect_min[302][0] = (mid_1[2431:2424] < top_0[2423:2416]) ? 1 : 0;
assign detect_min[302][1] = (mid_1[2431:2424] < top_0[2431:2424]) ? 1 : 0;
assign detect_min[302][2] = (mid_1[2431:2424] < top_0[2439:2432]) ? 1 : 0;
assign detect_min[302][3] = (mid_1[2431:2424] < top_1[2423:2416]) ? 1 : 0;
assign detect_min[302][4] = (mid_1[2431:2424] < top_1[2431:2424]) ? 1 : 0;
assign detect_min[302][5] = (mid_1[2431:2424] < top_1[2439:2432]) ? 1 : 0;
assign detect_min[302][6] = (mid_1[2431:2424] < top_2[2423:2416]) ? 1 : 0;
assign detect_min[302][7] = (mid_1[2431:2424] < top_2[2431:2424]) ? 1 : 0;
assign detect_min[302][8] = (mid_1[2431:2424] < top_2[2439:2432]) ? 1 : 0;
assign detect_min[302][9] = (mid_1[2431:2424] < mid_0[2423:2416]) ? 1 : 0;
assign detect_min[302][10] = (mid_1[2431:2424] < mid_0[2431:2424]) ? 1 : 0;
assign detect_min[302][11] = (mid_1[2431:2424] < mid_0[2439:2432]) ? 1 : 0;
assign detect_min[302][12] = (mid_1[2431:2424] < mid_1[2423:2416]) ? 1 : 0;
assign detect_min[302][13] = (mid_1[2431:2424] < mid_1[2439:2432]) ? 1 : 0;
assign detect_min[302][14] = (mid_1[2431:2424] < mid_2[2423:2416]) ? 1 : 0;
assign detect_min[302][15] = (mid_1[2431:2424] < mid_2[2431:2424]) ? 1 : 0;
assign detect_min[302][16] = (mid_1[2431:2424] < mid_2[2439:2432]) ? 1 : 0;
assign detect_min[302][17] = (mid_1[2431:2424] < btm_0[2423:2416]) ? 1 : 0;
assign detect_min[302][18] = (mid_1[2431:2424] < btm_0[2431:2424]) ? 1 : 0;
assign detect_min[302][19] = (mid_1[2431:2424] < btm_0[2439:2432]) ? 1 : 0;
assign detect_min[302][20] = (mid_1[2431:2424] < btm_1[2423:2416]) ? 1 : 0;
assign detect_min[302][21] = (mid_1[2431:2424] < btm_1[2431:2424]) ? 1 : 0;
assign detect_min[302][22] = (mid_1[2431:2424] < btm_1[2439:2432]) ? 1 : 0;
assign detect_min[302][23] = (mid_1[2431:2424] < btm_2[2423:2416]) ? 1 : 0;
assign detect_min[302][24] = (mid_1[2431:2424] < btm_2[2431:2424]) ? 1 : 0;
assign detect_min[302][25] = (mid_1[2431:2424] < btm_2[2439:2432]) ? 1 : 0;

assign detect_min[303][0] = (mid_1[2439:2432] < top_0[2431:2424]) ? 1 : 0;
assign detect_min[303][1] = (mid_1[2439:2432] < top_0[2439:2432]) ? 1 : 0;
assign detect_min[303][2] = (mid_1[2439:2432] < top_0[2447:2440]) ? 1 : 0;
assign detect_min[303][3] = (mid_1[2439:2432] < top_1[2431:2424]) ? 1 : 0;
assign detect_min[303][4] = (mid_1[2439:2432] < top_1[2439:2432]) ? 1 : 0;
assign detect_min[303][5] = (mid_1[2439:2432] < top_1[2447:2440]) ? 1 : 0;
assign detect_min[303][6] = (mid_1[2439:2432] < top_2[2431:2424]) ? 1 : 0;
assign detect_min[303][7] = (mid_1[2439:2432] < top_2[2439:2432]) ? 1 : 0;
assign detect_min[303][8] = (mid_1[2439:2432] < top_2[2447:2440]) ? 1 : 0;
assign detect_min[303][9] = (mid_1[2439:2432] < mid_0[2431:2424]) ? 1 : 0;
assign detect_min[303][10] = (mid_1[2439:2432] < mid_0[2439:2432]) ? 1 : 0;
assign detect_min[303][11] = (mid_1[2439:2432] < mid_0[2447:2440]) ? 1 : 0;
assign detect_min[303][12] = (mid_1[2439:2432] < mid_1[2431:2424]) ? 1 : 0;
assign detect_min[303][13] = (mid_1[2439:2432] < mid_1[2447:2440]) ? 1 : 0;
assign detect_min[303][14] = (mid_1[2439:2432] < mid_2[2431:2424]) ? 1 : 0;
assign detect_min[303][15] = (mid_1[2439:2432] < mid_2[2439:2432]) ? 1 : 0;
assign detect_min[303][16] = (mid_1[2439:2432] < mid_2[2447:2440]) ? 1 : 0;
assign detect_min[303][17] = (mid_1[2439:2432] < btm_0[2431:2424]) ? 1 : 0;
assign detect_min[303][18] = (mid_1[2439:2432] < btm_0[2439:2432]) ? 1 : 0;
assign detect_min[303][19] = (mid_1[2439:2432] < btm_0[2447:2440]) ? 1 : 0;
assign detect_min[303][20] = (mid_1[2439:2432] < btm_1[2431:2424]) ? 1 : 0;
assign detect_min[303][21] = (mid_1[2439:2432] < btm_1[2439:2432]) ? 1 : 0;
assign detect_min[303][22] = (mid_1[2439:2432] < btm_1[2447:2440]) ? 1 : 0;
assign detect_min[303][23] = (mid_1[2439:2432] < btm_2[2431:2424]) ? 1 : 0;
assign detect_min[303][24] = (mid_1[2439:2432] < btm_2[2439:2432]) ? 1 : 0;
assign detect_min[303][25] = (mid_1[2439:2432] < btm_2[2447:2440]) ? 1 : 0;

assign detect_min[304][0] = (mid_1[2447:2440] < top_0[2439:2432]) ? 1 : 0;
assign detect_min[304][1] = (mid_1[2447:2440] < top_0[2447:2440]) ? 1 : 0;
assign detect_min[304][2] = (mid_1[2447:2440] < top_0[2455:2448]) ? 1 : 0;
assign detect_min[304][3] = (mid_1[2447:2440] < top_1[2439:2432]) ? 1 : 0;
assign detect_min[304][4] = (mid_1[2447:2440] < top_1[2447:2440]) ? 1 : 0;
assign detect_min[304][5] = (mid_1[2447:2440] < top_1[2455:2448]) ? 1 : 0;
assign detect_min[304][6] = (mid_1[2447:2440] < top_2[2439:2432]) ? 1 : 0;
assign detect_min[304][7] = (mid_1[2447:2440] < top_2[2447:2440]) ? 1 : 0;
assign detect_min[304][8] = (mid_1[2447:2440] < top_2[2455:2448]) ? 1 : 0;
assign detect_min[304][9] = (mid_1[2447:2440] < mid_0[2439:2432]) ? 1 : 0;
assign detect_min[304][10] = (mid_1[2447:2440] < mid_0[2447:2440]) ? 1 : 0;
assign detect_min[304][11] = (mid_1[2447:2440] < mid_0[2455:2448]) ? 1 : 0;
assign detect_min[304][12] = (mid_1[2447:2440] < mid_1[2439:2432]) ? 1 : 0;
assign detect_min[304][13] = (mid_1[2447:2440] < mid_1[2455:2448]) ? 1 : 0;
assign detect_min[304][14] = (mid_1[2447:2440] < mid_2[2439:2432]) ? 1 : 0;
assign detect_min[304][15] = (mid_1[2447:2440] < mid_2[2447:2440]) ? 1 : 0;
assign detect_min[304][16] = (mid_1[2447:2440] < mid_2[2455:2448]) ? 1 : 0;
assign detect_min[304][17] = (mid_1[2447:2440] < btm_0[2439:2432]) ? 1 : 0;
assign detect_min[304][18] = (mid_1[2447:2440] < btm_0[2447:2440]) ? 1 : 0;
assign detect_min[304][19] = (mid_1[2447:2440] < btm_0[2455:2448]) ? 1 : 0;
assign detect_min[304][20] = (mid_1[2447:2440] < btm_1[2439:2432]) ? 1 : 0;
assign detect_min[304][21] = (mid_1[2447:2440] < btm_1[2447:2440]) ? 1 : 0;
assign detect_min[304][22] = (mid_1[2447:2440] < btm_1[2455:2448]) ? 1 : 0;
assign detect_min[304][23] = (mid_1[2447:2440] < btm_2[2439:2432]) ? 1 : 0;
assign detect_min[304][24] = (mid_1[2447:2440] < btm_2[2447:2440]) ? 1 : 0;
assign detect_min[304][25] = (mid_1[2447:2440] < btm_2[2455:2448]) ? 1 : 0;

assign detect_min[305][0] = (mid_1[2455:2448] < top_0[2447:2440]) ? 1 : 0;
assign detect_min[305][1] = (mid_1[2455:2448] < top_0[2455:2448]) ? 1 : 0;
assign detect_min[305][2] = (mid_1[2455:2448] < top_0[2463:2456]) ? 1 : 0;
assign detect_min[305][3] = (mid_1[2455:2448] < top_1[2447:2440]) ? 1 : 0;
assign detect_min[305][4] = (mid_1[2455:2448] < top_1[2455:2448]) ? 1 : 0;
assign detect_min[305][5] = (mid_1[2455:2448] < top_1[2463:2456]) ? 1 : 0;
assign detect_min[305][6] = (mid_1[2455:2448] < top_2[2447:2440]) ? 1 : 0;
assign detect_min[305][7] = (mid_1[2455:2448] < top_2[2455:2448]) ? 1 : 0;
assign detect_min[305][8] = (mid_1[2455:2448] < top_2[2463:2456]) ? 1 : 0;
assign detect_min[305][9] = (mid_1[2455:2448] < mid_0[2447:2440]) ? 1 : 0;
assign detect_min[305][10] = (mid_1[2455:2448] < mid_0[2455:2448]) ? 1 : 0;
assign detect_min[305][11] = (mid_1[2455:2448] < mid_0[2463:2456]) ? 1 : 0;
assign detect_min[305][12] = (mid_1[2455:2448] < mid_1[2447:2440]) ? 1 : 0;
assign detect_min[305][13] = (mid_1[2455:2448] < mid_1[2463:2456]) ? 1 : 0;
assign detect_min[305][14] = (mid_1[2455:2448] < mid_2[2447:2440]) ? 1 : 0;
assign detect_min[305][15] = (mid_1[2455:2448] < mid_2[2455:2448]) ? 1 : 0;
assign detect_min[305][16] = (mid_1[2455:2448] < mid_2[2463:2456]) ? 1 : 0;
assign detect_min[305][17] = (mid_1[2455:2448] < btm_0[2447:2440]) ? 1 : 0;
assign detect_min[305][18] = (mid_1[2455:2448] < btm_0[2455:2448]) ? 1 : 0;
assign detect_min[305][19] = (mid_1[2455:2448] < btm_0[2463:2456]) ? 1 : 0;
assign detect_min[305][20] = (mid_1[2455:2448] < btm_1[2447:2440]) ? 1 : 0;
assign detect_min[305][21] = (mid_1[2455:2448] < btm_1[2455:2448]) ? 1 : 0;
assign detect_min[305][22] = (mid_1[2455:2448] < btm_1[2463:2456]) ? 1 : 0;
assign detect_min[305][23] = (mid_1[2455:2448] < btm_2[2447:2440]) ? 1 : 0;
assign detect_min[305][24] = (mid_1[2455:2448] < btm_2[2455:2448]) ? 1 : 0;
assign detect_min[305][25] = (mid_1[2455:2448] < btm_2[2463:2456]) ? 1 : 0;

assign detect_min[306][0] = (mid_1[2463:2456] < top_0[2455:2448]) ? 1 : 0;
assign detect_min[306][1] = (mid_1[2463:2456] < top_0[2463:2456]) ? 1 : 0;
assign detect_min[306][2] = (mid_1[2463:2456] < top_0[2471:2464]) ? 1 : 0;
assign detect_min[306][3] = (mid_1[2463:2456] < top_1[2455:2448]) ? 1 : 0;
assign detect_min[306][4] = (mid_1[2463:2456] < top_1[2463:2456]) ? 1 : 0;
assign detect_min[306][5] = (mid_1[2463:2456] < top_1[2471:2464]) ? 1 : 0;
assign detect_min[306][6] = (mid_1[2463:2456] < top_2[2455:2448]) ? 1 : 0;
assign detect_min[306][7] = (mid_1[2463:2456] < top_2[2463:2456]) ? 1 : 0;
assign detect_min[306][8] = (mid_1[2463:2456] < top_2[2471:2464]) ? 1 : 0;
assign detect_min[306][9] = (mid_1[2463:2456] < mid_0[2455:2448]) ? 1 : 0;
assign detect_min[306][10] = (mid_1[2463:2456] < mid_0[2463:2456]) ? 1 : 0;
assign detect_min[306][11] = (mid_1[2463:2456] < mid_0[2471:2464]) ? 1 : 0;
assign detect_min[306][12] = (mid_1[2463:2456] < mid_1[2455:2448]) ? 1 : 0;
assign detect_min[306][13] = (mid_1[2463:2456] < mid_1[2471:2464]) ? 1 : 0;
assign detect_min[306][14] = (mid_1[2463:2456] < mid_2[2455:2448]) ? 1 : 0;
assign detect_min[306][15] = (mid_1[2463:2456] < mid_2[2463:2456]) ? 1 : 0;
assign detect_min[306][16] = (mid_1[2463:2456] < mid_2[2471:2464]) ? 1 : 0;
assign detect_min[306][17] = (mid_1[2463:2456] < btm_0[2455:2448]) ? 1 : 0;
assign detect_min[306][18] = (mid_1[2463:2456] < btm_0[2463:2456]) ? 1 : 0;
assign detect_min[306][19] = (mid_1[2463:2456] < btm_0[2471:2464]) ? 1 : 0;
assign detect_min[306][20] = (mid_1[2463:2456] < btm_1[2455:2448]) ? 1 : 0;
assign detect_min[306][21] = (mid_1[2463:2456] < btm_1[2463:2456]) ? 1 : 0;
assign detect_min[306][22] = (mid_1[2463:2456] < btm_1[2471:2464]) ? 1 : 0;
assign detect_min[306][23] = (mid_1[2463:2456] < btm_2[2455:2448]) ? 1 : 0;
assign detect_min[306][24] = (mid_1[2463:2456] < btm_2[2463:2456]) ? 1 : 0;
assign detect_min[306][25] = (mid_1[2463:2456] < btm_2[2471:2464]) ? 1 : 0;

assign detect_min[307][0] = (mid_1[2471:2464] < top_0[2463:2456]) ? 1 : 0;
assign detect_min[307][1] = (mid_1[2471:2464] < top_0[2471:2464]) ? 1 : 0;
assign detect_min[307][2] = (mid_1[2471:2464] < top_0[2479:2472]) ? 1 : 0;
assign detect_min[307][3] = (mid_1[2471:2464] < top_1[2463:2456]) ? 1 : 0;
assign detect_min[307][4] = (mid_1[2471:2464] < top_1[2471:2464]) ? 1 : 0;
assign detect_min[307][5] = (mid_1[2471:2464] < top_1[2479:2472]) ? 1 : 0;
assign detect_min[307][6] = (mid_1[2471:2464] < top_2[2463:2456]) ? 1 : 0;
assign detect_min[307][7] = (mid_1[2471:2464] < top_2[2471:2464]) ? 1 : 0;
assign detect_min[307][8] = (mid_1[2471:2464] < top_2[2479:2472]) ? 1 : 0;
assign detect_min[307][9] = (mid_1[2471:2464] < mid_0[2463:2456]) ? 1 : 0;
assign detect_min[307][10] = (mid_1[2471:2464] < mid_0[2471:2464]) ? 1 : 0;
assign detect_min[307][11] = (mid_1[2471:2464] < mid_0[2479:2472]) ? 1 : 0;
assign detect_min[307][12] = (mid_1[2471:2464] < mid_1[2463:2456]) ? 1 : 0;
assign detect_min[307][13] = (mid_1[2471:2464] < mid_1[2479:2472]) ? 1 : 0;
assign detect_min[307][14] = (mid_1[2471:2464] < mid_2[2463:2456]) ? 1 : 0;
assign detect_min[307][15] = (mid_1[2471:2464] < mid_2[2471:2464]) ? 1 : 0;
assign detect_min[307][16] = (mid_1[2471:2464] < mid_2[2479:2472]) ? 1 : 0;
assign detect_min[307][17] = (mid_1[2471:2464] < btm_0[2463:2456]) ? 1 : 0;
assign detect_min[307][18] = (mid_1[2471:2464] < btm_0[2471:2464]) ? 1 : 0;
assign detect_min[307][19] = (mid_1[2471:2464] < btm_0[2479:2472]) ? 1 : 0;
assign detect_min[307][20] = (mid_1[2471:2464] < btm_1[2463:2456]) ? 1 : 0;
assign detect_min[307][21] = (mid_1[2471:2464] < btm_1[2471:2464]) ? 1 : 0;
assign detect_min[307][22] = (mid_1[2471:2464] < btm_1[2479:2472]) ? 1 : 0;
assign detect_min[307][23] = (mid_1[2471:2464] < btm_2[2463:2456]) ? 1 : 0;
assign detect_min[307][24] = (mid_1[2471:2464] < btm_2[2471:2464]) ? 1 : 0;
assign detect_min[307][25] = (mid_1[2471:2464] < btm_2[2479:2472]) ? 1 : 0;

assign detect_min[308][0] = (mid_1[2479:2472] < top_0[2471:2464]) ? 1 : 0;
assign detect_min[308][1] = (mid_1[2479:2472] < top_0[2479:2472]) ? 1 : 0;
assign detect_min[308][2] = (mid_1[2479:2472] < top_0[2487:2480]) ? 1 : 0;
assign detect_min[308][3] = (mid_1[2479:2472] < top_1[2471:2464]) ? 1 : 0;
assign detect_min[308][4] = (mid_1[2479:2472] < top_1[2479:2472]) ? 1 : 0;
assign detect_min[308][5] = (mid_1[2479:2472] < top_1[2487:2480]) ? 1 : 0;
assign detect_min[308][6] = (mid_1[2479:2472] < top_2[2471:2464]) ? 1 : 0;
assign detect_min[308][7] = (mid_1[2479:2472] < top_2[2479:2472]) ? 1 : 0;
assign detect_min[308][8] = (mid_1[2479:2472] < top_2[2487:2480]) ? 1 : 0;
assign detect_min[308][9] = (mid_1[2479:2472] < mid_0[2471:2464]) ? 1 : 0;
assign detect_min[308][10] = (mid_1[2479:2472] < mid_0[2479:2472]) ? 1 : 0;
assign detect_min[308][11] = (mid_1[2479:2472] < mid_0[2487:2480]) ? 1 : 0;
assign detect_min[308][12] = (mid_1[2479:2472] < mid_1[2471:2464]) ? 1 : 0;
assign detect_min[308][13] = (mid_1[2479:2472] < mid_1[2487:2480]) ? 1 : 0;
assign detect_min[308][14] = (mid_1[2479:2472] < mid_2[2471:2464]) ? 1 : 0;
assign detect_min[308][15] = (mid_1[2479:2472] < mid_2[2479:2472]) ? 1 : 0;
assign detect_min[308][16] = (mid_1[2479:2472] < mid_2[2487:2480]) ? 1 : 0;
assign detect_min[308][17] = (mid_1[2479:2472] < btm_0[2471:2464]) ? 1 : 0;
assign detect_min[308][18] = (mid_1[2479:2472] < btm_0[2479:2472]) ? 1 : 0;
assign detect_min[308][19] = (mid_1[2479:2472] < btm_0[2487:2480]) ? 1 : 0;
assign detect_min[308][20] = (mid_1[2479:2472] < btm_1[2471:2464]) ? 1 : 0;
assign detect_min[308][21] = (mid_1[2479:2472] < btm_1[2479:2472]) ? 1 : 0;
assign detect_min[308][22] = (mid_1[2479:2472] < btm_1[2487:2480]) ? 1 : 0;
assign detect_min[308][23] = (mid_1[2479:2472] < btm_2[2471:2464]) ? 1 : 0;
assign detect_min[308][24] = (mid_1[2479:2472] < btm_2[2479:2472]) ? 1 : 0;
assign detect_min[308][25] = (mid_1[2479:2472] < btm_2[2487:2480]) ? 1 : 0;

assign detect_min[309][0] = (mid_1[2487:2480] < top_0[2479:2472]) ? 1 : 0;
assign detect_min[309][1] = (mid_1[2487:2480] < top_0[2487:2480]) ? 1 : 0;
assign detect_min[309][2] = (mid_1[2487:2480] < top_0[2495:2488]) ? 1 : 0;
assign detect_min[309][3] = (mid_1[2487:2480] < top_1[2479:2472]) ? 1 : 0;
assign detect_min[309][4] = (mid_1[2487:2480] < top_1[2487:2480]) ? 1 : 0;
assign detect_min[309][5] = (mid_1[2487:2480] < top_1[2495:2488]) ? 1 : 0;
assign detect_min[309][6] = (mid_1[2487:2480] < top_2[2479:2472]) ? 1 : 0;
assign detect_min[309][7] = (mid_1[2487:2480] < top_2[2487:2480]) ? 1 : 0;
assign detect_min[309][8] = (mid_1[2487:2480] < top_2[2495:2488]) ? 1 : 0;
assign detect_min[309][9] = (mid_1[2487:2480] < mid_0[2479:2472]) ? 1 : 0;
assign detect_min[309][10] = (mid_1[2487:2480] < mid_0[2487:2480]) ? 1 : 0;
assign detect_min[309][11] = (mid_1[2487:2480] < mid_0[2495:2488]) ? 1 : 0;
assign detect_min[309][12] = (mid_1[2487:2480] < mid_1[2479:2472]) ? 1 : 0;
assign detect_min[309][13] = (mid_1[2487:2480] < mid_1[2495:2488]) ? 1 : 0;
assign detect_min[309][14] = (mid_1[2487:2480] < mid_2[2479:2472]) ? 1 : 0;
assign detect_min[309][15] = (mid_1[2487:2480] < mid_2[2487:2480]) ? 1 : 0;
assign detect_min[309][16] = (mid_1[2487:2480] < mid_2[2495:2488]) ? 1 : 0;
assign detect_min[309][17] = (mid_1[2487:2480] < btm_0[2479:2472]) ? 1 : 0;
assign detect_min[309][18] = (mid_1[2487:2480] < btm_0[2487:2480]) ? 1 : 0;
assign detect_min[309][19] = (mid_1[2487:2480] < btm_0[2495:2488]) ? 1 : 0;
assign detect_min[309][20] = (mid_1[2487:2480] < btm_1[2479:2472]) ? 1 : 0;
assign detect_min[309][21] = (mid_1[2487:2480] < btm_1[2487:2480]) ? 1 : 0;
assign detect_min[309][22] = (mid_1[2487:2480] < btm_1[2495:2488]) ? 1 : 0;
assign detect_min[309][23] = (mid_1[2487:2480] < btm_2[2479:2472]) ? 1 : 0;
assign detect_min[309][24] = (mid_1[2487:2480] < btm_2[2487:2480]) ? 1 : 0;
assign detect_min[309][25] = (mid_1[2487:2480] < btm_2[2495:2488]) ? 1 : 0;

assign detect_min[310][0] = (mid_1[2495:2488] < top_0[2487:2480]) ? 1 : 0;
assign detect_min[310][1] = (mid_1[2495:2488] < top_0[2495:2488]) ? 1 : 0;
assign detect_min[310][2] = (mid_1[2495:2488] < top_0[2503:2496]) ? 1 : 0;
assign detect_min[310][3] = (mid_1[2495:2488] < top_1[2487:2480]) ? 1 : 0;
assign detect_min[310][4] = (mid_1[2495:2488] < top_1[2495:2488]) ? 1 : 0;
assign detect_min[310][5] = (mid_1[2495:2488] < top_1[2503:2496]) ? 1 : 0;
assign detect_min[310][6] = (mid_1[2495:2488] < top_2[2487:2480]) ? 1 : 0;
assign detect_min[310][7] = (mid_1[2495:2488] < top_2[2495:2488]) ? 1 : 0;
assign detect_min[310][8] = (mid_1[2495:2488] < top_2[2503:2496]) ? 1 : 0;
assign detect_min[310][9] = (mid_1[2495:2488] < mid_0[2487:2480]) ? 1 : 0;
assign detect_min[310][10] = (mid_1[2495:2488] < mid_0[2495:2488]) ? 1 : 0;
assign detect_min[310][11] = (mid_1[2495:2488] < mid_0[2503:2496]) ? 1 : 0;
assign detect_min[310][12] = (mid_1[2495:2488] < mid_1[2487:2480]) ? 1 : 0;
assign detect_min[310][13] = (mid_1[2495:2488] < mid_1[2503:2496]) ? 1 : 0;
assign detect_min[310][14] = (mid_1[2495:2488] < mid_2[2487:2480]) ? 1 : 0;
assign detect_min[310][15] = (mid_1[2495:2488] < mid_2[2495:2488]) ? 1 : 0;
assign detect_min[310][16] = (mid_1[2495:2488] < mid_2[2503:2496]) ? 1 : 0;
assign detect_min[310][17] = (mid_1[2495:2488] < btm_0[2487:2480]) ? 1 : 0;
assign detect_min[310][18] = (mid_1[2495:2488] < btm_0[2495:2488]) ? 1 : 0;
assign detect_min[310][19] = (mid_1[2495:2488] < btm_0[2503:2496]) ? 1 : 0;
assign detect_min[310][20] = (mid_1[2495:2488] < btm_1[2487:2480]) ? 1 : 0;
assign detect_min[310][21] = (mid_1[2495:2488] < btm_1[2495:2488]) ? 1 : 0;
assign detect_min[310][22] = (mid_1[2495:2488] < btm_1[2503:2496]) ? 1 : 0;
assign detect_min[310][23] = (mid_1[2495:2488] < btm_2[2487:2480]) ? 1 : 0;
assign detect_min[310][24] = (mid_1[2495:2488] < btm_2[2495:2488]) ? 1 : 0;
assign detect_min[310][25] = (mid_1[2495:2488] < btm_2[2503:2496]) ? 1 : 0;

assign detect_min[311][0] = (mid_1[2503:2496] < top_0[2495:2488]) ? 1 : 0;
assign detect_min[311][1] = (mid_1[2503:2496] < top_0[2503:2496]) ? 1 : 0;
assign detect_min[311][2] = (mid_1[2503:2496] < top_0[2511:2504]) ? 1 : 0;
assign detect_min[311][3] = (mid_1[2503:2496] < top_1[2495:2488]) ? 1 : 0;
assign detect_min[311][4] = (mid_1[2503:2496] < top_1[2503:2496]) ? 1 : 0;
assign detect_min[311][5] = (mid_1[2503:2496] < top_1[2511:2504]) ? 1 : 0;
assign detect_min[311][6] = (mid_1[2503:2496] < top_2[2495:2488]) ? 1 : 0;
assign detect_min[311][7] = (mid_1[2503:2496] < top_2[2503:2496]) ? 1 : 0;
assign detect_min[311][8] = (mid_1[2503:2496] < top_2[2511:2504]) ? 1 : 0;
assign detect_min[311][9] = (mid_1[2503:2496] < mid_0[2495:2488]) ? 1 : 0;
assign detect_min[311][10] = (mid_1[2503:2496] < mid_0[2503:2496]) ? 1 : 0;
assign detect_min[311][11] = (mid_1[2503:2496] < mid_0[2511:2504]) ? 1 : 0;
assign detect_min[311][12] = (mid_1[2503:2496] < mid_1[2495:2488]) ? 1 : 0;
assign detect_min[311][13] = (mid_1[2503:2496] < mid_1[2511:2504]) ? 1 : 0;
assign detect_min[311][14] = (mid_1[2503:2496] < mid_2[2495:2488]) ? 1 : 0;
assign detect_min[311][15] = (mid_1[2503:2496] < mid_2[2503:2496]) ? 1 : 0;
assign detect_min[311][16] = (mid_1[2503:2496] < mid_2[2511:2504]) ? 1 : 0;
assign detect_min[311][17] = (mid_1[2503:2496] < btm_0[2495:2488]) ? 1 : 0;
assign detect_min[311][18] = (mid_1[2503:2496] < btm_0[2503:2496]) ? 1 : 0;
assign detect_min[311][19] = (mid_1[2503:2496] < btm_0[2511:2504]) ? 1 : 0;
assign detect_min[311][20] = (mid_1[2503:2496] < btm_1[2495:2488]) ? 1 : 0;
assign detect_min[311][21] = (mid_1[2503:2496] < btm_1[2503:2496]) ? 1 : 0;
assign detect_min[311][22] = (mid_1[2503:2496] < btm_1[2511:2504]) ? 1 : 0;
assign detect_min[311][23] = (mid_1[2503:2496] < btm_2[2495:2488]) ? 1 : 0;
assign detect_min[311][24] = (mid_1[2503:2496] < btm_2[2503:2496]) ? 1 : 0;
assign detect_min[311][25] = (mid_1[2503:2496] < btm_2[2511:2504]) ? 1 : 0;

assign detect_min[312][0] = (mid_1[2511:2504] < top_0[2503:2496]) ? 1 : 0;
assign detect_min[312][1] = (mid_1[2511:2504] < top_0[2511:2504]) ? 1 : 0;
assign detect_min[312][2] = (mid_1[2511:2504] < top_0[2519:2512]) ? 1 : 0;
assign detect_min[312][3] = (mid_1[2511:2504] < top_1[2503:2496]) ? 1 : 0;
assign detect_min[312][4] = (mid_1[2511:2504] < top_1[2511:2504]) ? 1 : 0;
assign detect_min[312][5] = (mid_1[2511:2504] < top_1[2519:2512]) ? 1 : 0;
assign detect_min[312][6] = (mid_1[2511:2504] < top_2[2503:2496]) ? 1 : 0;
assign detect_min[312][7] = (mid_1[2511:2504] < top_2[2511:2504]) ? 1 : 0;
assign detect_min[312][8] = (mid_1[2511:2504] < top_2[2519:2512]) ? 1 : 0;
assign detect_min[312][9] = (mid_1[2511:2504] < mid_0[2503:2496]) ? 1 : 0;
assign detect_min[312][10] = (mid_1[2511:2504] < mid_0[2511:2504]) ? 1 : 0;
assign detect_min[312][11] = (mid_1[2511:2504] < mid_0[2519:2512]) ? 1 : 0;
assign detect_min[312][12] = (mid_1[2511:2504] < mid_1[2503:2496]) ? 1 : 0;
assign detect_min[312][13] = (mid_1[2511:2504] < mid_1[2519:2512]) ? 1 : 0;
assign detect_min[312][14] = (mid_1[2511:2504] < mid_2[2503:2496]) ? 1 : 0;
assign detect_min[312][15] = (mid_1[2511:2504] < mid_2[2511:2504]) ? 1 : 0;
assign detect_min[312][16] = (mid_1[2511:2504] < mid_2[2519:2512]) ? 1 : 0;
assign detect_min[312][17] = (mid_1[2511:2504] < btm_0[2503:2496]) ? 1 : 0;
assign detect_min[312][18] = (mid_1[2511:2504] < btm_0[2511:2504]) ? 1 : 0;
assign detect_min[312][19] = (mid_1[2511:2504] < btm_0[2519:2512]) ? 1 : 0;
assign detect_min[312][20] = (mid_1[2511:2504] < btm_1[2503:2496]) ? 1 : 0;
assign detect_min[312][21] = (mid_1[2511:2504] < btm_1[2511:2504]) ? 1 : 0;
assign detect_min[312][22] = (mid_1[2511:2504] < btm_1[2519:2512]) ? 1 : 0;
assign detect_min[312][23] = (mid_1[2511:2504] < btm_2[2503:2496]) ? 1 : 0;
assign detect_min[312][24] = (mid_1[2511:2504] < btm_2[2511:2504]) ? 1 : 0;
assign detect_min[312][25] = (mid_1[2511:2504] < btm_2[2519:2512]) ? 1 : 0;

assign detect_min[313][0] = (mid_1[2519:2512] < top_0[2511:2504]) ? 1 : 0;
assign detect_min[313][1] = (mid_1[2519:2512] < top_0[2519:2512]) ? 1 : 0;
assign detect_min[313][2] = (mid_1[2519:2512] < top_0[2527:2520]) ? 1 : 0;
assign detect_min[313][3] = (mid_1[2519:2512] < top_1[2511:2504]) ? 1 : 0;
assign detect_min[313][4] = (mid_1[2519:2512] < top_1[2519:2512]) ? 1 : 0;
assign detect_min[313][5] = (mid_1[2519:2512] < top_1[2527:2520]) ? 1 : 0;
assign detect_min[313][6] = (mid_1[2519:2512] < top_2[2511:2504]) ? 1 : 0;
assign detect_min[313][7] = (mid_1[2519:2512] < top_2[2519:2512]) ? 1 : 0;
assign detect_min[313][8] = (mid_1[2519:2512] < top_2[2527:2520]) ? 1 : 0;
assign detect_min[313][9] = (mid_1[2519:2512] < mid_0[2511:2504]) ? 1 : 0;
assign detect_min[313][10] = (mid_1[2519:2512] < mid_0[2519:2512]) ? 1 : 0;
assign detect_min[313][11] = (mid_1[2519:2512] < mid_0[2527:2520]) ? 1 : 0;
assign detect_min[313][12] = (mid_1[2519:2512] < mid_1[2511:2504]) ? 1 : 0;
assign detect_min[313][13] = (mid_1[2519:2512] < mid_1[2527:2520]) ? 1 : 0;
assign detect_min[313][14] = (mid_1[2519:2512] < mid_2[2511:2504]) ? 1 : 0;
assign detect_min[313][15] = (mid_1[2519:2512] < mid_2[2519:2512]) ? 1 : 0;
assign detect_min[313][16] = (mid_1[2519:2512] < mid_2[2527:2520]) ? 1 : 0;
assign detect_min[313][17] = (mid_1[2519:2512] < btm_0[2511:2504]) ? 1 : 0;
assign detect_min[313][18] = (mid_1[2519:2512] < btm_0[2519:2512]) ? 1 : 0;
assign detect_min[313][19] = (mid_1[2519:2512] < btm_0[2527:2520]) ? 1 : 0;
assign detect_min[313][20] = (mid_1[2519:2512] < btm_1[2511:2504]) ? 1 : 0;
assign detect_min[313][21] = (mid_1[2519:2512] < btm_1[2519:2512]) ? 1 : 0;
assign detect_min[313][22] = (mid_1[2519:2512] < btm_1[2527:2520]) ? 1 : 0;
assign detect_min[313][23] = (mid_1[2519:2512] < btm_2[2511:2504]) ? 1 : 0;
assign detect_min[313][24] = (mid_1[2519:2512] < btm_2[2519:2512]) ? 1 : 0;
assign detect_min[313][25] = (mid_1[2519:2512] < btm_2[2527:2520]) ? 1 : 0;

assign detect_min[314][0] = (mid_1[2527:2520] < top_0[2519:2512]) ? 1 : 0;
assign detect_min[314][1] = (mid_1[2527:2520] < top_0[2527:2520]) ? 1 : 0;
assign detect_min[314][2] = (mid_1[2527:2520] < top_0[2535:2528]) ? 1 : 0;
assign detect_min[314][3] = (mid_1[2527:2520] < top_1[2519:2512]) ? 1 : 0;
assign detect_min[314][4] = (mid_1[2527:2520] < top_1[2527:2520]) ? 1 : 0;
assign detect_min[314][5] = (mid_1[2527:2520] < top_1[2535:2528]) ? 1 : 0;
assign detect_min[314][6] = (mid_1[2527:2520] < top_2[2519:2512]) ? 1 : 0;
assign detect_min[314][7] = (mid_1[2527:2520] < top_2[2527:2520]) ? 1 : 0;
assign detect_min[314][8] = (mid_1[2527:2520] < top_2[2535:2528]) ? 1 : 0;
assign detect_min[314][9] = (mid_1[2527:2520] < mid_0[2519:2512]) ? 1 : 0;
assign detect_min[314][10] = (mid_1[2527:2520] < mid_0[2527:2520]) ? 1 : 0;
assign detect_min[314][11] = (mid_1[2527:2520] < mid_0[2535:2528]) ? 1 : 0;
assign detect_min[314][12] = (mid_1[2527:2520] < mid_1[2519:2512]) ? 1 : 0;
assign detect_min[314][13] = (mid_1[2527:2520] < mid_1[2535:2528]) ? 1 : 0;
assign detect_min[314][14] = (mid_1[2527:2520] < mid_2[2519:2512]) ? 1 : 0;
assign detect_min[314][15] = (mid_1[2527:2520] < mid_2[2527:2520]) ? 1 : 0;
assign detect_min[314][16] = (mid_1[2527:2520] < mid_2[2535:2528]) ? 1 : 0;
assign detect_min[314][17] = (mid_1[2527:2520] < btm_0[2519:2512]) ? 1 : 0;
assign detect_min[314][18] = (mid_1[2527:2520] < btm_0[2527:2520]) ? 1 : 0;
assign detect_min[314][19] = (mid_1[2527:2520] < btm_0[2535:2528]) ? 1 : 0;
assign detect_min[314][20] = (mid_1[2527:2520] < btm_1[2519:2512]) ? 1 : 0;
assign detect_min[314][21] = (mid_1[2527:2520] < btm_1[2527:2520]) ? 1 : 0;
assign detect_min[314][22] = (mid_1[2527:2520] < btm_1[2535:2528]) ? 1 : 0;
assign detect_min[314][23] = (mid_1[2527:2520] < btm_2[2519:2512]) ? 1 : 0;
assign detect_min[314][24] = (mid_1[2527:2520] < btm_2[2527:2520]) ? 1 : 0;
assign detect_min[314][25] = (mid_1[2527:2520] < btm_2[2535:2528]) ? 1 : 0;

assign detect_min[315][0] = (mid_1[2535:2528] < top_0[2527:2520]) ? 1 : 0;
assign detect_min[315][1] = (mid_1[2535:2528] < top_0[2535:2528]) ? 1 : 0;
assign detect_min[315][2] = (mid_1[2535:2528] < top_0[2543:2536]) ? 1 : 0;
assign detect_min[315][3] = (mid_1[2535:2528] < top_1[2527:2520]) ? 1 : 0;
assign detect_min[315][4] = (mid_1[2535:2528] < top_1[2535:2528]) ? 1 : 0;
assign detect_min[315][5] = (mid_1[2535:2528] < top_1[2543:2536]) ? 1 : 0;
assign detect_min[315][6] = (mid_1[2535:2528] < top_2[2527:2520]) ? 1 : 0;
assign detect_min[315][7] = (mid_1[2535:2528] < top_2[2535:2528]) ? 1 : 0;
assign detect_min[315][8] = (mid_1[2535:2528] < top_2[2543:2536]) ? 1 : 0;
assign detect_min[315][9] = (mid_1[2535:2528] < mid_0[2527:2520]) ? 1 : 0;
assign detect_min[315][10] = (mid_1[2535:2528] < mid_0[2535:2528]) ? 1 : 0;
assign detect_min[315][11] = (mid_1[2535:2528] < mid_0[2543:2536]) ? 1 : 0;
assign detect_min[315][12] = (mid_1[2535:2528] < mid_1[2527:2520]) ? 1 : 0;
assign detect_min[315][13] = (mid_1[2535:2528] < mid_1[2543:2536]) ? 1 : 0;
assign detect_min[315][14] = (mid_1[2535:2528] < mid_2[2527:2520]) ? 1 : 0;
assign detect_min[315][15] = (mid_1[2535:2528] < mid_2[2535:2528]) ? 1 : 0;
assign detect_min[315][16] = (mid_1[2535:2528] < mid_2[2543:2536]) ? 1 : 0;
assign detect_min[315][17] = (mid_1[2535:2528] < btm_0[2527:2520]) ? 1 : 0;
assign detect_min[315][18] = (mid_1[2535:2528] < btm_0[2535:2528]) ? 1 : 0;
assign detect_min[315][19] = (mid_1[2535:2528] < btm_0[2543:2536]) ? 1 : 0;
assign detect_min[315][20] = (mid_1[2535:2528] < btm_1[2527:2520]) ? 1 : 0;
assign detect_min[315][21] = (mid_1[2535:2528] < btm_1[2535:2528]) ? 1 : 0;
assign detect_min[315][22] = (mid_1[2535:2528] < btm_1[2543:2536]) ? 1 : 0;
assign detect_min[315][23] = (mid_1[2535:2528] < btm_2[2527:2520]) ? 1 : 0;
assign detect_min[315][24] = (mid_1[2535:2528] < btm_2[2535:2528]) ? 1 : 0;
assign detect_min[315][25] = (mid_1[2535:2528] < btm_2[2543:2536]) ? 1 : 0;

assign detect_min[316][0] = (mid_1[2543:2536] < top_0[2535:2528]) ? 1 : 0;
assign detect_min[316][1] = (mid_1[2543:2536] < top_0[2543:2536]) ? 1 : 0;
assign detect_min[316][2] = (mid_1[2543:2536] < top_0[2551:2544]) ? 1 : 0;
assign detect_min[316][3] = (mid_1[2543:2536] < top_1[2535:2528]) ? 1 : 0;
assign detect_min[316][4] = (mid_1[2543:2536] < top_1[2543:2536]) ? 1 : 0;
assign detect_min[316][5] = (mid_1[2543:2536] < top_1[2551:2544]) ? 1 : 0;
assign detect_min[316][6] = (mid_1[2543:2536] < top_2[2535:2528]) ? 1 : 0;
assign detect_min[316][7] = (mid_1[2543:2536] < top_2[2543:2536]) ? 1 : 0;
assign detect_min[316][8] = (mid_1[2543:2536] < top_2[2551:2544]) ? 1 : 0;
assign detect_min[316][9] = (mid_1[2543:2536] < mid_0[2535:2528]) ? 1 : 0;
assign detect_min[316][10] = (mid_1[2543:2536] < mid_0[2543:2536]) ? 1 : 0;
assign detect_min[316][11] = (mid_1[2543:2536] < mid_0[2551:2544]) ? 1 : 0;
assign detect_min[316][12] = (mid_1[2543:2536] < mid_1[2535:2528]) ? 1 : 0;
assign detect_min[316][13] = (mid_1[2543:2536] < mid_1[2551:2544]) ? 1 : 0;
assign detect_min[316][14] = (mid_1[2543:2536] < mid_2[2535:2528]) ? 1 : 0;
assign detect_min[316][15] = (mid_1[2543:2536] < mid_2[2543:2536]) ? 1 : 0;
assign detect_min[316][16] = (mid_1[2543:2536] < mid_2[2551:2544]) ? 1 : 0;
assign detect_min[316][17] = (mid_1[2543:2536] < btm_0[2535:2528]) ? 1 : 0;
assign detect_min[316][18] = (mid_1[2543:2536] < btm_0[2543:2536]) ? 1 : 0;
assign detect_min[316][19] = (mid_1[2543:2536] < btm_0[2551:2544]) ? 1 : 0;
assign detect_min[316][20] = (mid_1[2543:2536] < btm_1[2535:2528]) ? 1 : 0;
assign detect_min[316][21] = (mid_1[2543:2536] < btm_1[2543:2536]) ? 1 : 0;
assign detect_min[316][22] = (mid_1[2543:2536] < btm_1[2551:2544]) ? 1 : 0;
assign detect_min[316][23] = (mid_1[2543:2536] < btm_2[2535:2528]) ? 1 : 0;
assign detect_min[316][24] = (mid_1[2543:2536] < btm_2[2543:2536]) ? 1 : 0;
assign detect_min[316][25] = (mid_1[2543:2536] < btm_2[2551:2544]) ? 1 : 0;

assign detect_min[317][0] = (mid_1[2551:2544] < top_0[2543:2536]) ? 1 : 0;
assign detect_min[317][1] = (mid_1[2551:2544] < top_0[2551:2544]) ? 1 : 0;
assign detect_min[317][2] = (mid_1[2551:2544] < top_0[2559:2552]) ? 1 : 0;
assign detect_min[317][3] = (mid_1[2551:2544] < top_1[2543:2536]) ? 1 : 0;
assign detect_min[317][4] = (mid_1[2551:2544] < top_1[2551:2544]) ? 1 : 0;
assign detect_min[317][5] = (mid_1[2551:2544] < top_1[2559:2552]) ? 1 : 0;
assign detect_min[317][6] = (mid_1[2551:2544] < top_2[2543:2536]) ? 1 : 0;
assign detect_min[317][7] = (mid_1[2551:2544] < top_2[2551:2544]) ? 1 : 0;
assign detect_min[317][8] = (mid_1[2551:2544] < top_2[2559:2552]) ? 1 : 0;
assign detect_min[317][9] = (mid_1[2551:2544] < mid_0[2543:2536]) ? 1 : 0;
assign detect_min[317][10] = (mid_1[2551:2544] < mid_0[2551:2544]) ? 1 : 0;
assign detect_min[317][11] = (mid_1[2551:2544] < mid_0[2559:2552]) ? 1 : 0;
assign detect_min[317][12] = (mid_1[2551:2544] < mid_1[2543:2536]) ? 1 : 0;
assign detect_min[317][13] = (mid_1[2551:2544] < mid_1[2559:2552]) ? 1 : 0;
assign detect_min[317][14] = (mid_1[2551:2544] < mid_2[2543:2536]) ? 1 : 0;
assign detect_min[317][15] = (mid_1[2551:2544] < mid_2[2551:2544]) ? 1 : 0;
assign detect_min[317][16] = (mid_1[2551:2544] < mid_2[2559:2552]) ? 1 : 0;
assign detect_min[317][17] = (mid_1[2551:2544] < btm_0[2543:2536]) ? 1 : 0;
assign detect_min[317][18] = (mid_1[2551:2544] < btm_0[2551:2544]) ? 1 : 0;
assign detect_min[317][19] = (mid_1[2551:2544] < btm_0[2559:2552]) ? 1 : 0;
assign detect_min[317][20] = (mid_1[2551:2544] < btm_1[2543:2536]) ? 1 : 0;
assign detect_min[317][21] = (mid_1[2551:2544] < btm_1[2551:2544]) ? 1 : 0;
assign detect_min[317][22] = (mid_1[2551:2544] < btm_1[2559:2552]) ? 1 : 0;
assign detect_min[317][23] = (mid_1[2551:2544] < btm_2[2543:2536]) ? 1 : 0;
assign detect_min[317][24] = (mid_1[2551:2544] < btm_2[2551:2544]) ? 1 : 0;
assign detect_min[317][25] = (mid_1[2551:2544] < btm_2[2559:2552]) ? 1 : 0;

assign detect_min[318][0] = (mid_1[2559:2552] < top_0[2551:2544]) ? 1 : 0;
assign detect_min[318][1] = (mid_1[2559:2552] < top_0[2559:2552]) ? 1 : 0;
assign detect_min[318][2] = (mid_1[2559:2552] < top_0[2567:2560]) ? 1 : 0;
assign detect_min[318][3] = (mid_1[2559:2552] < top_1[2551:2544]) ? 1 : 0;
assign detect_min[318][4] = (mid_1[2559:2552] < top_1[2559:2552]) ? 1 : 0;
assign detect_min[318][5] = (mid_1[2559:2552] < top_1[2567:2560]) ? 1 : 0;
assign detect_min[318][6] = (mid_1[2559:2552] < top_2[2551:2544]) ? 1 : 0;
assign detect_min[318][7] = (mid_1[2559:2552] < top_2[2559:2552]) ? 1 : 0;
assign detect_min[318][8] = (mid_1[2559:2552] < top_2[2567:2560]) ? 1 : 0;
assign detect_min[318][9] = (mid_1[2559:2552] < mid_0[2551:2544]) ? 1 : 0;
assign detect_min[318][10] = (mid_1[2559:2552] < mid_0[2559:2552]) ? 1 : 0;
assign detect_min[318][11] = (mid_1[2559:2552] < mid_0[2567:2560]) ? 1 : 0;
assign detect_min[318][12] = (mid_1[2559:2552] < mid_1[2551:2544]) ? 1 : 0;
assign detect_min[318][13] = (mid_1[2559:2552] < mid_1[2567:2560]) ? 1 : 0;
assign detect_min[318][14] = (mid_1[2559:2552] < mid_2[2551:2544]) ? 1 : 0;
assign detect_min[318][15] = (mid_1[2559:2552] < mid_2[2559:2552]) ? 1 : 0;
assign detect_min[318][16] = (mid_1[2559:2552] < mid_2[2567:2560]) ? 1 : 0;
assign detect_min[318][17] = (mid_1[2559:2552] < btm_0[2551:2544]) ? 1 : 0;
assign detect_min[318][18] = (mid_1[2559:2552] < btm_0[2559:2552]) ? 1 : 0;
assign detect_min[318][19] = (mid_1[2559:2552] < btm_0[2567:2560]) ? 1 : 0;
assign detect_min[318][20] = (mid_1[2559:2552] < btm_1[2551:2544]) ? 1 : 0;
assign detect_min[318][21] = (mid_1[2559:2552] < btm_1[2559:2552]) ? 1 : 0;
assign detect_min[318][22] = (mid_1[2559:2552] < btm_1[2567:2560]) ? 1 : 0;
assign detect_min[318][23] = (mid_1[2559:2552] < btm_2[2551:2544]) ? 1 : 0;
assign detect_min[318][24] = (mid_1[2559:2552] < btm_2[2559:2552]) ? 1 : 0;
assign detect_min[318][25] = (mid_1[2559:2552] < btm_2[2567:2560]) ? 1 : 0;

assign detect_min[319][0] = (mid_1[2567:2560] < top_0[2559:2552]) ? 1 : 0;
assign detect_min[319][1] = (mid_1[2567:2560] < top_0[2567:2560]) ? 1 : 0;
assign detect_min[319][2] = (mid_1[2567:2560] < top_0[2575:2568]) ? 1 : 0;
assign detect_min[319][3] = (mid_1[2567:2560] < top_1[2559:2552]) ? 1 : 0;
assign detect_min[319][4] = (mid_1[2567:2560] < top_1[2567:2560]) ? 1 : 0;
assign detect_min[319][5] = (mid_1[2567:2560] < top_1[2575:2568]) ? 1 : 0;
assign detect_min[319][6] = (mid_1[2567:2560] < top_2[2559:2552]) ? 1 : 0;
assign detect_min[319][7] = (mid_1[2567:2560] < top_2[2567:2560]) ? 1 : 0;
assign detect_min[319][8] = (mid_1[2567:2560] < top_2[2575:2568]) ? 1 : 0;
assign detect_min[319][9] = (mid_1[2567:2560] < mid_0[2559:2552]) ? 1 : 0;
assign detect_min[319][10] = (mid_1[2567:2560] < mid_0[2567:2560]) ? 1 : 0;
assign detect_min[319][11] = (mid_1[2567:2560] < mid_0[2575:2568]) ? 1 : 0;
assign detect_min[319][12] = (mid_1[2567:2560] < mid_1[2559:2552]) ? 1 : 0;
assign detect_min[319][13] = (mid_1[2567:2560] < mid_1[2575:2568]) ? 1 : 0;
assign detect_min[319][14] = (mid_1[2567:2560] < mid_2[2559:2552]) ? 1 : 0;
assign detect_min[319][15] = (mid_1[2567:2560] < mid_2[2567:2560]) ? 1 : 0;
assign detect_min[319][16] = (mid_1[2567:2560] < mid_2[2575:2568]) ? 1 : 0;
assign detect_min[319][17] = (mid_1[2567:2560] < btm_0[2559:2552]) ? 1 : 0;
assign detect_min[319][18] = (mid_1[2567:2560] < btm_0[2567:2560]) ? 1 : 0;
assign detect_min[319][19] = (mid_1[2567:2560] < btm_0[2575:2568]) ? 1 : 0;
assign detect_min[319][20] = (mid_1[2567:2560] < btm_1[2559:2552]) ? 1 : 0;
assign detect_min[319][21] = (mid_1[2567:2560] < btm_1[2567:2560]) ? 1 : 0;
assign detect_min[319][22] = (mid_1[2567:2560] < btm_1[2575:2568]) ? 1 : 0;
assign detect_min[319][23] = (mid_1[2567:2560] < btm_2[2559:2552]) ? 1 : 0;
assign detect_min[319][24] = (mid_1[2567:2560] < btm_2[2567:2560]) ? 1 : 0;
assign detect_min[319][25] = (mid_1[2567:2560] < btm_2[2575:2568]) ? 1 : 0;

assign detect_min[320][0] = (mid_1[2575:2568] < top_0[2567:2560]) ? 1 : 0;
assign detect_min[320][1] = (mid_1[2575:2568] < top_0[2575:2568]) ? 1 : 0;
assign detect_min[320][2] = (mid_1[2575:2568] < top_0[2583:2576]) ? 1 : 0;
assign detect_min[320][3] = (mid_1[2575:2568] < top_1[2567:2560]) ? 1 : 0;
assign detect_min[320][4] = (mid_1[2575:2568] < top_1[2575:2568]) ? 1 : 0;
assign detect_min[320][5] = (mid_1[2575:2568] < top_1[2583:2576]) ? 1 : 0;
assign detect_min[320][6] = (mid_1[2575:2568] < top_2[2567:2560]) ? 1 : 0;
assign detect_min[320][7] = (mid_1[2575:2568] < top_2[2575:2568]) ? 1 : 0;
assign detect_min[320][8] = (mid_1[2575:2568] < top_2[2583:2576]) ? 1 : 0;
assign detect_min[320][9] = (mid_1[2575:2568] < mid_0[2567:2560]) ? 1 : 0;
assign detect_min[320][10] = (mid_1[2575:2568] < mid_0[2575:2568]) ? 1 : 0;
assign detect_min[320][11] = (mid_1[2575:2568] < mid_0[2583:2576]) ? 1 : 0;
assign detect_min[320][12] = (mid_1[2575:2568] < mid_1[2567:2560]) ? 1 : 0;
assign detect_min[320][13] = (mid_1[2575:2568] < mid_1[2583:2576]) ? 1 : 0;
assign detect_min[320][14] = (mid_1[2575:2568] < mid_2[2567:2560]) ? 1 : 0;
assign detect_min[320][15] = (mid_1[2575:2568] < mid_2[2575:2568]) ? 1 : 0;
assign detect_min[320][16] = (mid_1[2575:2568] < mid_2[2583:2576]) ? 1 : 0;
assign detect_min[320][17] = (mid_1[2575:2568] < btm_0[2567:2560]) ? 1 : 0;
assign detect_min[320][18] = (mid_1[2575:2568] < btm_0[2575:2568]) ? 1 : 0;
assign detect_min[320][19] = (mid_1[2575:2568] < btm_0[2583:2576]) ? 1 : 0;
assign detect_min[320][20] = (mid_1[2575:2568] < btm_1[2567:2560]) ? 1 : 0;
assign detect_min[320][21] = (mid_1[2575:2568] < btm_1[2575:2568]) ? 1 : 0;
assign detect_min[320][22] = (mid_1[2575:2568] < btm_1[2583:2576]) ? 1 : 0;
assign detect_min[320][23] = (mid_1[2575:2568] < btm_2[2567:2560]) ? 1 : 0;
assign detect_min[320][24] = (mid_1[2575:2568] < btm_2[2575:2568]) ? 1 : 0;
assign detect_min[320][25] = (mid_1[2575:2568] < btm_2[2583:2576]) ? 1 : 0;

assign detect_min[321][0] = (mid_1[2583:2576] < top_0[2575:2568]) ? 1 : 0;
assign detect_min[321][1] = (mid_1[2583:2576] < top_0[2583:2576]) ? 1 : 0;
assign detect_min[321][2] = (mid_1[2583:2576] < top_0[2591:2584]) ? 1 : 0;
assign detect_min[321][3] = (mid_1[2583:2576] < top_1[2575:2568]) ? 1 : 0;
assign detect_min[321][4] = (mid_1[2583:2576] < top_1[2583:2576]) ? 1 : 0;
assign detect_min[321][5] = (mid_1[2583:2576] < top_1[2591:2584]) ? 1 : 0;
assign detect_min[321][6] = (mid_1[2583:2576] < top_2[2575:2568]) ? 1 : 0;
assign detect_min[321][7] = (mid_1[2583:2576] < top_2[2583:2576]) ? 1 : 0;
assign detect_min[321][8] = (mid_1[2583:2576] < top_2[2591:2584]) ? 1 : 0;
assign detect_min[321][9] = (mid_1[2583:2576] < mid_0[2575:2568]) ? 1 : 0;
assign detect_min[321][10] = (mid_1[2583:2576] < mid_0[2583:2576]) ? 1 : 0;
assign detect_min[321][11] = (mid_1[2583:2576] < mid_0[2591:2584]) ? 1 : 0;
assign detect_min[321][12] = (mid_1[2583:2576] < mid_1[2575:2568]) ? 1 : 0;
assign detect_min[321][13] = (mid_1[2583:2576] < mid_1[2591:2584]) ? 1 : 0;
assign detect_min[321][14] = (mid_1[2583:2576] < mid_2[2575:2568]) ? 1 : 0;
assign detect_min[321][15] = (mid_1[2583:2576] < mid_2[2583:2576]) ? 1 : 0;
assign detect_min[321][16] = (mid_1[2583:2576] < mid_2[2591:2584]) ? 1 : 0;
assign detect_min[321][17] = (mid_1[2583:2576] < btm_0[2575:2568]) ? 1 : 0;
assign detect_min[321][18] = (mid_1[2583:2576] < btm_0[2583:2576]) ? 1 : 0;
assign detect_min[321][19] = (mid_1[2583:2576] < btm_0[2591:2584]) ? 1 : 0;
assign detect_min[321][20] = (mid_1[2583:2576] < btm_1[2575:2568]) ? 1 : 0;
assign detect_min[321][21] = (mid_1[2583:2576] < btm_1[2583:2576]) ? 1 : 0;
assign detect_min[321][22] = (mid_1[2583:2576] < btm_1[2591:2584]) ? 1 : 0;
assign detect_min[321][23] = (mid_1[2583:2576] < btm_2[2575:2568]) ? 1 : 0;
assign detect_min[321][24] = (mid_1[2583:2576] < btm_2[2583:2576]) ? 1 : 0;
assign detect_min[321][25] = (mid_1[2583:2576] < btm_2[2591:2584]) ? 1 : 0;

assign detect_min[322][0] = (mid_1[2591:2584] < top_0[2583:2576]) ? 1 : 0;
assign detect_min[322][1] = (mid_1[2591:2584] < top_0[2591:2584]) ? 1 : 0;
assign detect_min[322][2] = (mid_1[2591:2584] < top_0[2599:2592]) ? 1 : 0;
assign detect_min[322][3] = (mid_1[2591:2584] < top_1[2583:2576]) ? 1 : 0;
assign detect_min[322][4] = (mid_1[2591:2584] < top_1[2591:2584]) ? 1 : 0;
assign detect_min[322][5] = (mid_1[2591:2584] < top_1[2599:2592]) ? 1 : 0;
assign detect_min[322][6] = (mid_1[2591:2584] < top_2[2583:2576]) ? 1 : 0;
assign detect_min[322][7] = (mid_1[2591:2584] < top_2[2591:2584]) ? 1 : 0;
assign detect_min[322][8] = (mid_1[2591:2584] < top_2[2599:2592]) ? 1 : 0;
assign detect_min[322][9] = (mid_1[2591:2584] < mid_0[2583:2576]) ? 1 : 0;
assign detect_min[322][10] = (mid_1[2591:2584] < mid_0[2591:2584]) ? 1 : 0;
assign detect_min[322][11] = (mid_1[2591:2584] < mid_0[2599:2592]) ? 1 : 0;
assign detect_min[322][12] = (mid_1[2591:2584] < mid_1[2583:2576]) ? 1 : 0;
assign detect_min[322][13] = (mid_1[2591:2584] < mid_1[2599:2592]) ? 1 : 0;
assign detect_min[322][14] = (mid_1[2591:2584] < mid_2[2583:2576]) ? 1 : 0;
assign detect_min[322][15] = (mid_1[2591:2584] < mid_2[2591:2584]) ? 1 : 0;
assign detect_min[322][16] = (mid_1[2591:2584] < mid_2[2599:2592]) ? 1 : 0;
assign detect_min[322][17] = (mid_1[2591:2584] < btm_0[2583:2576]) ? 1 : 0;
assign detect_min[322][18] = (mid_1[2591:2584] < btm_0[2591:2584]) ? 1 : 0;
assign detect_min[322][19] = (mid_1[2591:2584] < btm_0[2599:2592]) ? 1 : 0;
assign detect_min[322][20] = (mid_1[2591:2584] < btm_1[2583:2576]) ? 1 : 0;
assign detect_min[322][21] = (mid_1[2591:2584] < btm_1[2591:2584]) ? 1 : 0;
assign detect_min[322][22] = (mid_1[2591:2584] < btm_1[2599:2592]) ? 1 : 0;
assign detect_min[322][23] = (mid_1[2591:2584] < btm_2[2583:2576]) ? 1 : 0;
assign detect_min[322][24] = (mid_1[2591:2584] < btm_2[2591:2584]) ? 1 : 0;
assign detect_min[322][25] = (mid_1[2591:2584] < btm_2[2599:2592]) ? 1 : 0;

assign detect_min[323][0] = (mid_1[2599:2592] < top_0[2591:2584]) ? 1 : 0;
assign detect_min[323][1] = (mid_1[2599:2592] < top_0[2599:2592]) ? 1 : 0;
assign detect_min[323][2] = (mid_1[2599:2592] < top_0[2607:2600]) ? 1 : 0;
assign detect_min[323][3] = (mid_1[2599:2592] < top_1[2591:2584]) ? 1 : 0;
assign detect_min[323][4] = (mid_1[2599:2592] < top_1[2599:2592]) ? 1 : 0;
assign detect_min[323][5] = (mid_1[2599:2592] < top_1[2607:2600]) ? 1 : 0;
assign detect_min[323][6] = (mid_1[2599:2592] < top_2[2591:2584]) ? 1 : 0;
assign detect_min[323][7] = (mid_1[2599:2592] < top_2[2599:2592]) ? 1 : 0;
assign detect_min[323][8] = (mid_1[2599:2592] < top_2[2607:2600]) ? 1 : 0;
assign detect_min[323][9] = (mid_1[2599:2592] < mid_0[2591:2584]) ? 1 : 0;
assign detect_min[323][10] = (mid_1[2599:2592] < mid_0[2599:2592]) ? 1 : 0;
assign detect_min[323][11] = (mid_1[2599:2592] < mid_0[2607:2600]) ? 1 : 0;
assign detect_min[323][12] = (mid_1[2599:2592] < mid_1[2591:2584]) ? 1 : 0;
assign detect_min[323][13] = (mid_1[2599:2592] < mid_1[2607:2600]) ? 1 : 0;
assign detect_min[323][14] = (mid_1[2599:2592] < mid_2[2591:2584]) ? 1 : 0;
assign detect_min[323][15] = (mid_1[2599:2592] < mid_2[2599:2592]) ? 1 : 0;
assign detect_min[323][16] = (mid_1[2599:2592] < mid_2[2607:2600]) ? 1 : 0;
assign detect_min[323][17] = (mid_1[2599:2592] < btm_0[2591:2584]) ? 1 : 0;
assign detect_min[323][18] = (mid_1[2599:2592] < btm_0[2599:2592]) ? 1 : 0;
assign detect_min[323][19] = (mid_1[2599:2592] < btm_0[2607:2600]) ? 1 : 0;
assign detect_min[323][20] = (mid_1[2599:2592] < btm_1[2591:2584]) ? 1 : 0;
assign detect_min[323][21] = (mid_1[2599:2592] < btm_1[2599:2592]) ? 1 : 0;
assign detect_min[323][22] = (mid_1[2599:2592] < btm_1[2607:2600]) ? 1 : 0;
assign detect_min[323][23] = (mid_1[2599:2592] < btm_2[2591:2584]) ? 1 : 0;
assign detect_min[323][24] = (mid_1[2599:2592] < btm_2[2599:2592]) ? 1 : 0;
assign detect_min[323][25] = (mid_1[2599:2592] < btm_2[2607:2600]) ? 1 : 0;

assign detect_min[324][0] = (mid_1[2607:2600] < top_0[2599:2592]) ? 1 : 0;
assign detect_min[324][1] = (mid_1[2607:2600] < top_0[2607:2600]) ? 1 : 0;
assign detect_min[324][2] = (mid_1[2607:2600] < top_0[2615:2608]) ? 1 : 0;
assign detect_min[324][3] = (mid_1[2607:2600] < top_1[2599:2592]) ? 1 : 0;
assign detect_min[324][4] = (mid_1[2607:2600] < top_1[2607:2600]) ? 1 : 0;
assign detect_min[324][5] = (mid_1[2607:2600] < top_1[2615:2608]) ? 1 : 0;
assign detect_min[324][6] = (mid_1[2607:2600] < top_2[2599:2592]) ? 1 : 0;
assign detect_min[324][7] = (mid_1[2607:2600] < top_2[2607:2600]) ? 1 : 0;
assign detect_min[324][8] = (mid_1[2607:2600] < top_2[2615:2608]) ? 1 : 0;
assign detect_min[324][9] = (mid_1[2607:2600] < mid_0[2599:2592]) ? 1 : 0;
assign detect_min[324][10] = (mid_1[2607:2600] < mid_0[2607:2600]) ? 1 : 0;
assign detect_min[324][11] = (mid_1[2607:2600] < mid_0[2615:2608]) ? 1 : 0;
assign detect_min[324][12] = (mid_1[2607:2600] < mid_1[2599:2592]) ? 1 : 0;
assign detect_min[324][13] = (mid_1[2607:2600] < mid_1[2615:2608]) ? 1 : 0;
assign detect_min[324][14] = (mid_1[2607:2600] < mid_2[2599:2592]) ? 1 : 0;
assign detect_min[324][15] = (mid_1[2607:2600] < mid_2[2607:2600]) ? 1 : 0;
assign detect_min[324][16] = (mid_1[2607:2600] < mid_2[2615:2608]) ? 1 : 0;
assign detect_min[324][17] = (mid_1[2607:2600] < btm_0[2599:2592]) ? 1 : 0;
assign detect_min[324][18] = (mid_1[2607:2600] < btm_0[2607:2600]) ? 1 : 0;
assign detect_min[324][19] = (mid_1[2607:2600] < btm_0[2615:2608]) ? 1 : 0;
assign detect_min[324][20] = (mid_1[2607:2600] < btm_1[2599:2592]) ? 1 : 0;
assign detect_min[324][21] = (mid_1[2607:2600] < btm_1[2607:2600]) ? 1 : 0;
assign detect_min[324][22] = (mid_1[2607:2600] < btm_1[2615:2608]) ? 1 : 0;
assign detect_min[324][23] = (mid_1[2607:2600] < btm_2[2599:2592]) ? 1 : 0;
assign detect_min[324][24] = (mid_1[2607:2600] < btm_2[2607:2600]) ? 1 : 0;
assign detect_min[324][25] = (mid_1[2607:2600] < btm_2[2615:2608]) ? 1 : 0;

assign detect_min[325][0] = (mid_1[2615:2608] < top_0[2607:2600]) ? 1 : 0;
assign detect_min[325][1] = (mid_1[2615:2608] < top_0[2615:2608]) ? 1 : 0;
assign detect_min[325][2] = (mid_1[2615:2608] < top_0[2623:2616]) ? 1 : 0;
assign detect_min[325][3] = (mid_1[2615:2608] < top_1[2607:2600]) ? 1 : 0;
assign detect_min[325][4] = (mid_1[2615:2608] < top_1[2615:2608]) ? 1 : 0;
assign detect_min[325][5] = (mid_1[2615:2608] < top_1[2623:2616]) ? 1 : 0;
assign detect_min[325][6] = (mid_1[2615:2608] < top_2[2607:2600]) ? 1 : 0;
assign detect_min[325][7] = (mid_1[2615:2608] < top_2[2615:2608]) ? 1 : 0;
assign detect_min[325][8] = (mid_1[2615:2608] < top_2[2623:2616]) ? 1 : 0;
assign detect_min[325][9] = (mid_1[2615:2608] < mid_0[2607:2600]) ? 1 : 0;
assign detect_min[325][10] = (mid_1[2615:2608] < mid_0[2615:2608]) ? 1 : 0;
assign detect_min[325][11] = (mid_1[2615:2608] < mid_0[2623:2616]) ? 1 : 0;
assign detect_min[325][12] = (mid_1[2615:2608] < mid_1[2607:2600]) ? 1 : 0;
assign detect_min[325][13] = (mid_1[2615:2608] < mid_1[2623:2616]) ? 1 : 0;
assign detect_min[325][14] = (mid_1[2615:2608] < mid_2[2607:2600]) ? 1 : 0;
assign detect_min[325][15] = (mid_1[2615:2608] < mid_2[2615:2608]) ? 1 : 0;
assign detect_min[325][16] = (mid_1[2615:2608] < mid_2[2623:2616]) ? 1 : 0;
assign detect_min[325][17] = (mid_1[2615:2608] < btm_0[2607:2600]) ? 1 : 0;
assign detect_min[325][18] = (mid_1[2615:2608] < btm_0[2615:2608]) ? 1 : 0;
assign detect_min[325][19] = (mid_1[2615:2608] < btm_0[2623:2616]) ? 1 : 0;
assign detect_min[325][20] = (mid_1[2615:2608] < btm_1[2607:2600]) ? 1 : 0;
assign detect_min[325][21] = (mid_1[2615:2608] < btm_1[2615:2608]) ? 1 : 0;
assign detect_min[325][22] = (mid_1[2615:2608] < btm_1[2623:2616]) ? 1 : 0;
assign detect_min[325][23] = (mid_1[2615:2608] < btm_2[2607:2600]) ? 1 : 0;
assign detect_min[325][24] = (mid_1[2615:2608] < btm_2[2615:2608]) ? 1 : 0;
assign detect_min[325][25] = (mid_1[2615:2608] < btm_2[2623:2616]) ? 1 : 0;

assign detect_min[326][0] = (mid_1[2623:2616] < top_0[2615:2608]) ? 1 : 0;
assign detect_min[326][1] = (mid_1[2623:2616] < top_0[2623:2616]) ? 1 : 0;
assign detect_min[326][2] = (mid_1[2623:2616] < top_0[2631:2624]) ? 1 : 0;
assign detect_min[326][3] = (mid_1[2623:2616] < top_1[2615:2608]) ? 1 : 0;
assign detect_min[326][4] = (mid_1[2623:2616] < top_1[2623:2616]) ? 1 : 0;
assign detect_min[326][5] = (mid_1[2623:2616] < top_1[2631:2624]) ? 1 : 0;
assign detect_min[326][6] = (mid_1[2623:2616] < top_2[2615:2608]) ? 1 : 0;
assign detect_min[326][7] = (mid_1[2623:2616] < top_2[2623:2616]) ? 1 : 0;
assign detect_min[326][8] = (mid_1[2623:2616] < top_2[2631:2624]) ? 1 : 0;
assign detect_min[326][9] = (mid_1[2623:2616] < mid_0[2615:2608]) ? 1 : 0;
assign detect_min[326][10] = (mid_1[2623:2616] < mid_0[2623:2616]) ? 1 : 0;
assign detect_min[326][11] = (mid_1[2623:2616] < mid_0[2631:2624]) ? 1 : 0;
assign detect_min[326][12] = (mid_1[2623:2616] < mid_1[2615:2608]) ? 1 : 0;
assign detect_min[326][13] = (mid_1[2623:2616] < mid_1[2631:2624]) ? 1 : 0;
assign detect_min[326][14] = (mid_1[2623:2616] < mid_2[2615:2608]) ? 1 : 0;
assign detect_min[326][15] = (mid_1[2623:2616] < mid_2[2623:2616]) ? 1 : 0;
assign detect_min[326][16] = (mid_1[2623:2616] < mid_2[2631:2624]) ? 1 : 0;
assign detect_min[326][17] = (mid_1[2623:2616] < btm_0[2615:2608]) ? 1 : 0;
assign detect_min[326][18] = (mid_1[2623:2616] < btm_0[2623:2616]) ? 1 : 0;
assign detect_min[326][19] = (mid_1[2623:2616] < btm_0[2631:2624]) ? 1 : 0;
assign detect_min[326][20] = (mid_1[2623:2616] < btm_1[2615:2608]) ? 1 : 0;
assign detect_min[326][21] = (mid_1[2623:2616] < btm_1[2623:2616]) ? 1 : 0;
assign detect_min[326][22] = (mid_1[2623:2616] < btm_1[2631:2624]) ? 1 : 0;
assign detect_min[326][23] = (mid_1[2623:2616] < btm_2[2615:2608]) ? 1 : 0;
assign detect_min[326][24] = (mid_1[2623:2616] < btm_2[2623:2616]) ? 1 : 0;
assign detect_min[326][25] = (mid_1[2623:2616] < btm_2[2631:2624]) ? 1 : 0;

assign detect_min[327][0] = (mid_1[2631:2624] < top_0[2623:2616]) ? 1 : 0;
assign detect_min[327][1] = (mid_1[2631:2624] < top_0[2631:2624]) ? 1 : 0;
assign detect_min[327][2] = (mid_1[2631:2624] < top_0[2639:2632]) ? 1 : 0;
assign detect_min[327][3] = (mid_1[2631:2624] < top_1[2623:2616]) ? 1 : 0;
assign detect_min[327][4] = (mid_1[2631:2624] < top_1[2631:2624]) ? 1 : 0;
assign detect_min[327][5] = (mid_1[2631:2624] < top_1[2639:2632]) ? 1 : 0;
assign detect_min[327][6] = (mid_1[2631:2624] < top_2[2623:2616]) ? 1 : 0;
assign detect_min[327][7] = (mid_1[2631:2624] < top_2[2631:2624]) ? 1 : 0;
assign detect_min[327][8] = (mid_1[2631:2624] < top_2[2639:2632]) ? 1 : 0;
assign detect_min[327][9] = (mid_1[2631:2624] < mid_0[2623:2616]) ? 1 : 0;
assign detect_min[327][10] = (mid_1[2631:2624] < mid_0[2631:2624]) ? 1 : 0;
assign detect_min[327][11] = (mid_1[2631:2624] < mid_0[2639:2632]) ? 1 : 0;
assign detect_min[327][12] = (mid_1[2631:2624] < mid_1[2623:2616]) ? 1 : 0;
assign detect_min[327][13] = (mid_1[2631:2624] < mid_1[2639:2632]) ? 1 : 0;
assign detect_min[327][14] = (mid_1[2631:2624] < mid_2[2623:2616]) ? 1 : 0;
assign detect_min[327][15] = (mid_1[2631:2624] < mid_2[2631:2624]) ? 1 : 0;
assign detect_min[327][16] = (mid_1[2631:2624] < mid_2[2639:2632]) ? 1 : 0;
assign detect_min[327][17] = (mid_1[2631:2624] < btm_0[2623:2616]) ? 1 : 0;
assign detect_min[327][18] = (mid_1[2631:2624] < btm_0[2631:2624]) ? 1 : 0;
assign detect_min[327][19] = (mid_1[2631:2624] < btm_0[2639:2632]) ? 1 : 0;
assign detect_min[327][20] = (mid_1[2631:2624] < btm_1[2623:2616]) ? 1 : 0;
assign detect_min[327][21] = (mid_1[2631:2624] < btm_1[2631:2624]) ? 1 : 0;
assign detect_min[327][22] = (mid_1[2631:2624] < btm_1[2639:2632]) ? 1 : 0;
assign detect_min[327][23] = (mid_1[2631:2624] < btm_2[2623:2616]) ? 1 : 0;
assign detect_min[327][24] = (mid_1[2631:2624] < btm_2[2631:2624]) ? 1 : 0;
assign detect_min[327][25] = (mid_1[2631:2624] < btm_2[2639:2632]) ? 1 : 0;

assign detect_min[328][0] = (mid_1[2639:2632] < top_0[2631:2624]) ? 1 : 0;
assign detect_min[328][1] = (mid_1[2639:2632] < top_0[2639:2632]) ? 1 : 0;
assign detect_min[328][2] = (mid_1[2639:2632] < top_0[2647:2640]) ? 1 : 0;
assign detect_min[328][3] = (mid_1[2639:2632] < top_1[2631:2624]) ? 1 : 0;
assign detect_min[328][4] = (mid_1[2639:2632] < top_1[2639:2632]) ? 1 : 0;
assign detect_min[328][5] = (mid_1[2639:2632] < top_1[2647:2640]) ? 1 : 0;
assign detect_min[328][6] = (mid_1[2639:2632] < top_2[2631:2624]) ? 1 : 0;
assign detect_min[328][7] = (mid_1[2639:2632] < top_2[2639:2632]) ? 1 : 0;
assign detect_min[328][8] = (mid_1[2639:2632] < top_2[2647:2640]) ? 1 : 0;
assign detect_min[328][9] = (mid_1[2639:2632] < mid_0[2631:2624]) ? 1 : 0;
assign detect_min[328][10] = (mid_1[2639:2632] < mid_0[2639:2632]) ? 1 : 0;
assign detect_min[328][11] = (mid_1[2639:2632] < mid_0[2647:2640]) ? 1 : 0;
assign detect_min[328][12] = (mid_1[2639:2632] < mid_1[2631:2624]) ? 1 : 0;
assign detect_min[328][13] = (mid_1[2639:2632] < mid_1[2647:2640]) ? 1 : 0;
assign detect_min[328][14] = (mid_1[2639:2632] < mid_2[2631:2624]) ? 1 : 0;
assign detect_min[328][15] = (mid_1[2639:2632] < mid_2[2639:2632]) ? 1 : 0;
assign detect_min[328][16] = (mid_1[2639:2632] < mid_2[2647:2640]) ? 1 : 0;
assign detect_min[328][17] = (mid_1[2639:2632] < btm_0[2631:2624]) ? 1 : 0;
assign detect_min[328][18] = (mid_1[2639:2632] < btm_0[2639:2632]) ? 1 : 0;
assign detect_min[328][19] = (mid_1[2639:2632] < btm_0[2647:2640]) ? 1 : 0;
assign detect_min[328][20] = (mid_1[2639:2632] < btm_1[2631:2624]) ? 1 : 0;
assign detect_min[328][21] = (mid_1[2639:2632] < btm_1[2639:2632]) ? 1 : 0;
assign detect_min[328][22] = (mid_1[2639:2632] < btm_1[2647:2640]) ? 1 : 0;
assign detect_min[328][23] = (mid_1[2639:2632] < btm_2[2631:2624]) ? 1 : 0;
assign detect_min[328][24] = (mid_1[2639:2632] < btm_2[2639:2632]) ? 1 : 0;
assign detect_min[328][25] = (mid_1[2639:2632] < btm_2[2647:2640]) ? 1 : 0;

assign detect_min[329][0] = (mid_1[2647:2640] < top_0[2639:2632]) ? 1 : 0;
assign detect_min[329][1] = (mid_1[2647:2640] < top_0[2647:2640]) ? 1 : 0;
assign detect_min[329][2] = (mid_1[2647:2640] < top_0[2655:2648]) ? 1 : 0;
assign detect_min[329][3] = (mid_1[2647:2640] < top_1[2639:2632]) ? 1 : 0;
assign detect_min[329][4] = (mid_1[2647:2640] < top_1[2647:2640]) ? 1 : 0;
assign detect_min[329][5] = (mid_1[2647:2640] < top_1[2655:2648]) ? 1 : 0;
assign detect_min[329][6] = (mid_1[2647:2640] < top_2[2639:2632]) ? 1 : 0;
assign detect_min[329][7] = (mid_1[2647:2640] < top_2[2647:2640]) ? 1 : 0;
assign detect_min[329][8] = (mid_1[2647:2640] < top_2[2655:2648]) ? 1 : 0;
assign detect_min[329][9] = (mid_1[2647:2640] < mid_0[2639:2632]) ? 1 : 0;
assign detect_min[329][10] = (mid_1[2647:2640] < mid_0[2647:2640]) ? 1 : 0;
assign detect_min[329][11] = (mid_1[2647:2640] < mid_0[2655:2648]) ? 1 : 0;
assign detect_min[329][12] = (mid_1[2647:2640] < mid_1[2639:2632]) ? 1 : 0;
assign detect_min[329][13] = (mid_1[2647:2640] < mid_1[2655:2648]) ? 1 : 0;
assign detect_min[329][14] = (mid_1[2647:2640] < mid_2[2639:2632]) ? 1 : 0;
assign detect_min[329][15] = (mid_1[2647:2640] < mid_2[2647:2640]) ? 1 : 0;
assign detect_min[329][16] = (mid_1[2647:2640] < mid_2[2655:2648]) ? 1 : 0;
assign detect_min[329][17] = (mid_1[2647:2640] < btm_0[2639:2632]) ? 1 : 0;
assign detect_min[329][18] = (mid_1[2647:2640] < btm_0[2647:2640]) ? 1 : 0;
assign detect_min[329][19] = (mid_1[2647:2640] < btm_0[2655:2648]) ? 1 : 0;
assign detect_min[329][20] = (mid_1[2647:2640] < btm_1[2639:2632]) ? 1 : 0;
assign detect_min[329][21] = (mid_1[2647:2640] < btm_1[2647:2640]) ? 1 : 0;
assign detect_min[329][22] = (mid_1[2647:2640] < btm_1[2655:2648]) ? 1 : 0;
assign detect_min[329][23] = (mid_1[2647:2640] < btm_2[2639:2632]) ? 1 : 0;
assign detect_min[329][24] = (mid_1[2647:2640] < btm_2[2647:2640]) ? 1 : 0;
assign detect_min[329][25] = (mid_1[2647:2640] < btm_2[2655:2648]) ? 1 : 0;

assign detect_min[330][0] = (mid_1[2655:2648] < top_0[2647:2640]) ? 1 : 0;
assign detect_min[330][1] = (mid_1[2655:2648] < top_0[2655:2648]) ? 1 : 0;
assign detect_min[330][2] = (mid_1[2655:2648] < top_0[2663:2656]) ? 1 : 0;
assign detect_min[330][3] = (mid_1[2655:2648] < top_1[2647:2640]) ? 1 : 0;
assign detect_min[330][4] = (mid_1[2655:2648] < top_1[2655:2648]) ? 1 : 0;
assign detect_min[330][5] = (mid_1[2655:2648] < top_1[2663:2656]) ? 1 : 0;
assign detect_min[330][6] = (mid_1[2655:2648] < top_2[2647:2640]) ? 1 : 0;
assign detect_min[330][7] = (mid_1[2655:2648] < top_2[2655:2648]) ? 1 : 0;
assign detect_min[330][8] = (mid_1[2655:2648] < top_2[2663:2656]) ? 1 : 0;
assign detect_min[330][9] = (mid_1[2655:2648] < mid_0[2647:2640]) ? 1 : 0;
assign detect_min[330][10] = (mid_1[2655:2648] < mid_0[2655:2648]) ? 1 : 0;
assign detect_min[330][11] = (mid_1[2655:2648] < mid_0[2663:2656]) ? 1 : 0;
assign detect_min[330][12] = (mid_1[2655:2648] < mid_1[2647:2640]) ? 1 : 0;
assign detect_min[330][13] = (mid_1[2655:2648] < mid_1[2663:2656]) ? 1 : 0;
assign detect_min[330][14] = (mid_1[2655:2648] < mid_2[2647:2640]) ? 1 : 0;
assign detect_min[330][15] = (mid_1[2655:2648] < mid_2[2655:2648]) ? 1 : 0;
assign detect_min[330][16] = (mid_1[2655:2648] < mid_2[2663:2656]) ? 1 : 0;
assign detect_min[330][17] = (mid_1[2655:2648] < btm_0[2647:2640]) ? 1 : 0;
assign detect_min[330][18] = (mid_1[2655:2648] < btm_0[2655:2648]) ? 1 : 0;
assign detect_min[330][19] = (mid_1[2655:2648] < btm_0[2663:2656]) ? 1 : 0;
assign detect_min[330][20] = (mid_1[2655:2648] < btm_1[2647:2640]) ? 1 : 0;
assign detect_min[330][21] = (mid_1[2655:2648] < btm_1[2655:2648]) ? 1 : 0;
assign detect_min[330][22] = (mid_1[2655:2648] < btm_1[2663:2656]) ? 1 : 0;
assign detect_min[330][23] = (mid_1[2655:2648] < btm_2[2647:2640]) ? 1 : 0;
assign detect_min[330][24] = (mid_1[2655:2648] < btm_2[2655:2648]) ? 1 : 0;
assign detect_min[330][25] = (mid_1[2655:2648] < btm_2[2663:2656]) ? 1 : 0;

assign detect_min[331][0] = (mid_1[2663:2656] < top_0[2655:2648]) ? 1 : 0;
assign detect_min[331][1] = (mid_1[2663:2656] < top_0[2663:2656]) ? 1 : 0;
assign detect_min[331][2] = (mid_1[2663:2656] < top_0[2671:2664]) ? 1 : 0;
assign detect_min[331][3] = (mid_1[2663:2656] < top_1[2655:2648]) ? 1 : 0;
assign detect_min[331][4] = (mid_1[2663:2656] < top_1[2663:2656]) ? 1 : 0;
assign detect_min[331][5] = (mid_1[2663:2656] < top_1[2671:2664]) ? 1 : 0;
assign detect_min[331][6] = (mid_1[2663:2656] < top_2[2655:2648]) ? 1 : 0;
assign detect_min[331][7] = (mid_1[2663:2656] < top_2[2663:2656]) ? 1 : 0;
assign detect_min[331][8] = (mid_1[2663:2656] < top_2[2671:2664]) ? 1 : 0;
assign detect_min[331][9] = (mid_1[2663:2656] < mid_0[2655:2648]) ? 1 : 0;
assign detect_min[331][10] = (mid_1[2663:2656] < mid_0[2663:2656]) ? 1 : 0;
assign detect_min[331][11] = (mid_1[2663:2656] < mid_0[2671:2664]) ? 1 : 0;
assign detect_min[331][12] = (mid_1[2663:2656] < mid_1[2655:2648]) ? 1 : 0;
assign detect_min[331][13] = (mid_1[2663:2656] < mid_1[2671:2664]) ? 1 : 0;
assign detect_min[331][14] = (mid_1[2663:2656] < mid_2[2655:2648]) ? 1 : 0;
assign detect_min[331][15] = (mid_1[2663:2656] < mid_2[2663:2656]) ? 1 : 0;
assign detect_min[331][16] = (mid_1[2663:2656] < mid_2[2671:2664]) ? 1 : 0;
assign detect_min[331][17] = (mid_1[2663:2656] < btm_0[2655:2648]) ? 1 : 0;
assign detect_min[331][18] = (mid_1[2663:2656] < btm_0[2663:2656]) ? 1 : 0;
assign detect_min[331][19] = (mid_1[2663:2656] < btm_0[2671:2664]) ? 1 : 0;
assign detect_min[331][20] = (mid_1[2663:2656] < btm_1[2655:2648]) ? 1 : 0;
assign detect_min[331][21] = (mid_1[2663:2656] < btm_1[2663:2656]) ? 1 : 0;
assign detect_min[331][22] = (mid_1[2663:2656] < btm_1[2671:2664]) ? 1 : 0;
assign detect_min[331][23] = (mid_1[2663:2656] < btm_2[2655:2648]) ? 1 : 0;
assign detect_min[331][24] = (mid_1[2663:2656] < btm_2[2663:2656]) ? 1 : 0;
assign detect_min[331][25] = (mid_1[2663:2656] < btm_2[2671:2664]) ? 1 : 0;

assign detect_min[332][0] = (mid_1[2671:2664] < top_0[2663:2656]) ? 1 : 0;
assign detect_min[332][1] = (mid_1[2671:2664] < top_0[2671:2664]) ? 1 : 0;
assign detect_min[332][2] = (mid_1[2671:2664] < top_0[2679:2672]) ? 1 : 0;
assign detect_min[332][3] = (mid_1[2671:2664] < top_1[2663:2656]) ? 1 : 0;
assign detect_min[332][4] = (mid_1[2671:2664] < top_1[2671:2664]) ? 1 : 0;
assign detect_min[332][5] = (mid_1[2671:2664] < top_1[2679:2672]) ? 1 : 0;
assign detect_min[332][6] = (mid_1[2671:2664] < top_2[2663:2656]) ? 1 : 0;
assign detect_min[332][7] = (mid_1[2671:2664] < top_2[2671:2664]) ? 1 : 0;
assign detect_min[332][8] = (mid_1[2671:2664] < top_2[2679:2672]) ? 1 : 0;
assign detect_min[332][9] = (mid_1[2671:2664] < mid_0[2663:2656]) ? 1 : 0;
assign detect_min[332][10] = (mid_1[2671:2664] < mid_0[2671:2664]) ? 1 : 0;
assign detect_min[332][11] = (mid_1[2671:2664] < mid_0[2679:2672]) ? 1 : 0;
assign detect_min[332][12] = (mid_1[2671:2664] < mid_1[2663:2656]) ? 1 : 0;
assign detect_min[332][13] = (mid_1[2671:2664] < mid_1[2679:2672]) ? 1 : 0;
assign detect_min[332][14] = (mid_1[2671:2664] < mid_2[2663:2656]) ? 1 : 0;
assign detect_min[332][15] = (mid_1[2671:2664] < mid_2[2671:2664]) ? 1 : 0;
assign detect_min[332][16] = (mid_1[2671:2664] < mid_2[2679:2672]) ? 1 : 0;
assign detect_min[332][17] = (mid_1[2671:2664] < btm_0[2663:2656]) ? 1 : 0;
assign detect_min[332][18] = (mid_1[2671:2664] < btm_0[2671:2664]) ? 1 : 0;
assign detect_min[332][19] = (mid_1[2671:2664] < btm_0[2679:2672]) ? 1 : 0;
assign detect_min[332][20] = (mid_1[2671:2664] < btm_1[2663:2656]) ? 1 : 0;
assign detect_min[332][21] = (mid_1[2671:2664] < btm_1[2671:2664]) ? 1 : 0;
assign detect_min[332][22] = (mid_1[2671:2664] < btm_1[2679:2672]) ? 1 : 0;
assign detect_min[332][23] = (mid_1[2671:2664] < btm_2[2663:2656]) ? 1 : 0;
assign detect_min[332][24] = (mid_1[2671:2664] < btm_2[2671:2664]) ? 1 : 0;
assign detect_min[332][25] = (mid_1[2671:2664] < btm_2[2679:2672]) ? 1 : 0;

assign detect_min[333][0] = (mid_1[2679:2672] < top_0[2671:2664]) ? 1 : 0;
assign detect_min[333][1] = (mid_1[2679:2672] < top_0[2679:2672]) ? 1 : 0;
assign detect_min[333][2] = (mid_1[2679:2672] < top_0[2687:2680]) ? 1 : 0;
assign detect_min[333][3] = (mid_1[2679:2672] < top_1[2671:2664]) ? 1 : 0;
assign detect_min[333][4] = (mid_1[2679:2672] < top_1[2679:2672]) ? 1 : 0;
assign detect_min[333][5] = (mid_1[2679:2672] < top_1[2687:2680]) ? 1 : 0;
assign detect_min[333][6] = (mid_1[2679:2672] < top_2[2671:2664]) ? 1 : 0;
assign detect_min[333][7] = (mid_1[2679:2672] < top_2[2679:2672]) ? 1 : 0;
assign detect_min[333][8] = (mid_1[2679:2672] < top_2[2687:2680]) ? 1 : 0;
assign detect_min[333][9] = (mid_1[2679:2672] < mid_0[2671:2664]) ? 1 : 0;
assign detect_min[333][10] = (mid_1[2679:2672] < mid_0[2679:2672]) ? 1 : 0;
assign detect_min[333][11] = (mid_1[2679:2672] < mid_0[2687:2680]) ? 1 : 0;
assign detect_min[333][12] = (mid_1[2679:2672] < mid_1[2671:2664]) ? 1 : 0;
assign detect_min[333][13] = (mid_1[2679:2672] < mid_1[2687:2680]) ? 1 : 0;
assign detect_min[333][14] = (mid_1[2679:2672] < mid_2[2671:2664]) ? 1 : 0;
assign detect_min[333][15] = (mid_1[2679:2672] < mid_2[2679:2672]) ? 1 : 0;
assign detect_min[333][16] = (mid_1[2679:2672] < mid_2[2687:2680]) ? 1 : 0;
assign detect_min[333][17] = (mid_1[2679:2672] < btm_0[2671:2664]) ? 1 : 0;
assign detect_min[333][18] = (mid_1[2679:2672] < btm_0[2679:2672]) ? 1 : 0;
assign detect_min[333][19] = (mid_1[2679:2672] < btm_0[2687:2680]) ? 1 : 0;
assign detect_min[333][20] = (mid_1[2679:2672] < btm_1[2671:2664]) ? 1 : 0;
assign detect_min[333][21] = (mid_1[2679:2672] < btm_1[2679:2672]) ? 1 : 0;
assign detect_min[333][22] = (mid_1[2679:2672] < btm_1[2687:2680]) ? 1 : 0;
assign detect_min[333][23] = (mid_1[2679:2672] < btm_2[2671:2664]) ? 1 : 0;
assign detect_min[333][24] = (mid_1[2679:2672] < btm_2[2679:2672]) ? 1 : 0;
assign detect_min[333][25] = (mid_1[2679:2672] < btm_2[2687:2680]) ? 1 : 0;

assign detect_min[334][0] = (mid_1[2687:2680] < top_0[2679:2672]) ? 1 : 0;
assign detect_min[334][1] = (mid_1[2687:2680] < top_0[2687:2680]) ? 1 : 0;
assign detect_min[334][2] = (mid_1[2687:2680] < top_0[2695:2688]) ? 1 : 0;
assign detect_min[334][3] = (mid_1[2687:2680] < top_1[2679:2672]) ? 1 : 0;
assign detect_min[334][4] = (mid_1[2687:2680] < top_1[2687:2680]) ? 1 : 0;
assign detect_min[334][5] = (mid_1[2687:2680] < top_1[2695:2688]) ? 1 : 0;
assign detect_min[334][6] = (mid_1[2687:2680] < top_2[2679:2672]) ? 1 : 0;
assign detect_min[334][7] = (mid_1[2687:2680] < top_2[2687:2680]) ? 1 : 0;
assign detect_min[334][8] = (mid_1[2687:2680] < top_2[2695:2688]) ? 1 : 0;
assign detect_min[334][9] = (mid_1[2687:2680] < mid_0[2679:2672]) ? 1 : 0;
assign detect_min[334][10] = (mid_1[2687:2680] < mid_0[2687:2680]) ? 1 : 0;
assign detect_min[334][11] = (mid_1[2687:2680] < mid_0[2695:2688]) ? 1 : 0;
assign detect_min[334][12] = (mid_1[2687:2680] < mid_1[2679:2672]) ? 1 : 0;
assign detect_min[334][13] = (mid_1[2687:2680] < mid_1[2695:2688]) ? 1 : 0;
assign detect_min[334][14] = (mid_1[2687:2680] < mid_2[2679:2672]) ? 1 : 0;
assign detect_min[334][15] = (mid_1[2687:2680] < mid_2[2687:2680]) ? 1 : 0;
assign detect_min[334][16] = (mid_1[2687:2680] < mid_2[2695:2688]) ? 1 : 0;
assign detect_min[334][17] = (mid_1[2687:2680] < btm_0[2679:2672]) ? 1 : 0;
assign detect_min[334][18] = (mid_1[2687:2680] < btm_0[2687:2680]) ? 1 : 0;
assign detect_min[334][19] = (mid_1[2687:2680] < btm_0[2695:2688]) ? 1 : 0;
assign detect_min[334][20] = (mid_1[2687:2680] < btm_1[2679:2672]) ? 1 : 0;
assign detect_min[334][21] = (mid_1[2687:2680] < btm_1[2687:2680]) ? 1 : 0;
assign detect_min[334][22] = (mid_1[2687:2680] < btm_1[2695:2688]) ? 1 : 0;
assign detect_min[334][23] = (mid_1[2687:2680] < btm_2[2679:2672]) ? 1 : 0;
assign detect_min[334][24] = (mid_1[2687:2680] < btm_2[2687:2680]) ? 1 : 0;
assign detect_min[334][25] = (mid_1[2687:2680] < btm_2[2695:2688]) ? 1 : 0;

assign detect_min[335][0] = (mid_1[2695:2688] < top_0[2687:2680]) ? 1 : 0;
assign detect_min[335][1] = (mid_1[2695:2688] < top_0[2695:2688]) ? 1 : 0;
assign detect_min[335][2] = (mid_1[2695:2688] < top_0[2703:2696]) ? 1 : 0;
assign detect_min[335][3] = (mid_1[2695:2688] < top_1[2687:2680]) ? 1 : 0;
assign detect_min[335][4] = (mid_1[2695:2688] < top_1[2695:2688]) ? 1 : 0;
assign detect_min[335][5] = (mid_1[2695:2688] < top_1[2703:2696]) ? 1 : 0;
assign detect_min[335][6] = (mid_1[2695:2688] < top_2[2687:2680]) ? 1 : 0;
assign detect_min[335][7] = (mid_1[2695:2688] < top_2[2695:2688]) ? 1 : 0;
assign detect_min[335][8] = (mid_1[2695:2688] < top_2[2703:2696]) ? 1 : 0;
assign detect_min[335][9] = (mid_1[2695:2688] < mid_0[2687:2680]) ? 1 : 0;
assign detect_min[335][10] = (mid_1[2695:2688] < mid_0[2695:2688]) ? 1 : 0;
assign detect_min[335][11] = (mid_1[2695:2688] < mid_0[2703:2696]) ? 1 : 0;
assign detect_min[335][12] = (mid_1[2695:2688] < mid_1[2687:2680]) ? 1 : 0;
assign detect_min[335][13] = (mid_1[2695:2688] < mid_1[2703:2696]) ? 1 : 0;
assign detect_min[335][14] = (mid_1[2695:2688] < mid_2[2687:2680]) ? 1 : 0;
assign detect_min[335][15] = (mid_1[2695:2688] < mid_2[2695:2688]) ? 1 : 0;
assign detect_min[335][16] = (mid_1[2695:2688] < mid_2[2703:2696]) ? 1 : 0;
assign detect_min[335][17] = (mid_1[2695:2688] < btm_0[2687:2680]) ? 1 : 0;
assign detect_min[335][18] = (mid_1[2695:2688] < btm_0[2695:2688]) ? 1 : 0;
assign detect_min[335][19] = (mid_1[2695:2688] < btm_0[2703:2696]) ? 1 : 0;
assign detect_min[335][20] = (mid_1[2695:2688] < btm_1[2687:2680]) ? 1 : 0;
assign detect_min[335][21] = (mid_1[2695:2688] < btm_1[2695:2688]) ? 1 : 0;
assign detect_min[335][22] = (mid_1[2695:2688] < btm_1[2703:2696]) ? 1 : 0;
assign detect_min[335][23] = (mid_1[2695:2688] < btm_2[2687:2680]) ? 1 : 0;
assign detect_min[335][24] = (mid_1[2695:2688] < btm_2[2695:2688]) ? 1 : 0;
assign detect_min[335][25] = (mid_1[2695:2688] < btm_2[2703:2696]) ? 1 : 0;

assign detect_min[336][0] = (mid_1[2703:2696] < top_0[2695:2688]) ? 1 : 0;
assign detect_min[336][1] = (mid_1[2703:2696] < top_0[2703:2696]) ? 1 : 0;
assign detect_min[336][2] = (mid_1[2703:2696] < top_0[2711:2704]) ? 1 : 0;
assign detect_min[336][3] = (mid_1[2703:2696] < top_1[2695:2688]) ? 1 : 0;
assign detect_min[336][4] = (mid_1[2703:2696] < top_1[2703:2696]) ? 1 : 0;
assign detect_min[336][5] = (mid_1[2703:2696] < top_1[2711:2704]) ? 1 : 0;
assign detect_min[336][6] = (mid_1[2703:2696] < top_2[2695:2688]) ? 1 : 0;
assign detect_min[336][7] = (mid_1[2703:2696] < top_2[2703:2696]) ? 1 : 0;
assign detect_min[336][8] = (mid_1[2703:2696] < top_2[2711:2704]) ? 1 : 0;
assign detect_min[336][9] = (mid_1[2703:2696] < mid_0[2695:2688]) ? 1 : 0;
assign detect_min[336][10] = (mid_1[2703:2696] < mid_0[2703:2696]) ? 1 : 0;
assign detect_min[336][11] = (mid_1[2703:2696] < mid_0[2711:2704]) ? 1 : 0;
assign detect_min[336][12] = (mid_1[2703:2696] < mid_1[2695:2688]) ? 1 : 0;
assign detect_min[336][13] = (mid_1[2703:2696] < mid_1[2711:2704]) ? 1 : 0;
assign detect_min[336][14] = (mid_1[2703:2696] < mid_2[2695:2688]) ? 1 : 0;
assign detect_min[336][15] = (mid_1[2703:2696] < mid_2[2703:2696]) ? 1 : 0;
assign detect_min[336][16] = (mid_1[2703:2696] < mid_2[2711:2704]) ? 1 : 0;
assign detect_min[336][17] = (mid_1[2703:2696] < btm_0[2695:2688]) ? 1 : 0;
assign detect_min[336][18] = (mid_1[2703:2696] < btm_0[2703:2696]) ? 1 : 0;
assign detect_min[336][19] = (mid_1[2703:2696] < btm_0[2711:2704]) ? 1 : 0;
assign detect_min[336][20] = (mid_1[2703:2696] < btm_1[2695:2688]) ? 1 : 0;
assign detect_min[336][21] = (mid_1[2703:2696] < btm_1[2703:2696]) ? 1 : 0;
assign detect_min[336][22] = (mid_1[2703:2696] < btm_1[2711:2704]) ? 1 : 0;
assign detect_min[336][23] = (mid_1[2703:2696] < btm_2[2695:2688]) ? 1 : 0;
assign detect_min[336][24] = (mid_1[2703:2696] < btm_2[2703:2696]) ? 1 : 0;
assign detect_min[336][25] = (mid_1[2703:2696] < btm_2[2711:2704]) ? 1 : 0;

assign detect_min[337][0] = (mid_1[2711:2704] < top_0[2703:2696]) ? 1 : 0;
assign detect_min[337][1] = (mid_1[2711:2704] < top_0[2711:2704]) ? 1 : 0;
assign detect_min[337][2] = (mid_1[2711:2704] < top_0[2719:2712]) ? 1 : 0;
assign detect_min[337][3] = (mid_1[2711:2704] < top_1[2703:2696]) ? 1 : 0;
assign detect_min[337][4] = (mid_1[2711:2704] < top_1[2711:2704]) ? 1 : 0;
assign detect_min[337][5] = (mid_1[2711:2704] < top_1[2719:2712]) ? 1 : 0;
assign detect_min[337][6] = (mid_1[2711:2704] < top_2[2703:2696]) ? 1 : 0;
assign detect_min[337][7] = (mid_1[2711:2704] < top_2[2711:2704]) ? 1 : 0;
assign detect_min[337][8] = (mid_1[2711:2704] < top_2[2719:2712]) ? 1 : 0;
assign detect_min[337][9] = (mid_1[2711:2704] < mid_0[2703:2696]) ? 1 : 0;
assign detect_min[337][10] = (mid_1[2711:2704] < mid_0[2711:2704]) ? 1 : 0;
assign detect_min[337][11] = (mid_1[2711:2704] < mid_0[2719:2712]) ? 1 : 0;
assign detect_min[337][12] = (mid_1[2711:2704] < mid_1[2703:2696]) ? 1 : 0;
assign detect_min[337][13] = (mid_1[2711:2704] < mid_1[2719:2712]) ? 1 : 0;
assign detect_min[337][14] = (mid_1[2711:2704] < mid_2[2703:2696]) ? 1 : 0;
assign detect_min[337][15] = (mid_1[2711:2704] < mid_2[2711:2704]) ? 1 : 0;
assign detect_min[337][16] = (mid_1[2711:2704] < mid_2[2719:2712]) ? 1 : 0;
assign detect_min[337][17] = (mid_1[2711:2704] < btm_0[2703:2696]) ? 1 : 0;
assign detect_min[337][18] = (mid_1[2711:2704] < btm_0[2711:2704]) ? 1 : 0;
assign detect_min[337][19] = (mid_1[2711:2704] < btm_0[2719:2712]) ? 1 : 0;
assign detect_min[337][20] = (mid_1[2711:2704] < btm_1[2703:2696]) ? 1 : 0;
assign detect_min[337][21] = (mid_1[2711:2704] < btm_1[2711:2704]) ? 1 : 0;
assign detect_min[337][22] = (mid_1[2711:2704] < btm_1[2719:2712]) ? 1 : 0;
assign detect_min[337][23] = (mid_1[2711:2704] < btm_2[2703:2696]) ? 1 : 0;
assign detect_min[337][24] = (mid_1[2711:2704] < btm_2[2711:2704]) ? 1 : 0;
assign detect_min[337][25] = (mid_1[2711:2704] < btm_2[2719:2712]) ? 1 : 0;

assign detect_min[338][0] = (mid_1[2719:2712] < top_0[2711:2704]) ? 1 : 0;
assign detect_min[338][1] = (mid_1[2719:2712] < top_0[2719:2712]) ? 1 : 0;
assign detect_min[338][2] = (mid_1[2719:2712] < top_0[2727:2720]) ? 1 : 0;
assign detect_min[338][3] = (mid_1[2719:2712] < top_1[2711:2704]) ? 1 : 0;
assign detect_min[338][4] = (mid_1[2719:2712] < top_1[2719:2712]) ? 1 : 0;
assign detect_min[338][5] = (mid_1[2719:2712] < top_1[2727:2720]) ? 1 : 0;
assign detect_min[338][6] = (mid_1[2719:2712] < top_2[2711:2704]) ? 1 : 0;
assign detect_min[338][7] = (mid_1[2719:2712] < top_2[2719:2712]) ? 1 : 0;
assign detect_min[338][8] = (mid_1[2719:2712] < top_2[2727:2720]) ? 1 : 0;
assign detect_min[338][9] = (mid_1[2719:2712] < mid_0[2711:2704]) ? 1 : 0;
assign detect_min[338][10] = (mid_1[2719:2712] < mid_0[2719:2712]) ? 1 : 0;
assign detect_min[338][11] = (mid_1[2719:2712] < mid_0[2727:2720]) ? 1 : 0;
assign detect_min[338][12] = (mid_1[2719:2712] < mid_1[2711:2704]) ? 1 : 0;
assign detect_min[338][13] = (mid_1[2719:2712] < mid_1[2727:2720]) ? 1 : 0;
assign detect_min[338][14] = (mid_1[2719:2712] < mid_2[2711:2704]) ? 1 : 0;
assign detect_min[338][15] = (mid_1[2719:2712] < mid_2[2719:2712]) ? 1 : 0;
assign detect_min[338][16] = (mid_1[2719:2712] < mid_2[2727:2720]) ? 1 : 0;
assign detect_min[338][17] = (mid_1[2719:2712] < btm_0[2711:2704]) ? 1 : 0;
assign detect_min[338][18] = (mid_1[2719:2712] < btm_0[2719:2712]) ? 1 : 0;
assign detect_min[338][19] = (mid_1[2719:2712] < btm_0[2727:2720]) ? 1 : 0;
assign detect_min[338][20] = (mid_1[2719:2712] < btm_1[2711:2704]) ? 1 : 0;
assign detect_min[338][21] = (mid_1[2719:2712] < btm_1[2719:2712]) ? 1 : 0;
assign detect_min[338][22] = (mid_1[2719:2712] < btm_1[2727:2720]) ? 1 : 0;
assign detect_min[338][23] = (mid_1[2719:2712] < btm_2[2711:2704]) ? 1 : 0;
assign detect_min[338][24] = (mid_1[2719:2712] < btm_2[2719:2712]) ? 1 : 0;
assign detect_min[338][25] = (mid_1[2719:2712] < btm_2[2727:2720]) ? 1 : 0;

assign detect_min[339][0] = (mid_1[2727:2720] < top_0[2719:2712]) ? 1 : 0;
assign detect_min[339][1] = (mid_1[2727:2720] < top_0[2727:2720]) ? 1 : 0;
assign detect_min[339][2] = (mid_1[2727:2720] < top_0[2735:2728]) ? 1 : 0;
assign detect_min[339][3] = (mid_1[2727:2720] < top_1[2719:2712]) ? 1 : 0;
assign detect_min[339][4] = (mid_1[2727:2720] < top_1[2727:2720]) ? 1 : 0;
assign detect_min[339][5] = (mid_1[2727:2720] < top_1[2735:2728]) ? 1 : 0;
assign detect_min[339][6] = (mid_1[2727:2720] < top_2[2719:2712]) ? 1 : 0;
assign detect_min[339][7] = (mid_1[2727:2720] < top_2[2727:2720]) ? 1 : 0;
assign detect_min[339][8] = (mid_1[2727:2720] < top_2[2735:2728]) ? 1 : 0;
assign detect_min[339][9] = (mid_1[2727:2720] < mid_0[2719:2712]) ? 1 : 0;
assign detect_min[339][10] = (mid_1[2727:2720] < mid_0[2727:2720]) ? 1 : 0;
assign detect_min[339][11] = (mid_1[2727:2720] < mid_0[2735:2728]) ? 1 : 0;
assign detect_min[339][12] = (mid_1[2727:2720] < mid_1[2719:2712]) ? 1 : 0;
assign detect_min[339][13] = (mid_1[2727:2720] < mid_1[2735:2728]) ? 1 : 0;
assign detect_min[339][14] = (mid_1[2727:2720] < mid_2[2719:2712]) ? 1 : 0;
assign detect_min[339][15] = (mid_1[2727:2720] < mid_2[2727:2720]) ? 1 : 0;
assign detect_min[339][16] = (mid_1[2727:2720] < mid_2[2735:2728]) ? 1 : 0;
assign detect_min[339][17] = (mid_1[2727:2720] < btm_0[2719:2712]) ? 1 : 0;
assign detect_min[339][18] = (mid_1[2727:2720] < btm_0[2727:2720]) ? 1 : 0;
assign detect_min[339][19] = (mid_1[2727:2720] < btm_0[2735:2728]) ? 1 : 0;
assign detect_min[339][20] = (mid_1[2727:2720] < btm_1[2719:2712]) ? 1 : 0;
assign detect_min[339][21] = (mid_1[2727:2720] < btm_1[2727:2720]) ? 1 : 0;
assign detect_min[339][22] = (mid_1[2727:2720] < btm_1[2735:2728]) ? 1 : 0;
assign detect_min[339][23] = (mid_1[2727:2720] < btm_2[2719:2712]) ? 1 : 0;
assign detect_min[339][24] = (mid_1[2727:2720] < btm_2[2727:2720]) ? 1 : 0;
assign detect_min[339][25] = (mid_1[2727:2720] < btm_2[2735:2728]) ? 1 : 0;

assign detect_min[340][0] = (mid_1[2735:2728] < top_0[2727:2720]) ? 1 : 0;
assign detect_min[340][1] = (mid_1[2735:2728] < top_0[2735:2728]) ? 1 : 0;
assign detect_min[340][2] = (mid_1[2735:2728] < top_0[2743:2736]) ? 1 : 0;
assign detect_min[340][3] = (mid_1[2735:2728] < top_1[2727:2720]) ? 1 : 0;
assign detect_min[340][4] = (mid_1[2735:2728] < top_1[2735:2728]) ? 1 : 0;
assign detect_min[340][5] = (mid_1[2735:2728] < top_1[2743:2736]) ? 1 : 0;
assign detect_min[340][6] = (mid_1[2735:2728] < top_2[2727:2720]) ? 1 : 0;
assign detect_min[340][7] = (mid_1[2735:2728] < top_2[2735:2728]) ? 1 : 0;
assign detect_min[340][8] = (mid_1[2735:2728] < top_2[2743:2736]) ? 1 : 0;
assign detect_min[340][9] = (mid_1[2735:2728] < mid_0[2727:2720]) ? 1 : 0;
assign detect_min[340][10] = (mid_1[2735:2728] < mid_0[2735:2728]) ? 1 : 0;
assign detect_min[340][11] = (mid_1[2735:2728] < mid_0[2743:2736]) ? 1 : 0;
assign detect_min[340][12] = (mid_1[2735:2728] < mid_1[2727:2720]) ? 1 : 0;
assign detect_min[340][13] = (mid_1[2735:2728] < mid_1[2743:2736]) ? 1 : 0;
assign detect_min[340][14] = (mid_1[2735:2728] < mid_2[2727:2720]) ? 1 : 0;
assign detect_min[340][15] = (mid_1[2735:2728] < mid_2[2735:2728]) ? 1 : 0;
assign detect_min[340][16] = (mid_1[2735:2728] < mid_2[2743:2736]) ? 1 : 0;
assign detect_min[340][17] = (mid_1[2735:2728] < btm_0[2727:2720]) ? 1 : 0;
assign detect_min[340][18] = (mid_1[2735:2728] < btm_0[2735:2728]) ? 1 : 0;
assign detect_min[340][19] = (mid_1[2735:2728] < btm_0[2743:2736]) ? 1 : 0;
assign detect_min[340][20] = (mid_1[2735:2728] < btm_1[2727:2720]) ? 1 : 0;
assign detect_min[340][21] = (mid_1[2735:2728] < btm_1[2735:2728]) ? 1 : 0;
assign detect_min[340][22] = (mid_1[2735:2728] < btm_1[2743:2736]) ? 1 : 0;
assign detect_min[340][23] = (mid_1[2735:2728] < btm_2[2727:2720]) ? 1 : 0;
assign detect_min[340][24] = (mid_1[2735:2728] < btm_2[2735:2728]) ? 1 : 0;
assign detect_min[340][25] = (mid_1[2735:2728] < btm_2[2743:2736]) ? 1 : 0;

assign detect_min[341][0] = (mid_1[2743:2736] < top_0[2735:2728]) ? 1 : 0;
assign detect_min[341][1] = (mid_1[2743:2736] < top_0[2743:2736]) ? 1 : 0;
assign detect_min[341][2] = (mid_1[2743:2736] < top_0[2751:2744]) ? 1 : 0;
assign detect_min[341][3] = (mid_1[2743:2736] < top_1[2735:2728]) ? 1 : 0;
assign detect_min[341][4] = (mid_1[2743:2736] < top_1[2743:2736]) ? 1 : 0;
assign detect_min[341][5] = (mid_1[2743:2736] < top_1[2751:2744]) ? 1 : 0;
assign detect_min[341][6] = (mid_1[2743:2736] < top_2[2735:2728]) ? 1 : 0;
assign detect_min[341][7] = (mid_1[2743:2736] < top_2[2743:2736]) ? 1 : 0;
assign detect_min[341][8] = (mid_1[2743:2736] < top_2[2751:2744]) ? 1 : 0;
assign detect_min[341][9] = (mid_1[2743:2736] < mid_0[2735:2728]) ? 1 : 0;
assign detect_min[341][10] = (mid_1[2743:2736] < mid_0[2743:2736]) ? 1 : 0;
assign detect_min[341][11] = (mid_1[2743:2736] < mid_0[2751:2744]) ? 1 : 0;
assign detect_min[341][12] = (mid_1[2743:2736] < mid_1[2735:2728]) ? 1 : 0;
assign detect_min[341][13] = (mid_1[2743:2736] < mid_1[2751:2744]) ? 1 : 0;
assign detect_min[341][14] = (mid_1[2743:2736] < mid_2[2735:2728]) ? 1 : 0;
assign detect_min[341][15] = (mid_1[2743:2736] < mid_2[2743:2736]) ? 1 : 0;
assign detect_min[341][16] = (mid_1[2743:2736] < mid_2[2751:2744]) ? 1 : 0;
assign detect_min[341][17] = (mid_1[2743:2736] < btm_0[2735:2728]) ? 1 : 0;
assign detect_min[341][18] = (mid_1[2743:2736] < btm_0[2743:2736]) ? 1 : 0;
assign detect_min[341][19] = (mid_1[2743:2736] < btm_0[2751:2744]) ? 1 : 0;
assign detect_min[341][20] = (mid_1[2743:2736] < btm_1[2735:2728]) ? 1 : 0;
assign detect_min[341][21] = (mid_1[2743:2736] < btm_1[2743:2736]) ? 1 : 0;
assign detect_min[341][22] = (mid_1[2743:2736] < btm_1[2751:2744]) ? 1 : 0;
assign detect_min[341][23] = (mid_1[2743:2736] < btm_2[2735:2728]) ? 1 : 0;
assign detect_min[341][24] = (mid_1[2743:2736] < btm_2[2743:2736]) ? 1 : 0;
assign detect_min[341][25] = (mid_1[2743:2736] < btm_2[2751:2744]) ? 1 : 0;

assign detect_min[342][0] = (mid_1[2751:2744] < top_0[2743:2736]) ? 1 : 0;
assign detect_min[342][1] = (mid_1[2751:2744] < top_0[2751:2744]) ? 1 : 0;
assign detect_min[342][2] = (mid_1[2751:2744] < top_0[2759:2752]) ? 1 : 0;
assign detect_min[342][3] = (mid_1[2751:2744] < top_1[2743:2736]) ? 1 : 0;
assign detect_min[342][4] = (mid_1[2751:2744] < top_1[2751:2744]) ? 1 : 0;
assign detect_min[342][5] = (mid_1[2751:2744] < top_1[2759:2752]) ? 1 : 0;
assign detect_min[342][6] = (mid_1[2751:2744] < top_2[2743:2736]) ? 1 : 0;
assign detect_min[342][7] = (mid_1[2751:2744] < top_2[2751:2744]) ? 1 : 0;
assign detect_min[342][8] = (mid_1[2751:2744] < top_2[2759:2752]) ? 1 : 0;
assign detect_min[342][9] = (mid_1[2751:2744] < mid_0[2743:2736]) ? 1 : 0;
assign detect_min[342][10] = (mid_1[2751:2744] < mid_0[2751:2744]) ? 1 : 0;
assign detect_min[342][11] = (mid_1[2751:2744] < mid_0[2759:2752]) ? 1 : 0;
assign detect_min[342][12] = (mid_1[2751:2744] < mid_1[2743:2736]) ? 1 : 0;
assign detect_min[342][13] = (mid_1[2751:2744] < mid_1[2759:2752]) ? 1 : 0;
assign detect_min[342][14] = (mid_1[2751:2744] < mid_2[2743:2736]) ? 1 : 0;
assign detect_min[342][15] = (mid_1[2751:2744] < mid_2[2751:2744]) ? 1 : 0;
assign detect_min[342][16] = (mid_1[2751:2744] < mid_2[2759:2752]) ? 1 : 0;
assign detect_min[342][17] = (mid_1[2751:2744] < btm_0[2743:2736]) ? 1 : 0;
assign detect_min[342][18] = (mid_1[2751:2744] < btm_0[2751:2744]) ? 1 : 0;
assign detect_min[342][19] = (mid_1[2751:2744] < btm_0[2759:2752]) ? 1 : 0;
assign detect_min[342][20] = (mid_1[2751:2744] < btm_1[2743:2736]) ? 1 : 0;
assign detect_min[342][21] = (mid_1[2751:2744] < btm_1[2751:2744]) ? 1 : 0;
assign detect_min[342][22] = (mid_1[2751:2744] < btm_1[2759:2752]) ? 1 : 0;
assign detect_min[342][23] = (mid_1[2751:2744] < btm_2[2743:2736]) ? 1 : 0;
assign detect_min[342][24] = (mid_1[2751:2744] < btm_2[2751:2744]) ? 1 : 0;
assign detect_min[342][25] = (mid_1[2751:2744] < btm_2[2759:2752]) ? 1 : 0;

assign detect_min[343][0] = (mid_1[2759:2752] < top_0[2751:2744]) ? 1 : 0;
assign detect_min[343][1] = (mid_1[2759:2752] < top_0[2759:2752]) ? 1 : 0;
assign detect_min[343][2] = (mid_1[2759:2752] < top_0[2767:2760]) ? 1 : 0;
assign detect_min[343][3] = (mid_1[2759:2752] < top_1[2751:2744]) ? 1 : 0;
assign detect_min[343][4] = (mid_1[2759:2752] < top_1[2759:2752]) ? 1 : 0;
assign detect_min[343][5] = (mid_1[2759:2752] < top_1[2767:2760]) ? 1 : 0;
assign detect_min[343][6] = (mid_1[2759:2752] < top_2[2751:2744]) ? 1 : 0;
assign detect_min[343][7] = (mid_1[2759:2752] < top_2[2759:2752]) ? 1 : 0;
assign detect_min[343][8] = (mid_1[2759:2752] < top_2[2767:2760]) ? 1 : 0;
assign detect_min[343][9] = (mid_1[2759:2752] < mid_0[2751:2744]) ? 1 : 0;
assign detect_min[343][10] = (mid_1[2759:2752] < mid_0[2759:2752]) ? 1 : 0;
assign detect_min[343][11] = (mid_1[2759:2752] < mid_0[2767:2760]) ? 1 : 0;
assign detect_min[343][12] = (mid_1[2759:2752] < mid_1[2751:2744]) ? 1 : 0;
assign detect_min[343][13] = (mid_1[2759:2752] < mid_1[2767:2760]) ? 1 : 0;
assign detect_min[343][14] = (mid_1[2759:2752] < mid_2[2751:2744]) ? 1 : 0;
assign detect_min[343][15] = (mid_1[2759:2752] < mid_2[2759:2752]) ? 1 : 0;
assign detect_min[343][16] = (mid_1[2759:2752] < mid_2[2767:2760]) ? 1 : 0;
assign detect_min[343][17] = (mid_1[2759:2752] < btm_0[2751:2744]) ? 1 : 0;
assign detect_min[343][18] = (mid_1[2759:2752] < btm_0[2759:2752]) ? 1 : 0;
assign detect_min[343][19] = (mid_1[2759:2752] < btm_0[2767:2760]) ? 1 : 0;
assign detect_min[343][20] = (mid_1[2759:2752] < btm_1[2751:2744]) ? 1 : 0;
assign detect_min[343][21] = (mid_1[2759:2752] < btm_1[2759:2752]) ? 1 : 0;
assign detect_min[343][22] = (mid_1[2759:2752] < btm_1[2767:2760]) ? 1 : 0;
assign detect_min[343][23] = (mid_1[2759:2752] < btm_2[2751:2744]) ? 1 : 0;
assign detect_min[343][24] = (mid_1[2759:2752] < btm_2[2759:2752]) ? 1 : 0;
assign detect_min[343][25] = (mid_1[2759:2752] < btm_2[2767:2760]) ? 1 : 0;

assign detect_min[344][0] = (mid_1[2767:2760] < top_0[2759:2752]) ? 1 : 0;
assign detect_min[344][1] = (mid_1[2767:2760] < top_0[2767:2760]) ? 1 : 0;
assign detect_min[344][2] = (mid_1[2767:2760] < top_0[2775:2768]) ? 1 : 0;
assign detect_min[344][3] = (mid_1[2767:2760] < top_1[2759:2752]) ? 1 : 0;
assign detect_min[344][4] = (mid_1[2767:2760] < top_1[2767:2760]) ? 1 : 0;
assign detect_min[344][5] = (mid_1[2767:2760] < top_1[2775:2768]) ? 1 : 0;
assign detect_min[344][6] = (mid_1[2767:2760] < top_2[2759:2752]) ? 1 : 0;
assign detect_min[344][7] = (mid_1[2767:2760] < top_2[2767:2760]) ? 1 : 0;
assign detect_min[344][8] = (mid_1[2767:2760] < top_2[2775:2768]) ? 1 : 0;
assign detect_min[344][9] = (mid_1[2767:2760] < mid_0[2759:2752]) ? 1 : 0;
assign detect_min[344][10] = (mid_1[2767:2760] < mid_0[2767:2760]) ? 1 : 0;
assign detect_min[344][11] = (mid_1[2767:2760] < mid_0[2775:2768]) ? 1 : 0;
assign detect_min[344][12] = (mid_1[2767:2760] < mid_1[2759:2752]) ? 1 : 0;
assign detect_min[344][13] = (mid_1[2767:2760] < mid_1[2775:2768]) ? 1 : 0;
assign detect_min[344][14] = (mid_1[2767:2760] < mid_2[2759:2752]) ? 1 : 0;
assign detect_min[344][15] = (mid_1[2767:2760] < mid_2[2767:2760]) ? 1 : 0;
assign detect_min[344][16] = (mid_1[2767:2760] < mid_2[2775:2768]) ? 1 : 0;
assign detect_min[344][17] = (mid_1[2767:2760] < btm_0[2759:2752]) ? 1 : 0;
assign detect_min[344][18] = (mid_1[2767:2760] < btm_0[2767:2760]) ? 1 : 0;
assign detect_min[344][19] = (mid_1[2767:2760] < btm_0[2775:2768]) ? 1 : 0;
assign detect_min[344][20] = (mid_1[2767:2760] < btm_1[2759:2752]) ? 1 : 0;
assign detect_min[344][21] = (mid_1[2767:2760] < btm_1[2767:2760]) ? 1 : 0;
assign detect_min[344][22] = (mid_1[2767:2760] < btm_1[2775:2768]) ? 1 : 0;
assign detect_min[344][23] = (mid_1[2767:2760] < btm_2[2759:2752]) ? 1 : 0;
assign detect_min[344][24] = (mid_1[2767:2760] < btm_2[2767:2760]) ? 1 : 0;
assign detect_min[344][25] = (mid_1[2767:2760] < btm_2[2775:2768]) ? 1 : 0;

assign detect_min[345][0] = (mid_1[2775:2768] < top_0[2767:2760]) ? 1 : 0;
assign detect_min[345][1] = (mid_1[2775:2768] < top_0[2775:2768]) ? 1 : 0;
assign detect_min[345][2] = (mid_1[2775:2768] < top_0[2783:2776]) ? 1 : 0;
assign detect_min[345][3] = (mid_1[2775:2768] < top_1[2767:2760]) ? 1 : 0;
assign detect_min[345][4] = (mid_1[2775:2768] < top_1[2775:2768]) ? 1 : 0;
assign detect_min[345][5] = (mid_1[2775:2768] < top_1[2783:2776]) ? 1 : 0;
assign detect_min[345][6] = (mid_1[2775:2768] < top_2[2767:2760]) ? 1 : 0;
assign detect_min[345][7] = (mid_1[2775:2768] < top_2[2775:2768]) ? 1 : 0;
assign detect_min[345][8] = (mid_1[2775:2768] < top_2[2783:2776]) ? 1 : 0;
assign detect_min[345][9] = (mid_1[2775:2768] < mid_0[2767:2760]) ? 1 : 0;
assign detect_min[345][10] = (mid_1[2775:2768] < mid_0[2775:2768]) ? 1 : 0;
assign detect_min[345][11] = (mid_1[2775:2768] < mid_0[2783:2776]) ? 1 : 0;
assign detect_min[345][12] = (mid_1[2775:2768] < mid_1[2767:2760]) ? 1 : 0;
assign detect_min[345][13] = (mid_1[2775:2768] < mid_1[2783:2776]) ? 1 : 0;
assign detect_min[345][14] = (mid_1[2775:2768] < mid_2[2767:2760]) ? 1 : 0;
assign detect_min[345][15] = (mid_1[2775:2768] < mid_2[2775:2768]) ? 1 : 0;
assign detect_min[345][16] = (mid_1[2775:2768] < mid_2[2783:2776]) ? 1 : 0;
assign detect_min[345][17] = (mid_1[2775:2768] < btm_0[2767:2760]) ? 1 : 0;
assign detect_min[345][18] = (mid_1[2775:2768] < btm_0[2775:2768]) ? 1 : 0;
assign detect_min[345][19] = (mid_1[2775:2768] < btm_0[2783:2776]) ? 1 : 0;
assign detect_min[345][20] = (mid_1[2775:2768] < btm_1[2767:2760]) ? 1 : 0;
assign detect_min[345][21] = (mid_1[2775:2768] < btm_1[2775:2768]) ? 1 : 0;
assign detect_min[345][22] = (mid_1[2775:2768] < btm_1[2783:2776]) ? 1 : 0;
assign detect_min[345][23] = (mid_1[2775:2768] < btm_2[2767:2760]) ? 1 : 0;
assign detect_min[345][24] = (mid_1[2775:2768] < btm_2[2775:2768]) ? 1 : 0;
assign detect_min[345][25] = (mid_1[2775:2768] < btm_2[2783:2776]) ? 1 : 0;

assign detect_min[346][0] = (mid_1[2783:2776] < top_0[2775:2768]) ? 1 : 0;
assign detect_min[346][1] = (mid_1[2783:2776] < top_0[2783:2776]) ? 1 : 0;
assign detect_min[346][2] = (mid_1[2783:2776] < top_0[2791:2784]) ? 1 : 0;
assign detect_min[346][3] = (mid_1[2783:2776] < top_1[2775:2768]) ? 1 : 0;
assign detect_min[346][4] = (mid_1[2783:2776] < top_1[2783:2776]) ? 1 : 0;
assign detect_min[346][5] = (mid_1[2783:2776] < top_1[2791:2784]) ? 1 : 0;
assign detect_min[346][6] = (mid_1[2783:2776] < top_2[2775:2768]) ? 1 : 0;
assign detect_min[346][7] = (mid_1[2783:2776] < top_2[2783:2776]) ? 1 : 0;
assign detect_min[346][8] = (mid_1[2783:2776] < top_2[2791:2784]) ? 1 : 0;
assign detect_min[346][9] = (mid_1[2783:2776] < mid_0[2775:2768]) ? 1 : 0;
assign detect_min[346][10] = (mid_1[2783:2776] < mid_0[2783:2776]) ? 1 : 0;
assign detect_min[346][11] = (mid_1[2783:2776] < mid_0[2791:2784]) ? 1 : 0;
assign detect_min[346][12] = (mid_1[2783:2776] < mid_1[2775:2768]) ? 1 : 0;
assign detect_min[346][13] = (mid_1[2783:2776] < mid_1[2791:2784]) ? 1 : 0;
assign detect_min[346][14] = (mid_1[2783:2776] < mid_2[2775:2768]) ? 1 : 0;
assign detect_min[346][15] = (mid_1[2783:2776] < mid_2[2783:2776]) ? 1 : 0;
assign detect_min[346][16] = (mid_1[2783:2776] < mid_2[2791:2784]) ? 1 : 0;
assign detect_min[346][17] = (mid_1[2783:2776] < btm_0[2775:2768]) ? 1 : 0;
assign detect_min[346][18] = (mid_1[2783:2776] < btm_0[2783:2776]) ? 1 : 0;
assign detect_min[346][19] = (mid_1[2783:2776] < btm_0[2791:2784]) ? 1 : 0;
assign detect_min[346][20] = (mid_1[2783:2776] < btm_1[2775:2768]) ? 1 : 0;
assign detect_min[346][21] = (mid_1[2783:2776] < btm_1[2783:2776]) ? 1 : 0;
assign detect_min[346][22] = (mid_1[2783:2776] < btm_1[2791:2784]) ? 1 : 0;
assign detect_min[346][23] = (mid_1[2783:2776] < btm_2[2775:2768]) ? 1 : 0;
assign detect_min[346][24] = (mid_1[2783:2776] < btm_2[2783:2776]) ? 1 : 0;
assign detect_min[346][25] = (mid_1[2783:2776] < btm_2[2791:2784]) ? 1 : 0;

assign detect_min[347][0] = (mid_1[2791:2784] < top_0[2783:2776]) ? 1 : 0;
assign detect_min[347][1] = (mid_1[2791:2784] < top_0[2791:2784]) ? 1 : 0;
assign detect_min[347][2] = (mid_1[2791:2784] < top_0[2799:2792]) ? 1 : 0;
assign detect_min[347][3] = (mid_1[2791:2784] < top_1[2783:2776]) ? 1 : 0;
assign detect_min[347][4] = (mid_1[2791:2784] < top_1[2791:2784]) ? 1 : 0;
assign detect_min[347][5] = (mid_1[2791:2784] < top_1[2799:2792]) ? 1 : 0;
assign detect_min[347][6] = (mid_1[2791:2784] < top_2[2783:2776]) ? 1 : 0;
assign detect_min[347][7] = (mid_1[2791:2784] < top_2[2791:2784]) ? 1 : 0;
assign detect_min[347][8] = (mid_1[2791:2784] < top_2[2799:2792]) ? 1 : 0;
assign detect_min[347][9] = (mid_1[2791:2784] < mid_0[2783:2776]) ? 1 : 0;
assign detect_min[347][10] = (mid_1[2791:2784] < mid_0[2791:2784]) ? 1 : 0;
assign detect_min[347][11] = (mid_1[2791:2784] < mid_0[2799:2792]) ? 1 : 0;
assign detect_min[347][12] = (mid_1[2791:2784] < mid_1[2783:2776]) ? 1 : 0;
assign detect_min[347][13] = (mid_1[2791:2784] < mid_1[2799:2792]) ? 1 : 0;
assign detect_min[347][14] = (mid_1[2791:2784] < mid_2[2783:2776]) ? 1 : 0;
assign detect_min[347][15] = (mid_1[2791:2784] < mid_2[2791:2784]) ? 1 : 0;
assign detect_min[347][16] = (mid_1[2791:2784] < mid_2[2799:2792]) ? 1 : 0;
assign detect_min[347][17] = (mid_1[2791:2784] < btm_0[2783:2776]) ? 1 : 0;
assign detect_min[347][18] = (mid_1[2791:2784] < btm_0[2791:2784]) ? 1 : 0;
assign detect_min[347][19] = (mid_1[2791:2784] < btm_0[2799:2792]) ? 1 : 0;
assign detect_min[347][20] = (mid_1[2791:2784] < btm_1[2783:2776]) ? 1 : 0;
assign detect_min[347][21] = (mid_1[2791:2784] < btm_1[2791:2784]) ? 1 : 0;
assign detect_min[347][22] = (mid_1[2791:2784] < btm_1[2799:2792]) ? 1 : 0;
assign detect_min[347][23] = (mid_1[2791:2784] < btm_2[2783:2776]) ? 1 : 0;
assign detect_min[347][24] = (mid_1[2791:2784] < btm_2[2791:2784]) ? 1 : 0;
assign detect_min[347][25] = (mid_1[2791:2784] < btm_2[2799:2792]) ? 1 : 0;

assign detect_min[348][0] = (mid_1[2799:2792] < top_0[2791:2784]) ? 1 : 0;
assign detect_min[348][1] = (mid_1[2799:2792] < top_0[2799:2792]) ? 1 : 0;
assign detect_min[348][2] = (mid_1[2799:2792] < top_0[2807:2800]) ? 1 : 0;
assign detect_min[348][3] = (mid_1[2799:2792] < top_1[2791:2784]) ? 1 : 0;
assign detect_min[348][4] = (mid_1[2799:2792] < top_1[2799:2792]) ? 1 : 0;
assign detect_min[348][5] = (mid_1[2799:2792] < top_1[2807:2800]) ? 1 : 0;
assign detect_min[348][6] = (mid_1[2799:2792] < top_2[2791:2784]) ? 1 : 0;
assign detect_min[348][7] = (mid_1[2799:2792] < top_2[2799:2792]) ? 1 : 0;
assign detect_min[348][8] = (mid_1[2799:2792] < top_2[2807:2800]) ? 1 : 0;
assign detect_min[348][9] = (mid_1[2799:2792] < mid_0[2791:2784]) ? 1 : 0;
assign detect_min[348][10] = (mid_1[2799:2792] < mid_0[2799:2792]) ? 1 : 0;
assign detect_min[348][11] = (mid_1[2799:2792] < mid_0[2807:2800]) ? 1 : 0;
assign detect_min[348][12] = (mid_1[2799:2792] < mid_1[2791:2784]) ? 1 : 0;
assign detect_min[348][13] = (mid_1[2799:2792] < mid_1[2807:2800]) ? 1 : 0;
assign detect_min[348][14] = (mid_1[2799:2792] < mid_2[2791:2784]) ? 1 : 0;
assign detect_min[348][15] = (mid_1[2799:2792] < mid_2[2799:2792]) ? 1 : 0;
assign detect_min[348][16] = (mid_1[2799:2792] < mid_2[2807:2800]) ? 1 : 0;
assign detect_min[348][17] = (mid_1[2799:2792] < btm_0[2791:2784]) ? 1 : 0;
assign detect_min[348][18] = (mid_1[2799:2792] < btm_0[2799:2792]) ? 1 : 0;
assign detect_min[348][19] = (mid_1[2799:2792] < btm_0[2807:2800]) ? 1 : 0;
assign detect_min[348][20] = (mid_1[2799:2792] < btm_1[2791:2784]) ? 1 : 0;
assign detect_min[348][21] = (mid_1[2799:2792] < btm_1[2799:2792]) ? 1 : 0;
assign detect_min[348][22] = (mid_1[2799:2792] < btm_1[2807:2800]) ? 1 : 0;
assign detect_min[348][23] = (mid_1[2799:2792] < btm_2[2791:2784]) ? 1 : 0;
assign detect_min[348][24] = (mid_1[2799:2792] < btm_2[2799:2792]) ? 1 : 0;
assign detect_min[348][25] = (mid_1[2799:2792] < btm_2[2807:2800]) ? 1 : 0;

assign detect_min[349][0] = (mid_1[2807:2800] < top_0[2799:2792]) ? 1 : 0;
assign detect_min[349][1] = (mid_1[2807:2800] < top_0[2807:2800]) ? 1 : 0;
assign detect_min[349][2] = (mid_1[2807:2800] < top_0[2815:2808]) ? 1 : 0;
assign detect_min[349][3] = (mid_1[2807:2800] < top_1[2799:2792]) ? 1 : 0;
assign detect_min[349][4] = (mid_1[2807:2800] < top_1[2807:2800]) ? 1 : 0;
assign detect_min[349][5] = (mid_1[2807:2800] < top_1[2815:2808]) ? 1 : 0;
assign detect_min[349][6] = (mid_1[2807:2800] < top_2[2799:2792]) ? 1 : 0;
assign detect_min[349][7] = (mid_1[2807:2800] < top_2[2807:2800]) ? 1 : 0;
assign detect_min[349][8] = (mid_1[2807:2800] < top_2[2815:2808]) ? 1 : 0;
assign detect_min[349][9] = (mid_1[2807:2800] < mid_0[2799:2792]) ? 1 : 0;
assign detect_min[349][10] = (mid_1[2807:2800] < mid_0[2807:2800]) ? 1 : 0;
assign detect_min[349][11] = (mid_1[2807:2800] < mid_0[2815:2808]) ? 1 : 0;
assign detect_min[349][12] = (mid_1[2807:2800] < mid_1[2799:2792]) ? 1 : 0;
assign detect_min[349][13] = (mid_1[2807:2800] < mid_1[2815:2808]) ? 1 : 0;
assign detect_min[349][14] = (mid_1[2807:2800] < mid_2[2799:2792]) ? 1 : 0;
assign detect_min[349][15] = (mid_1[2807:2800] < mid_2[2807:2800]) ? 1 : 0;
assign detect_min[349][16] = (mid_1[2807:2800] < mid_2[2815:2808]) ? 1 : 0;
assign detect_min[349][17] = (mid_1[2807:2800] < btm_0[2799:2792]) ? 1 : 0;
assign detect_min[349][18] = (mid_1[2807:2800] < btm_0[2807:2800]) ? 1 : 0;
assign detect_min[349][19] = (mid_1[2807:2800] < btm_0[2815:2808]) ? 1 : 0;
assign detect_min[349][20] = (mid_1[2807:2800] < btm_1[2799:2792]) ? 1 : 0;
assign detect_min[349][21] = (mid_1[2807:2800] < btm_1[2807:2800]) ? 1 : 0;
assign detect_min[349][22] = (mid_1[2807:2800] < btm_1[2815:2808]) ? 1 : 0;
assign detect_min[349][23] = (mid_1[2807:2800] < btm_2[2799:2792]) ? 1 : 0;
assign detect_min[349][24] = (mid_1[2807:2800] < btm_2[2807:2800]) ? 1 : 0;
assign detect_min[349][25] = (mid_1[2807:2800] < btm_2[2815:2808]) ? 1 : 0;

assign detect_min[350][0] = (mid_1[2815:2808] < top_0[2807:2800]) ? 1 : 0;
assign detect_min[350][1] = (mid_1[2815:2808] < top_0[2815:2808]) ? 1 : 0;
assign detect_min[350][2] = (mid_1[2815:2808] < top_0[2823:2816]) ? 1 : 0;
assign detect_min[350][3] = (mid_1[2815:2808] < top_1[2807:2800]) ? 1 : 0;
assign detect_min[350][4] = (mid_1[2815:2808] < top_1[2815:2808]) ? 1 : 0;
assign detect_min[350][5] = (mid_1[2815:2808] < top_1[2823:2816]) ? 1 : 0;
assign detect_min[350][6] = (mid_1[2815:2808] < top_2[2807:2800]) ? 1 : 0;
assign detect_min[350][7] = (mid_1[2815:2808] < top_2[2815:2808]) ? 1 : 0;
assign detect_min[350][8] = (mid_1[2815:2808] < top_2[2823:2816]) ? 1 : 0;
assign detect_min[350][9] = (mid_1[2815:2808] < mid_0[2807:2800]) ? 1 : 0;
assign detect_min[350][10] = (mid_1[2815:2808] < mid_0[2815:2808]) ? 1 : 0;
assign detect_min[350][11] = (mid_1[2815:2808] < mid_0[2823:2816]) ? 1 : 0;
assign detect_min[350][12] = (mid_1[2815:2808] < mid_1[2807:2800]) ? 1 : 0;
assign detect_min[350][13] = (mid_1[2815:2808] < mid_1[2823:2816]) ? 1 : 0;
assign detect_min[350][14] = (mid_1[2815:2808] < mid_2[2807:2800]) ? 1 : 0;
assign detect_min[350][15] = (mid_1[2815:2808] < mid_2[2815:2808]) ? 1 : 0;
assign detect_min[350][16] = (mid_1[2815:2808] < mid_2[2823:2816]) ? 1 : 0;
assign detect_min[350][17] = (mid_1[2815:2808] < btm_0[2807:2800]) ? 1 : 0;
assign detect_min[350][18] = (mid_1[2815:2808] < btm_0[2815:2808]) ? 1 : 0;
assign detect_min[350][19] = (mid_1[2815:2808] < btm_0[2823:2816]) ? 1 : 0;
assign detect_min[350][20] = (mid_1[2815:2808] < btm_1[2807:2800]) ? 1 : 0;
assign detect_min[350][21] = (mid_1[2815:2808] < btm_1[2815:2808]) ? 1 : 0;
assign detect_min[350][22] = (mid_1[2815:2808] < btm_1[2823:2816]) ? 1 : 0;
assign detect_min[350][23] = (mid_1[2815:2808] < btm_2[2807:2800]) ? 1 : 0;
assign detect_min[350][24] = (mid_1[2815:2808] < btm_2[2815:2808]) ? 1 : 0;
assign detect_min[350][25] = (mid_1[2815:2808] < btm_2[2823:2816]) ? 1 : 0;

assign detect_min[351][0] = (mid_1[2823:2816] < top_0[2815:2808]) ? 1 : 0;
assign detect_min[351][1] = (mid_1[2823:2816] < top_0[2823:2816]) ? 1 : 0;
assign detect_min[351][2] = (mid_1[2823:2816] < top_0[2831:2824]) ? 1 : 0;
assign detect_min[351][3] = (mid_1[2823:2816] < top_1[2815:2808]) ? 1 : 0;
assign detect_min[351][4] = (mid_1[2823:2816] < top_1[2823:2816]) ? 1 : 0;
assign detect_min[351][5] = (mid_1[2823:2816] < top_1[2831:2824]) ? 1 : 0;
assign detect_min[351][6] = (mid_1[2823:2816] < top_2[2815:2808]) ? 1 : 0;
assign detect_min[351][7] = (mid_1[2823:2816] < top_2[2823:2816]) ? 1 : 0;
assign detect_min[351][8] = (mid_1[2823:2816] < top_2[2831:2824]) ? 1 : 0;
assign detect_min[351][9] = (mid_1[2823:2816] < mid_0[2815:2808]) ? 1 : 0;
assign detect_min[351][10] = (mid_1[2823:2816] < mid_0[2823:2816]) ? 1 : 0;
assign detect_min[351][11] = (mid_1[2823:2816] < mid_0[2831:2824]) ? 1 : 0;
assign detect_min[351][12] = (mid_1[2823:2816] < mid_1[2815:2808]) ? 1 : 0;
assign detect_min[351][13] = (mid_1[2823:2816] < mid_1[2831:2824]) ? 1 : 0;
assign detect_min[351][14] = (mid_1[2823:2816] < mid_2[2815:2808]) ? 1 : 0;
assign detect_min[351][15] = (mid_1[2823:2816] < mid_2[2823:2816]) ? 1 : 0;
assign detect_min[351][16] = (mid_1[2823:2816] < mid_2[2831:2824]) ? 1 : 0;
assign detect_min[351][17] = (mid_1[2823:2816] < btm_0[2815:2808]) ? 1 : 0;
assign detect_min[351][18] = (mid_1[2823:2816] < btm_0[2823:2816]) ? 1 : 0;
assign detect_min[351][19] = (mid_1[2823:2816] < btm_0[2831:2824]) ? 1 : 0;
assign detect_min[351][20] = (mid_1[2823:2816] < btm_1[2815:2808]) ? 1 : 0;
assign detect_min[351][21] = (mid_1[2823:2816] < btm_1[2823:2816]) ? 1 : 0;
assign detect_min[351][22] = (mid_1[2823:2816] < btm_1[2831:2824]) ? 1 : 0;
assign detect_min[351][23] = (mid_1[2823:2816] < btm_2[2815:2808]) ? 1 : 0;
assign detect_min[351][24] = (mid_1[2823:2816] < btm_2[2823:2816]) ? 1 : 0;
assign detect_min[351][25] = (mid_1[2823:2816] < btm_2[2831:2824]) ? 1 : 0;

assign detect_min[352][0] = (mid_1[2831:2824] < top_0[2823:2816]) ? 1 : 0;
assign detect_min[352][1] = (mid_1[2831:2824] < top_0[2831:2824]) ? 1 : 0;
assign detect_min[352][2] = (mid_1[2831:2824] < top_0[2839:2832]) ? 1 : 0;
assign detect_min[352][3] = (mid_1[2831:2824] < top_1[2823:2816]) ? 1 : 0;
assign detect_min[352][4] = (mid_1[2831:2824] < top_1[2831:2824]) ? 1 : 0;
assign detect_min[352][5] = (mid_1[2831:2824] < top_1[2839:2832]) ? 1 : 0;
assign detect_min[352][6] = (mid_1[2831:2824] < top_2[2823:2816]) ? 1 : 0;
assign detect_min[352][7] = (mid_1[2831:2824] < top_2[2831:2824]) ? 1 : 0;
assign detect_min[352][8] = (mid_1[2831:2824] < top_2[2839:2832]) ? 1 : 0;
assign detect_min[352][9] = (mid_1[2831:2824] < mid_0[2823:2816]) ? 1 : 0;
assign detect_min[352][10] = (mid_1[2831:2824] < mid_0[2831:2824]) ? 1 : 0;
assign detect_min[352][11] = (mid_1[2831:2824] < mid_0[2839:2832]) ? 1 : 0;
assign detect_min[352][12] = (mid_1[2831:2824] < mid_1[2823:2816]) ? 1 : 0;
assign detect_min[352][13] = (mid_1[2831:2824] < mid_1[2839:2832]) ? 1 : 0;
assign detect_min[352][14] = (mid_1[2831:2824] < mid_2[2823:2816]) ? 1 : 0;
assign detect_min[352][15] = (mid_1[2831:2824] < mid_2[2831:2824]) ? 1 : 0;
assign detect_min[352][16] = (mid_1[2831:2824] < mid_2[2839:2832]) ? 1 : 0;
assign detect_min[352][17] = (mid_1[2831:2824] < btm_0[2823:2816]) ? 1 : 0;
assign detect_min[352][18] = (mid_1[2831:2824] < btm_0[2831:2824]) ? 1 : 0;
assign detect_min[352][19] = (mid_1[2831:2824] < btm_0[2839:2832]) ? 1 : 0;
assign detect_min[352][20] = (mid_1[2831:2824] < btm_1[2823:2816]) ? 1 : 0;
assign detect_min[352][21] = (mid_1[2831:2824] < btm_1[2831:2824]) ? 1 : 0;
assign detect_min[352][22] = (mid_1[2831:2824] < btm_1[2839:2832]) ? 1 : 0;
assign detect_min[352][23] = (mid_1[2831:2824] < btm_2[2823:2816]) ? 1 : 0;
assign detect_min[352][24] = (mid_1[2831:2824] < btm_2[2831:2824]) ? 1 : 0;
assign detect_min[352][25] = (mid_1[2831:2824] < btm_2[2839:2832]) ? 1 : 0;

assign detect_min[353][0] = (mid_1[2839:2832] < top_0[2831:2824]) ? 1 : 0;
assign detect_min[353][1] = (mid_1[2839:2832] < top_0[2839:2832]) ? 1 : 0;
assign detect_min[353][2] = (mid_1[2839:2832] < top_0[2847:2840]) ? 1 : 0;
assign detect_min[353][3] = (mid_1[2839:2832] < top_1[2831:2824]) ? 1 : 0;
assign detect_min[353][4] = (mid_1[2839:2832] < top_1[2839:2832]) ? 1 : 0;
assign detect_min[353][5] = (mid_1[2839:2832] < top_1[2847:2840]) ? 1 : 0;
assign detect_min[353][6] = (mid_1[2839:2832] < top_2[2831:2824]) ? 1 : 0;
assign detect_min[353][7] = (mid_1[2839:2832] < top_2[2839:2832]) ? 1 : 0;
assign detect_min[353][8] = (mid_1[2839:2832] < top_2[2847:2840]) ? 1 : 0;
assign detect_min[353][9] = (mid_1[2839:2832] < mid_0[2831:2824]) ? 1 : 0;
assign detect_min[353][10] = (mid_1[2839:2832] < mid_0[2839:2832]) ? 1 : 0;
assign detect_min[353][11] = (mid_1[2839:2832] < mid_0[2847:2840]) ? 1 : 0;
assign detect_min[353][12] = (mid_1[2839:2832] < mid_1[2831:2824]) ? 1 : 0;
assign detect_min[353][13] = (mid_1[2839:2832] < mid_1[2847:2840]) ? 1 : 0;
assign detect_min[353][14] = (mid_1[2839:2832] < mid_2[2831:2824]) ? 1 : 0;
assign detect_min[353][15] = (mid_1[2839:2832] < mid_2[2839:2832]) ? 1 : 0;
assign detect_min[353][16] = (mid_1[2839:2832] < mid_2[2847:2840]) ? 1 : 0;
assign detect_min[353][17] = (mid_1[2839:2832] < btm_0[2831:2824]) ? 1 : 0;
assign detect_min[353][18] = (mid_1[2839:2832] < btm_0[2839:2832]) ? 1 : 0;
assign detect_min[353][19] = (mid_1[2839:2832] < btm_0[2847:2840]) ? 1 : 0;
assign detect_min[353][20] = (mid_1[2839:2832] < btm_1[2831:2824]) ? 1 : 0;
assign detect_min[353][21] = (mid_1[2839:2832] < btm_1[2839:2832]) ? 1 : 0;
assign detect_min[353][22] = (mid_1[2839:2832] < btm_1[2847:2840]) ? 1 : 0;
assign detect_min[353][23] = (mid_1[2839:2832] < btm_2[2831:2824]) ? 1 : 0;
assign detect_min[353][24] = (mid_1[2839:2832] < btm_2[2839:2832]) ? 1 : 0;
assign detect_min[353][25] = (mid_1[2839:2832] < btm_2[2847:2840]) ? 1 : 0;

assign detect_min[354][0] = (mid_1[2847:2840] < top_0[2839:2832]) ? 1 : 0;
assign detect_min[354][1] = (mid_1[2847:2840] < top_0[2847:2840]) ? 1 : 0;
assign detect_min[354][2] = (mid_1[2847:2840] < top_0[2855:2848]) ? 1 : 0;
assign detect_min[354][3] = (mid_1[2847:2840] < top_1[2839:2832]) ? 1 : 0;
assign detect_min[354][4] = (mid_1[2847:2840] < top_1[2847:2840]) ? 1 : 0;
assign detect_min[354][5] = (mid_1[2847:2840] < top_1[2855:2848]) ? 1 : 0;
assign detect_min[354][6] = (mid_1[2847:2840] < top_2[2839:2832]) ? 1 : 0;
assign detect_min[354][7] = (mid_1[2847:2840] < top_2[2847:2840]) ? 1 : 0;
assign detect_min[354][8] = (mid_1[2847:2840] < top_2[2855:2848]) ? 1 : 0;
assign detect_min[354][9] = (mid_1[2847:2840] < mid_0[2839:2832]) ? 1 : 0;
assign detect_min[354][10] = (mid_1[2847:2840] < mid_0[2847:2840]) ? 1 : 0;
assign detect_min[354][11] = (mid_1[2847:2840] < mid_0[2855:2848]) ? 1 : 0;
assign detect_min[354][12] = (mid_1[2847:2840] < mid_1[2839:2832]) ? 1 : 0;
assign detect_min[354][13] = (mid_1[2847:2840] < mid_1[2855:2848]) ? 1 : 0;
assign detect_min[354][14] = (mid_1[2847:2840] < mid_2[2839:2832]) ? 1 : 0;
assign detect_min[354][15] = (mid_1[2847:2840] < mid_2[2847:2840]) ? 1 : 0;
assign detect_min[354][16] = (mid_1[2847:2840] < mid_2[2855:2848]) ? 1 : 0;
assign detect_min[354][17] = (mid_1[2847:2840] < btm_0[2839:2832]) ? 1 : 0;
assign detect_min[354][18] = (mid_1[2847:2840] < btm_0[2847:2840]) ? 1 : 0;
assign detect_min[354][19] = (mid_1[2847:2840] < btm_0[2855:2848]) ? 1 : 0;
assign detect_min[354][20] = (mid_1[2847:2840] < btm_1[2839:2832]) ? 1 : 0;
assign detect_min[354][21] = (mid_1[2847:2840] < btm_1[2847:2840]) ? 1 : 0;
assign detect_min[354][22] = (mid_1[2847:2840] < btm_1[2855:2848]) ? 1 : 0;
assign detect_min[354][23] = (mid_1[2847:2840] < btm_2[2839:2832]) ? 1 : 0;
assign detect_min[354][24] = (mid_1[2847:2840] < btm_2[2847:2840]) ? 1 : 0;
assign detect_min[354][25] = (mid_1[2847:2840] < btm_2[2855:2848]) ? 1 : 0;

assign detect_min[355][0] = (mid_1[2855:2848] < top_0[2847:2840]) ? 1 : 0;
assign detect_min[355][1] = (mid_1[2855:2848] < top_0[2855:2848]) ? 1 : 0;
assign detect_min[355][2] = (mid_1[2855:2848] < top_0[2863:2856]) ? 1 : 0;
assign detect_min[355][3] = (mid_1[2855:2848] < top_1[2847:2840]) ? 1 : 0;
assign detect_min[355][4] = (mid_1[2855:2848] < top_1[2855:2848]) ? 1 : 0;
assign detect_min[355][5] = (mid_1[2855:2848] < top_1[2863:2856]) ? 1 : 0;
assign detect_min[355][6] = (mid_1[2855:2848] < top_2[2847:2840]) ? 1 : 0;
assign detect_min[355][7] = (mid_1[2855:2848] < top_2[2855:2848]) ? 1 : 0;
assign detect_min[355][8] = (mid_1[2855:2848] < top_2[2863:2856]) ? 1 : 0;
assign detect_min[355][9] = (mid_1[2855:2848] < mid_0[2847:2840]) ? 1 : 0;
assign detect_min[355][10] = (mid_1[2855:2848] < mid_0[2855:2848]) ? 1 : 0;
assign detect_min[355][11] = (mid_1[2855:2848] < mid_0[2863:2856]) ? 1 : 0;
assign detect_min[355][12] = (mid_1[2855:2848] < mid_1[2847:2840]) ? 1 : 0;
assign detect_min[355][13] = (mid_1[2855:2848] < mid_1[2863:2856]) ? 1 : 0;
assign detect_min[355][14] = (mid_1[2855:2848] < mid_2[2847:2840]) ? 1 : 0;
assign detect_min[355][15] = (mid_1[2855:2848] < mid_2[2855:2848]) ? 1 : 0;
assign detect_min[355][16] = (mid_1[2855:2848] < mid_2[2863:2856]) ? 1 : 0;
assign detect_min[355][17] = (mid_1[2855:2848] < btm_0[2847:2840]) ? 1 : 0;
assign detect_min[355][18] = (mid_1[2855:2848] < btm_0[2855:2848]) ? 1 : 0;
assign detect_min[355][19] = (mid_1[2855:2848] < btm_0[2863:2856]) ? 1 : 0;
assign detect_min[355][20] = (mid_1[2855:2848] < btm_1[2847:2840]) ? 1 : 0;
assign detect_min[355][21] = (mid_1[2855:2848] < btm_1[2855:2848]) ? 1 : 0;
assign detect_min[355][22] = (mid_1[2855:2848] < btm_1[2863:2856]) ? 1 : 0;
assign detect_min[355][23] = (mid_1[2855:2848] < btm_2[2847:2840]) ? 1 : 0;
assign detect_min[355][24] = (mid_1[2855:2848] < btm_2[2855:2848]) ? 1 : 0;
assign detect_min[355][25] = (mid_1[2855:2848] < btm_2[2863:2856]) ? 1 : 0;

assign detect_min[356][0] = (mid_1[2863:2856] < top_0[2855:2848]) ? 1 : 0;
assign detect_min[356][1] = (mid_1[2863:2856] < top_0[2863:2856]) ? 1 : 0;
assign detect_min[356][2] = (mid_1[2863:2856] < top_0[2871:2864]) ? 1 : 0;
assign detect_min[356][3] = (mid_1[2863:2856] < top_1[2855:2848]) ? 1 : 0;
assign detect_min[356][4] = (mid_1[2863:2856] < top_1[2863:2856]) ? 1 : 0;
assign detect_min[356][5] = (mid_1[2863:2856] < top_1[2871:2864]) ? 1 : 0;
assign detect_min[356][6] = (mid_1[2863:2856] < top_2[2855:2848]) ? 1 : 0;
assign detect_min[356][7] = (mid_1[2863:2856] < top_2[2863:2856]) ? 1 : 0;
assign detect_min[356][8] = (mid_1[2863:2856] < top_2[2871:2864]) ? 1 : 0;
assign detect_min[356][9] = (mid_1[2863:2856] < mid_0[2855:2848]) ? 1 : 0;
assign detect_min[356][10] = (mid_1[2863:2856] < mid_0[2863:2856]) ? 1 : 0;
assign detect_min[356][11] = (mid_1[2863:2856] < mid_0[2871:2864]) ? 1 : 0;
assign detect_min[356][12] = (mid_1[2863:2856] < mid_1[2855:2848]) ? 1 : 0;
assign detect_min[356][13] = (mid_1[2863:2856] < mid_1[2871:2864]) ? 1 : 0;
assign detect_min[356][14] = (mid_1[2863:2856] < mid_2[2855:2848]) ? 1 : 0;
assign detect_min[356][15] = (mid_1[2863:2856] < mid_2[2863:2856]) ? 1 : 0;
assign detect_min[356][16] = (mid_1[2863:2856] < mid_2[2871:2864]) ? 1 : 0;
assign detect_min[356][17] = (mid_1[2863:2856] < btm_0[2855:2848]) ? 1 : 0;
assign detect_min[356][18] = (mid_1[2863:2856] < btm_0[2863:2856]) ? 1 : 0;
assign detect_min[356][19] = (mid_1[2863:2856] < btm_0[2871:2864]) ? 1 : 0;
assign detect_min[356][20] = (mid_1[2863:2856] < btm_1[2855:2848]) ? 1 : 0;
assign detect_min[356][21] = (mid_1[2863:2856] < btm_1[2863:2856]) ? 1 : 0;
assign detect_min[356][22] = (mid_1[2863:2856] < btm_1[2871:2864]) ? 1 : 0;
assign detect_min[356][23] = (mid_1[2863:2856] < btm_2[2855:2848]) ? 1 : 0;
assign detect_min[356][24] = (mid_1[2863:2856] < btm_2[2863:2856]) ? 1 : 0;
assign detect_min[356][25] = (mid_1[2863:2856] < btm_2[2871:2864]) ? 1 : 0;

assign detect_min[357][0] = (mid_1[2871:2864] < top_0[2863:2856]) ? 1 : 0;
assign detect_min[357][1] = (mid_1[2871:2864] < top_0[2871:2864]) ? 1 : 0;
assign detect_min[357][2] = (mid_1[2871:2864] < top_0[2879:2872]) ? 1 : 0;
assign detect_min[357][3] = (mid_1[2871:2864] < top_1[2863:2856]) ? 1 : 0;
assign detect_min[357][4] = (mid_1[2871:2864] < top_1[2871:2864]) ? 1 : 0;
assign detect_min[357][5] = (mid_1[2871:2864] < top_1[2879:2872]) ? 1 : 0;
assign detect_min[357][6] = (mid_1[2871:2864] < top_2[2863:2856]) ? 1 : 0;
assign detect_min[357][7] = (mid_1[2871:2864] < top_2[2871:2864]) ? 1 : 0;
assign detect_min[357][8] = (mid_1[2871:2864] < top_2[2879:2872]) ? 1 : 0;
assign detect_min[357][9] = (mid_1[2871:2864] < mid_0[2863:2856]) ? 1 : 0;
assign detect_min[357][10] = (mid_1[2871:2864] < mid_0[2871:2864]) ? 1 : 0;
assign detect_min[357][11] = (mid_1[2871:2864] < mid_0[2879:2872]) ? 1 : 0;
assign detect_min[357][12] = (mid_1[2871:2864] < mid_1[2863:2856]) ? 1 : 0;
assign detect_min[357][13] = (mid_1[2871:2864] < mid_1[2879:2872]) ? 1 : 0;
assign detect_min[357][14] = (mid_1[2871:2864] < mid_2[2863:2856]) ? 1 : 0;
assign detect_min[357][15] = (mid_1[2871:2864] < mid_2[2871:2864]) ? 1 : 0;
assign detect_min[357][16] = (mid_1[2871:2864] < mid_2[2879:2872]) ? 1 : 0;
assign detect_min[357][17] = (mid_1[2871:2864] < btm_0[2863:2856]) ? 1 : 0;
assign detect_min[357][18] = (mid_1[2871:2864] < btm_0[2871:2864]) ? 1 : 0;
assign detect_min[357][19] = (mid_1[2871:2864] < btm_0[2879:2872]) ? 1 : 0;
assign detect_min[357][20] = (mid_1[2871:2864] < btm_1[2863:2856]) ? 1 : 0;
assign detect_min[357][21] = (mid_1[2871:2864] < btm_1[2871:2864]) ? 1 : 0;
assign detect_min[357][22] = (mid_1[2871:2864] < btm_1[2879:2872]) ? 1 : 0;
assign detect_min[357][23] = (mid_1[2871:2864] < btm_2[2863:2856]) ? 1 : 0;
assign detect_min[357][24] = (mid_1[2871:2864] < btm_2[2871:2864]) ? 1 : 0;
assign detect_min[357][25] = (mid_1[2871:2864] < btm_2[2879:2872]) ? 1 : 0;

assign detect_min[358][0] = (mid_1[2879:2872] < top_0[2871:2864]) ? 1 : 0;
assign detect_min[358][1] = (mid_1[2879:2872] < top_0[2879:2872]) ? 1 : 0;
assign detect_min[358][2] = (mid_1[2879:2872] < top_0[2887:2880]) ? 1 : 0;
assign detect_min[358][3] = (mid_1[2879:2872] < top_1[2871:2864]) ? 1 : 0;
assign detect_min[358][4] = (mid_1[2879:2872] < top_1[2879:2872]) ? 1 : 0;
assign detect_min[358][5] = (mid_1[2879:2872] < top_1[2887:2880]) ? 1 : 0;
assign detect_min[358][6] = (mid_1[2879:2872] < top_2[2871:2864]) ? 1 : 0;
assign detect_min[358][7] = (mid_1[2879:2872] < top_2[2879:2872]) ? 1 : 0;
assign detect_min[358][8] = (mid_1[2879:2872] < top_2[2887:2880]) ? 1 : 0;
assign detect_min[358][9] = (mid_1[2879:2872] < mid_0[2871:2864]) ? 1 : 0;
assign detect_min[358][10] = (mid_1[2879:2872] < mid_0[2879:2872]) ? 1 : 0;
assign detect_min[358][11] = (mid_1[2879:2872] < mid_0[2887:2880]) ? 1 : 0;
assign detect_min[358][12] = (mid_1[2879:2872] < mid_1[2871:2864]) ? 1 : 0;
assign detect_min[358][13] = (mid_1[2879:2872] < mid_1[2887:2880]) ? 1 : 0;
assign detect_min[358][14] = (mid_1[2879:2872] < mid_2[2871:2864]) ? 1 : 0;
assign detect_min[358][15] = (mid_1[2879:2872] < mid_2[2879:2872]) ? 1 : 0;
assign detect_min[358][16] = (mid_1[2879:2872] < mid_2[2887:2880]) ? 1 : 0;
assign detect_min[358][17] = (mid_1[2879:2872] < btm_0[2871:2864]) ? 1 : 0;
assign detect_min[358][18] = (mid_1[2879:2872] < btm_0[2879:2872]) ? 1 : 0;
assign detect_min[358][19] = (mid_1[2879:2872] < btm_0[2887:2880]) ? 1 : 0;
assign detect_min[358][20] = (mid_1[2879:2872] < btm_1[2871:2864]) ? 1 : 0;
assign detect_min[358][21] = (mid_1[2879:2872] < btm_1[2879:2872]) ? 1 : 0;
assign detect_min[358][22] = (mid_1[2879:2872] < btm_1[2887:2880]) ? 1 : 0;
assign detect_min[358][23] = (mid_1[2879:2872] < btm_2[2871:2864]) ? 1 : 0;
assign detect_min[358][24] = (mid_1[2879:2872] < btm_2[2879:2872]) ? 1 : 0;
assign detect_min[358][25] = (mid_1[2879:2872] < btm_2[2887:2880]) ? 1 : 0;

assign detect_min[359][0] = (mid_1[2887:2880] < top_0[2879:2872]) ? 1 : 0;
assign detect_min[359][1] = (mid_1[2887:2880] < top_0[2887:2880]) ? 1 : 0;
assign detect_min[359][2] = (mid_1[2887:2880] < top_0[2895:2888]) ? 1 : 0;
assign detect_min[359][3] = (mid_1[2887:2880] < top_1[2879:2872]) ? 1 : 0;
assign detect_min[359][4] = (mid_1[2887:2880] < top_1[2887:2880]) ? 1 : 0;
assign detect_min[359][5] = (mid_1[2887:2880] < top_1[2895:2888]) ? 1 : 0;
assign detect_min[359][6] = (mid_1[2887:2880] < top_2[2879:2872]) ? 1 : 0;
assign detect_min[359][7] = (mid_1[2887:2880] < top_2[2887:2880]) ? 1 : 0;
assign detect_min[359][8] = (mid_1[2887:2880] < top_2[2895:2888]) ? 1 : 0;
assign detect_min[359][9] = (mid_1[2887:2880] < mid_0[2879:2872]) ? 1 : 0;
assign detect_min[359][10] = (mid_1[2887:2880] < mid_0[2887:2880]) ? 1 : 0;
assign detect_min[359][11] = (mid_1[2887:2880] < mid_0[2895:2888]) ? 1 : 0;
assign detect_min[359][12] = (mid_1[2887:2880] < mid_1[2879:2872]) ? 1 : 0;
assign detect_min[359][13] = (mid_1[2887:2880] < mid_1[2895:2888]) ? 1 : 0;
assign detect_min[359][14] = (mid_1[2887:2880] < mid_2[2879:2872]) ? 1 : 0;
assign detect_min[359][15] = (mid_1[2887:2880] < mid_2[2887:2880]) ? 1 : 0;
assign detect_min[359][16] = (mid_1[2887:2880] < mid_2[2895:2888]) ? 1 : 0;
assign detect_min[359][17] = (mid_1[2887:2880] < btm_0[2879:2872]) ? 1 : 0;
assign detect_min[359][18] = (mid_1[2887:2880] < btm_0[2887:2880]) ? 1 : 0;
assign detect_min[359][19] = (mid_1[2887:2880] < btm_0[2895:2888]) ? 1 : 0;
assign detect_min[359][20] = (mid_1[2887:2880] < btm_1[2879:2872]) ? 1 : 0;
assign detect_min[359][21] = (mid_1[2887:2880] < btm_1[2887:2880]) ? 1 : 0;
assign detect_min[359][22] = (mid_1[2887:2880] < btm_1[2895:2888]) ? 1 : 0;
assign detect_min[359][23] = (mid_1[2887:2880] < btm_2[2879:2872]) ? 1 : 0;
assign detect_min[359][24] = (mid_1[2887:2880] < btm_2[2887:2880]) ? 1 : 0;
assign detect_min[359][25] = (mid_1[2887:2880] < btm_2[2895:2888]) ? 1 : 0;

assign detect_min[360][0] = (mid_1[2895:2888] < top_0[2887:2880]) ? 1 : 0;
assign detect_min[360][1] = (mid_1[2895:2888] < top_0[2895:2888]) ? 1 : 0;
assign detect_min[360][2] = (mid_1[2895:2888] < top_0[2903:2896]) ? 1 : 0;
assign detect_min[360][3] = (mid_1[2895:2888] < top_1[2887:2880]) ? 1 : 0;
assign detect_min[360][4] = (mid_1[2895:2888] < top_1[2895:2888]) ? 1 : 0;
assign detect_min[360][5] = (mid_1[2895:2888] < top_1[2903:2896]) ? 1 : 0;
assign detect_min[360][6] = (mid_1[2895:2888] < top_2[2887:2880]) ? 1 : 0;
assign detect_min[360][7] = (mid_1[2895:2888] < top_2[2895:2888]) ? 1 : 0;
assign detect_min[360][8] = (mid_1[2895:2888] < top_2[2903:2896]) ? 1 : 0;
assign detect_min[360][9] = (mid_1[2895:2888] < mid_0[2887:2880]) ? 1 : 0;
assign detect_min[360][10] = (mid_1[2895:2888] < mid_0[2895:2888]) ? 1 : 0;
assign detect_min[360][11] = (mid_1[2895:2888] < mid_0[2903:2896]) ? 1 : 0;
assign detect_min[360][12] = (mid_1[2895:2888] < mid_1[2887:2880]) ? 1 : 0;
assign detect_min[360][13] = (mid_1[2895:2888] < mid_1[2903:2896]) ? 1 : 0;
assign detect_min[360][14] = (mid_1[2895:2888] < mid_2[2887:2880]) ? 1 : 0;
assign detect_min[360][15] = (mid_1[2895:2888] < mid_2[2895:2888]) ? 1 : 0;
assign detect_min[360][16] = (mid_1[2895:2888] < mid_2[2903:2896]) ? 1 : 0;
assign detect_min[360][17] = (mid_1[2895:2888] < btm_0[2887:2880]) ? 1 : 0;
assign detect_min[360][18] = (mid_1[2895:2888] < btm_0[2895:2888]) ? 1 : 0;
assign detect_min[360][19] = (mid_1[2895:2888] < btm_0[2903:2896]) ? 1 : 0;
assign detect_min[360][20] = (mid_1[2895:2888] < btm_1[2887:2880]) ? 1 : 0;
assign detect_min[360][21] = (mid_1[2895:2888] < btm_1[2895:2888]) ? 1 : 0;
assign detect_min[360][22] = (mid_1[2895:2888] < btm_1[2903:2896]) ? 1 : 0;
assign detect_min[360][23] = (mid_1[2895:2888] < btm_2[2887:2880]) ? 1 : 0;
assign detect_min[360][24] = (mid_1[2895:2888] < btm_2[2895:2888]) ? 1 : 0;
assign detect_min[360][25] = (mid_1[2895:2888] < btm_2[2903:2896]) ? 1 : 0;

assign detect_min[361][0] = (mid_1[2903:2896] < top_0[2895:2888]) ? 1 : 0;
assign detect_min[361][1] = (mid_1[2903:2896] < top_0[2903:2896]) ? 1 : 0;
assign detect_min[361][2] = (mid_1[2903:2896] < top_0[2911:2904]) ? 1 : 0;
assign detect_min[361][3] = (mid_1[2903:2896] < top_1[2895:2888]) ? 1 : 0;
assign detect_min[361][4] = (mid_1[2903:2896] < top_1[2903:2896]) ? 1 : 0;
assign detect_min[361][5] = (mid_1[2903:2896] < top_1[2911:2904]) ? 1 : 0;
assign detect_min[361][6] = (mid_1[2903:2896] < top_2[2895:2888]) ? 1 : 0;
assign detect_min[361][7] = (mid_1[2903:2896] < top_2[2903:2896]) ? 1 : 0;
assign detect_min[361][8] = (mid_1[2903:2896] < top_2[2911:2904]) ? 1 : 0;
assign detect_min[361][9] = (mid_1[2903:2896] < mid_0[2895:2888]) ? 1 : 0;
assign detect_min[361][10] = (mid_1[2903:2896] < mid_0[2903:2896]) ? 1 : 0;
assign detect_min[361][11] = (mid_1[2903:2896] < mid_0[2911:2904]) ? 1 : 0;
assign detect_min[361][12] = (mid_1[2903:2896] < mid_1[2895:2888]) ? 1 : 0;
assign detect_min[361][13] = (mid_1[2903:2896] < mid_1[2911:2904]) ? 1 : 0;
assign detect_min[361][14] = (mid_1[2903:2896] < mid_2[2895:2888]) ? 1 : 0;
assign detect_min[361][15] = (mid_1[2903:2896] < mid_2[2903:2896]) ? 1 : 0;
assign detect_min[361][16] = (mid_1[2903:2896] < mid_2[2911:2904]) ? 1 : 0;
assign detect_min[361][17] = (mid_1[2903:2896] < btm_0[2895:2888]) ? 1 : 0;
assign detect_min[361][18] = (mid_1[2903:2896] < btm_0[2903:2896]) ? 1 : 0;
assign detect_min[361][19] = (mid_1[2903:2896] < btm_0[2911:2904]) ? 1 : 0;
assign detect_min[361][20] = (mid_1[2903:2896] < btm_1[2895:2888]) ? 1 : 0;
assign detect_min[361][21] = (mid_1[2903:2896] < btm_1[2903:2896]) ? 1 : 0;
assign detect_min[361][22] = (mid_1[2903:2896] < btm_1[2911:2904]) ? 1 : 0;
assign detect_min[361][23] = (mid_1[2903:2896] < btm_2[2895:2888]) ? 1 : 0;
assign detect_min[361][24] = (mid_1[2903:2896] < btm_2[2903:2896]) ? 1 : 0;
assign detect_min[361][25] = (mid_1[2903:2896] < btm_2[2911:2904]) ? 1 : 0;

assign detect_min[362][0] = (mid_1[2911:2904] < top_0[2903:2896]) ? 1 : 0;
assign detect_min[362][1] = (mid_1[2911:2904] < top_0[2911:2904]) ? 1 : 0;
assign detect_min[362][2] = (mid_1[2911:2904] < top_0[2919:2912]) ? 1 : 0;
assign detect_min[362][3] = (mid_1[2911:2904] < top_1[2903:2896]) ? 1 : 0;
assign detect_min[362][4] = (mid_1[2911:2904] < top_1[2911:2904]) ? 1 : 0;
assign detect_min[362][5] = (mid_1[2911:2904] < top_1[2919:2912]) ? 1 : 0;
assign detect_min[362][6] = (mid_1[2911:2904] < top_2[2903:2896]) ? 1 : 0;
assign detect_min[362][7] = (mid_1[2911:2904] < top_2[2911:2904]) ? 1 : 0;
assign detect_min[362][8] = (mid_1[2911:2904] < top_2[2919:2912]) ? 1 : 0;
assign detect_min[362][9] = (mid_1[2911:2904] < mid_0[2903:2896]) ? 1 : 0;
assign detect_min[362][10] = (mid_1[2911:2904] < mid_0[2911:2904]) ? 1 : 0;
assign detect_min[362][11] = (mid_1[2911:2904] < mid_0[2919:2912]) ? 1 : 0;
assign detect_min[362][12] = (mid_1[2911:2904] < mid_1[2903:2896]) ? 1 : 0;
assign detect_min[362][13] = (mid_1[2911:2904] < mid_1[2919:2912]) ? 1 : 0;
assign detect_min[362][14] = (mid_1[2911:2904] < mid_2[2903:2896]) ? 1 : 0;
assign detect_min[362][15] = (mid_1[2911:2904] < mid_2[2911:2904]) ? 1 : 0;
assign detect_min[362][16] = (mid_1[2911:2904] < mid_2[2919:2912]) ? 1 : 0;
assign detect_min[362][17] = (mid_1[2911:2904] < btm_0[2903:2896]) ? 1 : 0;
assign detect_min[362][18] = (mid_1[2911:2904] < btm_0[2911:2904]) ? 1 : 0;
assign detect_min[362][19] = (mid_1[2911:2904] < btm_0[2919:2912]) ? 1 : 0;
assign detect_min[362][20] = (mid_1[2911:2904] < btm_1[2903:2896]) ? 1 : 0;
assign detect_min[362][21] = (mid_1[2911:2904] < btm_1[2911:2904]) ? 1 : 0;
assign detect_min[362][22] = (mid_1[2911:2904] < btm_1[2919:2912]) ? 1 : 0;
assign detect_min[362][23] = (mid_1[2911:2904] < btm_2[2903:2896]) ? 1 : 0;
assign detect_min[362][24] = (mid_1[2911:2904] < btm_2[2911:2904]) ? 1 : 0;
assign detect_min[362][25] = (mid_1[2911:2904] < btm_2[2919:2912]) ? 1 : 0;

assign detect_min[363][0] = (mid_1[2919:2912] < top_0[2911:2904]) ? 1 : 0;
assign detect_min[363][1] = (mid_1[2919:2912] < top_0[2919:2912]) ? 1 : 0;
assign detect_min[363][2] = (mid_1[2919:2912] < top_0[2927:2920]) ? 1 : 0;
assign detect_min[363][3] = (mid_1[2919:2912] < top_1[2911:2904]) ? 1 : 0;
assign detect_min[363][4] = (mid_1[2919:2912] < top_1[2919:2912]) ? 1 : 0;
assign detect_min[363][5] = (mid_1[2919:2912] < top_1[2927:2920]) ? 1 : 0;
assign detect_min[363][6] = (mid_1[2919:2912] < top_2[2911:2904]) ? 1 : 0;
assign detect_min[363][7] = (mid_1[2919:2912] < top_2[2919:2912]) ? 1 : 0;
assign detect_min[363][8] = (mid_1[2919:2912] < top_2[2927:2920]) ? 1 : 0;
assign detect_min[363][9] = (mid_1[2919:2912] < mid_0[2911:2904]) ? 1 : 0;
assign detect_min[363][10] = (mid_1[2919:2912] < mid_0[2919:2912]) ? 1 : 0;
assign detect_min[363][11] = (mid_1[2919:2912] < mid_0[2927:2920]) ? 1 : 0;
assign detect_min[363][12] = (mid_1[2919:2912] < mid_1[2911:2904]) ? 1 : 0;
assign detect_min[363][13] = (mid_1[2919:2912] < mid_1[2927:2920]) ? 1 : 0;
assign detect_min[363][14] = (mid_1[2919:2912] < mid_2[2911:2904]) ? 1 : 0;
assign detect_min[363][15] = (mid_1[2919:2912] < mid_2[2919:2912]) ? 1 : 0;
assign detect_min[363][16] = (mid_1[2919:2912] < mid_2[2927:2920]) ? 1 : 0;
assign detect_min[363][17] = (mid_1[2919:2912] < btm_0[2911:2904]) ? 1 : 0;
assign detect_min[363][18] = (mid_1[2919:2912] < btm_0[2919:2912]) ? 1 : 0;
assign detect_min[363][19] = (mid_1[2919:2912] < btm_0[2927:2920]) ? 1 : 0;
assign detect_min[363][20] = (mid_1[2919:2912] < btm_1[2911:2904]) ? 1 : 0;
assign detect_min[363][21] = (mid_1[2919:2912] < btm_1[2919:2912]) ? 1 : 0;
assign detect_min[363][22] = (mid_1[2919:2912] < btm_1[2927:2920]) ? 1 : 0;
assign detect_min[363][23] = (mid_1[2919:2912] < btm_2[2911:2904]) ? 1 : 0;
assign detect_min[363][24] = (mid_1[2919:2912] < btm_2[2919:2912]) ? 1 : 0;
assign detect_min[363][25] = (mid_1[2919:2912] < btm_2[2927:2920]) ? 1 : 0;

assign detect_min[364][0] = (mid_1[2927:2920] < top_0[2919:2912]) ? 1 : 0;
assign detect_min[364][1] = (mid_1[2927:2920] < top_0[2927:2920]) ? 1 : 0;
assign detect_min[364][2] = (mid_1[2927:2920] < top_0[2935:2928]) ? 1 : 0;
assign detect_min[364][3] = (mid_1[2927:2920] < top_1[2919:2912]) ? 1 : 0;
assign detect_min[364][4] = (mid_1[2927:2920] < top_1[2927:2920]) ? 1 : 0;
assign detect_min[364][5] = (mid_1[2927:2920] < top_1[2935:2928]) ? 1 : 0;
assign detect_min[364][6] = (mid_1[2927:2920] < top_2[2919:2912]) ? 1 : 0;
assign detect_min[364][7] = (mid_1[2927:2920] < top_2[2927:2920]) ? 1 : 0;
assign detect_min[364][8] = (mid_1[2927:2920] < top_2[2935:2928]) ? 1 : 0;
assign detect_min[364][9] = (mid_1[2927:2920] < mid_0[2919:2912]) ? 1 : 0;
assign detect_min[364][10] = (mid_1[2927:2920] < mid_0[2927:2920]) ? 1 : 0;
assign detect_min[364][11] = (mid_1[2927:2920] < mid_0[2935:2928]) ? 1 : 0;
assign detect_min[364][12] = (mid_1[2927:2920] < mid_1[2919:2912]) ? 1 : 0;
assign detect_min[364][13] = (mid_1[2927:2920] < mid_1[2935:2928]) ? 1 : 0;
assign detect_min[364][14] = (mid_1[2927:2920] < mid_2[2919:2912]) ? 1 : 0;
assign detect_min[364][15] = (mid_1[2927:2920] < mid_2[2927:2920]) ? 1 : 0;
assign detect_min[364][16] = (mid_1[2927:2920] < mid_2[2935:2928]) ? 1 : 0;
assign detect_min[364][17] = (mid_1[2927:2920] < btm_0[2919:2912]) ? 1 : 0;
assign detect_min[364][18] = (mid_1[2927:2920] < btm_0[2927:2920]) ? 1 : 0;
assign detect_min[364][19] = (mid_1[2927:2920] < btm_0[2935:2928]) ? 1 : 0;
assign detect_min[364][20] = (mid_1[2927:2920] < btm_1[2919:2912]) ? 1 : 0;
assign detect_min[364][21] = (mid_1[2927:2920] < btm_1[2927:2920]) ? 1 : 0;
assign detect_min[364][22] = (mid_1[2927:2920] < btm_1[2935:2928]) ? 1 : 0;
assign detect_min[364][23] = (mid_1[2927:2920] < btm_2[2919:2912]) ? 1 : 0;
assign detect_min[364][24] = (mid_1[2927:2920] < btm_2[2927:2920]) ? 1 : 0;
assign detect_min[364][25] = (mid_1[2927:2920] < btm_2[2935:2928]) ? 1 : 0;

assign detect_min[365][0] = (mid_1[2935:2928] < top_0[2927:2920]) ? 1 : 0;
assign detect_min[365][1] = (mid_1[2935:2928] < top_0[2935:2928]) ? 1 : 0;
assign detect_min[365][2] = (mid_1[2935:2928] < top_0[2943:2936]) ? 1 : 0;
assign detect_min[365][3] = (mid_1[2935:2928] < top_1[2927:2920]) ? 1 : 0;
assign detect_min[365][4] = (mid_1[2935:2928] < top_1[2935:2928]) ? 1 : 0;
assign detect_min[365][5] = (mid_1[2935:2928] < top_1[2943:2936]) ? 1 : 0;
assign detect_min[365][6] = (mid_1[2935:2928] < top_2[2927:2920]) ? 1 : 0;
assign detect_min[365][7] = (mid_1[2935:2928] < top_2[2935:2928]) ? 1 : 0;
assign detect_min[365][8] = (mid_1[2935:2928] < top_2[2943:2936]) ? 1 : 0;
assign detect_min[365][9] = (mid_1[2935:2928] < mid_0[2927:2920]) ? 1 : 0;
assign detect_min[365][10] = (mid_1[2935:2928] < mid_0[2935:2928]) ? 1 : 0;
assign detect_min[365][11] = (mid_1[2935:2928] < mid_0[2943:2936]) ? 1 : 0;
assign detect_min[365][12] = (mid_1[2935:2928] < mid_1[2927:2920]) ? 1 : 0;
assign detect_min[365][13] = (mid_1[2935:2928] < mid_1[2943:2936]) ? 1 : 0;
assign detect_min[365][14] = (mid_1[2935:2928] < mid_2[2927:2920]) ? 1 : 0;
assign detect_min[365][15] = (mid_1[2935:2928] < mid_2[2935:2928]) ? 1 : 0;
assign detect_min[365][16] = (mid_1[2935:2928] < mid_2[2943:2936]) ? 1 : 0;
assign detect_min[365][17] = (mid_1[2935:2928] < btm_0[2927:2920]) ? 1 : 0;
assign detect_min[365][18] = (mid_1[2935:2928] < btm_0[2935:2928]) ? 1 : 0;
assign detect_min[365][19] = (mid_1[2935:2928] < btm_0[2943:2936]) ? 1 : 0;
assign detect_min[365][20] = (mid_1[2935:2928] < btm_1[2927:2920]) ? 1 : 0;
assign detect_min[365][21] = (mid_1[2935:2928] < btm_1[2935:2928]) ? 1 : 0;
assign detect_min[365][22] = (mid_1[2935:2928] < btm_1[2943:2936]) ? 1 : 0;
assign detect_min[365][23] = (mid_1[2935:2928] < btm_2[2927:2920]) ? 1 : 0;
assign detect_min[365][24] = (mid_1[2935:2928] < btm_2[2935:2928]) ? 1 : 0;
assign detect_min[365][25] = (mid_1[2935:2928] < btm_2[2943:2936]) ? 1 : 0;

assign detect_min[366][0] = (mid_1[2943:2936] < top_0[2935:2928]) ? 1 : 0;
assign detect_min[366][1] = (mid_1[2943:2936] < top_0[2943:2936]) ? 1 : 0;
assign detect_min[366][2] = (mid_1[2943:2936] < top_0[2951:2944]) ? 1 : 0;
assign detect_min[366][3] = (mid_1[2943:2936] < top_1[2935:2928]) ? 1 : 0;
assign detect_min[366][4] = (mid_1[2943:2936] < top_1[2943:2936]) ? 1 : 0;
assign detect_min[366][5] = (mid_1[2943:2936] < top_1[2951:2944]) ? 1 : 0;
assign detect_min[366][6] = (mid_1[2943:2936] < top_2[2935:2928]) ? 1 : 0;
assign detect_min[366][7] = (mid_1[2943:2936] < top_2[2943:2936]) ? 1 : 0;
assign detect_min[366][8] = (mid_1[2943:2936] < top_2[2951:2944]) ? 1 : 0;
assign detect_min[366][9] = (mid_1[2943:2936] < mid_0[2935:2928]) ? 1 : 0;
assign detect_min[366][10] = (mid_1[2943:2936] < mid_0[2943:2936]) ? 1 : 0;
assign detect_min[366][11] = (mid_1[2943:2936] < mid_0[2951:2944]) ? 1 : 0;
assign detect_min[366][12] = (mid_1[2943:2936] < mid_1[2935:2928]) ? 1 : 0;
assign detect_min[366][13] = (mid_1[2943:2936] < mid_1[2951:2944]) ? 1 : 0;
assign detect_min[366][14] = (mid_1[2943:2936] < mid_2[2935:2928]) ? 1 : 0;
assign detect_min[366][15] = (mid_1[2943:2936] < mid_2[2943:2936]) ? 1 : 0;
assign detect_min[366][16] = (mid_1[2943:2936] < mid_2[2951:2944]) ? 1 : 0;
assign detect_min[366][17] = (mid_1[2943:2936] < btm_0[2935:2928]) ? 1 : 0;
assign detect_min[366][18] = (mid_1[2943:2936] < btm_0[2943:2936]) ? 1 : 0;
assign detect_min[366][19] = (mid_1[2943:2936] < btm_0[2951:2944]) ? 1 : 0;
assign detect_min[366][20] = (mid_1[2943:2936] < btm_1[2935:2928]) ? 1 : 0;
assign detect_min[366][21] = (mid_1[2943:2936] < btm_1[2943:2936]) ? 1 : 0;
assign detect_min[366][22] = (mid_1[2943:2936] < btm_1[2951:2944]) ? 1 : 0;
assign detect_min[366][23] = (mid_1[2943:2936] < btm_2[2935:2928]) ? 1 : 0;
assign detect_min[366][24] = (mid_1[2943:2936] < btm_2[2943:2936]) ? 1 : 0;
assign detect_min[366][25] = (mid_1[2943:2936] < btm_2[2951:2944]) ? 1 : 0;

assign detect_min[367][0] = (mid_1[2951:2944] < top_0[2943:2936]) ? 1 : 0;
assign detect_min[367][1] = (mid_1[2951:2944] < top_0[2951:2944]) ? 1 : 0;
assign detect_min[367][2] = (mid_1[2951:2944] < top_0[2959:2952]) ? 1 : 0;
assign detect_min[367][3] = (mid_1[2951:2944] < top_1[2943:2936]) ? 1 : 0;
assign detect_min[367][4] = (mid_1[2951:2944] < top_1[2951:2944]) ? 1 : 0;
assign detect_min[367][5] = (mid_1[2951:2944] < top_1[2959:2952]) ? 1 : 0;
assign detect_min[367][6] = (mid_1[2951:2944] < top_2[2943:2936]) ? 1 : 0;
assign detect_min[367][7] = (mid_1[2951:2944] < top_2[2951:2944]) ? 1 : 0;
assign detect_min[367][8] = (mid_1[2951:2944] < top_2[2959:2952]) ? 1 : 0;
assign detect_min[367][9] = (mid_1[2951:2944] < mid_0[2943:2936]) ? 1 : 0;
assign detect_min[367][10] = (mid_1[2951:2944] < mid_0[2951:2944]) ? 1 : 0;
assign detect_min[367][11] = (mid_1[2951:2944] < mid_0[2959:2952]) ? 1 : 0;
assign detect_min[367][12] = (mid_1[2951:2944] < mid_1[2943:2936]) ? 1 : 0;
assign detect_min[367][13] = (mid_1[2951:2944] < mid_1[2959:2952]) ? 1 : 0;
assign detect_min[367][14] = (mid_1[2951:2944] < mid_2[2943:2936]) ? 1 : 0;
assign detect_min[367][15] = (mid_1[2951:2944] < mid_2[2951:2944]) ? 1 : 0;
assign detect_min[367][16] = (mid_1[2951:2944] < mid_2[2959:2952]) ? 1 : 0;
assign detect_min[367][17] = (mid_1[2951:2944] < btm_0[2943:2936]) ? 1 : 0;
assign detect_min[367][18] = (mid_1[2951:2944] < btm_0[2951:2944]) ? 1 : 0;
assign detect_min[367][19] = (mid_1[2951:2944] < btm_0[2959:2952]) ? 1 : 0;
assign detect_min[367][20] = (mid_1[2951:2944] < btm_1[2943:2936]) ? 1 : 0;
assign detect_min[367][21] = (mid_1[2951:2944] < btm_1[2951:2944]) ? 1 : 0;
assign detect_min[367][22] = (mid_1[2951:2944] < btm_1[2959:2952]) ? 1 : 0;
assign detect_min[367][23] = (mid_1[2951:2944] < btm_2[2943:2936]) ? 1 : 0;
assign detect_min[367][24] = (mid_1[2951:2944] < btm_2[2951:2944]) ? 1 : 0;
assign detect_min[367][25] = (mid_1[2951:2944] < btm_2[2959:2952]) ? 1 : 0;

assign detect_min[368][0] = (mid_1[2959:2952] < top_0[2951:2944]) ? 1 : 0;
assign detect_min[368][1] = (mid_1[2959:2952] < top_0[2959:2952]) ? 1 : 0;
assign detect_min[368][2] = (mid_1[2959:2952] < top_0[2967:2960]) ? 1 : 0;
assign detect_min[368][3] = (mid_1[2959:2952] < top_1[2951:2944]) ? 1 : 0;
assign detect_min[368][4] = (mid_1[2959:2952] < top_1[2959:2952]) ? 1 : 0;
assign detect_min[368][5] = (mid_1[2959:2952] < top_1[2967:2960]) ? 1 : 0;
assign detect_min[368][6] = (mid_1[2959:2952] < top_2[2951:2944]) ? 1 : 0;
assign detect_min[368][7] = (mid_1[2959:2952] < top_2[2959:2952]) ? 1 : 0;
assign detect_min[368][8] = (mid_1[2959:2952] < top_2[2967:2960]) ? 1 : 0;
assign detect_min[368][9] = (mid_1[2959:2952] < mid_0[2951:2944]) ? 1 : 0;
assign detect_min[368][10] = (mid_1[2959:2952] < mid_0[2959:2952]) ? 1 : 0;
assign detect_min[368][11] = (mid_1[2959:2952] < mid_0[2967:2960]) ? 1 : 0;
assign detect_min[368][12] = (mid_1[2959:2952] < mid_1[2951:2944]) ? 1 : 0;
assign detect_min[368][13] = (mid_1[2959:2952] < mid_1[2967:2960]) ? 1 : 0;
assign detect_min[368][14] = (mid_1[2959:2952] < mid_2[2951:2944]) ? 1 : 0;
assign detect_min[368][15] = (mid_1[2959:2952] < mid_2[2959:2952]) ? 1 : 0;
assign detect_min[368][16] = (mid_1[2959:2952] < mid_2[2967:2960]) ? 1 : 0;
assign detect_min[368][17] = (mid_1[2959:2952] < btm_0[2951:2944]) ? 1 : 0;
assign detect_min[368][18] = (mid_1[2959:2952] < btm_0[2959:2952]) ? 1 : 0;
assign detect_min[368][19] = (mid_1[2959:2952] < btm_0[2967:2960]) ? 1 : 0;
assign detect_min[368][20] = (mid_1[2959:2952] < btm_1[2951:2944]) ? 1 : 0;
assign detect_min[368][21] = (mid_1[2959:2952] < btm_1[2959:2952]) ? 1 : 0;
assign detect_min[368][22] = (mid_1[2959:2952] < btm_1[2967:2960]) ? 1 : 0;
assign detect_min[368][23] = (mid_1[2959:2952] < btm_2[2951:2944]) ? 1 : 0;
assign detect_min[368][24] = (mid_1[2959:2952] < btm_2[2959:2952]) ? 1 : 0;
assign detect_min[368][25] = (mid_1[2959:2952] < btm_2[2967:2960]) ? 1 : 0;

assign detect_min[369][0] = (mid_1[2967:2960] < top_0[2959:2952]) ? 1 : 0;
assign detect_min[369][1] = (mid_1[2967:2960] < top_0[2967:2960]) ? 1 : 0;
assign detect_min[369][2] = (mid_1[2967:2960] < top_0[2975:2968]) ? 1 : 0;
assign detect_min[369][3] = (mid_1[2967:2960] < top_1[2959:2952]) ? 1 : 0;
assign detect_min[369][4] = (mid_1[2967:2960] < top_1[2967:2960]) ? 1 : 0;
assign detect_min[369][5] = (mid_1[2967:2960] < top_1[2975:2968]) ? 1 : 0;
assign detect_min[369][6] = (mid_1[2967:2960] < top_2[2959:2952]) ? 1 : 0;
assign detect_min[369][7] = (mid_1[2967:2960] < top_2[2967:2960]) ? 1 : 0;
assign detect_min[369][8] = (mid_1[2967:2960] < top_2[2975:2968]) ? 1 : 0;
assign detect_min[369][9] = (mid_1[2967:2960] < mid_0[2959:2952]) ? 1 : 0;
assign detect_min[369][10] = (mid_1[2967:2960] < mid_0[2967:2960]) ? 1 : 0;
assign detect_min[369][11] = (mid_1[2967:2960] < mid_0[2975:2968]) ? 1 : 0;
assign detect_min[369][12] = (mid_1[2967:2960] < mid_1[2959:2952]) ? 1 : 0;
assign detect_min[369][13] = (mid_1[2967:2960] < mid_1[2975:2968]) ? 1 : 0;
assign detect_min[369][14] = (mid_1[2967:2960] < mid_2[2959:2952]) ? 1 : 0;
assign detect_min[369][15] = (mid_1[2967:2960] < mid_2[2967:2960]) ? 1 : 0;
assign detect_min[369][16] = (mid_1[2967:2960] < mid_2[2975:2968]) ? 1 : 0;
assign detect_min[369][17] = (mid_1[2967:2960] < btm_0[2959:2952]) ? 1 : 0;
assign detect_min[369][18] = (mid_1[2967:2960] < btm_0[2967:2960]) ? 1 : 0;
assign detect_min[369][19] = (mid_1[2967:2960] < btm_0[2975:2968]) ? 1 : 0;
assign detect_min[369][20] = (mid_1[2967:2960] < btm_1[2959:2952]) ? 1 : 0;
assign detect_min[369][21] = (mid_1[2967:2960] < btm_1[2967:2960]) ? 1 : 0;
assign detect_min[369][22] = (mid_1[2967:2960] < btm_1[2975:2968]) ? 1 : 0;
assign detect_min[369][23] = (mid_1[2967:2960] < btm_2[2959:2952]) ? 1 : 0;
assign detect_min[369][24] = (mid_1[2967:2960] < btm_2[2967:2960]) ? 1 : 0;
assign detect_min[369][25] = (mid_1[2967:2960] < btm_2[2975:2968]) ? 1 : 0;

assign detect_min[370][0] = (mid_1[2975:2968] < top_0[2967:2960]) ? 1 : 0;
assign detect_min[370][1] = (mid_1[2975:2968] < top_0[2975:2968]) ? 1 : 0;
assign detect_min[370][2] = (mid_1[2975:2968] < top_0[2983:2976]) ? 1 : 0;
assign detect_min[370][3] = (mid_1[2975:2968] < top_1[2967:2960]) ? 1 : 0;
assign detect_min[370][4] = (mid_1[2975:2968] < top_1[2975:2968]) ? 1 : 0;
assign detect_min[370][5] = (mid_1[2975:2968] < top_1[2983:2976]) ? 1 : 0;
assign detect_min[370][6] = (mid_1[2975:2968] < top_2[2967:2960]) ? 1 : 0;
assign detect_min[370][7] = (mid_1[2975:2968] < top_2[2975:2968]) ? 1 : 0;
assign detect_min[370][8] = (mid_1[2975:2968] < top_2[2983:2976]) ? 1 : 0;
assign detect_min[370][9] = (mid_1[2975:2968] < mid_0[2967:2960]) ? 1 : 0;
assign detect_min[370][10] = (mid_1[2975:2968] < mid_0[2975:2968]) ? 1 : 0;
assign detect_min[370][11] = (mid_1[2975:2968] < mid_0[2983:2976]) ? 1 : 0;
assign detect_min[370][12] = (mid_1[2975:2968] < mid_1[2967:2960]) ? 1 : 0;
assign detect_min[370][13] = (mid_1[2975:2968] < mid_1[2983:2976]) ? 1 : 0;
assign detect_min[370][14] = (mid_1[2975:2968] < mid_2[2967:2960]) ? 1 : 0;
assign detect_min[370][15] = (mid_1[2975:2968] < mid_2[2975:2968]) ? 1 : 0;
assign detect_min[370][16] = (mid_1[2975:2968] < mid_2[2983:2976]) ? 1 : 0;
assign detect_min[370][17] = (mid_1[2975:2968] < btm_0[2967:2960]) ? 1 : 0;
assign detect_min[370][18] = (mid_1[2975:2968] < btm_0[2975:2968]) ? 1 : 0;
assign detect_min[370][19] = (mid_1[2975:2968] < btm_0[2983:2976]) ? 1 : 0;
assign detect_min[370][20] = (mid_1[2975:2968] < btm_1[2967:2960]) ? 1 : 0;
assign detect_min[370][21] = (mid_1[2975:2968] < btm_1[2975:2968]) ? 1 : 0;
assign detect_min[370][22] = (mid_1[2975:2968] < btm_1[2983:2976]) ? 1 : 0;
assign detect_min[370][23] = (mid_1[2975:2968] < btm_2[2967:2960]) ? 1 : 0;
assign detect_min[370][24] = (mid_1[2975:2968] < btm_2[2975:2968]) ? 1 : 0;
assign detect_min[370][25] = (mid_1[2975:2968] < btm_2[2983:2976]) ? 1 : 0;

assign detect_min[371][0] = (mid_1[2983:2976] < top_0[2975:2968]) ? 1 : 0;
assign detect_min[371][1] = (mid_1[2983:2976] < top_0[2983:2976]) ? 1 : 0;
assign detect_min[371][2] = (mid_1[2983:2976] < top_0[2991:2984]) ? 1 : 0;
assign detect_min[371][3] = (mid_1[2983:2976] < top_1[2975:2968]) ? 1 : 0;
assign detect_min[371][4] = (mid_1[2983:2976] < top_1[2983:2976]) ? 1 : 0;
assign detect_min[371][5] = (mid_1[2983:2976] < top_1[2991:2984]) ? 1 : 0;
assign detect_min[371][6] = (mid_1[2983:2976] < top_2[2975:2968]) ? 1 : 0;
assign detect_min[371][7] = (mid_1[2983:2976] < top_2[2983:2976]) ? 1 : 0;
assign detect_min[371][8] = (mid_1[2983:2976] < top_2[2991:2984]) ? 1 : 0;
assign detect_min[371][9] = (mid_1[2983:2976] < mid_0[2975:2968]) ? 1 : 0;
assign detect_min[371][10] = (mid_1[2983:2976] < mid_0[2983:2976]) ? 1 : 0;
assign detect_min[371][11] = (mid_1[2983:2976] < mid_0[2991:2984]) ? 1 : 0;
assign detect_min[371][12] = (mid_1[2983:2976] < mid_1[2975:2968]) ? 1 : 0;
assign detect_min[371][13] = (mid_1[2983:2976] < mid_1[2991:2984]) ? 1 : 0;
assign detect_min[371][14] = (mid_1[2983:2976] < mid_2[2975:2968]) ? 1 : 0;
assign detect_min[371][15] = (mid_1[2983:2976] < mid_2[2983:2976]) ? 1 : 0;
assign detect_min[371][16] = (mid_1[2983:2976] < mid_2[2991:2984]) ? 1 : 0;
assign detect_min[371][17] = (mid_1[2983:2976] < btm_0[2975:2968]) ? 1 : 0;
assign detect_min[371][18] = (mid_1[2983:2976] < btm_0[2983:2976]) ? 1 : 0;
assign detect_min[371][19] = (mid_1[2983:2976] < btm_0[2991:2984]) ? 1 : 0;
assign detect_min[371][20] = (mid_1[2983:2976] < btm_1[2975:2968]) ? 1 : 0;
assign detect_min[371][21] = (mid_1[2983:2976] < btm_1[2983:2976]) ? 1 : 0;
assign detect_min[371][22] = (mid_1[2983:2976] < btm_1[2991:2984]) ? 1 : 0;
assign detect_min[371][23] = (mid_1[2983:2976] < btm_2[2975:2968]) ? 1 : 0;
assign detect_min[371][24] = (mid_1[2983:2976] < btm_2[2983:2976]) ? 1 : 0;
assign detect_min[371][25] = (mid_1[2983:2976] < btm_2[2991:2984]) ? 1 : 0;

assign detect_min[372][0] = (mid_1[2991:2984] < top_0[2983:2976]) ? 1 : 0;
assign detect_min[372][1] = (mid_1[2991:2984] < top_0[2991:2984]) ? 1 : 0;
assign detect_min[372][2] = (mid_1[2991:2984] < top_0[2999:2992]) ? 1 : 0;
assign detect_min[372][3] = (mid_1[2991:2984] < top_1[2983:2976]) ? 1 : 0;
assign detect_min[372][4] = (mid_1[2991:2984] < top_1[2991:2984]) ? 1 : 0;
assign detect_min[372][5] = (mid_1[2991:2984] < top_1[2999:2992]) ? 1 : 0;
assign detect_min[372][6] = (mid_1[2991:2984] < top_2[2983:2976]) ? 1 : 0;
assign detect_min[372][7] = (mid_1[2991:2984] < top_2[2991:2984]) ? 1 : 0;
assign detect_min[372][8] = (mid_1[2991:2984] < top_2[2999:2992]) ? 1 : 0;
assign detect_min[372][9] = (mid_1[2991:2984] < mid_0[2983:2976]) ? 1 : 0;
assign detect_min[372][10] = (mid_1[2991:2984] < mid_0[2991:2984]) ? 1 : 0;
assign detect_min[372][11] = (mid_1[2991:2984] < mid_0[2999:2992]) ? 1 : 0;
assign detect_min[372][12] = (mid_1[2991:2984] < mid_1[2983:2976]) ? 1 : 0;
assign detect_min[372][13] = (mid_1[2991:2984] < mid_1[2999:2992]) ? 1 : 0;
assign detect_min[372][14] = (mid_1[2991:2984] < mid_2[2983:2976]) ? 1 : 0;
assign detect_min[372][15] = (mid_1[2991:2984] < mid_2[2991:2984]) ? 1 : 0;
assign detect_min[372][16] = (mid_1[2991:2984] < mid_2[2999:2992]) ? 1 : 0;
assign detect_min[372][17] = (mid_1[2991:2984] < btm_0[2983:2976]) ? 1 : 0;
assign detect_min[372][18] = (mid_1[2991:2984] < btm_0[2991:2984]) ? 1 : 0;
assign detect_min[372][19] = (mid_1[2991:2984] < btm_0[2999:2992]) ? 1 : 0;
assign detect_min[372][20] = (mid_1[2991:2984] < btm_1[2983:2976]) ? 1 : 0;
assign detect_min[372][21] = (mid_1[2991:2984] < btm_1[2991:2984]) ? 1 : 0;
assign detect_min[372][22] = (mid_1[2991:2984] < btm_1[2999:2992]) ? 1 : 0;
assign detect_min[372][23] = (mid_1[2991:2984] < btm_2[2983:2976]) ? 1 : 0;
assign detect_min[372][24] = (mid_1[2991:2984] < btm_2[2991:2984]) ? 1 : 0;
assign detect_min[372][25] = (mid_1[2991:2984] < btm_2[2999:2992]) ? 1 : 0;

assign detect_min[373][0] = (mid_1[2999:2992] < top_0[2991:2984]) ? 1 : 0;
assign detect_min[373][1] = (mid_1[2999:2992] < top_0[2999:2992]) ? 1 : 0;
assign detect_min[373][2] = (mid_1[2999:2992] < top_0[3007:3000]) ? 1 : 0;
assign detect_min[373][3] = (mid_1[2999:2992] < top_1[2991:2984]) ? 1 : 0;
assign detect_min[373][4] = (mid_1[2999:2992] < top_1[2999:2992]) ? 1 : 0;
assign detect_min[373][5] = (mid_1[2999:2992] < top_1[3007:3000]) ? 1 : 0;
assign detect_min[373][6] = (mid_1[2999:2992] < top_2[2991:2984]) ? 1 : 0;
assign detect_min[373][7] = (mid_1[2999:2992] < top_2[2999:2992]) ? 1 : 0;
assign detect_min[373][8] = (mid_1[2999:2992] < top_2[3007:3000]) ? 1 : 0;
assign detect_min[373][9] = (mid_1[2999:2992] < mid_0[2991:2984]) ? 1 : 0;
assign detect_min[373][10] = (mid_1[2999:2992] < mid_0[2999:2992]) ? 1 : 0;
assign detect_min[373][11] = (mid_1[2999:2992] < mid_0[3007:3000]) ? 1 : 0;
assign detect_min[373][12] = (mid_1[2999:2992] < mid_1[2991:2984]) ? 1 : 0;
assign detect_min[373][13] = (mid_1[2999:2992] < mid_1[3007:3000]) ? 1 : 0;
assign detect_min[373][14] = (mid_1[2999:2992] < mid_2[2991:2984]) ? 1 : 0;
assign detect_min[373][15] = (mid_1[2999:2992] < mid_2[2999:2992]) ? 1 : 0;
assign detect_min[373][16] = (mid_1[2999:2992] < mid_2[3007:3000]) ? 1 : 0;
assign detect_min[373][17] = (mid_1[2999:2992] < btm_0[2991:2984]) ? 1 : 0;
assign detect_min[373][18] = (mid_1[2999:2992] < btm_0[2999:2992]) ? 1 : 0;
assign detect_min[373][19] = (mid_1[2999:2992] < btm_0[3007:3000]) ? 1 : 0;
assign detect_min[373][20] = (mid_1[2999:2992] < btm_1[2991:2984]) ? 1 : 0;
assign detect_min[373][21] = (mid_1[2999:2992] < btm_1[2999:2992]) ? 1 : 0;
assign detect_min[373][22] = (mid_1[2999:2992] < btm_1[3007:3000]) ? 1 : 0;
assign detect_min[373][23] = (mid_1[2999:2992] < btm_2[2991:2984]) ? 1 : 0;
assign detect_min[373][24] = (mid_1[2999:2992] < btm_2[2999:2992]) ? 1 : 0;
assign detect_min[373][25] = (mid_1[2999:2992] < btm_2[3007:3000]) ? 1 : 0;

assign detect_min[374][0] = (mid_1[3007:3000] < top_0[2999:2992]) ? 1 : 0;
assign detect_min[374][1] = (mid_1[3007:3000] < top_0[3007:3000]) ? 1 : 0;
assign detect_min[374][2] = (mid_1[3007:3000] < top_0[3015:3008]) ? 1 : 0;
assign detect_min[374][3] = (mid_1[3007:3000] < top_1[2999:2992]) ? 1 : 0;
assign detect_min[374][4] = (mid_1[3007:3000] < top_1[3007:3000]) ? 1 : 0;
assign detect_min[374][5] = (mid_1[3007:3000] < top_1[3015:3008]) ? 1 : 0;
assign detect_min[374][6] = (mid_1[3007:3000] < top_2[2999:2992]) ? 1 : 0;
assign detect_min[374][7] = (mid_1[3007:3000] < top_2[3007:3000]) ? 1 : 0;
assign detect_min[374][8] = (mid_1[3007:3000] < top_2[3015:3008]) ? 1 : 0;
assign detect_min[374][9] = (mid_1[3007:3000] < mid_0[2999:2992]) ? 1 : 0;
assign detect_min[374][10] = (mid_1[3007:3000] < mid_0[3007:3000]) ? 1 : 0;
assign detect_min[374][11] = (mid_1[3007:3000] < mid_0[3015:3008]) ? 1 : 0;
assign detect_min[374][12] = (mid_1[3007:3000] < mid_1[2999:2992]) ? 1 : 0;
assign detect_min[374][13] = (mid_1[3007:3000] < mid_1[3015:3008]) ? 1 : 0;
assign detect_min[374][14] = (mid_1[3007:3000] < mid_2[2999:2992]) ? 1 : 0;
assign detect_min[374][15] = (mid_1[3007:3000] < mid_2[3007:3000]) ? 1 : 0;
assign detect_min[374][16] = (mid_1[3007:3000] < mid_2[3015:3008]) ? 1 : 0;
assign detect_min[374][17] = (mid_1[3007:3000] < btm_0[2999:2992]) ? 1 : 0;
assign detect_min[374][18] = (mid_1[3007:3000] < btm_0[3007:3000]) ? 1 : 0;
assign detect_min[374][19] = (mid_1[3007:3000] < btm_0[3015:3008]) ? 1 : 0;
assign detect_min[374][20] = (mid_1[3007:3000] < btm_1[2999:2992]) ? 1 : 0;
assign detect_min[374][21] = (mid_1[3007:3000] < btm_1[3007:3000]) ? 1 : 0;
assign detect_min[374][22] = (mid_1[3007:3000] < btm_1[3015:3008]) ? 1 : 0;
assign detect_min[374][23] = (mid_1[3007:3000] < btm_2[2999:2992]) ? 1 : 0;
assign detect_min[374][24] = (mid_1[3007:3000] < btm_2[3007:3000]) ? 1 : 0;
assign detect_min[374][25] = (mid_1[3007:3000] < btm_2[3015:3008]) ? 1 : 0;

assign detect_min[375][0] = (mid_1[3015:3008] < top_0[3007:3000]) ? 1 : 0;
assign detect_min[375][1] = (mid_1[3015:3008] < top_0[3015:3008]) ? 1 : 0;
assign detect_min[375][2] = (mid_1[3015:3008] < top_0[3023:3016]) ? 1 : 0;
assign detect_min[375][3] = (mid_1[3015:3008] < top_1[3007:3000]) ? 1 : 0;
assign detect_min[375][4] = (mid_1[3015:3008] < top_1[3015:3008]) ? 1 : 0;
assign detect_min[375][5] = (mid_1[3015:3008] < top_1[3023:3016]) ? 1 : 0;
assign detect_min[375][6] = (mid_1[3015:3008] < top_2[3007:3000]) ? 1 : 0;
assign detect_min[375][7] = (mid_1[3015:3008] < top_2[3015:3008]) ? 1 : 0;
assign detect_min[375][8] = (mid_1[3015:3008] < top_2[3023:3016]) ? 1 : 0;
assign detect_min[375][9] = (mid_1[3015:3008] < mid_0[3007:3000]) ? 1 : 0;
assign detect_min[375][10] = (mid_1[3015:3008] < mid_0[3015:3008]) ? 1 : 0;
assign detect_min[375][11] = (mid_1[3015:3008] < mid_0[3023:3016]) ? 1 : 0;
assign detect_min[375][12] = (mid_1[3015:3008] < mid_1[3007:3000]) ? 1 : 0;
assign detect_min[375][13] = (mid_1[3015:3008] < mid_1[3023:3016]) ? 1 : 0;
assign detect_min[375][14] = (mid_1[3015:3008] < mid_2[3007:3000]) ? 1 : 0;
assign detect_min[375][15] = (mid_1[3015:3008] < mid_2[3015:3008]) ? 1 : 0;
assign detect_min[375][16] = (mid_1[3015:3008] < mid_2[3023:3016]) ? 1 : 0;
assign detect_min[375][17] = (mid_1[3015:3008] < btm_0[3007:3000]) ? 1 : 0;
assign detect_min[375][18] = (mid_1[3015:3008] < btm_0[3015:3008]) ? 1 : 0;
assign detect_min[375][19] = (mid_1[3015:3008] < btm_0[3023:3016]) ? 1 : 0;
assign detect_min[375][20] = (mid_1[3015:3008] < btm_1[3007:3000]) ? 1 : 0;
assign detect_min[375][21] = (mid_1[3015:3008] < btm_1[3015:3008]) ? 1 : 0;
assign detect_min[375][22] = (mid_1[3015:3008] < btm_1[3023:3016]) ? 1 : 0;
assign detect_min[375][23] = (mid_1[3015:3008] < btm_2[3007:3000]) ? 1 : 0;
assign detect_min[375][24] = (mid_1[3015:3008] < btm_2[3015:3008]) ? 1 : 0;
assign detect_min[375][25] = (mid_1[3015:3008] < btm_2[3023:3016]) ? 1 : 0;

assign detect_min[376][0] = (mid_1[3023:3016] < top_0[3015:3008]) ? 1 : 0;
assign detect_min[376][1] = (mid_1[3023:3016] < top_0[3023:3016]) ? 1 : 0;
assign detect_min[376][2] = (mid_1[3023:3016] < top_0[3031:3024]) ? 1 : 0;
assign detect_min[376][3] = (mid_1[3023:3016] < top_1[3015:3008]) ? 1 : 0;
assign detect_min[376][4] = (mid_1[3023:3016] < top_1[3023:3016]) ? 1 : 0;
assign detect_min[376][5] = (mid_1[3023:3016] < top_1[3031:3024]) ? 1 : 0;
assign detect_min[376][6] = (mid_1[3023:3016] < top_2[3015:3008]) ? 1 : 0;
assign detect_min[376][7] = (mid_1[3023:3016] < top_2[3023:3016]) ? 1 : 0;
assign detect_min[376][8] = (mid_1[3023:3016] < top_2[3031:3024]) ? 1 : 0;
assign detect_min[376][9] = (mid_1[3023:3016] < mid_0[3015:3008]) ? 1 : 0;
assign detect_min[376][10] = (mid_1[3023:3016] < mid_0[3023:3016]) ? 1 : 0;
assign detect_min[376][11] = (mid_1[3023:3016] < mid_0[3031:3024]) ? 1 : 0;
assign detect_min[376][12] = (mid_1[3023:3016] < mid_1[3015:3008]) ? 1 : 0;
assign detect_min[376][13] = (mid_1[3023:3016] < mid_1[3031:3024]) ? 1 : 0;
assign detect_min[376][14] = (mid_1[3023:3016] < mid_2[3015:3008]) ? 1 : 0;
assign detect_min[376][15] = (mid_1[3023:3016] < mid_2[3023:3016]) ? 1 : 0;
assign detect_min[376][16] = (mid_1[3023:3016] < mid_2[3031:3024]) ? 1 : 0;
assign detect_min[376][17] = (mid_1[3023:3016] < btm_0[3015:3008]) ? 1 : 0;
assign detect_min[376][18] = (mid_1[3023:3016] < btm_0[3023:3016]) ? 1 : 0;
assign detect_min[376][19] = (mid_1[3023:3016] < btm_0[3031:3024]) ? 1 : 0;
assign detect_min[376][20] = (mid_1[3023:3016] < btm_1[3015:3008]) ? 1 : 0;
assign detect_min[376][21] = (mid_1[3023:3016] < btm_1[3023:3016]) ? 1 : 0;
assign detect_min[376][22] = (mid_1[3023:3016] < btm_1[3031:3024]) ? 1 : 0;
assign detect_min[376][23] = (mid_1[3023:3016] < btm_2[3015:3008]) ? 1 : 0;
assign detect_min[376][24] = (mid_1[3023:3016] < btm_2[3023:3016]) ? 1 : 0;
assign detect_min[376][25] = (mid_1[3023:3016] < btm_2[3031:3024]) ? 1 : 0;

assign detect_min[377][0] = (mid_1[3031:3024] < top_0[3023:3016]) ? 1 : 0;
assign detect_min[377][1] = (mid_1[3031:3024] < top_0[3031:3024]) ? 1 : 0;
assign detect_min[377][2] = (mid_1[3031:3024] < top_0[3039:3032]) ? 1 : 0;
assign detect_min[377][3] = (mid_1[3031:3024] < top_1[3023:3016]) ? 1 : 0;
assign detect_min[377][4] = (mid_1[3031:3024] < top_1[3031:3024]) ? 1 : 0;
assign detect_min[377][5] = (mid_1[3031:3024] < top_1[3039:3032]) ? 1 : 0;
assign detect_min[377][6] = (mid_1[3031:3024] < top_2[3023:3016]) ? 1 : 0;
assign detect_min[377][7] = (mid_1[3031:3024] < top_2[3031:3024]) ? 1 : 0;
assign detect_min[377][8] = (mid_1[3031:3024] < top_2[3039:3032]) ? 1 : 0;
assign detect_min[377][9] = (mid_1[3031:3024] < mid_0[3023:3016]) ? 1 : 0;
assign detect_min[377][10] = (mid_1[3031:3024] < mid_0[3031:3024]) ? 1 : 0;
assign detect_min[377][11] = (mid_1[3031:3024] < mid_0[3039:3032]) ? 1 : 0;
assign detect_min[377][12] = (mid_1[3031:3024] < mid_1[3023:3016]) ? 1 : 0;
assign detect_min[377][13] = (mid_1[3031:3024] < mid_1[3039:3032]) ? 1 : 0;
assign detect_min[377][14] = (mid_1[3031:3024] < mid_2[3023:3016]) ? 1 : 0;
assign detect_min[377][15] = (mid_1[3031:3024] < mid_2[3031:3024]) ? 1 : 0;
assign detect_min[377][16] = (mid_1[3031:3024] < mid_2[3039:3032]) ? 1 : 0;
assign detect_min[377][17] = (mid_1[3031:3024] < btm_0[3023:3016]) ? 1 : 0;
assign detect_min[377][18] = (mid_1[3031:3024] < btm_0[3031:3024]) ? 1 : 0;
assign detect_min[377][19] = (mid_1[3031:3024] < btm_0[3039:3032]) ? 1 : 0;
assign detect_min[377][20] = (mid_1[3031:3024] < btm_1[3023:3016]) ? 1 : 0;
assign detect_min[377][21] = (mid_1[3031:3024] < btm_1[3031:3024]) ? 1 : 0;
assign detect_min[377][22] = (mid_1[3031:3024] < btm_1[3039:3032]) ? 1 : 0;
assign detect_min[377][23] = (mid_1[3031:3024] < btm_2[3023:3016]) ? 1 : 0;
assign detect_min[377][24] = (mid_1[3031:3024] < btm_2[3031:3024]) ? 1 : 0;
assign detect_min[377][25] = (mid_1[3031:3024] < btm_2[3039:3032]) ? 1 : 0;

assign detect_min[378][0] = (mid_1[3039:3032] < top_0[3031:3024]) ? 1 : 0;
assign detect_min[378][1] = (mid_1[3039:3032] < top_0[3039:3032]) ? 1 : 0;
assign detect_min[378][2] = (mid_1[3039:3032] < top_0[3047:3040]) ? 1 : 0;
assign detect_min[378][3] = (mid_1[3039:3032] < top_1[3031:3024]) ? 1 : 0;
assign detect_min[378][4] = (mid_1[3039:3032] < top_1[3039:3032]) ? 1 : 0;
assign detect_min[378][5] = (mid_1[3039:3032] < top_1[3047:3040]) ? 1 : 0;
assign detect_min[378][6] = (mid_1[3039:3032] < top_2[3031:3024]) ? 1 : 0;
assign detect_min[378][7] = (mid_1[3039:3032] < top_2[3039:3032]) ? 1 : 0;
assign detect_min[378][8] = (mid_1[3039:3032] < top_2[3047:3040]) ? 1 : 0;
assign detect_min[378][9] = (mid_1[3039:3032] < mid_0[3031:3024]) ? 1 : 0;
assign detect_min[378][10] = (mid_1[3039:3032] < mid_0[3039:3032]) ? 1 : 0;
assign detect_min[378][11] = (mid_1[3039:3032] < mid_0[3047:3040]) ? 1 : 0;
assign detect_min[378][12] = (mid_1[3039:3032] < mid_1[3031:3024]) ? 1 : 0;
assign detect_min[378][13] = (mid_1[3039:3032] < mid_1[3047:3040]) ? 1 : 0;
assign detect_min[378][14] = (mid_1[3039:3032] < mid_2[3031:3024]) ? 1 : 0;
assign detect_min[378][15] = (mid_1[3039:3032] < mid_2[3039:3032]) ? 1 : 0;
assign detect_min[378][16] = (mid_1[3039:3032] < mid_2[3047:3040]) ? 1 : 0;
assign detect_min[378][17] = (mid_1[3039:3032] < btm_0[3031:3024]) ? 1 : 0;
assign detect_min[378][18] = (mid_1[3039:3032] < btm_0[3039:3032]) ? 1 : 0;
assign detect_min[378][19] = (mid_1[3039:3032] < btm_0[3047:3040]) ? 1 : 0;
assign detect_min[378][20] = (mid_1[3039:3032] < btm_1[3031:3024]) ? 1 : 0;
assign detect_min[378][21] = (mid_1[3039:3032] < btm_1[3039:3032]) ? 1 : 0;
assign detect_min[378][22] = (mid_1[3039:3032] < btm_1[3047:3040]) ? 1 : 0;
assign detect_min[378][23] = (mid_1[3039:3032] < btm_2[3031:3024]) ? 1 : 0;
assign detect_min[378][24] = (mid_1[3039:3032] < btm_2[3039:3032]) ? 1 : 0;
assign detect_min[378][25] = (mid_1[3039:3032] < btm_2[3047:3040]) ? 1 : 0;

assign detect_min[379][0] = (mid_1[3047:3040] < top_0[3039:3032]) ? 1 : 0;
assign detect_min[379][1] = (mid_1[3047:3040] < top_0[3047:3040]) ? 1 : 0;
assign detect_min[379][2] = (mid_1[3047:3040] < top_0[3055:3048]) ? 1 : 0;
assign detect_min[379][3] = (mid_1[3047:3040] < top_1[3039:3032]) ? 1 : 0;
assign detect_min[379][4] = (mid_1[3047:3040] < top_1[3047:3040]) ? 1 : 0;
assign detect_min[379][5] = (mid_1[3047:3040] < top_1[3055:3048]) ? 1 : 0;
assign detect_min[379][6] = (mid_1[3047:3040] < top_2[3039:3032]) ? 1 : 0;
assign detect_min[379][7] = (mid_1[3047:3040] < top_2[3047:3040]) ? 1 : 0;
assign detect_min[379][8] = (mid_1[3047:3040] < top_2[3055:3048]) ? 1 : 0;
assign detect_min[379][9] = (mid_1[3047:3040] < mid_0[3039:3032]) ? 1 : 0;
assign detect_min[379][10] = (mid_1[3047:3040] < mid_0[3047:3040]) ? 1 : 0;
assign detect_min[379][11] = (mid_1[3047:3040] < mid_0[3055:3048]) ? 1 : 0;
assign detect_min[379][12] = (mid_1[3047:3040] < mid_1[3039:3032]) ? 1 : 0;
assign detect_min[379][13] = (mid_1[3047:3040] < mid_1[3055:3048]) ? 1 : 0;
assign detect_min[379][14] = (mid_1[3047:3040] < mid_2[3039:3032]) ? 1 : 0;
assign detect_min[379][15] = (mid_1[3047:3040] < mid_2[3047:3040]) ? 1 : 0;
assign detect_min[379][16] = (mid_1[3047:3040] < mid_2[3055:3048]) ? 1 : 0;
assign detect_min[379][17] = (mid_1[3047:3040] < btm_0[3039:3032]) ? 1 : 0;
assign detect_min[379][18] = (mid_1[3047:3040] < btm_0[3047:3040]) ? 1 : 0;
assign detect_min[379][19] = (mid_1[3047:3040] < btm_0[3055:3048]) ? 1 : 0;
assign detect_min[379][20] = (mid_1[3047:3040] < btm_1[3039:3032]) ? 1 : 0;
assign detect_min[379][21] = (mid_1[3047:3040] < btm_1[3047:3040]) ? 1 : 0;
assign detect_min[379][22] = (mid_1[3047:3040] < btm_1[3055:3048]) ? 1 : 0;
assign detect_min[379][23] = (mid_1[3047:3040] < btm_2[3039:3032]) ? 1 : 0;
assign detect_min[379][24] = (mid_1[3047:3040] < btm_2[3047:3040]) ? 1 : 0;
assign detect_min[379][25] = (mid_1[3047:3040] < btm_2[3055:3048]) ? 1 : 0;

assign detect_min[380][0] = (mid_1[3055:3048] < top_0[3047:3040]) ? 1 : 0;
assign detect_min[380][1] = (mid_1[3055:3048] < top_0[3055:3048]) ? 1 : 0;
assign detect_min[380][2] = (mid_1[3055:3048] < top_0[3063:3056]) ? 1 : 0;
assign detect_min[380][3] = (mid_1[3055:3048] < top_1[3047:3040]) ? 1 : 0;
assign detect_min[380][4] = (mid_1[3055:3048] < top_1[3055:3048]) ? 1 : 0;
assign detect_min[380][5] = (mid_1[3055:3048] < top_1[3063:3056]) ? 1 : 0;
assign detect_min[380][6] = (mid_1[3055:3048] < top_2[3047:3040]) ? 1 : 0;
assign detect_min[380][7] = (mid_1[3055:3048] < top_2[3055:3048]) ? 1 : 0;
assign detect_min[380][8] = (mid_1[3055:3048] < top_2[3063:3056]) ? 1 : 0;
assign detect_min[380][9] = (mid_1[3055:3048] < mid_0[3047:3040]) ? 1 : 0;
assign detect_min[380][10] = (mid_1[3055:3048] < mid_0[3055:3048]) ? 1 : 0;
assign detect_min[380][11] = (mid_1[3055:3048] < mid_0[3063:3056]) ? 1 : 0;
assign detect_min[380][12] = (mid_1[3055:3048] < mid_1[3047:3040]) ? 1 : 0;
assign detect_min[380][13] = (mid_1[3055:3048] < mid_1[3063:3056]) ? 1 : 0;
assign detect_min[380][14] = (mid_1[3055:3048] < mid_2[3047:3040]) ? 1 : 0;
assign detect_min[380][15] = (mid_1[3055:3048] < mid_2[3055:3048]) ? 1 : 0;
assign detect_min[380][16] = (mid_1[3055:3048] < mid_2[3063:3056]) ? 1 : 0;
assign detect_min[380][17] = (mid_1[3055:3048] < btm_0[3047:3040]) ? 1 : 0;
assign detect_min[380][18] = (mid_1[3055:3048] < btm_0[3055:3048]) ? 1 : 0;
assign detect_min[380][19] = (mid_1[3055:3048] < btm_0[3063:3056]) ? 1 : 0;
assign detect_min[380][20] = (mid_1[3055:3048] < btm_1[3047:3040]) ? 1 : 0;
assign detect_min[380][21] = (mid_1[3055:3048] < btm_1[3055:3048]) ? 1 : 0;
assign detect_min[380][22] = (mid_1[3055:3048] < btm_1[3063:3056]) ? 1 : 0;
assign detect_min[380][23] = (mid_1[3055:3048] < btm_2[3047:3040]) ? 1 : 0;
assign detect_min[380][24] = (mid_1[3055:3048] < btm_2[3055:3048]) ? 1 : 0;
assign detect_min[380][25] = (mid_1[3055:3048] < btm_2[3063:3056]) ? 1 : 0;

assign detect_min[381][0] = (mid_1[3063:3056] < top_0[3055:3048]) ? 1 : 0;
assign detect_min[381][1] = (mid_1[3063:3056] < top_0[3063:3056]) ? 1 : 0;
assign detect_min[381][2] = (mid_1[3063:3056] < top_0[3071:3064]) ? 1 : 0;
assign detect_min[381][3] = (mid_1[3063:3056] < top_1[3055:3048]) ? 1 : 0;
assign detect_min[381][4] = (mid_1[3063:3056] < top_1[3063:3056]) ? 1 : 0;
assign detect_min[381][5] = (mid_1[3063:3056] < top_1[3071:3064]) ? 1 : 0;
assign detect_min[381][6] = (mid_1[3063:3056] < top_2[3055:3048]) ? 1 : 0;
assign detect_min[381][7] = (mid_1[3063:3056] < top_2[3063:3056]) ? 1 : 0;
assign detect_min[381][8] = (mid_1[3063:3056] < top_2[3071:3064]) ? 1 : 0;
assign detect_min[381][9] = (mid_1[3063:3056] < mid_0[3055:3048]) ? 1 : 0;
assign detect_min[381][10] = (mid_1[3063:3056] < mid_0[3063:3056]) ? 1 : 0;
assign detect_min[381][11] = (mid_1[3063:3056] < mid_0[3071:3064]) ? 1 : 0;
assign detect_min[381][12] = (mid_1[3063:3056] < mid_1[3055:3048]) ? 1 : 0;
assign detect_min[381][13] = (mid_1[3063:3056] < mid_1[3071:3064]) ? 1 : 0;
assign detect_min[381][14] = (mid_1[3063:3056] < mid_2[3055:3048]) ? 1 : 0;
assign detect_min[381][15] = (mid_1[3063:3056] < mid_2[3063:3056]) ? 1 : 0;
assign detect_min[381][16] = (mid_1[3063:3056] < mid_2[3071:3064]) ? 1 : 0;
assign detect_min[381][17] = (mid_1[3063:3056] < btm_0[3055:3048]) ? 1 : 0;
assign detect_min[381][18] = (mid_1[3063:3056] < btm_0[3063:3056]) ? 1 : 0;
assign detect_min[381][19] = (mid_1[3063:3056] < btm_0[3071:3064]) ? 1 : 0;
assign detect_min[381][20] = (mid_1[3063:3056] < btm_1[3055:3048]) ? 1 : 0;
assign detect_min[381][21] = (mid_1[3063:3056] < btm_1[3063:3056]) ? 1 : 0;
assign detect_min[381][22] = (mid_1[3063:3056] < btm_1[3071:3064]) ? 1 : 0;
assign detect_min[381][23] = (mid_1[3063:3056] < btm_2[3055:3048]) ? 1 : 0;
assign detect_min[381][24] = (mid_1[3063:3056] < btm_2[3063:3056]) ? 1 : 0;
assign detect_min[381][25] = (mid_1[3063:3056] < btm_2[3071:3064]) ? 1 : 0;

assign detect_min[382][0] = (mid_1[3071:3064] < top_0[3063:3056]) ? 1 : 0;
assign detect_min[382][1] = (mid_1[3071:3064] < top_0[3071:3064]) ? 1 : 0;
assign detect_min[382][2] = (mid_1[3071:3064] < top_0[3079:3072]) ? 1 : 0;
assign detect_min[382][3] = (mid_1[3071:3064] < top_1[3063:3056]) ? 1 : 0;
assign detect_min[382][4] = (mid_1[3071:3064] < top_1[3071:3064]) ? 1 : 0;
assign detect_min[382][5] = (mid_1[3071:3064] < top_1[3079:3072]) ? 1 : 0;
assign detect_min[382][6] = (mid_1[3071:3064] < top_2[3063:3056]) ? 1 : 0;
assign detect_min[382][7] = (mid_1[3071:3064] < top_2[3071:3064]) ? 1 : 0;
assign detect_min[382][8] = (mid_1[3071:3064] < top_2[3079:3072]) ? 1 : 0;
assign detect_min[382][9] = (mid_1[3071:3064] < mid_0[3063:3056]) ? 1 : 0;
assign detect_min[382][10] = (mid_1[3071:3064] < mid_0[3071:3064]) ? 1 : 0;
assign detect_min[382][11] = (mid_1[3071:3064] < mid_0[3079:3072]) ? 1 : 0;
assign detect_min[382][12] = (mid_1[3071:3064] < mid_1[3063:3056]) ? 1 : 0;
assign detect_min[382][13] = (mid_1[3071:3064] < mid_1[3079:3072]) ? 1 : 0;
assign detect_min[382][14] = (mid_1[3071:3064] < mid_2[3063:3056]) ? 1 : 0;
assign detect_min[382][15] = (mid_1[3071:3064] < mid_2[3071:3064]) ? 1 : 0;
assign detect_min[382][16] = (mid_1[3071:3064] < mid_2[3079:3072]) ? 1 : 0;
assign detect_min[382][17] = (mid_1[3071:3064] < btm_0[3063:3056]) ? 1 : 0;
assign detect_min[382][18] = (mid_1[3071:3064] < btm_0[3071:3064]) ? 1 : 0;
assign detect_min[382][19] = (mid_1[3071:3064] < btm_0[3079:3072]) ? 1 : 0;
assign detect_min[382][20] = (mid_1[3071:3064] < btm_1[3063:3056]) ? 1 : 0;
assign detect_min[382][21] = (mid_1[3071:3064] < btm_1[3071:3064]) ? 1 : 0;
assign detect_min[382][22] = (mid_1[3071:3064] < btm_1[3079:3072]) ? 1 : 0;
assign detect_min[382][23] = (mid_1[3071:3064] < btm_2[3063:3056]) ? 1 : 0;
assign detect_min[382][24] = (mid_1[3071:3064] < btm_2[3071:3064]) ? 1 : 0;
assign detect_min[382][25] = (mid_1[3071:3064] < btm_2[3079:3072]) ? 1 : 0;

assign detect_min[383][0] = (mid_1[3079:3072] < top_0[3071:3064]) ? 1 : 0;
assign detect_min[383][1] = (mid_1[3079:3072] < top_0[3079:3072]) ? 1 : 0;
assign detect_min[383][2] = (mid_1[3079:3072] < top_0[3087:3080]) ? 1 : 0;
assign detect_min[383][3] = (mid_1[3079:3072] < top_1[3071:3064]) ? 1 : 0;
assign detect_min[383][4] = (mid_1[3079:3072] < top_1[3079:3072]) ? 1 : 0;
assign detect_min[383][5] = (mid_1[3079:3072] < top_1[3087:3080]) ? 1 : 0;
assign detect_min[383][6] = (mid_1[3079:3072] < top_2[3071:3064]) ? 1 : 0;
assign detect_min[383][7] = (mid_1[3079:3072] < top_2[3079:3072]) ? 1 : 0;
assign detect_min[383][8] = (mid_1[3079:3072] < top_2[3087:3080]) ? 1 : 0;
assign detect_min[383][9] = (mid_1[3079:3072] < mid_0[3071:3064]) ? 1 : 0;
assign detect_min[383][10] = (mid_1[3079:3072] < mid_0[3079:3072]) ? 1 : 0;
assign detect_min[383][11] = (mid_1[3079:3072] < mid_0[3087:3080]) ? 1 : 0;
assign detect_min[383][12] = (mid_1[3079:3072] < mid_1[3071:3064]) ? 1 : 0;
assign detect_min[383][13] = (mid_1[3079:3072] < mid_1[3087:3080]) ? 1 : 0;
assign detect_min[383][14] = (mid_1[3079:3072] < mid_2[3071:3064]) ? 1 : 0;
assign detect_min[383][15] = (mid_1[3079:3072] < mid_2[3079:3072]) ? 1 : 0;
assign detect_min[383][16] = (mid_1[3079:3072] < mid_2[3087:3080]) ? 1 : 0;
assign detect_min[383][17] = (mid_1[3079:3072] < btm_0[3071:3064]) ? 1 : 0;
assign detect_min[383][18] = (mid_1[3079:3072] < btm_0[3079:3072]) ? 1 : 0;
assign detect_min[383][19] = (mid_1[3079:3072] < btm_0[3087:3080]) ? 1 : 0;
assign detect_min[383][20] = (mid_1[3079:3072] < btm_1[3071:3064]) ? 1 : 0;
assign detect_min[383][21] = (mid_1[3079:3072] < btm_1[3079:3072]) ? 1 : 0;
assign detect_min[383][22] = (mid_1[3079:3072] < btm_1[3087:3080]) ? 1 : 0;
assign detect_min[383][23] = (mid_1[3079:3072] < btm_2[3071:3064]) ? 1 : 0;
assign detect_min[383][24] = (mid_1[3079:3072] < btm_2[3079:3072]) ? 1 : 0;
assign detect_min[383][25] = (mid_1[3079:3072] < btm_2[3087:3080]) ? 1 : 0;

assign detect_min[384][0] = (mid_1[3087:3080] < top_0[3079:3072]) ? 1 : 0;
assign detect_min[384][1] = (mid_1[3087:3080] < top_0[3087:3080]) ? 1 : 0;
assign detect_min[384][2] = (mid_1[3087:3080] < top_0[3095:3088]) ? 1 : 0;
assign detect_min[384][3] = (mid_1[3087:3080] < top_1[3079:3072]) ? 1 : 0;
assign detect_min[384][4] = (mid_1[3087:3080] < top_1[3087:3080]) ? 1 : 0;
assign detect_min[384][5] = (mid_1[3087:3080] < top_1[3095:3088]) ? 1 : 0;
assign detect_min[384][6] = (mid_1[3087:3080] < top_2[3079:3072]) ? 1 : 0;
assign detect_min[384][7] = (mid_1[3087:3080] < top_2[3087:3080]) ? 1 : 0;
assign detect_min[384][8] = (mid_1[3087:3080] < top_2[3095:3088]) ? 1 : 0;
assign detect_min[384][9] = (mid_1[3087:3080] < mid_0[3079:3072]) ? 1 : 0;
assign detect_min[384][10] = (mid_1[3087:3080] < mid_0[3087:3080]) ? 1 : 0;
assign detect_min[384][11] = (mid_1[3087:3080] < mid_0[3095:3088]) ? 1 : 0;
assign detect_min[384][12] = (mid_1[3087:3080] < mid_1[3079:3072]) ? 1 : 0;
assign detect_min[384][13] = (mid_1[3087:3080] < mid_1[3095:3088]) ? 1 : 0;
assign detect_min[384][14] = (mid_1[3087:3080] < mid_2[3079:3072]) ? 1 : 0;
assign detect_min[384][15] = (mid_1[3087:3080] < mid_2[3087:3080]) ? 1 : 0;
assign detect_min[384][16] = (mid_1[3087:3080] < mid_2[3095:3088]) ? 1 : 0;
assign detect_min[384][17] = (mid_1[3087:3080] < btm_0[3079:3072]) ? 1 : 0;
assign detect_min[384][18] = (mid_1[3087:3080] < btm_0[3087:3080]) ? 1 : 0;
assign detect_min[384][19] = (mid_1[3087:3080] < btm_0[3095:3088]) ? 1 : 0;
assign detect_min[384][20] = (mid_1[3087:3080] < btm_1[3079:3072]) ? 1 : 0;
assign detect_min[384][21] = (mid_1[3087:3080] < btm_1[3087:3080]) ? 1 : 0;
assign detect_min[384][22] = (mid_1[3087:3080] < btm_1[3095:3088]) ? 1 : 0;
assign detect_min[384][23] = (mid_1[3087:3080] < btm_2[3079:3072]) ? 1 : 0;
assign detect_min[384][24] = (mid_1[3087:3080] < btm_2[3087:3080]) ? 1 : 0;
assign detect_min[384][25] = (mid_1[3087:3080] < btm_2[3095:3088]) ? 1 : 0;

assign detect_min[385][0] = (mid_1[3095:3088] < top_0[3087:3080]) ? 1 : 0;
assign detect_min[385][1] = (mid_1[3095:3088] < top_0[3095:3088]) ? 1 : 0;
assign detect_min[385][2] = (mid_1[3095:3088] < top_0[3103:3096]) ? 1 : 0;
assign detect_min[385][3] = (mid_1[3095:3088] < top_1[3087:3080]) ? 1 : 0;
assign detect_min[385][4] = (mid_1[3095:3088] < top_1[3095:3088]) ? 1 : 0;
assign detect_min[385][5] = (mid_1[3095:3088] < top_1[3103:3096]) ? 1 : 0;
assign detect_min[385][6] = (mid_1[3095:3088] < top_2[3087:3080]) ? 1 : 0;
assign detect_min[385][7] = (mid_1[3095:3088] < top_2[3095:3088]) ? 1 : 0;
assign detect_min[385][8] = (mid_1[3095:3088] < top_2[3103:3096]) ? 1 : 0;
assign detect_min[385][9] = (mid_1[3095:3088] < mid_0[3087:3080]) ? 1 : 0;
assign detect_min[385][10] = (mid_1[3095:3088] < mid_0[3095:3088]) ? 1 : 0;
assign detect_min[385][11] = (mid_1[3095:3088] < mid_0[3103:3096]) ? 1 : 0;
assign detect_min[385][12] = (mid_1[3095:3088] < mid_1[3087:3080]) ? 1 : 0;
assign detect_min[385][13] = (mid_1[3095:3088] < mid_1[3103:3096]) ? 1 : 0;
assign detect_min[385][14] = (mid_1[3095:3088] < mid_2[3087:3080]) ? 1 : 0;
assign detect_min[385][15] = (mid_1[3095:3088] < mid_2[3095:3088]) ? 1 : 0;
assign detect_min[385][16] = (mid_1[3095:3088] < mid_2[3103:3096]) ? 1 : 0;
assign detect_min[385][17] = (mid_1[3095:3088] < btm_0[3087:3080]) ? 1 : 0;
assign detect_min[385][18] = (mid_1[3095:3088] < btm_0[3095:3088]) ? 1 : 0;
assign detect_min[385][19] = (mid_1[3095:3088] < btm_0[3103:3096]) ? 1 : 0;
assign detect_min[385][20] = (mid_1[3095:3088] < btm_1[3087:3080]) ? 1 : 0;
assign detect_min[385][21] = (mid_1[3095:3088] < btm_1[3095:3088]) ? 1 : 0;
assign detect_min[385][22] = (mid_1[3095:3088] < btm_1[3103:3096]) ? 1 : 0;
assign detect_min[385][23] = (mid_1[3095:3088] < btm_2[3087:3080]) ? 1 : 0;
assign detect_min[385][24] = (mid_1[3095:3088] < btm_2[3095:3088]) ? 1 : 0;
assign detect_min[385][25] = (mid_1[3095:3088] < btm_2[3103:3096]) ? 1 : 0;

assign detect_min[386][0] = (mid_1[3103:3096] < top_0[3095:3088]) ? 1 : 0;
assign detect_min[386][1] = (mid_1[3103:3096] < top_0[3103:3096]) ? 1 : 0;
assign detect_min[386][2] = (mid_1[3103:3096] < top_0[3111:3104]) ? 1 : 0;
assign detect_min[386][3] = (mid_1[3103:3096] < top_1[3095:3088]) ? 1 : 0;
assign detect_min[386][4] = (mid_1[3103:3096] < top_1[3103:3096]) ? 1 : 0;
assign detect_min[386][5] = (mid_1[3103:3096] < top_1[3111:3104]) ? 1 : 0;
assign detect_min[386][6] = (mid_1[3103:3096] < top_2[3095:3088]) ? 1 : 0;
assign detect_min[386][7] = (mid_1[3103:3096] < top_2[3103:3096]) ? 1 : 0;
assign detect_min[386][8] = (mid_1[3103:3096] < top_2[3111:3104]) ? 1 : 0;
assign detect_min[386][9] = (mid_1[3103:3096] < mid_0[3095:3088]) ? 1 : 0;
assign detect_min[386][10] = (mid_1[3103:3096] < mid_0[3103:3096]) ? 1 : 0;
assign detect_min[386][11] = (mid_1[3103:3096] < mid_0[3111:3104]) ? 1 : 0;
assign detect_min[386][12] = (mid_1[3103:3096] < mid_1[3095:3088]) ? 1 : 0;
assign detect_min[386][13] = (mid_1[3103:3096] < mid_1[3111:3104]) ? 1 : 0;
assign detect_min[386][14] = (mid_1[3103:3096] < mid_2[3095:3088]) ? 1 : 0;
assign detect_min[386][15] = (mid_1[3103:3096] < mid_2[3103:3096]) ? 1 : 0;
assign detect_min[386][16] = (mid_1[3103:3096] < mid_2[3111:3104]) ? 1 : 0;
assign detect_min[386][17] = (mid_1[3103:3096] < btm_0[3095:3088]) ? 1 : 0;
assign detect_min[386][18] = (mid_1[3103:3096] < btm_0[3103:3096]) ? 1 : 0;
assign detect_min[386][19] = (mid_1[3103:3096] < btm_0[3111:3104]) ? 1 : 0;
assign detect_min[386][20] = (mid_1[3103:3096] < btm_1[3095:3088]) ? 1 : 0;
assign detect_min[386][21] = (mid_1[3103:3096] < btm_1[3103:3096]) ? 1 : 0;
assign detect_min[386][22] = (mid_1[3103:3096] < btm_1[3111:3104]) ? 1 : 0;
assign detect_min[386][23] = (mid_1[3103:3096] < btm_2[3095:3088]) ? 1 : 0;
assign detect_min[386][24] = (mid_1[3103:3096] < btm_2[3103:3096]) ? 1 : 0;
assign detect_min[386][25] = (mid_1[3103:3096] < btm_2[3111:3104]) ? 1 : 0;

assign detect_min[387][0] = (mid_1[3111:3104] < top_0[3103:3096]) ? 1 : 0;
assign detect_min[387][1] = (mid_1[3111:3104] < top_0[3111:3104]) ? 1 : 0;
assign detect_min[387][2] = (mid_1[3111:3104] < top_0[3119:3112]) ? 1 : 0;
assign detect_min[387][3] = (mid_1[3111:3104] < top_1[3103:3096]) ? 1 : 0;
assign detect_min[387][4] = (mid_1[3111:3104] < top_1[3111:3104]) ? 1 : 0;
assign detect_min[387][5] = (mid_1[3111:3104] < top_1[3119:3112]) ? 1 : 0;
assign detect_min[387][6] = (mid_1[3111:3104] < top_2[3103:3096]) ? 1 : 0;
assign detect_min[387][7] = (mid_1[3111:3104] < top_2[3111:3104]) ? 1 : 0;
assign detect_min[387][8] = (mid_1[3111:3104] < top_2[3119:3112]) ? 1 : 0;
assign detect_min[387][9] = (mid_1[3111:3104] < mid_0[3103:3096]) ? 1 : 0;
assign detect_min[387][10] = (mid_1[3111:3104] < mid_0[3111:3104]) ? 1 : 0;
assign detect_min[387][11] = (mid_1[3111:3104] < mid_0[3119:3112]) ? 1 : 0;
assign detect_min[387][12] = (mid_1[3111:3104] < mid_1[3103:3096]) ? 1 : 0;
assign detect_min[387][13] = (mid_1[3111:3104] < mid_1[3119:3112]) ? 1 : 0;
assign detect_min[387][14] = (mid_1[3111:3104] < mid_2[3103:3096]) ? 1 : 0;
assign detect_min[387][15] = (mid_1[3111:3104] < mid_2[3111:3104]) ? 1 : 0;
assign detect_min[387][16] = (mid_1[3111:3104] < mid_2[3119:3112]) ? 1 : 0;
assign detect_min[387][17] = (mid_1[3111:3104] < btm_0[3103:3096]) ? 1 : 0;
assign detect_min[387][18] = (mid_1[3111:3104] < btm_0[3111:3104]) ? 1 : 0;
assign detect_min[387][19] = (mid_1[3111:3104] < btm_0[3119:3112]) ? 1 : 0;
assign detect_min[387][20] = (mid_1[3111:3104] < btm_1[3103:3096]) ? 1 : 0;
assign detect_min[387][21] = (mid_1[3111:3104] < btm_1[3111:3104]) ? 1 : 0;
assign detect_min[387][22] = (mid_1[3111:3104] < btm_1[3119:3112]) ? 1 : 0;
assign detect_min[387][23] = (mid_1[3111:3104] < btm_2[3103:3096]) ? 1 : 0;
assign detect_min[387][24] = (mid_1[3111:3104] < btm_2[3111:3104]) ? 1 : 0;
assign detect_min[387][25] = (mid_1[3111:3104] < btm_2[3119:3112]) ? 1 : 0;

assign detect_min[388][0] = (mid_1[3119:3112] < top_0[3111:3104]) ? 1 : 0;
assign detect_min[388][1] = (mid_1[3119:3112] < top_0[3119:3112]) ? 1 : 0;
assign detect_min[388][2] = (mid_1[3119:3112] < top_0[3127:3120]) ? 1 : 0;
assign detect_min[388][3] = (mid_1[3119:3112] < top_1[3111:3104]) ? 1 : 0;
assign detect_min[388][4] = (mid_1[3119:3112] < top_1[3119:3112]) ? 1 : 0;
assign detect_min[388][5] = (mid_1[3119:3112] < top_1[3127:3120]) ? 1 : 0;
assign detect_min[388][6] = (mid_1[3119:3112] < top_2[3111:3104]) ? 1 : 0;
assign detect_min[388][7] = (mid_1[3119:3112] < top_2[3119:3112]) ? 1 : 0;
assign detect_min[388][8] = (mid_1[3119:3112] < top_2[3127:3120]) ? 1 : 0;
assign detect_min[388][9] = (mid_1[3119:3112] < mid_0[3111:3104]) ? 1 : 0;
assign detect_min[388][10] = (mid_1[3119:3112] < mid_0[3119:3112]) ? 1 : 0;
assign detect_min[388][11] = (mid_1[3119:3112] < mid_0[3127:3120]) ? 1 : 0;
assign detect_min[388][12] = (mid_1[3119:3112] < mid_1[3111:3104]) ? 1 : 0;
assign detect_min[388][13] = (mid_1[3119:3112] < mid_1[3127:3120]) ? 1 : 0;
assign detect_min[388][14] = (mid_1[3119:3112] < mid_2[3111:3104]) ? 1 : 0;
assign detect_min[388][15] = (mid_1[3119:3112] < mid_2[3119:3112]) ? 1 : 0;
assign detect_min[388][16] = (mid_1[3119:3112] < mid_2[3127:3120]) ? 1 : 0;
assign detect_min[388][17] = (mid_1[3119:3112] < btm_0[3111:3104]) ? 1 : 0;
assign detect_min[388][18] = (mid_1[3119:3112] < btm_0[3119:3112]) ? 1 : 0;
assign detect_min[388][19] = (mid_1[3119:3112] < btm_0[3127:3120]) ? 1 : 0;
assign detect_min[388][20] = (mid_1[3119:3112] < btm_1[3111:3104]) ? 1 : 0;
assign detect_min[388][21] = (mid_1[3119:3112] < btm_1[3119:3112]) ? 1 : 0;
assign detect_min[388][22] = (mid_1[3119:3112] < btm_1[3127:3120]) ? 1 : 0;
assign detect_min[388][23] = (mid_1[3119:3112] < btm_2[3111:3104]) ? 1 : 0;
assign detect_min[388][24] = (mid_1[3119:3112] < btm_2[3119:3112]) ? 1 : 0;
assign detect_min[388][25] = (mid_1[3119:3112] < btm_2[3127:3120]) ? 1 : 0;

assign detect_min[389][0] = (mid_1[3127:3120] < top_0[3119:3112]) ? 1 : 0;
assign detect_min[389][1] = (mid_1[3127:3120] < top_0[3127:3120]) ? 1 : 0;
assign detect_min[389][2] = (mid_1[3127:3120] < top_0[3135:3128]) ? 1 : 0;
assign detect_min[389][3] = (mid_1[3127:3120] < top_1[3119:3112]) ? 1 : 0;
assign detect_min[389][4] = (mid_1[3127:3120] < top_1[3127:3120]) ? 1 : 0;
assign detect_min[389][5] = (mid_1[3127:3120] < top_1[3135:3128]) ? 1 : 0;
assign detect_min[389][6] = (mid_1[3127:3120] < top_2[3119:3112]) ? 1 : 0;
assign detect_min[389][7] = (mid_1[3127:3120] < top_2[3127:3120]) ? 1 : 0;
assign detect_min[389][8] = (mid_1[3127:3120] < top_2[3135:3128]) ? 1 : 0;
assign detect_min[389][9] = (mid_1[3127:3120] < mid_0[3119:3112]) ? 1 : 0;
assign detect_min[389][10] = (mid_1[3127:3120] < mid_0[3127:3120]) ? 1 : 0;
assign detect_min[389][11] = (mid_1[3127:3120] < mid_0[3135:3128]) ? 1 : 0;
assign detect_min[389][12] = (mid_1[3127:3120] < mid_1[3119:3112]) ? 1 : 0;
assign detect_min[389][13] = (mid_1[3127:3120] < mid_1[3135:3128]) ? 1 : 0;
assign detect_min[389][14] = (mid_1[3127:3120] < mid_2[3119:3112]) ? 1 : 0;
assign detect_min[389][15] = (mid_1[3127:3120] < mid_2[3127:3120]) ? 1 : 0;
assign detect_min[389][16] = (mid_1[3127:3120] < mid_2[3135:3128]) ? 1 : 0;
assign detect_min[389][17] = (mid_1[3127:3120] < btm_0[3119:3112]) ? 1 : 0;
assign detect_min[389][18] = (mid_1[3127:3120] < btm_0[3127:3120]) ? 1 : 0;
assign detect_min[389][19] = (mid_1[3127:3120] < btm_0[3135:3128]) ? 1 : 0;
assign detect_min[389][20] = (mid_1[3127:3120] < btm_1[3119:3112]) ? 1 : 0;
assign detect_min[389][21] = (mid_1[3127:3120] < btm_1[3127:3120]) ? 1 : 0;
assign detect_min[389][22] = (mid_1[3127:3120] < btm_1[3135:3128]) ? 1 : 0;
assign detect_min[389][23] = (mid_1[3127:3120] < btm_2[3119:3112]) ? 1 : 0;
assign detect_min[389][24] = (mid_1[3127:3120] < btm_2[3127:3120]) ? 1 : 0;
assign detect_min[389][25] = (mid_1[3127:3120] < btm_2[3135:3128]) ? 1 : 0;

assign detect_min[390][0] = (mid_1[3135:3128] < top_0[3127:3120]) ? 1 : 0;
assign detect_min[390][1] = (mid_1[3135:3128] < top_0[3135:3128]) ? 1 : 0;
assign detect_min[390][2] = (mid_1[3135:3128] < top_0[3143:3136]) ? 1 : 0;
assign detect_min[390][3] = (mid_1[3135:3128] < top_1[3127:3120]) ? 1 : 0;
assign detect_min[390][4] = (mid_1[3135:3128] < top_1[3135:3128]) ? 1 : 0;
assign detect_min[390][5] = (mid_1[3135:3128] < top_1[3143:3136]) ? 1 : 0;
assign detect_min[390][6] = (mid_1[3135:3128] < top_2[3127:3120]) ? 1 : 0;
assign detect_min[390][7] = (mid_1[3135:3128] < top_2[3135:3128]) ? 1 : 0;
assign detect_min[390][8] = (mid_1[3135:3128] < top_2[3143:3136]) ? 1 : 0;
assign detect_min[390][9] = (mid_1[3135:3128] < mid_0[3127:3120]) ? 1 : 0;
assign detect_min[390][10] = (mid_1[3135:3128] < mid_0[3135:3128]) ? 1 : 0;
assign detect_min[390][11] = (mid_1[3135:3128] < mid_0[3143:3136]) ? 1 : 0;
assign detect_min[390][12] = (mid_1[3135:3128] < mid_1[3127:3120]) ? 1 : 0;
assign detect_min[390][13] = (mid_1[3135:3128] < mid_1[3143:3136]) ? 1 : 0;
assign detect_min[390][14] = (mid_1[3135:3128] < mid_2[3127:3120]) ? 1 : 0;
assign detect_min[390][15] = (mid_1[3135:3128] < mid_2[3135:3128]) ? 1 : 0;
assign detect_min[390][16] = (mid_1[3135:3128] < mid_2[3143:3136]) ? 1 : 0;
assign detect_min[390][17] = (mid_1[3135:3128] < btm_0[3127:3120]) ? 1 : 0;
assign detect_min[390][18] = (mid_1[3135:3128] < btm_0[3135:3128]) ? 1 : 0;
assign detect_min[390][19] = (mid_1[3135:3128] < btm_0[3143:3136]) ? 1 : 0;
assign detect_min[390][20] = (mid_1[3135:3128] < btm_1[3127:3120]) ? 1 : 0;
assign detect_min[390][21] = (mid_1[3135:3128] < btm_1[3135:3128]) ? 1 : 0;
assign detect_min[390][22] = (mid_1[3135:3128] < btm_1[3143:3136]) ? 1 : 0;
assign detect_min[390][23] = (mid_1[3135:3128] < btm_2[3127:3120]) ? 1 : 0;
assign detect_min[390][24] = (mid_1[3135:3128] < btm_2[3135:3128]) ? 1 : 0;
assign detect_min[390][25] = (mid_1[3135:3128] < btm_2[3143:3136]) ? 1 : 0;

assign detect_min[391][0] = (mid_1[3143:3136] < top_0[3135:3128]) ? 1 : 0;
assign detect_min[391][1] = (mid_1[3143:3136] < top_0[3143:3136]) ? 1 : 0;
assign detect_min[391][2] = (mid_1[3143:3136] < top_0[3151:3144]) ? 1 : 0;
assign detect_min[391][3] = (mid_1[3143:3136] < top_1[3135:3128]) ? 1 : 0;
assign detect_min[391][4] = (mid_1[3143:3136] < top_1[3143:3136]) ? 1 : 0;
assign detect_min[391][5] = (mid_1[3143:3136] < top_1[3151:3144]) ? 1 : 0;
assign detect_min[391][6] = (mid_1[3143:3136] < top_2[3135:3128]) ? 1 : 0;
assign detect_min[391][7] = (mid_1[3143:3136] < top_2[3143:3136]) ? 1 : 0;
assign detect_min[391][8] = (mid_1[3143:3136] < top_2[3151:3144]) ? 1 : 0;
assign detect_min[391][9] = (mid_1[3143:3136] < mid_0[3135:3128]) ? 1 : 0;
assign detect_min[391][10] = (mid_1[3143:3136] < mid_0[3143:3136]) ? 1 : 0;
assign detect_min[391][11] = (mid_1[3143:3136] < mid_0[3151:3144]) ? 1 : 0;
assign detect_min[391][12] = (mid_1[3143:3136] < mid_1[3135:3128]) ? 1 : 0;
assign detect_min[391][13] = (mid_1[3143:3136] < mid_1[3151:3144]) ? 1 : 0;
assign detect_min[391][14] = (mid_1[3143:3136] < mid_2[3135:3128]) ? 1 : 0;
assign detect_min[391][15] = (mid_1[3143:3136] < mid_2[3143:3136]) ? 1 : 0;
assign detect_min[391][16] = (mid_1[3143:3136] < mid_2[3151:3144]) ? 1 : 0;
assign detect_min[391][17] = (mid_1[3143:3136] < btm_0[3135:3128]) ? 1 : 0;
assign detect_min[391][18] = (mid_1[3143:3136] < btm_0[3143:3136]) ? 1 : 0;
assign detect_min[391][19] = (mid_1[3143:3136] < btm_0[3151:3144]) ? 1 : 0;
assign detect_min[391][20] = (mid_1[3143:3136] < btm_1[3135:3128]) ? 1 : 0;
assign detect_min[391][21] = (mid_1[3143:3136] < btm_1[3143:3136]) ? 1 : 0;
assign detect_min[391][22] = (mid_1[3143:3136] < btm_1[3151:3144]) ? 1 : 0;
assign detect_min[391][23] = (mid_1[3143:3136] < btm_2[3135:3128]) ? 1 : 0;
assign detect_min[391][24] = (mid_1[3143:3136] < btm_2[3143:3136]) ? 1 : 0;
assign detect_min[391][25] = (mid_1[3143:3136] < btm_2[3151:3144]) ? 1 : 0;

assign detect_min[392][0] = (mid_1[3151:3144] < top_0[3143:3136]) ? 1 : 0;
assign detect_min[392][1] = (mid_1[3151:3144] < top_0[3151:3144]) ? 1 : 0;
assign detect_min[392][2] = (mid_1[3151:3144] < top_0[3159:3152]) ? 1 : 0;
assign detect_min[392][3] = (mid_1[3151:3144] < top_1[3143:3136]) ? 1 : 0;
assign detect_min[392][4] = (mid_1[3151:3144] < top_1[3151:3144]) ? 1 : 0;
assign detect_min[392][5] = (mid_1[3151:3144] < top_1[3159:3152]) ? 1 : 0;
assign detect_min[392][6] = (mid_1[3151:3144] < top_2[3143:3136]) ? 1 : 0;
assign detect_min[392][7] = (mid_1[3151:3144] < top_2[3151:3144]) ? 1 : 0;
assign detect_min[392][8] = (mid_1[3151:3144] < top_2[3159:3152]) ? 1 : 0;
assign detect_min[392][9] = (mid_1[3151:3144] < mid_0[3143:3136]) ? 1 : 0;
assign detect_min[392][10] = (mid_1[3151:3144] < mid_0[3151:3144]) ? 1 : 0;
assign detect_min[392][11] = (mid_1[3151:3144] < mid_0[3159:3152]) ? 1 : 0;
assign detect_min[392][12] = (mid_1[3151:3144] < mid_1[3143:3136]) ? 1 : 0;
assign detect_min[392][13] = (mid_1[3151:3144] < mid_1[3159:3152]) ? 1 : 0;
assign detect_min[392][14] = (mid_1[3151:3144] < mid_2[3143:3136]) ? 1 : 0;
assign detect_min[392][15] = (mid_1[3151:3144] < mid_2[3151:3144]) ? 1 : 0;
assign detect_min[392][16] = (mid_1[3151:3144] < mid_2[3159:3152]) ? 1 : 0;
assign detect_min[392][17] = (mid_1[3151:3144] < btm_0[3143:3136]) ? 1 : 0;
assign detect_min[392][18] = (mid_1[3151:3144] < btm_0[3151:3144]) ? 1 : 0;
assign detect_min[392][19] = (mid_1[3151:3144] < btm_0[3159:3152]) ? 1 : 0;
assign detect_min[392][20] = (mid_1[3151:3144] < btm_1[3143:3136]) ? 1 : 0;
assign detect_min[392][21] = (mid_1[3151:3144] < btm_1[3151:3144]) ? 1 : 0;
assign detect_min[392][22] = (mid_1[3151:3144] < btm_1[3159:3152]) ? 1 : 0;
assign detect_min[392][23] = (mid_1[3151:3144] < btm_2[3143:3136]) ? 1 : 0;
assign detect_min[392][24] = (mid_1[3151:3144] < btm_2[3151:3144]) ? 1 : 0;
assign detect_min[392][25] = (mid_1[3151:3144] < btm_2[3159:3152]) ? 1 : 0;

assign detect_min[393][0] = (mid_1[3159:3152] < top_0[3151:3144]) ? 1 : 0;
assign detect_min[393][1] = (mid_1[3159:3152] < top_0[3159:3152]) ? 1 : 0;
assign detect_min[393][2] = (mid_1[3159:3152] < top_0[3167:3160]) ? 1 : 0;
assign detect_min[393][3] = (mid_1[3159:3152] < top_1[3151:3144]) ? 1 : 0;
assign detect_min[393][4] = (mid_1[3159:3152] < top_1[3159:3152]) ? 1 : 0;
assign detect_min[393][5] = (mid_1[3159:3152] < top_1[3167:3160]) ? 1 : 0;
assign detect_min[393][6] = (mid_1[3159:3152] < top_2[3151:3144]) ? 1 : 0;
assign detect_min[393][7] = (mid_1[3159:3152] < top_2[3159:3152]) ? 1 : 0;
assign detect_min[393][8] = (mid_1[3159:3152] < top_2[3167:3160]) ? 1 : 0;
assign detect_min[393][9] = (mid_1[3159:3152] < mid_0[3151:3144]) ? 1 : 0;
assign detect_min[393][10] = (mid_1[3159:3152] < mid_0[3159:3152]) ? 1 : 0;
assign detect_min[393][11] = (mid_1[3159:3152] < mid_0[3167:3160]) ? 1 : 0;
assign detect_min[393][12] = (mid_1[3159:3152] < mid_1[3151:3144]) ? 1 : 0;
assign detect_min[393][13] = (mid_1[3159:3152] < mid_1[3167:3160]) ? 1 : 0;
assign detect_min[393][14] = (mid_1[3159:3152] < mid_2[3151:3144]) ? 1 : 0;
assign detect_min[393][15] = (mid_1[3159:3152] < mid_2[3159:3152]) ? 1 : 0;
assign detect_min[393][16] = (mid_1[3159:3152] < mid_2[3167:3160]) ? 1 : 0;
assign detect_min[393][17] = (mid_1[3159:3152] < btm_0[3151:3144]) ? 1 : 0;
assign detect_min[393][18] = (mid_1[3159:3152] < btm_0[3159:3152]) ? 1 : 0;
assign detect_min[393][19] = (mid_1[3159:3152] < btm_0[3167:3160]) ? 1 : 0;
assign detect_min[393][20] = (mid_1[3159:3152] < btm_1[3151:3144]) ? 1 : 0;
assign detect_min[393][21] = (mid_1[3159:3152] < btm_1[3159:3152]) ? 1 : 0;
assign detect_min[393][22] = (mid_1[3159:3152] < btm_1[3167:3160]) ? 1 : 0;
assign detect_min[393][23] = (mid_1[3159:3152] < btm_2[3151:3144]) ? 1 : 0;
assign detect_min[393][24] = (mid_1[3159:3152] < btm_2[3159:3152]) ? 1 : 0;
assign detect_min[393][25] = (mid_1[3159:3152] < btm_2[3167:3160]) ? 1 : 0;

assign detect_min[394][0] = (mid_1[3167:3160] < top_0[3159:3152]) ? 1 : 0;
assign detect_min[394][1] = (mid_1[3167:3160] < top_0[3167:3160]) ? 1 : 0;
assign detect_min[394][2] = (mid_1[3167:3160] < top_0[3175:3168]) ? 1 : 0;
assign detect_min[394][3] = (mid_1[3167:3160] < top_1[3159:3152]) ? 1 : 0;
assign detect_min[394][4] = (mid_1[3167:3160] < top_1[3167:3160]) ? 1 : 0;
assign detect_min[394][5] = (mid_1[3167:3160] < top_1[3175:3168]) ? 1 : 0;
assign detect_min[394][6] = (mid_1[3167:3160] < top_2[3159:3152]) ? 1 : 0;
assign detect_min[394][7] = (mid_1[3167:3160] < top_2[3167:3160]) ? 1 : 0;
assign detect_min[394][8] = (mid_1[3167:3160] < top_2[3175:3168]) ? 1 : 0;
assign detect_min[394][9] = (mid_1[3167:3160] < mid_0[3159:3152]) ? 1 : 0;
assign detect_min[394][10] = (mid_1[3167:3160] < mid_0[3167:3160]) ? 1 : 0;
assign detect_min[394][11] = (mid_1[3167:3160] < mid_0[3175:3168]) ? 1 : 0;
assign detect_min[394][12] = (mid_1[3167:3160] < mid_1[3159:3152]) ? 1 : 0;
assign detect_min[394][13] = (mid_1[3167:3160] < mid_1[3175:3168]) ? 1 : 0;
assign detect_min[394][14] = (mid_1[3167:3160] < mid_2[3159:3152]) ? 1 : 0;
assign detect_min[394][15] = (mid_1[3167:3160] < mid_2[3167:3160]) ? 1 : 0;
assign detect_min[394][16] = (mid_1[3167:3160] < mid_2[3175:3168]) ? 1 : 0;
assign detect_min[394][17] = (mid_1[3167:3160] < btm_0[3159:3152]) ? 1 : 0;
assign detect_min[394][18] = (mid_1[3167:3160] < btm_0[3167:3160]) ? 1 : 0;
assign detect_min[394][19] = (mid_1[3167:3160] < btm_0[3175:3168]) ? 1 : 0;
assign detect_min[394][20] = (mid_1[3167:3160] < btm_1[3159:3152]) ? 1 : 0;
assign detect_min[394][21] = (mid_1[3167:3160] < btm_1[3167:3160]) ? 1 : 0;
assign detect_min[394][22] = (mid_1[3167:3160] < btm_1[3175:3168]) ? 1 : 0;
assign detect_min[394][23] = (mid_1[3167:3160] < btm_2[3159:3152]) ? 1 : 0;
assign detect_min[394][24] = (mid_1[3167:3160] < btm_2[3167:3160]) ? 1 : 0;
assign detect_min[394][25] = (mid_1[3167:3160] < btm_2[3175:3168]) ? 1 : 0;

assign detect_min[395][0] = (mid_1[3175:3168] < top_0[3167:3160]) ? 1 : 0;
assign detect_min[395][1] = (mid_1[3175:3168] < top_0[3175:3168]) ? 1 : 0;
assign detect_min[395][2] = (mid_1[3175:3168] < top_0[3183:3176]) ? 1 : 0;
assign detect_min[395][3] = (mid_1[3175:3168] < top_1[3167:3160]) ? 1 : 0;
assign detect_min[395][4] = (mid_1[3175:3168] < top_1[3175:3168]) ? 1 : 0;
assign detect_min[395][5] = (mid_1[3175:3168] < top_1[3183:3176]) ? 1 : 0;
assign detect_min[395][6] = (mid_1[3175:3168] < top_2[3167:3160]) ? 1 : 0;
assign detect_min[395][7] = (mid_1[3175:3168] < top_2[3175:3168]) ? 1 : 0;
assign detect_min[395][8] = (mid_1[3175:3168] < top_2[3183:3176]) ? 1 : 0;
assign detect_min[395][9] = (mid_1[3175:3168] < mid_0[3167:3160]) ? 1 : 0;
assign detect_min[395][10] = (mid_1[3175:3168] < mid_0[3175:3168]) ? 1 : 0;
assign detect_min[395][11] = (mid_1[3175:3168] < mid_0[3183:3176]) ? 1 : 0;
assign detect_min[395][12] = (mid_1[3175:3168] < mid_1[3167:3160]) ? 1 : 0;
assign detect_min[395][13] = (mid_1[3175:3168] < mid_1[3183:3176]) ? 1 : 0;
assign detect_min[395][14] = (mid_1[3175:3168] < mid_2[3167:3160]) ? 1 : 0;
assign detect_min[395][15] = (mid_1[3175:3168] < mid_2[3175:3168]) ? 1 : 0;
assign detect_min[395][16] = (mid_1[3175:3168] < mid_2[3183:3176]) ? 1 : 0;
assign detect_min[395][17] = (mid_1[3175:3168] < btm_0[3167:3160]) ? 1 : 0;
assign detect_min[395][18] = (mid_1[3175:3168] < btm_0[3175:3168]) ? 1 : 0;
assign detect_min[395][19] = (mid_1[3175:3168] < btm_0[3183:3176]) ? 1 : 0;
assign detect_min[395][20] = (mid_1[3175:3168] < btm_1[3167:3160]) ? 1 : 0;
assign detect_min[395][21] = (mid_1[3175:3168] < btm_1[3175:3168]) ? 1 : 0;
assign detect_min[395][22] = (mid_1[3175:3168] < btm_1[3183:3176]) ? 1 : 0;
assign detect_min[395][23] = (mid_1[3175:3168] < btm_2[3167:3160]) ? 1 : 0;
assign detect_min[395][24] = (mid_1[3175:3168] < btm_2[3175:3168]) ? 1 : 0;
assign detect_min[395][25] = (mid_1[3175:3168] < btm_2[3183:3176]) ? 1 : 0;

assign detect_min[396][0] = (mid_1[3183:3176] < top_0[3175:3168]) ? 1 : 0;
assign detect_min[396][1] = (mid_1[3183:3176] < top_0[3183:3176]) ? 1 : 0;
assign detect_min[396][2] = (mid_1[3183:3176] < top_0[3191:3184]) ? 1 : 0;
assign detect_min[396][3] = (mid_1[3183:3176] < top_1[3175:3168]) ? 1 : 0;
assign detect_min[396][4] = (mid_1[3183:3176] < top_1[3183:3176]) ? 1 : 0;
assign detect_min[396][5] = (mid_1[3183:3176] < top_1[3191:3184]) ? 1 : 0;
assign detect_min[396][6] = (mid_1[3183:3176] < top_2[3175:3168]) ? 1 : 0;
assign detect_min[396][7] = (mid_1[3183:3176] < top_2[3183:3176]) ? 1 : 0;
assign detect_min[396][8] = (mid_1[3183:3176] < top_2[3191:3184]) ? 1 : 0;
assign detect_min[396][9] = (mid_1[3183:3176] < mid_0[3175:3168]) ? 1 : 0;
assign detect_min[396][10] = (mid_1[3183:3176] < mid_0[3183:3176]) ? 1 : 0;
assign detect_min[396][11] = (mid_1[3183:3176] < mid_0[3191:3184]) ? 1 : 0;
assign detect_min[396][12] = (mid_1[3183:3176] < mid_1[3175:3168]) ? 1 : 0;
assign detect_min[396][13] = (mid_1[3183:3176] < mid_1[3191:3184]) ? 1 : 0;
assign detect_min[396][14] = (mid_1[3183:3176] < mid_2[3175:3168]) ? 1 : 0;
assign detect_min[396][15] = (mid_1[3183:3176] < mid_2[3183:3176]) ? 1 : 0;
assign detect_min[396][16] = (mid_1[3183:3176] < mid_2[3191:3184]) ? 1 : 0;
assign detect_min[396][17] = (mid_1[3183:3176] < btm_0[3175:3168]) ? 1 : 0;
assign detect_min[396][18] = (mid_1[3183:3176] < btm_0[3183:3176]) ? 1 : 0;
assign detect_min[396][19] = (mid_1[3183:3176] < btm_0[3191:3184]) ? 1 : 0;
assign detect_min[396][20] = (mid_1[3183:3176] < btm_1[3175:3168]) ? 1 : 0;
assign detect_min[396][21] = (mid_1[3183:3176] < btm_1[3183:3176]) ? 1 : 0;
assign detect_min[396][22] = (mid_1[3183:3176] < btm_1[3191:3184]) ? 1 : 0;
assign detect_min[396][23] = (mid_1[3183:3176] < btm_2[3175:3168]) ? 1 : 0;
assign detect_min[396][24] = (mid_1[3183:3176] < btm_2[3183:3176]) ? 1 : 0;
assign detect_min[396][25] = (mid_1[3183:3176] < btm_2[3191:3184]) ? 1 : 0;

assign detect_min[397][0] = (mid_1[3191:3184] < top_0[3183:3176]) ? 1 : 0;
assign detect_min[397][1] = (mid_1[3191:3184] < top_0[3191:3184]) ? 1 : 0;
assign detect_min[397][2] = (mid_1[3191:3184] < top_0[3199:3192]) ? 1 : 0;
assign detect_min[397][3] = (mid_1[3191:3184] < top_1[3183:3176]) ? 1 : 0;
assign detect_min[397][4] = (mid_1[3191:3184] < top_1[3191:3184]) ? 1 : 0;
assign detect_min[397][5] = (mid_1[3191:3184] < top_1[3199:3192]) ? 1 : 0;
assign detect_min[397][6] = (mid_1[3191:3184] < top_2[3183:3176]) ? 1 : 0;
assign detect_min[397][7] = (mid_1[3191:3184] < top_2[3191:3184]) ? 1 : 0;
assign detect_min[397][8] = (mid_1[3191:3184] < top_2[3199:3192]) ? 1 : 0;
assign detect_min[397][9] = (mid_1[3191:3184] < mid_0[3183:3176]) ? 1 : 0;
assign detect_min[397][10] = (mid_1[3191:3184] < mid_0[3191:3184]) ? 1 : 0;
assign detect_min[397][11] = (mid_1[3191:3184] < mid_0[3199:3192]) ? 1 : 0;
assign detect_min[397][12] = (mid_1[3191:3184] < mid_1[3183:3176]) ? 1 : 0;
assign detect_min[397][13] = (mid_1[3191:3184] < mid_1[3199:3192]) ? 1 : 0;
assign detect_min[397][14] = (mid_1[3191:3184] < mid_2[3183:3176]) ? 1 : 0;
assign detect_min[397][15] = (mid_1[3191:3184] < mid_2[3191:3184]) ? 1 : 0;
assign detect_min[397][16] = (mid_1[3191:3184] < mid_2[3199:3192]) ? 1 : 0;
assign detect_min[397][17] = (mid_1[3191:3184] < btm_0[3183:3176]) ? 1 : 0;
assign detect_min[397][18] = (mid_1[3191:3184] < btm_0[3191:3184]) ? 1 : 0;
assign detect_min[397][19] = (mid_1[3191:3184] < btm_0[3199:3192]) ? 1 : 0;
assign detect_min[397][20] = (mid_1[3191:3184] < btm_1[3183:3176]) ? 1 : 0;
assign detect_min[397][21] = (mid_1[3191:3184] < btm_1[3191:3184]) ? 1 : 0;
assign detect_min[397][22] = (mid_1[3191:3184] < btm_1[3199:3192]) ? 1 : 0;
assign detect_min[397][23] = (mid_1[3191:3184] < btm_2[3183:3176]) ? 1 : 0;
assign detect_min[397][24] = (mid_1[3191:3184] < btm_2[3191:3184]) ? 1 : 0;
assign detect_min[397][25] = (mid_1[3191:3184] < btm_2[3199:3192]) ? 1 : 0;

assign detect_min[398][0] = (mid_1[3199:3192] < top_0[3191:3184]) ? 1 : 0;
assign detect_min[398][1] = (mid_1[3199:3192] < top_0[3199:3192]) ? 1 : 0;
assign detect_min[398][2] = (mid_1[3199:3192] < top_0[3207:3200]) ? 1 : 0;
assign detect_min[398][3] = (mid_1[3199:3192] < top_1[3191:3184]) ? 1 : 0;
assign detect_min[398][4] = (mid_1[3199:3192] < top_1[3199:3192]) ? 1 : 0;
assign detect_min[398][5] = (mid_1[3199:3192] < top_1[3207:3200]) ? 1 : 0;
assign detect_min[398][6] = (mid_1[3199:3192] < top_2[3191:3184]) ? 1 : 0;
assign detect_min[398][7] = (mid_1[3199:3192] < top_2[3199:3192]) ? 1 : 0;
assign detect_min[398][8] = (mid_1[3199:3192] < top_2[3207:3200]) ? 1 : 0;
assign detect_min[398][9] = (mid_1[3199:3192] < mid_0[3191:3184]) ? 1 : 0;
assign detect_min[398][10] = (mid_1[3199:3192] < mid_0[3199:3192]) ? 1 : 0;
assign detect_min[398][11] = (mid_1[3199:3192] < mid_0[3207:3200]) ? 1 : 0;
assign detect_min[398][12] = (mid_1[3199:3192] < mid_1[3191:3184]) ? 1 : 0;
assign detect_min[398][13] = (mid_1[3199:3192] < mid_1[3207:3200]) ? 1 : 0;
assign detect_min[398][14] = (mid_1[3199:3192] < mid_2[3191:3184]) ? 1 : 0;
assign detect_min[398][15] = (mid_1[3199:3192] < mid_2[3199:3192]) ? 1 : 0;
assign detect_min[398][16] = (mid_1[3199:3192] < mid_2[3207:3200]) ? 1 : 0;
assign detect_min[398][17] = (mid_1[3199:3192] < btm_0[3191:3184]) ? 1 : 0;
assign detect_min[398][18] = (mid_1[3199:3192] < btm_0[3199:3192]) ? 1 : 0;
assign detect_min[398][19] = (mid_1[3199:3192] < btm_0[3207:3200]) ? 1 : 0;
assign detect_min[398][20] = (mid_1[3199:3192] < btm_1[3191:3184]) ? 1 : 0;
assign detect_min[398][21] = (mid_1[3199:3192] < btm_1[3199:3192]) ? 1 : 0;
assign detect_min[398][22] = (mid_1[3199:3192] < btm_1[3207:3200]) ? 1 : 0;
assign detect_min[398][23] = (mid_1[3199:3192] < btm_2[3191:3184]) ? 1 : 0;
assign detect_min[398][24] = (mid_1[3199:3192] < btm_2[3199:3192]) ? 1 : 0;
assign detect_min[398][25] = (mid_1[3199:3192] < btm_2[3207:3200]) ? 1 : 0;

assign detect_min[399][0] = (mid_1[3207:3200] < top_0[3199:3192]) ? 1 : 0;
assign detect_min[399][1] = (mid_1[3207:3200] < top_0[3207:3200]) ? 1 : 0;
assign detect_min[399][2] = (mid_1[3207:3200] < top_0[3215:3208]) ? 1 : 0;
assign detect_min[399][3] = (mid_1[3207:3200] < top_1[3199:3192]) ? 1 : 0;
assign detect_min[399][4] = (mid_1[3207:3200] < top_1[3207:3200]) ? 1 : 0;
assign detect_min[399][5] = (mid_1[3207:3200] < top_1[3215:3208]) ? 1 : 0;
assign detect_min[399][6] = (mid_1[3207:3200] < top_2[3199:3192]) ? 1 : 0;
assign detect_min[399][7] = (mid_1[3207:3200] < top_2[3207:3200]) ? 1 : 0;
assign detect_min[399][8] = (mid_1[3207:3200] < top_2[3215:3208]) ? 1 : 0;
assign detect_min[399][9] = (mid_1[3207:3200] < mid_0[3199:3192]) ? 1 : 0;
assign detect_min[399][10] = (mid_1[3207:3200] < mid_0[3207:3200]) ? 1 : 0;
assign detect_min[399][11] = (mid_1[3207:3200] < mid_0[3215:3208]) ? 1 : 0;
assign detect_min[399][12] = (mid_1[3207:3200] < mid_1[3199:3192]) ? 1 : 0;
assign detect_min[399][13] = (mid_1[3207:3200] < mid_1[3215:3208]) ? 1 : 0;
assign detect_min[399][14] = (mid_1[3207:3200] < mid_2[3199:3192]) ? 1 : 0;
assign detect_min[399][15] = (mid_1[3207:3200] < mid_2[3207:3200]) ? 1 : 0;
assign detect_min[399][16] = (mid_1[3207:3200] < mid_2[3215:3208]) ? 1 : 0;
assign detect_min[399][17] = (mid_1[3207:3200] < btm_0[3199:3192]) ? 1 : 0;
assign detect_min[399][18] = (mid_1[3207:3200] < btm_0[3207:3200]) ? 1 : 0;
assign detect_min[399][19] = (mid_1[3207:3200] < btm_0[3215:3208]) ? 1 : 0;
assign detect_min[399][20] = (mid_1[3207:3200] < btm_1[3199:3192]) ? 1 : 0;
assign detect_min[399][21] = (mid_1[3207:3200] < btm_1[3207:3200]) ? 1 : 0;
assign detect_min[399][22] = (mid_1[3207:3200] < btm_1[3215:3208]) ? 1 : 0;
assign detect_min[399][23] = (mid_1[3207:3200] < btm_2[3199:3192]) ? 1 : 0;
assign detect_min[399][24] = (mid_1[3207:3200] < btm_2[3207:3200]) ? 1 : 0;
assign detect_min[399][25] = (mid_1[3207:3200] < btm_2[3215:3208]) ? 1 : 0;

assign detect_min[400][0] = (mid_1[3215:3208] < top_0[3207:3200]) ? 1 : 0;
assign detect_min[400][1] = (mid_1[3215:3208] < top_0[3215:3208]) ? 1 : 0;
assign detect_min[400][2] = (mid_1[3215:3208] < top_0[3223:3216]) ? 1 : 0;
assign detect_min[400][3] = (mid_1[3215:3208] < top_1[3207:3200]) ? 1 : 0;
assign detect_min[400][4] = (mid_1[3215:3208] < top_1[3215:3208]) ? 1 : 0;
assign detect_min[400][5] = (mid_1[3215:3208] < top_1[3223:3216]) ? 1 : 0;
assign detect_min[400][6] = (mid_1[3215:3208] < top_2[3207:3200]) ? 1 : 0;
assign detect_min[400][7] = (mid_1[3215:3208] < top_2[3215:3208]) ? 1 : 0;
assign detect_min[400][8] = (mid_1[3215:3208] < top_2[3223:3216]) ? 1 : 0;
assign detect_min[400][9] = (mid_1[3215:3208] < mid_0[3207:3200]) ? 1 : 0;
assign detect_min[400][10] = (mid_1[3215:3208] < mid_0[3215:3208]) ? 1 : 0;
assign detect_min[400][11] = (mid_1[3215:3208] < mid_0[3223:3216]) ? 1 : 0;
assign detect_min[400][12] = (mid_1[3215:3208] < mid_1[3207:3200]) ? 1 : 0;
assign detect_min[400][13] = (mid_1[3215:3208] < mid_1[3223:3216]) ? 1 : 0;
assign detect_min[400][14] = (mid_1[3215:3208] < mid_2[3207:3200]) ? 1 : 0;
assign detect_min[400][15] = (mid_1[3215:3208] < mid_2[3215:3208]) ? 1 : 0;
assign detect_min[400][16] = (mid_1[3215:3208] < mid_2[3223:3216]) ? 1 : 0;
assign detect_min[400][17] = (mid_1[3215:3208] < btm_0[3207:3200]) ? 1 : 0;
assign detect_min[400][18] = (mid_1[3215:3208] < btm_0[3215:3208]) ? 1 : 0;
assign detect_min[400][19] = (mid_1[3215:3208] < btm_0[3223:3216]) ? 1 : 0;
assign detect_min[400][20] = (mid_1[3215:3208] < btm_1[3207:3200]) ? 1 : 0;
assign detect_min[400][21] = (mid_1[3215:3208] < btm_1[3215:3208]) ? 1 : 0;
assign detect_min[400][22] = (mid_1[3215:3208] < btm_1[3223:3216]) ? 1 : 0;
assign detect_min[400][23] = (mid_1[3215:3208] < btm_2[3207:3200]) ? 1 : 0;
assign detect_min[400][24] = (mid_1[3215:3208] < btm_2[3215:3208]) ? 1 : 0;
assign detect_min[400][25] = (mid_1[3215:3208] < btm_2[3223:3216]) ? 1 : 0;

assign detect_min[401][0] = (mid_1[3223:3216] < top_0[3215:3208]) ? 1 : 0;
assign detect_min[401][1] = (mid_1[3223:3216] < top_0[3223:3216]) ? 1 : 0;
assign detect_min[401][2] = (mid_1[3223:3216] < top_0[3231:3224]) ? 1 : 0;
assign detect_min[401][3] = (mid_1[3223:3216] < top_1[3215:3208]) ? 1 : 0;
assign detect_min[401][4] = (mid_1[3223:3216] < top_1[3223:3216]) ? 1 : 0;
assign detect_min[401][5] = (mid_1[3223:3216] < top_1[3231:3224]) ? 1 : 0;
assign detect_min[401][6] = (mid_1[3223:3216] < top_2[3215:3208]) ? 1 : 0;
assign detect_min[401][7] = (mid_1[3223:3216] < top_2[3223:3216]) ? 1 : 0;
assign detect_min[401][8] = (mid_1[3223:3216] < top_2[3231:3224]) ? 1 : 0;
assign detect_min[401][9] = (mid_1[3223:3216] < mid_0[3215:3208]) ? 1 : 0;
assign detect_min[401][10] = (mid_1[3223:3216] < mid_0[3223:3216]) ? 1 : 0;
assign detect_min[401][11] = (mid_1[3223:3216] < mid_0[3231:3224]) ? 1 : 0;
assign detect_min[401][12] = (mid_1[3223:3216] < mid_1[3215:3208]) ? 1 : 0;
assign detect_min[401][13] = (mid_1[3223:3216] < mid_1[3231:3224]) ? 1 : 0;
assign detect_min[401][14] = (mid_1[3223:3216] < mid_2[3215:3208]) ? 1 : 0;
assign detect_min[401][15] = (mid_1[3223:3216] < mid_2[3223:3216]) ? 1 : 0;
assign detect_min[401][16] = (mid_1[3223:3216] < mid_2[3231:3224]) ? 1 : 0;
assign detect_min[401][17] = (mid_1[3223:3216] < btm_0[3215:3208]) ? 1 : 0;
assign detect_min[401][18] = (mid_1[3223:3216] < btm_0[3223:3216]) ? 1 : 0;
assign detect_min[401][19] = (mid_1[3223:3216] < btm_0[3231:3224]) ? 1 : 0;
assign detect_min[401][20] = (mid_1[3223:3216] < btm_1[3215:3208]) ? 1 : 0;
assign detect_min[401][21] = (mid_1[3223:3216] < btm_1[3223:3216]) ? 1 : 0;
assign detect_min[401][22] = (mid_1[3223:3216] < btm_1[3231:3224]) ? 1 : 0;
assign detect_min[401][23] = (mid_1[3223:3216] < btm_2[3215:3208]) ? 1 : 0;
assign detect_min[401][24] = (mid_1[3223:3216] < btm_2[3223:3216]) ? 1 : 0;
assign detect_min[401][25] = (mid_1[3223:3216] < btm_2[3231:3224]) ? 1 : 0;

assign detect_min[402][0] = (mid_1[3231:3224] < top_0[3223:3216]) ? 1 : 0;
assign detect_min[402][1] = (mid_1[3231:3224] < top_0[3231:3224]) ? 1 : 0;
assign detect_min[402][2] = (mid_1[3231:3224] < top_0[3239:3232]) ? 1 : 0;
assign detect_min[402][3] = (mid_1[3231:3224] < top_1[3223:3216]) ? 1 : 0;
assign detect_min[402][4] = (mid_1[3231:3224] < top_1[3231:3224]) ? 1 : 0;
assign detect_min[402][5] = (mid_1[3231:3224] < top_1[3239:3232]) ? 1 : 0;
assign detect_min[402][6] = (mid_1[3231:3224] < top_2[3223:3216]) ? 1 : 0;
assign detect_min[402][7] = (mid_1[3231:3224] < top_2[3231:3224]) ? 1 : 0;
assign detect_min[402][8] = (mid_1[3231:3224] < top_2[3239:3232]) ? 1 : 0;
assign detect_min[402][9] = (mid_1[3231:3224] < mid_0[3223:3216]) ? 1 : 0;
assign detect_min[402][10] = (mid_1[3231:3224] < mid_0[3231:3224]) ? 1 : 0;
assign detect_min[402][11] = (mid_1[3231:3224] < mid_0[3239:3232]) ? 1 : 0;
assign detect_min[402][12] = (mid_1[3231:3224] < mid_1[3223:3216]) ? 1 : 0;
assign detect_min[402][13] = (mid_1[3231:3224] < mid_1[3239:3232]) ? 1 : 0;
assign detect_min[402][14] = (mid_1[3231:3224] < mid_2[3223:3216]) ? 1 : 0;
assign detect_min[402][15] = (mid_1[3231:3224] < mid_2[3231:3224]) ? 1 : 0;
assign detect_min[402][16] = (mid_1[3231:3224] < mid_2[3239:3232]) ? 1 : 0;
assign detect_min[402][17] = (mid_1[3231:3224] < btm_0[3223:3216]) ? 1 : 0;
assign detect_min[402][18] = (mid_1[3231:3224] < btm_0[3231:3224]) ? 1 : 0;
assign detect_min[402][19] = (mid_1[3231:3224] < btm_0[3239:3232]) ? 1 : 0;
assign detect_min[402][20] = (mid_1[3231:3224] < btm_1[3223:3216]) ? 1 : 0;
assign detect_min[402][21] = (mid_1[3231:3224] < btm_1[3231:3224]) ? 1 : 0;
assign detect_min[402][22] = (mid_1[3231:3224] < btm_1[3239:3232]) ? 1 : 0;
assign detect_min[402][23] = (mid_1[3231:3224] < btm_2[3223:3216]) ? 1 : 0;
assign detect_min[402][24] = (mid_1[3231:3224] < btm_2[3231:3224]) ? 1 : 0;
assign detect_min[402][25] = (mid_1[3231:3224] < btm_2[3239:3232]) ? 1 : 0;

assign detect_min[403][0] = (mid_1[3239:3232] < top_0[3231:3224]) ? 1 : 0;
assign detect_min[403][1] = (mid_1[3239:3232] < top_0[3239:3232]) ? 1 : 0;
assign detect_min[403][2] = (mid_1[3239:3232] < top_0[3247:3240]) ? 1 : 0;
assign detect_min[403][3] = (mid_1[3239:3232] < top_1[3231:3224]) ? 1 : 0;
assign detect_min[403][4] = (mid_1[3239:3232] < top_1[3239:3232]) ? 1 : 0;
assign detect_min[403][5] = (mid_1[3239:3232] < top_1[3247:3240]) ? 1 : 0;
assign detect_min[403][6] = (mid_1[3239:3232] < top_2[3231:3224]) ? 1 : 0;
assign detect_min[403][7] = (mid_1[3239:3232] < top_2[3239:3232]) ? 1 : 0;
assign detect_min[403][8] = (mid_1[3239:3232] < top_2[3247:3240]) ? 1 : 0;
assign detect_min[403][9] = (mid_1[3239:3232] < mid_0[3231:3224]) ? 1 : 0;
assign detect_min[403][10] = (mid_1[3239:3232] < mid_0[3239:3232]) ? 1 : 0;
assign detect_min[403][11] = (mid_1[3239:3232] < mid_0[3247:3240]) ? 1 : 0;
assign detect_min[403][12] = (mid_1[3239:3232] < mid_1[3231:3224]) ? 1 : 0;
assign detect_min[403][13] = (mid_1[3239:3232] < mid_1[3247:3240]) ? 1 : 0;
assign detect_min[403][14] = (mid_1[3239:3232] < mid_2[3231:3224]) ? 1 : 0;
assign detect_min[403][15] = (mid_1[3239:3232] < mid_2[3239:3232]) ? 1 : 0;
assign detect_min[403][16] = (mid_1[3239:3232] < mid_2[3247:3240]) ? 1 : 0;
assign detect_min[403][17] = (mid_1[3239:3232] < btm_0[3231:3224]) ? 1 : 0;
assign detect_min[403][18] = (mid_1[3239:3232] < btm_0[3239:3232]) ? 1 : 0;
assign detect_min[403][19] = (mid_1[3239:3232] < btm_0[3247:3240]) ? 1 : 0;
assign detect_min[403][20] = (mid_1[3239:3232] < btm_1[3231:3224]) ? 1 : 0;
assign detect_min[403][21] = (mid_1[3239:3232] < btm_1[3239:3232]) ? 1 : 0;
assign detect_min[403][22] = (mid_1[3239:3232] < btm_1[3247:3240]) ? 1 : 0;
assign detect_min[403][23] = (mid_1[3239:3232] < btm_2[3231:3224]) ? 1 : 0;
assign detect_min[403][24] = (mid_1[3239:3232] < btm_2[3239:3232]) ? 1 : 0;
assign detect_min[403][25] = (mid_1[3239:3232] < btm_2[3247:3240]) ? 1 : 0;

assign detect_min[404][0] = (mid_1[3247:3240] < top_0[3239:3232]) ? 1 : 0;
assign detect_min[404][1] = (mid_1[3247:3240] < top_0[3247:3240]) ? 1 : 0;
assign detect_min[404][2] = (mid_1[3247:3240] < top_0[3255:3248]) ? 1 : 0;
assign detect_min[404][3] = (mid_1[3247:3240] < top_1[3239:3232]) ? 1 : 0;
assign detect_min[404][4] = (mid_1[3247:3240] < top_1[3247:3240]) ? 1 : 0;
assign detect_min[404][5] = (mid_1[3247:3240] < top_1[3255:3248]) ? 1 : 0;
assign detect_min[404][6] = (mid_1[3247:3240] < top_2[3239:3232]) ? 1 : 0;
assign detect_min[404][7] = (mid_1[3247:3240] < top_2[3247:3240]) ? 1 : 0;
assign detect_min[404][8] = (mid_1[3247:3240] < top_2[3255:3248]) ? 1 : 0;
assign detect_min[404][9] = (mid_1[3247:3240] < mid_0[3239:3232]) ? 1 : 0;
assign detect_min[404][10] = (mid_1[3247:3240] < mid_0[3247:3240]) ? 1 : 0;
assign detect_min[404][11] = (mid_1[3247:3240] < mid_0[3255:3248]) ? 1 : 0;
assign detect_min[404][12] = (mid_1[3247:3240] < mid_1[3239:3232]) ? 1 : 0;
assign detect_min[404][13] = (mid_1[3247:3240] < mid_1[3255:3248]) ? 1 : 0;
assign detect_min[404][14] = (mid_1[3247:3240] < mid_2[3239:3232]) ? 1 : 0;
assign detect_min[404][15] = (mid_1[3247:3240] < mid_2[3247:3240]) ? 1 : 0;
assign detect_min[404][16] = (mid_1[3247:3240] < mid_2[3255:3248]) ? 1 : 0;
assign detect_min[404][17] = (mid_1[3247:3240] < btm_0[3239:3232]) ? 1 : 0;
assign detect_min[404][18] = (mid_1[3247:3240] < btm_0[3247:3240]) ? 1 : 0;
assign detect_min[404][19] = (mid_1[3247:3240] < btm_0[3255:3248]) ? 1 : 0;
assign detect_min[404][20] = (mid_1[3247:3240] < btm_1[3239:3232]) ? 1 : 0;
assign detect_min[404][21] = (mid_1[3247:3240] < btm_1[3247:3240]) ? 1 : 0;
assign detect_min[404][22] = (mid_1[3247:3240] < btm_1[3255:3248]) ? 1 : 0;
assign detect_min[404][23] = (mid_1[3247:3240] < btm_2[3239:3232]) ? 1 : 0;
assign detect_min[404][24] = (mid_1[3247:3240] < btm_2[3247:3240]) ? 1 : 0;
assign detect_min[404][25] = (mid_1[3247:3240] < btm_2[3255:3248]) ? 1 : 0;

assign detect_min[405][0] = (mid_1[3255:3248] < top_0[3247:3240]) ? 1 : 0;
assign detect_min[405][1] = (mid_1[3255:3248] < top_0[3255:3248]) ? 1 : 0;
assign detect_min[405][2] = (mid_1[3255:3248] < top_0[3263:3256]) ? 1 : 0;
assign detect_min[405][3] = (mid_1[3255:3248] < top_1[3247:3240]) ? 1 : 0;
assign detect_min[405][4] = (mid_1[3255:3248] < top_1[3255:3248]) ? 1 : 0;
assign detect_min[405][5] = (mid_1[3255:3248] < top_1[3263:3256]) ? 1 : 0;
assign detect_min[405][6] = (mid_1[3255:3248] < top_2[3247:3240]) ? 1 : 0;
assign detect_min[405][7] = (mid_1[3255:3248] < top_2[3255:3248]) ? 1 : 0;
assign detect_min[405][8] = (mid_1[3255:3248] < top_2[3263:3256]) ? 1 : 0;
assign detect_min[405][9] = (mid_1[3255:3248] < mid_0[3247:3240]) ? 1 : 0;
assign detect_min[405][10] = (mid_1[3255:3248] < mid_0[3255:3248]) ? 1 : 0;
assign detect_min[405][11] = (mid_1[3255:3248] < mid_0[3263:3256]) ? 1 : 0;
assign detect_min[405][12] = (mid_1[3255:3248] < mid_1[3247:3240]) ? 1 : 0;
assign detect_min[405][13] = (mid_1[3255:3248] < mid_1[3263:3256]) ? 1 : 0;
assign detect_min[405][14] = (mid_1[3255:3248] < mid_2[3247:3240]) ? 1 : 0;
assign detect_min[405][15] = (mid_1[3255:3248] < mid_2[3255:3248]) ? 1 : 0;
assign detect_min[405][16] = (mid_1[3255:3248] < mid_2[3263:3256]) ? 1 : 0;
assign detect_min[405][17] = (mid_1[3255:3248] < btm_0[3247:3240]) ? 1 : 0;
assign detect_min[405][18] = (mid_1[3255:3248] < btm_0[3255:3248]) ? 1 : 0;
assign detect_min[405][19] = (mid_1[3255:3248] < btm_0[3263:3256]) ? 1 : 0;
assign detect_min[405][20] = (mid_1[3255:3248] < btm_1[3247:3240]) ? 1 : 0;
assign detect_min[405][21] = (mid_1[3255:3248] < btm_1[3255:3248]) ? 1 : 0;
assign detect_min[405][22] = (mid_1[3255:3248] < btm_1[3263:3256]) ? 1 : 0;
assign detect_min[405][23] = (mid_1[3255:3248] < btm_2[3247:3240]) ? 1 : 0;
assign detect_min[405][24] = (mid_1[3255:3248] < btm_2[3255:3248]) ? 1 : 0;
assign detect_min[405][25] = (mid_1[3255:3248] < btm_2[3263:3256]) ? 1 : 0;

assign detect_min[406][0] = (mid_1[3263:3256] < top_0[3255:3248]) ? 1 : 0;
assign detect_min[406][1] = (mid_1[3263:3256] < top_0[3263:3256]) ? 1 : 0;
assign detect_min[406][2] = (mid_1[3263:3256] < top_0[3271:3264]) ? 1 : 0;
assign detect_min[406][3] = (mid_1[3263:3256] < top_1[3255:3248]) ? 1 : 0;
assign detect_min[406][4] = (mid_1[3263:3256] < top_1[3263:3256]) ? 1 : 0;
assign detect_min[406][5] = (mid_1[3263:3256] < top_1[3271:3264]) ? 1 : 0;
assign detect_min[406][6] = (mid_1[3263:3256] < top_2[3255:3248]) ? 1 : 0;
assign detect_min[406][7] = (mid_1[3263:3256] < top_2[3263:3256]) ? 1 : 0;
assign detect_min[406][8] = (mid_1[3263:3256] < top_2[3271:3264]) ? 1 : 0;
assign detect_min[406][9] = (mid_1[3263:3256] < mid_0[3255:3248]) ? 1 : 0;
assign detect_min[406][10] = (mid_1[3263:3256] < mid_0[3263:3256]) ? 1 : 0;
assign detect_min[406][11] = (mid_1[3263:3256] < mid_0[3271:3264]) ? 1 : 0;
assign detect_min[406][12] = (mid_1[3263:3256] < mid_1[3255:3248]) ? 1 : 0;
assign detect_min[406][13] = (mid_1[3263:3256] < mid_1[3271:3264]) ? 1 : 0;
assign detect_min[406][14] = (mid_1[3263:3256] < mid_2[3255:3248]) ? 1 : 0;
assign detect_min[406][15] = (mid_1[3263:3256] < mid_2[3263:3256]) ? 1 : 0;
assign detect_min[406][16] = (mid_1[3263:3256] < mid_2[3271:3264]) ? 1 : 0;
assign detect_min[406][17] = (mid_1[3263:3256] < btm_0[3255:3248]) ? 1 : 0;
assign detect_min[406][18] = (mid_1[3263:3256] < btm_0[3263:3256]) ? 1 : 0;
assign detect_min[406][19] = (mid_1[3263:3256] < btm_0[3271:3264]) ? 1 : 0;
assign detect_min[406][20] = (mid_1[3263:3256] < btm_1[3255:3248]) ? 1 : 0;
assign detect_min[406][21] = (mid_1[3263:3256] < btm_1[3263:3256]) ? 1 : 0;
assign detect_min[406][22] = (mid_1[3263:3256] < btm_1[3271:3264]) ? 1 : 0;
assign detect_min[406][23] = (mid_1[3263:3256] < btm_2[3255:3248]) ? 1 : 0;
assign detect_min[406][24] = (mid_1[3263:3256] < btm_2[3263:3256]) ? 1 : 0;
assign detect_min[406][25] = (mid_1[3263:3256] < btm_2[3271:3264]) ? 1 : 0;

assign detect_min[407][0] = (mid_1[3271:3264] < top_0[3263:3256]) ? 1 : 0;
assign detect_min[407][1] = (mid_1[3271:3264] < top_0[3271:3264]) ? 1 : 0;
assign detect_min[407][2] = (mid_1[3271:3264] < top_0[3279:3272]) ? 1 : 0;
assign detect_min[407][3] = (mid_1[3271:3264] < top_1[3263:3256]) ? 1 : 0;
assign detect_min[407][4] = (mid_1[3271:3264] < top_1[3271:3264]) ? 1 : 0;
assign detect_min[407][5] = (mid_1[3271:3264] < top_1[3279:3272]) ? 1 : 0;
assign detect_min[407][6] = (mid_1[3271:3264] < top_2[3263:3256]) ? 1 : 0;
assign detect_min[407][7] = (mid_1[3271:3264] < top_2[3271:3264]) ? 1 : 0;
assign detect_min[407][8] = (mid_1[3271:3264] < top_2[3279:3272]) ? 1 : 0;
assign detect_min[407][9] = (mid_1[3271:3264] < mid_0[3263:3256]) ? 1 : 0;
assign detect_min[407][10] = (mid_1[3271:3264] < mid_0[3271:3264]) ? 1 : 0;
assign detect_min[407][11] = (mid_1[3271:3264] < mid_0[3279:3272]) ? 1 : 0;
assign detect_min[407][12] = (mid_1[3271:3264] < mid_1[3263:3256]) ? 1 : 0;
assign detect_min[407][13] = (mid_1[3271:3264] < mid_1[3279:3272]) ? 1 : 0;
assign detect_min[407][14] = (mid_1[3271:3264] < mid_2[3263:3256]) ? 1 : 0;
assign detect_min[407][15] = (mid_1[3271:3264] < mid_2[3271:3264]) ? 1 : 0;
assign detect_min[407][16] = (mid_1[3271:3264] < mid_2[3279:3272]) ? 1 : 0;
assign detect_min[407][17] = (mid_1[3271:3264] < btm_0[3263:3256]) ? 1 : 0;
assign detect_min[407][18] = (mid_1[3271:3264] < btm_0[3271:3264]) ? 1 : 0;
assign detect_min[407][19] = (mid_1[3271:3264] < btm_0[3279:3272]) ? 1 : 0;
assign detect_min[407][20] = (mid_1[3271:3264] < btm_1[3263:3256]) ? 1 : 0;
assign detect_min[407][21] = (mid_1[3271:3264] < btm_1[3271:3264]) ? 1 : 0;
assign detect_min[407][22] = (mid_1[3271:3264] < btm_1[3279:3272]) ? 1 : 0;
assign detect_min[407][23] = (mid_1[3271:3264] < btm_2[3263:3256]) ? 1 : 0;
assign detect_min[407][24] = (mid_1[3271:3264] < btm_2[3271:3264]) ? 1 : 0;
assign detect_min[407][25] = (mid_1[3271:3264] < btm_2[3279:3272]) ? 1 : 0;

assign detect_min[408][0] = (mid_1[3279:3272] < top_0[3271:3264]) ? 1 : 0;
assign detect_min[408][1] = (mid_1[3279:3272] < top_0[3279:3272]) ? 1 : 0;
assign detect_min[408][2] = (mid_1[3279:3272] < top_0[3287:3280]) ? 1 : 0;
assign detect_min[408][3] = (mid_1[3279:3272] < top_1[3271:3264]) ? 1 : 0;
assign detect_min[408][4] = (mid_1[3279:3272] < top_1[3279:3272]) ? 1 : 0;
assign detect_min[408][5] = (mid_1[3279:3272] < top_1[3287:3280]) ? 1 : 0;
assign detect_min[408][6] = (mid_1[3279:3272] < top_2[3271:3264]) ? 1 : 0;
assign detect_min[408][7] = (mid_1[3279:3272] < top_2[3279:3272]) ? 1 : 0;
assign detect_min[408][8] = (mid_1[3279:3272] < top_2[3287:3280]) ? 1 : 0;
assign detect_min[408][9] = (mid_1[3279:3272] < mid_0[3271:3264]) ? 1 : 0;
assign detect_min[408][10] = (mid_1[3279:3272] < mid_0[3279:3272]) ? 1 : 0;
assign detect_min[408][11] = (mid_1[3279:3272] < mid_0[3287:3280]) ? 1 : 0;
assign detect_min[408][12] = (mid_1[3279:3272] < mid_1[3271:3264]) ? 1 : 0;
assign detect_min[408][13] = (mid_1[3279:3272] < mid_1[3287:3280]) ? 1 : 0;
assign detect_min[408][14] = (mid_1[3279:3272] < mid_2[3271:3264]) ? 1 : 0;
assign detect_min[408][15] = (mid_1[3279:3272] < mid_2[3279:3272]) ? 1 : 0;
assign detect_min[408][16] = (mid_1[3279:3272] < mid_2[3287:3280]) ? 1 : 0;
assign detect_min[408][17] = (mid_1[3279:3272] < btm_0[3271:3264]) ? 1 : 0;
assign detect_min[408][18] = (mid_1[3279:3272] < btm_0[3279:3272]) ? 1 : 0;
assign detect_min[408][19] = (mid_1[3279:3272] < btm_0[3287:3280]) ? 1 : 0;
assign detect_min[408][20] = (mid_1[3279:3272] < btm_1[3271:3264]) ? 1 : 0;
assign detect_min[408][21] = (mid_1[3279:3272] < btm_1[3279:3272]) ? 1 : 0;
assign detect_min[408][22] = (mid_1[3279:3272] < btm_1[3287:3280]) ? 1 : 0;
assign detect_min[408][23] = (mid_1[3279:3272] < btm_2[3271:3264]) ? 1 : 0;
assign detect_min[408][24] = (mid_1[3279:3272] < btm_2[3279:3272]) ? 1 : 0;
assign detect_min[408][25] = (mid_1[3279:3272] < btm_2[3287:3280]) ? 1 : 0;

assign detect_min[409][0] = (mid_1[3287:3280] < top_0[3279:3272]) ? 1 : 0;
assign detect_min[409][1] = (mid_1[3287:3280] < top_0[3287:3280]) ? 1 : 0;
assign detect_min[409][2] = (mid_1[3287:3280] < top_0[3295:3288]) ? 1 : 0;
assign detect_min[409][3] = (mid_1[3287:3280] < top_1[3279:3272]) ? 1 : 0;
assign detect_min[409][4] = (mid_1[3287:3280] < top_1[3287:3280]) ? 1 : 0;
assign detect_min[409][5] = (mid_1[3287:3280] < top_1[3295:3288]) ? 1 : 0;
assign detect_min[409][6] = (mid_1[3287:3280] < top_2[3279:3272]) ? 1 : 0;
assign detect_min[409][7] = (mid_1[3287:3280] < top_2[3287:3280]) ? 1 : 0;
assign detect_min[409][8] = (mid_1[3287:3280] < top_2[3295:3288]) ? 1 : 0;
assign detect_min[409][9] = (mid_1[3287:3280] < mid_0[3279:3272]) ? 1 : 0;
assign detect_min[409][10] = (mid_1[3287:3280] < mid_0[3287:3280]) ? 1 : 0;
assign detect_min[409][11] = (mid_1[3287:3280] < mid_0[3295:3288]) ? 1 : 0;
assign detect_min[409][12] = (mid_1[3287:3280] < mid_1[3279:3272]) ? 1 : 0;
assign detect_min[409][13] = (mid_1[3287:3280] < mid_1[3295:3288]) ? 1 : 0;
assign detect_min[409][14] = (mid_1[3287:3280] < mid_2[3279:3272]) ? 1 : 0;
assign detect_min[409][15] = (mid_1[3287:3280] < mid_2[3287:3280]) ? 1 : 0;
assign detect_min[409][16] = (mid_1[3287:3280] < mid_2[3295:3288]) ? 1 : 0;
assign detect_min[409][17] = (mid_1[3287:3280] < btm_0[3279:3272]) ? 1 : 0;
assign detect_min[409][18] = (mid_1[3287:3280] < btm_0[3287:3280]) ? 1 : 0;
assign detect_min[409][19] = (mid_1[3287:3280] < btm_0[3295:3288]) ? 1 : 0;
assign detect_min[409][20] = (mid_1[3287:3280] < btm_1[3279:3272]) ? 1 : 0;
assign detect_min[409][21] = (mid_1[3287:3280] < btm_1[3287:3280]) ? 1 : 0;
assign detect_min[409][22] = (mid_1[3287:3280] < btm_1[3295:3288]) ? 1 : 0;
assign detect_min[409][23] = (mid_1[3287:3280] < btm_2[3279:3272]) ? 1 : 0;
assign detect_min[409][24] = (mid_1[3287:3280] < btm_2[3287:3280]) ? 1 : 0;
assign detect_min[409][25] = (mid_1[3287:3280] < btm_2[3295:3288]) ? 1 : 0;

assign detect_min[410][0] = (mid_1[3295:3288] < top_0[3287:3280]) ? 1 : 0;
assign detect_min[410][1] = (mid_1[3295:3288] < top_0[3295:3288]) ? 1 : 0;
assign detect_min[410][2] = (mid_1[3295:3288] < top_0[3303:3296]) ? 1 : 0;
assign detect_min[410][3] = (mid_1[3295:3288] < top_1[3287:3280]) ? 1 : 0;
assign detect_min[410][4] = (mid_1[3295:3288] < top_1[3295:3288]) ? 1 : 0;
assign detect_min[410][5] = (mid_1[3295:3288] < top_1[3303:3296]) ? 1 : 0;
assign detect_min[410][6] = (mid_1[3295:3288] < top_2[3287:3280]) ? 1 : 0;
assign detect_min[410][7] = (mid_1[3295:3288] < top_2[3295:3288]) ? 1 : 0;
assign detect_min[410][8] = (mid_1[3295:3288] < top_2[3303:3296]) ? 1 : 0;
assign detect_min[410][9] = (mid_1[3295:3288] < mid_0[3287:3280]) ? 1 : 0;
assign detect_min[410][10] = (mid_1[3295:3288] < mid_0[3295:3288]) ? 1 : 0;
assign detect_min[410][11] = (mid_1[3295:3288] < mid_0[3303:3296]) ? 1 : 0;
assign detect_min[410][12] = (mid_1[3295:3288] < mid_1[3287:3280]) ? 1 : 0;
assign detect_min[410][13] = (mid_1[3295:3288] < mid_1[3303:3296]) ? 1 : 0;
assign detect_min[410][14] = (mid_1[3295:3288] < mid_2[3287:3280]) ? 1 : 0;
assign detect_min[410][15] = (mid_1[3295:3288] < mid_2[3295:3288]) ? 1 : 0;
assign detect_min[410][16] = (mid_1[3295:3288] < mid_2[3303:3296]) ? 1 : 0;
assign detect_min[410][17] = (mid_1[3295:3288] < btm_0[3287:3280]) ? 1 : 0;
assign detect_min[410][18] = (mid_1[3295:3288] < btm_0[3295:3288]) ? 1 : 0;
assign detect_min[410][19] = (mid_1[3295:3288] < btm_0[3303:3296]) ? 1 : 0;
assign detect_min[410][20] = (mid_1[3295:3288] < btm_1[3287:3280]) ? 1 : 0;
assign detect_min[410][21] = (mid_1[3295:3288] < btm_1[3295:3288]) ? 1 : 0;
assign detect_min[410][22] = (mid_1[3295:3288] < btm_1[3303:3296]) ? 1 : 0;
assign detect_min[410][23] = (mid_1[3295:3288] < btm_2[3287:3280]) ? 1 : 0;
assign detect_min[410][24] = (mid_1[3295:3288] < btm_2[3295:3288]) ? 1 : 0;
assign detect_min[410][25] = (mid_1[3295:3288] < btm_2[3303:3296]) ? 1 : 0;

assign detect_min[411][0] = (mid_1[3303:3296] < top_0[3295:3288]) ? 1 : 0;
assign detect_min[411][1] = (mid_1[3303:3296] < top_0[3303:3296]) ? 1 : 0;
assign detect_min[411][2] = (mid_1[3303:3296] < top_0[3311:3304]) ? 1 : 0;
assign detect_min[411][3] = (mid_1[3303:3296] < top_1[3295:3288]) ? 1 : 0;
assign detect_min[411][4] = (mid_1[3303:3296] < top_1[3303:3296]) ? 1 : 0;
assign detect_min[411][5] = (mid_1[3303:3296] < top_1[3311:3304]) ? 1 : 0;
assign detect_min[411][6] = (mid_1[3303:3296] < top_2[3295:3288]) ? 1 : 0;
assign detect_min[411][7] = (mid_1[3303:3296] < top_2[3303:3296]) ? 1 : 0;
assign detect_min[411][8] = (mid_1[3303:3296] < top_2[3311:3304]) ? 1 : 0;
assign detect_min[411][9] = (mid_1[3303:3296] < mid_0[3295:3288]) ? 1 : 0;
assign detect_min[411][10] = (mid_1[3303:3296] < mid_0[3303:3296]) ? 1 : 0;
assign detect_min[411][11] = (mid_1[3303:3296] < mid_0[3311:3304]) ? 1 : 0;
assign detect_min[411][12] = (mid_1[3303:3296] < mid_1[3295:3288]) ? 1 : 0;
assign detect_min[411][13] = (mid_1[3303:3296] < mid_1[3311:3304]) ? 1 : 0;
assign detect_min[411][14] = (mid_1[3303:3296] < mid_2[3295:3288]) ? 1 : 0;
assign detect_min[411][15] = (mid_1[3303:3296] < mid_2[3303:3296]) ? 1 : 0;
assign detect_min[411][16] = (mid_1[3303:3296] < mid_2[3311:3304]) ? 1 : 0;
assign detect_min[411][17] = (mid_1[3303:3296] < btm_0[3295:3288]) ? 1 : 0;
assign detect_min[411][18] = (mid_1[3303:3296] < btm_0[3303:3296]) ? 1 : 0;
assign detect_min[411][19] = (mid_1[3303:3296] < btm_0[3311:3304]) ? 1 : 0;
assign detect_min[411][20] = (mid_1[3303:3296] < btm_1[3295:3288]) ? 1 : 0;
assign detect_min[411][21] = (mid_1[3303:3296] < btm_1[3303:3296]) ? 1 : 0;
assign detect_min[411][22] = (mid_1[3303:3296] < btm_1[3311:3304]) ? 1 : 0;
assign detect_min[411][23] = (mid_1[3303:3296] < btm_2[3295:3288]) ? 1 : 0;
assign detect_min[411][24] = (mid_1[3303:3296] < btm_2[3303:3296]) ? 1 : 0;
assign detect_min[411][25] = (mid_1[3303:3296] < btm_2[3311:3304]) ? 1 : 0;

assign detect_min[412][0] = (mid_1[3311:3304] < top_0[3303:3296]) ? 1 : 0;
assign detect_min[412][1] = (mid_1[3311:3304] < top_0[3311:3304]) ? 1 : 0;
assign detect_min[412][2] = (mid_1[3311:3304] < top_0[3319:3312]) ? 1 : 0;
assign detect_min[412][3] = (mid_1[3311:3304] < top_1[3303:3296]) ? 1 : 0;
assign detect_min[412][4] = (mid_1[3311:3304] < top_1[3311:3304]) ? 1 : 0;
assign detect_min[412][5] = (mid_1[3311:3304] < top_1[3319:3312]) ? 1 : 0;
assign detect_min[412][6] = (mid_1[3311:3304] < top_2[3303:3296]) ? 1 : 0;
assign detect_min[412][7] = (mid_1[3311:3304] < top_2[3311:3304]) ? 1 : 0;
assign detect_min[412][8] = (mid_1[3311:3304] < top_2[3319:3312]) ? 1 : 0;
assign detect_min[412][9] = (mid_1[3311:3304] < mid_0[3303:3296]) ? 1 : 0;
assign detect_min[412][10] = (mid_1[3311:3304] < mid_0[3311:3304]) ? 1 : 0;
assign detect_min[412][11] = (mid_1[3311:3304] < mid_0[3319:3312]) ? 1 : 0;
assign detect_min[412][12] = (mid_1[3311:3304] < mid_1[3303:3296]) ? 1 : 0;
assign detect_min[412][13] = (mid_1[3311:3304] < mid_1[3319:3312]) ? 1 : 0;
assign detect_min[412][14] = (mid_1[3311:3304] < mid_2[3303:3296]) ? 1 : 0;
assign detect_min[412][15] = (mid_1[3311:3304] < mid_2[3311:3304]) ? 1 : 0;
assign detect_min[412][16] = (mid_1[3311:3304] < mid_2[3319:3312]) ? 1 : 0;
assign detect_min[412][17] = (mid_1[3311:3304] < btm_0[3303:3296]) ? 1 : 0;
assign detect_min[412][18] = (mid_1[3311:3304] < btm_0[3311:3304]) ? 1 : 0;
assign detect_min[412][19] = (mid_1[3311:3304] < btm_0[3319:3312]) ? 1 : 0;
assign detect_min[412][20] = (mid_1[3311:3304] < btm_1[3303:3296]) ? 1 : 0;
assign detect_min[412][21] = (mid_1[3311:3304] < btm_1[3311:3304]) ? 1 : 0;
assign detect_min[412][22] = (mid_1[3311:3304] < btm_1[3319:3312]) ? 1 : 0;
assign detect_min[412][23] = (mid_1[3311:3304] < btm_2[3303:3296]) ? 1 : 0;
assign detect_min[412][24] = (mid_1[3311:3304] < btm_2[3311:3304]) ? 1 : 0;
assign detect_min[412][25] = (mid_1[3311:3304] < btm_2[3319:3312]) ? 1 : 0;

assign detect_min[413][0] = (mid_1[3319:3312] < top_0[3311:3304]) ? 1 : 0;
assign detect_min[413][1] = (mid_1[3319:3312] < top_0[3319:3312]) ? 1 : 0;
assign detect_min[413][2] = (mid_1[3319:3312] < top_0[3327:3320]) ? 1 : 0;
assign detect_min[413][3] = (mid_1[3319:3312] < top_1[3311:3304]) ? 1 : 0;
assign detect_min[413][4] = (mid_1[3319:3312] < top_1[3319:3312]) ? 1 : 0;
assign detect_min[413][5] = (mid_1[3319:3312] < top_1[3327:3320]) ? 1 : 0;
assign detect_min[413][6] = (mid_1[3319:3312] < top_2[3311:3304]) ? 1 : 0;
assign detect_min[413][7] = (mid_1[3319:3312] < top_2[3319:3312]) ? 1 : 0;
assign detect_min[413][8] = (mid_1[3319:3312] < top_2[3327:3320]) ? 1 : 0;
assign detect_min[413][9] = (mid_1[3319:3312] < mid_0[3311:3304]) ? 1 : 0;
assign detect_min[413][10] = (mid_1[3319:3312] < mid_0[3319:3312]) ? 1 : 0;
assign detect_min[413][11] = (mid_1[3319:3312] < mid_0[3327:3320]) ? 1 : 0;
assign detect_min[413][12] = (mid_1[3319:3312] < mid_1[3311:3304]) ? 1 : 0;
assign detect_min[413][13] = (mid_1[3319:3312] < mid_1[3327:3320]) ? 1 : 0;
assign detect_min[413][14] = (mid_1[3319:3312] < mid_2[3311:3304]) ? 1 : 0;
assign detect_min[413][15] = (mid_1[3319:3312] < mid_2[3319:3312]) ? 1 : 0;
assign detect_min[413][16] = (mid_1[3319:3312] < mid_2[3327:3320]) ? 1 : 0;
assign detect_min[413][17] = (mid_1[3319:3312] < btm_0[3311:3304]) ? 1 : 0;
assign detect_min[413][18] = (mid_1[3319:3312] < btm_0[3319:3312]) ? 1 : 0;
assign detect_min[413][19] = (mid_1[3319:3312] < btm_0[3327:3320]) ? 1 : 0;
assign detect_min[413][20] = (mid_1[3319:3312] < btm_1[3311:3304]) ? 1 : 0;
assign detect_min[413][21] = (mid_1[3319:3312] < btm_1[3319:3312]) ? 1 : 0;
assign detect_min[413][22] = (mid_1[3319:3312] < btm_1[3327:3320]) ? 1 : 0;
assign detect_min[413][23] = (mid_1[3319:3312] < btm_2[3311:3304]) ? 1 : 0;
assign detect_min[413][24] = (mid_1[3319:3312] < btm_2[3319:3312]) ? 1 : 0;
assign detect_min[413][25] = (mid_1[3319:3312] < btm_2[3327:3320]) ? 1 : 0;

assign detect_min[414][0] = (mid_1[3327:3320] < top_0[3319:3312]) ? 1 : 0;
assign detect_min[414][1] = (mid_1[3327:3320] < top_0[3327:3320]) ? 1 : 0;
assign detect_min[414][2] = (mid_1[3327:3320] < top_0[3335:3328]) ? 1 : 0;
assign detect_min[414][3] = (mid_1[3327:3320] < top_1[3319:3312]) ? 1 : 0;
assign detect_min[414][4] = (mid_1[3327:3320] < top_1[3327:3320]) ? 1 : 0;
assign detect_min[414][5] = (mid_1[3327:3320] < top_1[3335:3328]) ? 1 : 0;
assign detect_min[414][6] = (mid_1[3327:3320] < top_2[3319:3312]) ? 1 : 0;
assign detect_min[414][7] = (mid_1[3327:3320] < top_2[3327:3320]) ? 1 : 0;
assign detect_min[414][8] = (mid_1[3327:3320] < top_2[3335:3328]) ? 1 : 0;
assign detect_min[414][9] = (mid_1[3327:3320] < mid_0[3319:3312]) ? 1 : 0;
assign detect_min[414][10] = (mid_1[3327:3320] < mid_0[3327:3320]) ? 1 : 0;
assign detect_min[414][11] = (mid_1[3327:3320] < mid_0[3335:3328]) ? 1 : 0;
assign detect_min[414][12] = (mid_1[3327:3320] < mid_1[3319:3312]) ? 1 : 0;
assign detect_min[414][13] = (mid_1[3327:3320] < mid_1[3335:3328]) ? 1 : 0;
assign detect_min[414][14] = (mid_1[3327:3320] < mid_2[3319:3312]) ? 1 : 0;
assign detect_min[414][15] = (mid_1[3327:3320] < mid_2[3327:3320]) ? 1 : 0;
assign detect_min[414][16] = (mid_1[3327:3320] < mid_2[3335:3328]) ? 1 : 0;
assign detect_min[414][17] = (mid_1[3327:3320] < btm_0[3319:3312]) ? 1 : 0;
assign detect_min[414][18] = (mid_1[3327:3320] < btm_0[3327:3320]) ? 1 : 0;
assign detect_min[414][19] = (mid_1[3327:3320] < btm_0[3335:3328]) ? 1 : 0;
assign detect_min[414][20] = (mid_1[3327:3320] < btm_1[3319:3312]) ? 1 : 0;
assign detect_min[414][21] = (mid_1[3327:3320] < btm_1[3327:3320]) ? 1 : 0;
assign detect_min[414][22] = (mid_1[3327:3320] < btm_1[3335:3328]) ? 1 : 0;
assign detect_min[414][23] = (mid_1[3327:3320] < btm_2[3319:3312]) ? 1 : 0;
assign detect_min[414][24] = (mid_1[3327:3320] < btm_2[3327:3320]) ? 1 : 0;
assign detect_min[414][25] = (mid_1[3327:3320] < btm_2[3335:3328]) ? 1 : 0;

assign detect_min[415][0] = (mid_1[3335:3328] < top_0[3327:3320]) ? 1 : 0;
assign detect_min[415][1] = (mid_1[3335:3328] < top_0[3335:3328]) ? 1 : 0;
assign detect_min[415][2] = (mid_1[3335:3328] < top_0[3343:3336]) ? 1 : 0;
assign detect_min[415][3] = (mid_1[3335:3328] < top_1[3327:3320]) ? 1 : 0;
assign detect_min[415][4] = (mid_1[3335:3328] < top_1[3335:3328]) ? 1 : 0;
assign detect_min[415][5] = (mid_1[3335:3328] < top_1[3343:3336]) ? 1 : 0;
assign detect_min[415][6] = (mid_1[3335:3328] < top_2[3327:3320]) ? 1 : 0;
assign detect_min[415][7] = (mid_1[3335:3328] < top_2[3335:3328]) ? 1 : 0;
assign detect_min[415][8] = (mid_1[3335:3328] < top_2[3343:3336]) ? 1 : 0;
assign detect_min[415][9] = (mid_1[3335:3328] < mid_0[3327:3320]) ? 1 : 0;
assign detect_min[415][10] = (mid_1[3335:3328] < mid_0[3335:3328]) ? 1 : 0;
assign detect_min[415][11] = (mid_1[3335:3328] < mid_0[3343:3336]) ? 1 : 0;
assign detect_min[415][12] = (mid_1[3335:3328] < mid_1[3327:3320]) ? 1 : 0;
assign detect_min[415][13] = (mid_1[3335:3328] < mid_1[3343:3336]) ? 1 : 0;
assign detect_min[415][14] = (mid_1[3335:3328] < mid_2[3327:3320]) ? 1 : 0;
assign detect_min[415][15] = (mid_1[3335:3328] < mid_2[3335:3328]) ? 1 : 0;
assign detect_min[415][16] = (mid_1[3335:3328] < mid_2[3343:3336]) ? 1 : 0;
assign detect_min[415][17] = (mid_1[3335:3328] < btm_0[3327:3320]) ? 1 : 0;
assign detect_min[415][18] = (mid_1[3335:3328] < btm_0[3335:3328]) ? 1 : 0;
assign detect_min[415][19] = (mid_1[3335:3328] < btm_0[3343:3336]) ? 1 : 0;
assign detect_min[415][20] = (mid_1[3335:3328] < btm_1[3327:3320]) ? 1 : 0;
assign detect_min[415][21] = (mid_1[3335:3328] < btm_1[3335:3328]) ? 1 : 0;
assign detect_min[415][22] = (mid_1[3335:3328] < btm_1[3343:3336]) ? 1 : 0;
assign detect_min[415][23] = (mid_1[3335:3328] < btm_2[3327:3320]) ? 1 : 0;
assign detect_min[415][24] = (mid_1[3335:3328] < btm_2[3335:3328]) ? 1 : 0;
assign detect_min[415][25] = (mid_1[3335:3328] < btm_2[3343:3336]) ? 1 : 0;

assign detect_min[416][0] = (mid_1[3343:3336] < top_0[3335:3328]) ? 1 : 0;
assign detect_min[416][1] = (mid_1[3343:3336] < top_0[3343:3336]) ? 1 : 0;
assign detect_min[416][2] = (mid_1[3343:3336] < top_0[3351:3344]) ? 1 : 0;
assign detect_min[416][3] = (mid_1[3343:3336] < top_1[3335:3328]) ? 1 : 0;
assign detect_min[416][4] = (mid_1[3343:3336] < top_1[3343:3336]) ? 1 : 0;
assign detect_min[416][5] = (mid_1[3343:3336] < top_1[3351:3344]) ? 1 : 0;
assign detect_min[416][6] = (mid_1[3343:3336] < top_2[3335:3328]) ? 1 : 0;
assign detect_min[416][7] = (mid_1[3343:3336] < top_2[3343:3336]) ? 1 : 0;
assign detect_min[416][8] = (mid_1[3343:3336] < top_2[3351:3344]) ? 1 : 0;
assign detect_min[416][9] = (mid_1[3343:3336] < mid_0[3335:3328]) ? 1 : 0;
assign detect_min[416][10] = (mid_1[3343:3336] < mid_0[3343:3336]) ? 1 : 0;
assign detect_min[416][11] = (mid_1[3343:3336] < mid_0[3351:3344]) ? 1 : 0;
assign detect_min[416][12] = (mid_1[3343:3336] < mid_1[3335:3328]) ? 1 : 0;
assign detect_min[416][13] = (mid_1[3343:3336] < mid_1[3351:3344]) ? 1 : 0;
assign detect_min[416][14] = (mid_1[3343:3336] < mid_2[3335:3328]) ? 1 : 0;
assign detect_min[416][15] = (mid_1[3343:3336] < mid_2[3343:3336]) ? 1 : 0;
assign detect_min[416][16] = (mid_1[3343:3336] < mid_2[3351:3344]) ? 1 : 0;
assign detect_min[416][17] = (mid_1[3343:3336] < btm_0[3335:3328]) ? 1 : 0;
assign detect_min[416][18] = (mid_1[3343:3336] < btm_0[3343:3336]) ? 1 : 0;
assign detect_min[416][19] = (mid_1[3343:3336] < btm_0[3351:3344]) ? 1 : 0;
assign detect_min[416][20] = (mid_1[3343:3336] < btm_1[3335:3328]) ? 1 : 0;
assign detect_min[416][21] = (mid_1[3343:3336] < btm_1[3343:3336]) ? 1 : 0;
assign detect_min[416][22] = (mid_1[3343:3336] < btm_1[3351:3344]) ? 1 : 0;
assign detect_min[416][23] = (mid_1[3343:3336] < btm_2[3335:3328]) ? 1 : 0;
assign detect_min[416][24] = (mid_1[3343:3336] < btm_2[3343:3336]) ? 1 : 0;
assign detect_min[416][25] = (mid_1[3343:3336] < btm_2[3351:3344]) ? 1 : 0;

assign detect_min[417][0] = (mid_1[3351:3344] < top_0[3343:3336]) ? 1 : 0;
assign detect_min[417][1] = (mid_1[3351:3344] < top_0[3351:3344]) ? 1 : 0;
assign detect_min[417][2] = (mid_1[3351:3344] < top_0[3359:3352]) ? 1 : 0;
assign detect_min[417][3] = (mid_1[3351:3344] < top_1[3343:3336]) ? 1 : 0;
assign detect_min[417][4] = (mid_1[3351:3344] < top_1[3351:3344]) ? 1 : 0;
assign detect_min[417][5] = (mid_1[3351:3344] < top_1[3359:3352]) ? 1 : 0;
assign detect_min[417][6] = (mid_1[3351:3344] < top_2[3343:3336]) ? 1 : 0;
assign detect_min[417][7] = (mid_1[3351:3344] < top_2[3351:3344]) ? 1 : 0;
assign detect_min[417][8] = (mid_1[3351:3344] < top_2[3359:3352]) ? 1 : 0;
assign detect_min[417][9] = (mid_1[3351:3344] < mid_0[3343:3336]) ? 1 : 0;
assign detect_min[417][10] = (mid_1[3351:3344] < mid_0[3351:3344]) ? 1 : 0;
assign detect_min[417][11] = (mid_1[3351:3344] < mid_0[3359:3352]) ? 1 : 0;
assign detect_min[417][12] = (mid_1[3351:3344] < mid_1[3343:3336]) ? 1 : 0;
assign detect_min[417][13] = (mid_1[3351:3344] < mid_1[3359:3352]) ? 1 : 0;
assign detect_min[417][14] = (mid_1[3351:3344] < mid_2[3343:3336]) ? 1 : 0;
assign detect_min[417][15] = (mid_1[3351:3344] < mid_2[3351:3344]) ? 1 : 0;
assign detect_min[417][16] = (mid_1[3351:3344] < mid_2[3359:3352]) ? 1 : 0;
assign detect_min[417][17] = (mid_1[3351:3344] < btm_0[3343:3336]) ? 1 : 0;
assign detect_min[417][18] = (mid_1[3351:3344] < btm_0[3351:3344]) ? 1 : 0;
assign detect_min[417][19] = (mid_1[3351:3344] < btm_0[3359:3352]) ? 1 : 0;
assign detect_min[417][20] = (mid_1[3351:3344] < btm_1[3343:3336]) ? 1 : 0;
assign detect_min[417][21] = (mid_1[3351:3344] < btm_1[3351:3344]) ? 1 : 0;
assign detect_min[417][22] = (mid_1[3351:3344] < btm_1[3359:3352]) ? 1 : 0;
assign detect_min[417][23] = (mid_1[3351:3344] < btm_2[3343:3336]) ? 1 : 0;
assign detect_min[417][24] = (mid_1[3351:3344] < btm_2[3351:3344]) ? 1 : 0;
assign detect_min[417][25] = (mid_1[3351:3344] < btm_2[3359:3352]) ? 1 : 0;

assign detect_min[418][0] = (mid_1[3359:3352] < top_0[3351:3344]) ? 1 : 0;
assign detect_min[418][1] = (mid_1[3359:3352] < top_0[3359:3352]) ? 1 : 0;
assign detect_min[418][2] = (mid_1[3359:3352] < top_0[3367:3360]) ? 1 : 0;
assign detect_min[418][3] = (mid_1[3359:3352] < top_1[3351:3344]) ? 1 : 0;
assign detect_min[418][4] = (mid_1[3359:3352] < top_1[3359:3352]) ? 1 : 0;
assign detect_min[418][5] = (mid_1[3359:3352] < top_1[3367:3360]) ? 1 : 0;
assign detect_min[418][6] = (mid_1[3359:3352] < top_2[3351:3344]) ? 1 : 0;
assign detect_min[418][7] = (mid_1[3359:3352] < top_2[3359:3352]) ? 1 : 0;
assign detect_min[418][8] = (mid_1[3359:3352] < top_2[3367:3360]) ? 1 : 0;
assign detect_min[418][9] = (mid_1[3359:3352] < mid_0[3351:3344]) ? 1 : 0;
assign detect_min[418][10] = (mid_1[3359:3352] < mid_0[3359:3352]) ? 1 : 0;
assign detect_min[418][11] = (mid_1[3359:3352] < mid_0[3367:3360]) ? 1 : 0;
assign detect_min[418][12] = (mid_1[3359:3352] < mid_1[3351:3344]) ? 1 : 0;
assign detect_min[418][13] = (mid_1[3359:3352] < mid_1[3367:3360]) ? 1 : 0;
assign detect_min[418][14] = (mid_1[3359:3352] < mid_2[3351:3344]) ? 1 : 0;
assign detect_min[418][15] = (mid_1[3359:3352] < mid_2[3359:3352]) ? 1 : 0;
assign detect_min[418][16] = (mid_1[3359:3352] < mid_2[3367:3360]) ? 1 : 0;
assign detect_min[418][17] = (mid_1[3359:3352] < btm_0[3351:3344]) ? 1 : 0;
assign detect_min[418][18] = (mid_1[3359:3352] < btm_0[3359:3352]) ? 1 : 0;
assign detect_min[418][19] = (mid_1[3359:3352] < btm_0[3367:3360]) ? 1 : 0;
assign detect_min[418][20] = (mid_1[3359:3352] < btm_1[3351:3344]) ? 1 : 0;
assign detect_min[418][21] = (mid_1[3359:3352] < btm_1[3359:3352]) ? 1 : 0;
assign detect_min[418][22] = (mid_1[3359:3352] < btm_1[3367:3360]) ? 1 : 0;
assign detect_min[418][23] = (mid_1[3359:3352] < btm_2[3351:3344]) ? 1 : 0;
assign detect_min[418][24] = (mid_1[3359:3352] < btm_2[3359:3352]) ? 1 : 0;
assign detect_min[418][25] = (mid_1[3359:3352] < btm_2[3367:3360]) ? 1 : 0;

assign detect_min[419][0] = (mid_1[3367:3360] < top_0[3359:3352]) ? 1 : 0;
assign detect_min[419][1] = (mid_1[3367:3360] < top_0[3367:3360]) ? 1 : 0;
assign detect_min[419][2] = (mid_1[3367:3360] < top_0[3375:3368]) ? 1 : 0;
assign detect_min[419][3] = (mid_1[3367:3360] < top_1[3359:3352]) ? 1 : 0;
assign detect_min[419][4] = (mid_1[3367:3360] < top_1[3367:3360]) ? 1 : 0;
assign detect_min[419][5] = (mid_1[3367:3360] < top_1[3375:3368]) ? 1 : 0;
assign detect_min[419][6] = (mid_1[3367:3360] < top_2[3359:3352]) ? 1 : 0;
assign detect_min[419][7] = (mid_1[3367:3360] < top_2[3367:3360]) ? 1 : 0;
assign detect_min[419][8] = (mid_1[3367:3360] < top_2[3375:3368]) ? 1 : 0;
assign detect_min[419][9] = (mid_1[3367:3360] < mid_0[3359:3352]) ? 1 : 0;
assign detect_min[419][10] = (mid_1[3367:3360] < mid_0[3367:3360]) ? 1 : 0;
assign detect_min[419][11] = (mid_1[3367:3360] < mid_0[3375:3368]) ? 1 : 0;
assign detect_min[419][12] = (mid_1[3367:3360] < mid_1[3359:3352]) ? 1 : 0;
assign detect_min[419][13] = (mid_1[3367:3360] < mid_1[3375:3368]) ? 1 : 0;
assign detect_min[419][14] = (mid_1[3367:3360] < mid_2[3359:3352]) ? 1 : 0;
assign detect_min[419][15] = (mid_1[3367:3360] < mid_2[3367:3360]) ? 1 : 0;
assign detect_min[419][16] = (mid_1[3367:3360] < mid_2[3375:3368]) ? 1 : 0;
assign detect_min[419][17] = (mid_1[3367:3360] < btm_0[3359:3352]) ? 1 : 0;
assign detect_min[419][18] = (mid_1[3367:3360] < btm_0[3367:3360]) ? 1 : 0;
assign detect_min[419][19] = (mid_1[3367:3360] < btm_0[3375:3368]) ? 1 : 0;
assign detect_min[419][20] = (mid_1[3367:3360] < btm_1[3359:3352]) ? 1 : 0;
assign detect_min[419][21] = (mid_1[3367:3360] < btm_1[3367:3360]) ? 1 : 0;
assign detect_min[419][22] = (mid_1[3367:3360] < btm_1[3375:3368]) ? 1 : 0;
assign detect_min[419][23] = (mid_1[3367:3360] < btm_2[3359:3352]) ? 1 : 0;
assign detect_min[419][24] = (mid_1[3367:3360] < btm_2[3367:3360]) ? 1 : 0;
assign detect_min[419][25] = (mid_1[3367:3360] < btm_2[3375:3368]) ? 1 : 0;

assign detect_min[420][0] = (mid_1[3375:3368] < top_0[3367:3360]) ? 1 : 0;
assign detect_min[420][1] = (mid_1[3375:3368] < top_0[3375:3368]) ? 1 : 0;
assign detect_min[420][2] = (mid_1[3375:3368] < top_0[3383:3376]) ? 1 : 0;
assign detect_min[420][3] = (mid_1[3375:3368] < top_1[3367:3360]) ? 1 : 0;
assign detect_min[420][4] = (mid_1[3375:3368] < top_1[3375:3368]) ? 1 : 0;
assign detect_min[420][5] = (mid_1[3375:3368] < top_1[3383:3376]) ? 1 : 0;
assign detect_min[420][6] = (mid_1[3375:3368] < top_2[3367:3360]) ? 1 : 0;
assign detect_min[420][7] = (mid_1[3375:3368] < top_2[3375:3368]) ? 1 : 0;
assign detect_min[420][8] = (mid_1[3375:3368] < top_2[3383:3376]) ? 1 : 0;
assign detect_min[420][9] = (mid_1[3375:3368] < mid_0[3367:3360]) ? 1 : 0;
assign detect_min[420][10] = (mid_1[3375:3368] < mid_0[3375:3368]) ? 1 : 0;
assign detect_min[420][11] = (mid_1[3375:3368] < mid_0[3383:3376]) ? 1 : 0;
assign detect_min[420][12] = (mid_1[3375:3368] < mid_1[3367:3360]) ? 1 : 0;
assign detect_min[420][13] = (mid_1[3375:3368] < mid_1[3383:3376]) ? 1 : 0;
assign detect_min[420][14] = (mid_1[3375:3368] < mid_2[3367:3360]) ? 1 : 0;
assign detect_min[420][15] = (mid_1[3375:3368] < mid_2[3375:3368]) ? 1 : 0;
assign detect_min[420][16] = (mid_1[3375:3368] < mid_2[3383:3376]) ? 1 : 0;
assign detect_min[420][17] = (mid_1[3375:3368] < btm_0[3367:3360]) ? 1 : 0;
assign detect_min[420][18] = (mid_1[3375:3368] < btm_0[3375:3368]) ? 1 : 0;
assign detect_min[420][19] = (mid_1[3375:3368] < btm_0[3383:3376]) ? 1 : 0;
assign detect_min[420][20] = (mid_1[3375:3368] < btm_1[3367:3360]) ? 1 : 0;
assign detect_min[420][21] = (mid_1[3375:3368] < btm_1[3375:3368]) ? 1 : 0;
assign detect_min[420][22] = (mid_1[3375:3368] < btm_1[3383:3376]) ? 1 : 0;
assign detect_min[420][23] = (mid_1[3375:3368] < btm_2[3367:3360]) ? 1 : 0;
assign detect_min[420][24] = (mid_1[3375:3368] < btm_2[3375:3368]) ? 1 : 0;
assign detect_min[420][25] = (mid_1[3375:3368] < btm_2[3383:3376]) ? 1 : 0;

assign detect_min[421][0] = (mid_1[3383:3376] < top_0[3375:3368]) ? 1 : 0;
assign detect_min[421][1] = (mid_1[3383:3376] < top_0[3383:3376]) ? 1 : 0;
assign detect_min[421][2] = (mid_1[3383:3376] < top_0[3391:3384]) ? 1 : 0;
assign detect_min[421][3] = (mid_1[3383:3376] < top_1[3375:3368]) ? 1 : 0;
assign detect_min[421][4] = (mid_1[3383:3376] < top_1[3383:3376]) ? 1 : 0;
assign detect_min[421][5] = (mid_1[3383:3376] < top_1[3391:3384]) ? 1 : 0;
assign detect_min[421][6] = (mid_1[3383:3376] < top_2[3375:3368]) ? 1 : 0;
assign detect_min[421][7] = (mid_1[3383:3376] < top_2[3383:3376]) ? 1 : 0;
assign detect_min[421][8] = (mid_1[3383:3376] < top_2[3391:3384]) ? 1 : 0;
assign detect_min[421][9] = (mid_1[3383:3376] < mid_0[3375:3368]) ? 1 : 0;
assign detect_min[421][10] = (mid_1[3383:3376] < mid_0[3383:3376]) ? 1 : 0;
assign detect_min[421][11] = (mid_1[3383:3376] < mid_0[3391:3384]) ? 1 : 0;
assign detect_min[421][12] = (mid_1[3383:3376] < mid_1[3375:3368]) ? 1 : 0;
assign detect_min[421][13] = (mid_1[3383:3376] < mid_1[3391:3384]) ? 1 : 0;
assign detect_min[421][14] = (mid_1[3383:3376] < mid_2[3375:3368]) ? 1 : 0;
assign detect_min[421][15] = (mid_1[3383:3376] < mid_2[3383:3376]) ? 1 : 0;
assign detect_min[421][16] = (mid_1[3383:3376] < mid_2[3391:3384]) ? 1 : 0;
assign detect_min[421][17] = (mid_1[3383:3376] < btm_0[3375:3368]) ? 1 : 0;
assign detect_min[421][18] = (mid_1[3383:3376] < btm_0[3383:3376]) ? 1 : 0;
assign detect_min[421][19] = (mid_1[3383:3376] < btm_0[3391:3384]) ? 1 : 0;
assign detect_min[421][20] = (mid_1[3383:3376] < btm_1[3375:3368]) ? 1 : 0;
assign detect_min[421][21] = (mid_1[3383:3376] < btm_1[3383:3376]) ? 1 : 0;
assign detect_min[421][22] = (mid_1[3383:3376] < btm_1[3391:3384]) ? 1 : 0;
assign detect_min[421][23] = (mid_1[3383:3376] < btm_2[3375:3368]) ? 1 : 0;
assign detect_min[421][24] = (mid_1[3383:3376] < btm_2[3383:3376]) ? 1 : 0;
assign detect_min[421][25] = (mid_1[3383:3376] < btm_2[3391:3384]) ? 1 : 0;

assign detect_min[422][0] = (mid_1[3391:3384] < top_0[3383:3376]) ? 1 : 0;
assign detect_min[422][1] = (mid_1[3391:3384] < top_0[3391:3384]) ? 1 : 0;
assign detect_min[422][2] = (mid_1[3391:3384] < top_0[3399:3392]) ? 1 : 0;
assign detect_min[422][3] = (mid_1[3391:3384] < top_1[3383:3376]) ? 1 : 0;
assign detect_min[422][4] = (mid_1[3391:3384] < top_1[3391:3384]) ? 1 : 0;
assign detect_min[422][5] = (mid_1[3391:3384] < top_1[3399:3392]) ? 1 : 0;
assign detect_min[422][6] = (mid_1[3391:3384] < top_2[3383:3376]) ? 1 : 0;
assign detect_min[422][7] = (mid_1[3391:3384] < top_2[3391:3384]) ? 1 : 0;
assign detect_min[422][8] = (mid_1[3391:3384] < top_2[3399:3392]) ? 1 : 0;
assign detect_min[422][9] = (mid_1[3391:3384] < mid_0[3383:3376]) ? 1 : 0;
assign detect_min[422][10] = (mid_1[3391:3384] < mid_0[3391:3384]) ? 1 : 0;
assign detect_min[422][11] = (mid_1[3391:3384] < mid_0[3399:3392]) ? 1 : 0;
assign detect_min[422][12] = (mid_1[3391:3384] < mid_1[3383:3376]) ? 1 : 0;
assign detect_min[422][13] = (mid_1[3391:3384] < mid_1[3399:3392]) ? 1 : 0;
assign detect_min[422][14] = (mid_1[3391:3384] < mid_2[3383:3376]) ? 1 : 0;
assign detect_min[422][15] = (mid_1[3391:3384] < mid_2[3391:3384]) ? 1 : 0;
assign detect_min[422][16] = (mid_1[3391:3384] < mid_2[3399:3392]) ? 1 : 0;
assign detect_min[422][17] = (mid_1[3391:3384] < btm_0[3383:3376]) ? 1 : 0;
assign detect_min[422][18] = (mid_1[3391:3384] < btm_0[3391:3384]) ? 1 : 0;
assign detect_min[422][19] = (mid_1[3391:3384] < btm_0[3399:3392]) ? 1 : 0;
assign detect_min[422][20] = (mid_1[3391:3384] < btm_1[3383:3376]) ? 1 : 0;
assign detect_min[422][21] = (mid_1[3391:3384] < btm_1[3391:3384]) ? 1 : 0;
assign detect_min[422][22] = (mid_1[3391:3384] < btm_1[3399:3392]) ? 1 : 0;
assign detect_min[422][23] = (mid_1[3391:3384] < btm_2[3383:3376]) ? 1 : 0;
assign detect_min[422][24] = (mid_1[3391:3384] < btm_2[3391:3384]) ? 1 : 0;
assign detect_min[422][25] = (mid_1[3391:3384] < btm_2[3399:3392]) ? 1 : 0;

assign detect_min[423][0] = (mid_1[3399:3392] < top_0[3391:3384]) ? 1 : 0;
assign detect_min[423][1] = (mid_1[3399:3392] < top_0[3399:3392]) ? 1 : 0;
assign detect_min[423][2] = (mid_1[3399:3392] < top_0[3407:3400]) ? 1 : 0;
assign detect_min[423][3] = (mid_1[3399:3392] < top_1[3391:3384]) ? 1 : 0;
assign detect_min[423][4] = (mid_1[3399:3392] < top_1[3399:3392]) ? 1 : 0;
assign detect_min[423][5] = (mid_1[3399:3392] < top_1[3407:3400]) ? 1 : 0;
assign detect_min[423][6] = (mid_1[3399:3392] < top_2[3391:3384]) ? 1 : 0;
assign detect_min[423][7] = (mid_1[3399:3392] < top_2[3399:3392]) ? 1 : 0;
assign detect_min[423][8] = (mid_1[3399:3392] < top_2[3407:3400]) ? 1 : 0;
assign detect_min[423][9] = (mid_1[3399:3392] < mid_0[3391:3384]) ? 1 : 0;
assign detect_min[423][10] = (mid_1[3399:3392] < mid_0[3399:3392]) ? 1 : 0;
assign detect_min[423][11] = (mid_1[3399:3392] < mid_0[3407:3400]) ? 1 : 0;
assign detect_min[423][12] = (mid_1[3399:3392] < mid_1[3391:3384]) ? 1 : 0;
assign detect_min[423][13] = (mid_1[3399:3392] < mid_1[3407:3400]) ? 1 : 0;
assign detect_min[423][14] = (mid_1[3399:3392] < mid_2[3391:3384]) ? 1 : 0;
assign detect_min[423][15] = (mid_1[3399:3392] < mid_2[3399:3392]) ? 1 : 0;
assign detect_min[423][16] = (mid_1[3399:3392] < mid_2[3407:3400]) ? 1 : 0;
assign detect_min[423][17] = (mid_1[3399:3392] < btm_0[3391:3384]) ? 1 : 0;
assign detect_min[423][18] = (mid_1[3399:3392] < btm_0[3399:3392]) ? 1 : 0;
assign detect_min[423][19] = (mid_1[3399:3392] < btm_0[3407:3400]) ? 1 : 0;
assign detect_min[423][20] = (mid_1[3399:3392] < btm_1[3391:3384]) ? 1 : 0;
assign detect_min[423][21] = (mid_1[3399:3392] < btm_1[3399:3392]) ? 1 : 0;
assign detect_min[423][22] = (mid_1[3399:3392] < btm_1[3407:3400]) ? 1 : 0;
assign detect_min[423][23] = (mid_1[3399:3392] < btm_2[3391:3384]) ? 1 : 0;
assign detect_min[423][24] = (mid_1[3399:3392] < btm_2[3399:3392]) ? 1 : 0;
assign detect_min[423][25] = (mid_1[3399:3392] < btm_2[3407:3400]) ? 1 : 0;

assign detect_min[424][0] = (mid_1[3407:3400] < top_0[3399:3392]) ? 1 : 0;
assign detect_min[424][1] = (mid_1[3407:3400] < top_0[3407:3400]) ? 1 : 0;
assign detect_min[424][2] = (mid_1[3407:3400] < top_0[3415:3408]) ? 1 : 0;
assign detect_min[424][3] = (mid_1[3407:3400] < top_1[3399:3392]) ? 1 : 0;
assign detect_min[424][4] = (mid_1[3407:3400] < top_1[3407:3400]) ? 1 : 0;
assign detect_min[424][5] = (mid_1[3407:3400] < top_1[3415:3408]) ? 1 : 0;
assign detect_min[424][6] = (mid_1[3407:3400] < top_2[3399:3392]) ? 1 : 0;
assign detect_min[424][7] = (mid_1[3407:3400] < top_2[3407:3400]) ? 1 : 0;
assign detect_min[424][8] = (mid_1[3407:3400] < top_2[3415:3408]) ? 1 : 0;
assign detect_min[424][9] = (mid_1[3407:3400] < mid_0[3399:3392]) ? 1 : 0;
assign detect_min[424][10] = (mid_1[3407:3400] < mid_0[3407:3400]) ? 1 : 0;
assign detect_min[424][11] = (mid_1[3407:3400] < mid_0[3415:3408]) ? 1 : 0;
assign detect_min[424][12] = (mid_1[3407:3400] < mid_1[3399:3392]) ? 1 : 0;
assign detect_min[424][13] = (mid_1[3407:3400] < mid_1[3415:3408]) ? 1 : 0;
assign detect_min[424][14] = (mid_1[3407:3400] < mid_2[3399:3392]) ? 1 : 0;
assign detect_min[424][15] = (mid_1[3407:3400] < mid_2[3407:3400]) ? 1 : 0;
assign detect_min[424][16] = (mid_1[3407:3400] < mid_2[3415:3408]) ? 1 : 0;
assign detect_min[424][17] = (mid_1[3407:3400] < btm_0[3399:3392]) ? 1 : 0;
assign detect_min[424][18] = (mid_1[3407:3400] < btm_0[3407:3400]) ? 1 : 0;
assign detect_min[424][19] = (mid_1[3407:3400] < btm_0[3415:3408]) ? 1 : 0;
assign detect_min[424][20] = (mid_1[3407:3400] < btm_1[3399:3392]) ? 1 : 0;
assign detect_min[424][21] = (mid_1[3407:3400] < btm_1[3407:3400]) ? 1 : 0;
assign detect_min[424][22] = (mid_1[3407:3400] < btm_1[3415:3408]) ? 1 : 0;
assign detect_min[424][23] = (mid_1[3407:3400] < btm_2[3399:3392]) ? 1 : 0;
assign detect_min[424][24] = (mid_1[3407:3400] < btm_2[3407:3400]) ? 1 : 0;
assign detect_min[424][25] = (mid_1[3407:3400] < btm_2[3415:3408]) ? 1 : 0;

assign detect_min[425][0] = (mid_1[3415:3408] < top_0[3407:3400]) ? 1 : 0;
assign detect_min[425][1] = (mid_1[3415:3408] < top_0[3415:3408]) ? 1 : 0;
assign detect_min[425][2] = (mid_1[3415:3408] < top_0[3423:3416]) ? 1 : 0;
assign detect_min[425][3] = (mid_1[3415:3408] < top_1[3407:3400]) ? 1 : 0;
assign detect_min[425][4] = (mid_1[3415:3408] < top_1[3415:3408]) ? 1 : 0;
assign detect_min[425][5] = (mid_1[3415:3408] < top_1[3423:3416]) ? 1 : 0;
assign detect_min[425][6] = (mid_1[3415:3408] < top_2[3407:3400]) ? 1 : 0;
assign detect_min[425][7] = (mid_1[3415:3408] < top_2[3415:3408]) ? 1 : 0;
assign detect_min[425][8] = (mid_1[3415:3408] < top_2[3423:3416]) ? 1 : 0;
assign detect_min[425][9] = (mid_1[3415:3408] < mid_0[3407:3400]) ? 1 : 0;
assign detect_min[425][10] = (mid_1[3415:3408] < mid_0[3415:3408]) ? 1 : 0;
assign detect_min[425][11] = (mid_1[3415:3408] < mid_0[3423:3416]) ? 1 : 0;
assign detect_min[425][12] = (mid_1[3415:3408] < mid_1[3407:3400]) ? 1 : 0;
assign detect_min[425][13] = (mid_1[3415:3408] < mid_1[3423:3416]) ? 1 : 0;
assign detect_min[425][14] = (mid_1[3415:3408] < mid_2[3407:3400]) ? 1 : 0;
assign detect_min[425][15] = (mid_1[3415:3408] < mid_2[3415:3408]) ? 1 : 0;
assign detect_min[425][16] = (mid_1[3415:3408] < mid_2[3423:3416]) ? 1 : 0;
assign detect_min[425][17] = (mid_1[3415:3408] < btm_0[3407:3400]) ? 1 : 0;
assign detect_min[425][18] = (mid_1[3415:3408] < btm_0[3415:3408]) ? 1 : 0;
assign detect_min[425][19] = (mid_1[3415:3408] < btm_0[3423:3416]) ? 1 : 0;
assign detect_min[425][20] = (mid_1[3415:3408] < btm_1[3407:3400]) ? 1 : 0;
assign detect_min[425][21] = (mid_1[3415:3408] < btm_1[3415:3408]) ? 1 : 0;
assign detect_min[425][22] = (mid_1[3415:3408] < btm_1[3423:3416]) ? 1 : 0;
assign detect_min[425][23] = (mid_1[3415:3408] < btm_2[3407:3400]) ? 1 : 0;
assign detect_min[425][24] = (mid_1[3415:3408] < btm_2[3415:3408]) ? 1 : 0;
assign detect_min[425][25] = (mid_1[3415:3408] < btm_2[3423:3416]) ? 1 : 0;

assign detect_min[426][0] = (mid_1[3423:3416] < top_0[3415:3408]) ? 1 : 0;
assign detect_min[426][1] = (mid_1[3423:3416] < top_0[3423:3416]) ? 1 : 0;
assign detect_min[426][2] = (mid_1[3423:3416] < top_0[3431:3424]) ? 1 : 0;
assign detect_min[426][3] = (mid_1[3423:3416] < top_1[3415:3408]) ? 1 : 0;
assign detect_min[426][4] = (mid_1[3423:3416] < top_1[3423:3416]) ? 1 : 0;
assign detect_min[426][5] = (mid_1[3423:3416] < top_1[3431:3424]) ? 1 : 0;
assign detect_min[426][6] = (mid_1[3423:3416] < top_2[3415:3408]) ? 1 : 0;
assign detect_min[426][7] = (mid_1[3423:3416] < top_2[3423:3416]) ? 1 : 0;
assign detect_min[426][8] = (mid_1[3423:3416] < top_2[3431:3424]) ? 1 : 0;
assign detect_min[426][9] = (mid_1[3423:3416] < mid_0[3415:3408]) ? 1 : 0;
assign detect_min[426][10] = (mid_1[3423:3416] < mid_0[3423:3416]) ? 1 : 0;
assign detect_min[426][11] = (mid_1[3423:3416] < mid_0[3431:3424]) ? 1 : 0;
assign detect_min[426][12] = (mid_1[3423:3416] < mid_1[3415:3408]) ? 1 : 0;
assign detect_min[426][13] = (mid_1[3423:3416] < mid_1[3431:3424]) ? 1 : 0;
assign detect_min[426][14] = (mid_1[3423:3416] < mid_2[3415:3408]) ? 1 : 0;
assign detect_min[426][15] = (mid_1[3423:3416] < mid_2[3423:3416]) ? 1 : 0;
assign detect_min[426][16] = (mid_1[3423:3416] < mid_2[3431:3424]) ? 1 : 0;
assign detect_min[426][17] = (mid_1[3423:3416] < btm_0[3415:3408]) ? 1 : 0;
assign detect_min[426][18] = (mid_1[3423:3416] < btm_0[3423:3416]) ? 1 : 0;
assign detect_min[426][19] = (mid_1[3423:3416] < btm_0[3431:3424]) ? 1 : 0;
assign detect_min[426][20] = (mid_1[3423:3416] < btm_1[3415:3408]) ? 1 : 0;
assign detect_min[426][21] = (mid_1[3423:3416] < btm_1[3423:3416]) ? 1 : 0;
assign detect_min[426][22] = (mid_1[3423:3416] < btm_1[3431:3424]) ? 1 : 0;
assign detect_min[426][23] = (mid_1[3423:3416] < btm_2[3415:3408]) ? 1 : 0;
assign detect_min[426][24] = (mid_1[3423:3416] < btm_2[3423:3416]) ? 1 : 0;
assign detect_min[426][25] = (mid_1[3423:3416] < btm_2[3431:3424]) ? 1 : 0;

assign detect_min[427][0] = (mid_1[3431:3424] < top_0[3423:3416]) ? 1 : 0;
assign detect_min[427][1] = (mid_1[3431:3424] < top_0[3431:3424]) ? 1 : 0;
assign detect_min[427][2] = (mid_1[3431:3424] < top_0[3439:3432]) ? 1 : 0;
assign detect_min[427][3] = (mid_1[3431:3424] < top_1[3423:3416]) ? 1 : 0;
assign detect_min[427][4] = (mid_1[3431:3424] < top_1[3431:3424]) ? 1 : 0;
assign detect_min[427][5] = (mid_1[3431:3424] < top_1[3439:3432]) ? 1 : 0;
assign detect_min[427][6] = (mid_1[3431:3424] < top_2[3423:3416]) ? 1 : 0;
assign detect_min[427][7] = (mid_1[3431:3424] < top_2[3431:3424]) ? 1 : 0;
assign detect_min[427][8] = (mid_1[3431:3424] < top_2[3439:3432]) ? 1 : 0;
assign detect_min[427][9] = (mid_1[3431:3424] < mid_0[3423:3416]) ? 1 : 0;
assign detect_min[427][10] = (mid_1[3431:3424] < mid_0[3431:3424]) ? 1 : 0;
assign detect_min[427][11] = (mid_1[3431:3424] < mid_0[3439:3432]) ? 1 : 0;
assign detect_min[427][12] = (mid_1[3431:3424] < mid_1[3423:3416]) ? 1 : 0;
assign detect_min[427][13] = (mid_1[3431:3424] < mid_1[3439:3432]) ? 1 : 0;
assign detect_min[427][14] = (mid_1[3431:3424] < mid_2[3423:3416]) ? 1 : 0;
assign detect_min[427][15] = (mid_1[3431:3424] < mid_2[3431:3424]) ? 1 : 0;
assign detect_min[427][16] = (mid_1[3431:3424] < mid_2[3439:3432]) ? 1 : 0;
assign detect_min[427][17] = (mid_1[3431:3424] < btm_0[3423:3416]) ? 1 : 0;
assign detect_min[427][18] = (mid_1[3431:3424] < btm_0[3431:3424]) ? 1 : 0;
assign detect_min[427][19] = (mid_1[3431:3424] < btm_0[3439:3432]) ? 1 : 0;
assign detect_min[427][20] = (mid_1[3431:3424] < btm_1[3423:3416]) ? 1 : 0;
assign detect_min[427][21] = (mid_1[3431:3424] < btm_1[3431:3424]) ? 1 : 0;
assign detect_min[427][22] = (mid_1[3431:3424] < btm_1[3439:3432]) ? 1 : 0;
assign detect_min[427][23] = (mid_1[3431:3424] < btm_2[3423:3416]) ? 1 : 0;
assign detect_min[427][24] = (mid_1[3431:3424] < btm_2[3431:3424]) ? 1 : 0;
assign detect_min[427][25] = (mid_1[3431:3424] < btm_2[3439:3432]) ? 1 : 0;

assign detect_min[428][0] = (mid_1[3439:3432] < top_0[3431:3424]) ? 1 : 0;
assign detect_min[428][1] = (mid_1[3439:3432] < top_0[3439:3432]) ? 1 : 0;
assign detect_min[428][2] = (mid_1[3439:3432] < top_0[3447:3440]) ? 1 : 0;
assign detect_min[428][3] = (mid_1[3439:3432] < top_1[3431:3424]) ? 1 : 0;
assign detect_min[428][4] = (mid_1[3439:3432] < top_1[3439:3432]) ? 1 : 0;
assign detect_min[428][5] = (mid_1[3439:3432] < top_1[3447:3440]) ? 1 : 0;
assign detect_min[428][6] = (mid_1[3439:3432] < top_2[3431:3424]) ? 1 : 0;
assign detect_min[428][7] = (mid_1[3439:3432] < top_2[3439:3432]) ? 1 : 0;
assign detect_min[428][8] = (mid_1[3439:3432] < top_2[3447:3440]) ? 1 : 0;
assign detect_min[428][9] = (mid_1[3439:3432] < mid_0[3431:3424]) ? 1 : 0;
assign detect_min[428][10] = (mid_1[3439:3432] < mid_0[3439:3432]) ? 1 : 0;
assign detect_min[428][11] = (mid_1[3439:3432] < mid_0[3447:3440]) ? 1 : 0;
assign detect_min[428][12] = (mid_1[3439:3432] < mid_1[3431:3424]) ? 1 : 0;
assign detect_min[428][13] = (mid_1[3439:3432] < mid_1[3447:3440]) ? 1 : 0;
assign detect_min[428][14] = (mid_1[3439:3432] < mid_2[3431:3424]) ? 1 : 0;
assign detect_min[428][15] = (mid_1[3439:3432] < mid_2[3439:3432]) ? 1 : 0;
assign detect_min[428][16] = (mid_1[3439:3432] < mid_2[3447:3440]) ? 1 : 0;
assign detect_min[428][17] = (mid_1[3439:3432] < btm_0[3431:3424]) ? 1 : 0;
assign detect_min[428][18] = (mid_1[3439:3432] < btm_0[3439:3432]) ? 1 : 0;
assign detect_min[428][19] = (mid_1[3439:3432] < btm_0[3447:3440]) ? 1 : 0;
assign detect_min[428][20] = (mid_1[3439:3432] < btm_1[3431:3424]) ? 1 : 0;
assign detect_min[428][21] = (mid_1[3439:3432] < btm_1[3439:3432]) ? 1 : 0;
assign detect_min[428][22] = (mid_1[3439:3432] < btm_1[3447:3440]) ? 1 : 0;
assign detect_min[428][23] = (mid_1[3439:3432] < btm_2[3431:3424]) ? 1 : 0;
assign detect_min[428][24] = (mid_1[3439:3432] < btm_2[3439:3432]) ? 1 : 0;
assign detect_min[428][25] = (mid_1[3439:3432] < btm_2[3447:3440]) ? 1 : 0;

assign detect_min[429][0] = (mid_1[3447:3440] < top_0[3439:3432]) ? 1 : 0;
assign detect_min[429][1] = (mid_1[3447:3440] < top_0[3447:3440]) ? 1 : 0;
assign detect_min[429][2] = (mid_1[3447:3440] < top_0[3455:3448]) ? 1 : 0;
assign detect_min[429][3] = (mid_1[3447:3440] < top_1[3439:3432]) ? 1 : 0;
assign detect_min[429][4] = (mid_1[3447:3440] < top_1[3447:3440]) ? 1 : 0;
assign detect_min[429][5] = (mid_1[3447:3440] < top_1[3455:3448]) ? 1 : 0;
assign detect_min[429][6] = (mid_1[3447:3440] < top_2[3439:3432]) ? 1 : 0;
assign detect_min[429][7] = (mid_1[3447:3440] < top_2[3447:3440]) ? 1 : 0;
assign detect_min[429][8] = (mid_1[3447:3440] < top_2[3455:3448]) ? 1 : 0;
assign detect_min[429][9] = (mid_1[3447:3440] < mid_0[3439:3432]) ? 1 : 0;
assign detect_min[429][10] = (mid_1[3447:3440] < mid_0[3447:3440]) ? 1 : 0;
assign detect_min[429][11] = (mid_1[3447:3440] < mid_0[3455:3448]) ? 1 : 0;
assign detect_min[429][12] = (mid_1[3447:3440] < mid_1[3439:3432]) ? 1 : 0;
assign detect_min[429][13] = (mid_1[3447:3440] < mid_1[3455:3448]) ? 1 : 0;
assign detect_min[429][14] = (mid_1[3447:3440] < mid_2[3439:3432]) ? 1 : 0;
assign detect_min[429][15] = (mid_1[3447:3440] < mid_2[3447:3440]) ? 1 : 0;
assign detect_min[429][16] = (mid_1[3447:3440] < mid_2[3455:3448]) ? 1 : 0;
assign detect_min[429][17] = (mid_1[3447:3440] < btm_0[3439:3432]) ? 1 : 0;
assign detect_min[429][18] = (mid_1[3447:3440] < btm_0[3447:3440]) ? 1 : 0;
assign detect_min[429][19] = (mid_1[3447:3440] < btm_0[3455:3448]) ? 1 : 0;
assign detect_min[429][20] = (mid_1[3447:3440] < btm_1[3439:3432]) ? 1 : 0;
assign detect_min[429][21] = (mid_1[3447:3440] < btm_1[3447:3440]) ? 1 : 0;
assign detect_min[429][22] = (mid_1[3447:3440] < btm_1[3455:3448]) ? 1 : 0;
assign detect_min[429][23] = (mid_1[3447:3440] < btm_2[3439:3432]) ? 1 : 0;
assign detect_min[429][24] = (mid_1[3447:3440] < btm_2[3447:3440]) ? 1 : 0;
assign detect_min[429][25] = (mid_1[3447:3440] < btm_2[3455:3448]) ? 1 : 0;

assign detect_min[430][0] = (mid_1[3455:3448] < top_0[3447:3440]) ? 1 : 0;
assign detect_min[430][1] = (mid_1[3455:3448] < top_0[3455:3448]) ? 1 : 0;
assign detect_min[430][2] = (mid_1[3455:3448] < top_0[3463:3456]) ? 1 : 0;
assign detect_min[430][3] = (mid_1[3455:3448] < top_1[3447:3440]) ? 1 : 0;
assign detect_min[430][4] = (mid_1[3455:3448] < top_1[3455:3448]) ? 1 : 0;
assign detect_min[430][5] = (mid_1[3455:3448] < top_1[3463:3456]) ? 1 : 0;
assign detect_min[430][6] = (mid_1[3455:3448] < top_2[3447:3440]) ? 1 : 0;
assign detect_min[430][7] = (mid_1[3455:3448] < top_2[3455:3448]) ? 1 : 0;
assign detect_min[430][8] = (mid_1[3455:3448] < top_2[3463:3456]) ? 1 : 0;
assign detect_min[430][9] = (mid_1[3455:3448] < mid_0[3447:3440]) ? 1 : 0;
assign detect_min[430][10] = (mid_1[3455:3448] < mid_0[3455:3448]) ? 1 : 0;
assign detect_min[430][11] = (mid_1[3455:3448] < mid_0[3463:3456]) ? 1 : 0;
assign detect_min[430][12] = (mid_1[3455:3448] < mid_1[3447:3440]) ? 1 : 0;
assign detect_min[430][13] = (mid_1[3455:3448] < mid_1[3463:3456]) ? 1 : 0;
assign detect_min[430][14] = (mid_1[3455:3448] < mid_2[3447:3440]) ? 1 : 0;
assign detect_min[430][15] = (mid_1[3455:3448] < mid_2[3455:3448]) ? 1 : 0;
assign detect_min[430][16] = (mid_1[3455:3448] < mid_2[3463:3456]) ? 1 : 0;
assign detect_min[430][17] = (mid_1[3455:3448] < btm_0[3447:3440]) ? 1 : 0;
assign detect_min[430][18] = (mid_1[3455:3448] < btm_0[3455:3448]) ? 1 : 0;
assign detect_min[430][19] = (mid_1[3455:3448] < btm_0[3463:3456]) ? 1 : 0;
assign detect_min[430][20] = (mid_1[3455:3448] < btm_1[3447:3440]) ? 1 : 0;
assign detect_min[430][21] = (mid_1[3455:3448] < btm_1[3455:3448]) ? 1 : 0;
assign detect_min[430][22] = (mid_1[3455:3448] < btm_1[3463:3456]) ? 1 : 0;
assign detect_min[430][23] = (mid_1[3455:3448] < btm_2[3447:3440]) ? 1 : 0;
assign detect_min[430][24] = (mid_1[3455:3448] < btm_2[3455:3448]) ? 1 : 0;
assign detect_min[430][25] = (mid_1[3455:3448] < btm_2[3463:3456]) ? 1 : 0;

assign detect_min[431][0] = (mid_1[3463:3456] < top_0[3455:3448]) ? 1 : 0;
assign detect_min[431][1] = (mid_1[3463:3456] < top_0[3463:3456]) ? 1 : 0;
assign detect_min[431][2] = (mid_1[3463:3456] < top_0[3471:3464]) ? 1 : 0;
assign detect_min[431][3] = (mid_1[3463:3456] < top_1[3455:3448]) ? 1 : 0;
assign detect_min[431][4] = (mid_1[3463:3456] < top_1[3463:3456]) ? 1 : 0;
assign detect_min[431][5] = (mid_1[3463:3456] < top_1[3471:3464]) ? 1 : 0;
assign detect_min[431][6] = (mid_1[3463:3456] < top_2[3455:3448]) ? 1 : 0;
assign detect_min[431][7] = (mid_1[3463:3456] < top_2[3463:3456]) ? 1 : 0;
assign detect_min[431][8] = (mid_1[3463:3456] < top_2[3471:3464]) ? 1 : 0;
assign detect_min[431][9] = (mid_1[3463:3456] < mid_0[3455:3448]) ? 1 : 0;
assign detect_min[431][10] = (mid_1[3463:3456] < mid_0[3463:3456]) ? 1 : 0;
assign detect_min[431][11] = (mid_1[3463:3456] < mid_0[3471:3464]) ? 1 : 0;
assign detect_min[431][12] = (mid_1[3463:3456] < mid_1[3455:3448]) ? 1 : 0;
assign detect_min[431][13] = (mid_1[3463:3456] < mid_1[3471:3464]) ? 1 : 0;
assign detect_min[431][14] = (mid_1[3463:3456] < mid_2[3455:3448]) ? 1 : 0;
assign detect_min[431][15] = (mid_1[3463:3456] < mid_2[3463:3456]) ? 1 : 0;
assign detect_min[431][16] = (mid_1[3463:3456] < mid_2[3471:3464]) ? 1 : 0;
assign detect_min[431][17] = (mid_1[3463:3456] < btm_0[3455:3448]) ? 1 : 0;
assign detect_min[431][18] = (mid_1[3463:3456] < btm_0[3463:3456]) ? 1 : 0;
assign detect_min[431][19] = (mid_1[3463:3456] < btm_0[3471:3464]) ? 1 : 0;
assign detect_min[431][20] = (mid_1[3463:3456] < btm_1[3455:3448]) ? 1 : 0;
assign detect_min[431][21] = (mid_1[3463:3456] < btm_1[3463:3456]) ? 1 : 0;
assign detect_min[431][22] = (mid_1[3463:3456] < btm_1[3471:3464]) ? 1 : 0;
assign detect_min[431][23] = (mid_1[3463:3456] < btm_2[3455:3448]) ? 1 : 0;
assign detect_min[431][24] = (mid_1[3463:3456] < btm_2[3463:3456]) ? 1 : 0;
assign detect_min[431][25] = (mid_1[3463:3456] < btm_2[3471:3464]) ? 1 : 0;

assign detect_min[432][0] = (mid_1[3471:3464] < top_0[3463:3456]) ? 1 : 0;
assign detect_min[432][1] = (mid_1[3471:3464] < top_0[3471:3464]) ? 1 : 0;
assign detect_min[432][2] = (mid_1[3471:3464] < top_0[3479:3472]) ? 1 : 0;
assign detect_min[432][3] = (mid_1[3471:3464] < top_1[3463:3456]) ? 1 : 0;
assign detect_min[432][4] = (mid_1[3471:3464] < top_1[3471:3464]) ? 1 : 0;
assign detect_min[432][5] = (mid_1[3471:3464] < top_1[3479:3472]) ? 1 : 0;
assign detect_min[432][6] = (mid_1[3471:3464] < top_2[3463:3456]) ? 1 : 0;
assign detect_min[432][7] = (mid_1[3471:3464] < top_2[3471:3464]) ? 1 : 0;
assign detect_min[432][8] = (mid_1[3471:3464] < top_2[3479:3472]) ? 1 : 0;
assign detect_min[432][9] = (mid_1[3471:3464] < mid_0[3463:3456]) ? 1 : 0;
assign detect_min[432][10] = (mid_1[3471:3464] < mid_0[3471:3464]) ? 1 : 0;
assign detect_min[432][11] = (mid_1[3471:3464] < mid_0[3479:3472]) ? 1 : 0;
assign detect_min[432][12] = (mid_1[3471:3464] < mid_1[3463:3456]) ? 1 : 0;
assign detect_min[432][13] = (mid_1[3471:3464] < mid_1[3479:3472]) ? 1 : 0;
assign detect_min[432][14] = (mid_1[3471:3464] < mid_2[3463:3456]) ? 1 : 0;
assign detect_min[432][15] = (mid_1[3471:3464] < mid_2[3471:3464]) ? 1 : 0;
assign detect_min[432][16] = (mid_1[3471:3464] < mid_2[3479:3472]) ? 1 : 0;
assign detect_min[432][17] = (mid_1[3471:3464] < btm_0[3463:3456]) ? 1 : 0;
assign detect_min[432][18] = (mid_1[3471:3464] < btm_0[3471:3464]) ? 1 : 0;
assign detect_min[432][19] = (mid_1[3471:3464] < btm_0[3479:3472]) ? 1 : 0;
assign detect_min[432][20] = (mid_1[3471:3464] < btm_1[3463:3456]) ? 1 : 0;
assign detect_min[432][21] = (mid_1[3471:3464] < btm_1[3471:3464]) ? 1 : 0;
assign detect_min[432][22] = (mid_1[3471:3464] < btm_1[3479:3472]) ? 1 : 0;
assign detect_min[432][23] = (mid_1[3471:3464] < btm_2[3463:3456]) ? 1 : 0;
assign detect_min[432][24] = (mid_1[3471:3464] < btm_2[3471:3464]) ? 1 : 0;
assign detect_min[432][25] = (mid_1[3471:3464] < btm_2[3479:3472]) ? 1 : 0;

assign detect_min[433][0] = (mid_1[3479:3472] < top_0[3471:3464]) ? 1 : 0;
assign detect_min[433][1] = (mid_1[3479:3472] < top_0[3479:3472]) ? 1 : 0;
assign detect_min[433][2] = (mid_1[3479:3472] < top_0[3487:3480]) ? 1 : 0;
assign detect_min[433][3] = (mid_1[3479:3472] < top_1[3471:3464]) ? 1 : 0;
assign detect_min[433][4] = (mid_1[3479:3472] < top_1[3479:3472]) ? 1 : 0;
assign detect_min[433][5] = (mid_1[3479:3472] < top_1[3487:3480]) ? 1 : 0;
assign detect_min[433][6] = (mid_1[3479:3472] < top_2[3471:3464]) ? 1 : 0;
assign detect_min[433][7] = (mid_1[3479:3472] < top_2[3479:3472]) ? 1 : 0;
assign detect_min[433][8] = (mid_1[3479:3472] < top_2[3487:3480]) ? 1 : 0;
assign detect_min[433][9] = (mid_1[3479:3472] < mid_0[3471:3464]) ? 1 : 0;
assign detect_min[433][10] = (mid_1[3479:3472] < mid_0[3479:3472]) ? 1 : 0;
assign detect_min[433][11] = (mid_1[3479:3472] < mid_0[3487:3480]) ? 1 : 0;
assign detect_min[433][12] = (mid_1[3479:3472] < mid_1[3471:3464]) ? 1 : 0;
assign detect_min[433][13] = (mid_1[3479:3472] < mid_1[3487:3480]) ? 1 : 0;
assign detect_min[433][14] = (mid_1[3479:3472] < mid_2[3471:3464]) ? 1 : 0;
assign detect_min[433][15] = (mid_1[3479:3472] < mid_2[3479:3472]) ? 1 : 0;
assign detect_min[433][16] = (mid_1[3479:3472] < mid_2[3487:3480]) ? 1 : 0;
assign detect_min[433][17] = (mid_1[3479:3472] < btm_0[3471:3464]) ? 1 : 0;
assign detect_min[433][18] = (mid_1[3479:3472] < btm_0[3479:3472]) ? 1 : 0;
assign detect_min[433][19] = (mid_1[3479:3472] < btm_0[3487:3480]) ? 1 : 0;
assign detect_min[433][20] = (mid_1[3479:3472] < btm_1[3471:3464]) ? 1 : 0;
assign detect_min[433][21] = (mid_1[3479:3472] < btm_1[3479:3472]) ? 1 : 0;
assign detect_min[433][22] = (mid_1[3479:3472] < btm_1[3487:3480]) ? 1 : 0;
assign detect_min[433][23] = (mid_1[3479:3472] < btm_2[3471:3464]) ? 1 : 0;
assign detect_min[433][24] = (mid_1[3479:3472] < btm_2[3479:3472]) ? 1 : 0;
assign detect_min[433][25] = (mid_1[3479:3472] < btm_2[3487:3480]) ? 1 : 0;

assign detect_min[434][0] = (mid_1[3487:3480] < top_0[3479:3472]) ? 1 : 0;
assign detect_min[434][1] = (mid_1[3487:3480] < top_0[3487:3480]) ? 1 : 0;
assign detect_min[434][2] = (mid_1[3487:3480] < top_0[3495:3488]) ? 1 : 0;
assign detect_min[434][3] = (mid_1[3487:3480] < top_1[3479:3472]) ? 1 : 0;
assign detect_min[434][4] = (mid_1[3487:3480] < top_1[3487:3480]) ? 1 : 0;
assign detect_min[434][5] = (mid_1[3487:3480] < top_1[3495:3488]) ? 1 : 0;
assign detect_min[434][6] = (mid_1[3487:3480] < top_2[3479:3472]) ? 1 : 0;
assign detect_min[434][7] = (mid_1[3487:3480] < top_2[3487:3480]) ? 1 : 0;
assign detect_min[434][8] = (mid_1[3487:3480] < top_2[3495:3488]) ? 1 : 0;
assign detect_min[434][9] = (mid_1[3487:3480] < mid_0[3479:3472]) ? 1 : 0;
assign detect_min[434][10] = (mid_1[3487:3480] < mid_0[3487:3480]) ? 1 : 0;
assign detect_min[434][11] = (mid_1[3487:3480] < mid_0[3495:3488]) ? 1 : 0;
assign detect_min[434][12] = (mid_1[3487:3480] < mid_1[3479:3472]) ? 1 : 0;
assign detect_min[434][13] = (mid_1[3487:3480] < mid_1[3495:3488]) ? 1 : 0;
assign detect_min[434][14] = (mid_1[3487:3480] < mid_2[3479:3472]) ? 1 : 0;
assign detect_min[434][15] = (mid_1[3487:3480] < mid_2[3487:3480]) ? 1 : 0;
assign detect_min[434][16] = (mid_1[3487:3480] < mid_2[3495:3488]) ? 1 : 0;
assign detect_min[434][17] = (mid_1[3487:3480] < btm_0[3479:3472]) ? 1 : 0;
assign detect_min[434][18] = (mid_1[3487:3480] < btm_0[3487:3480]) ? 1 : 0;
assign detect_min[434][19] = (mid_1[3487:3480] < btm_0[3495:3488]) ? 1 : 0;
assign detect_min[434][20] = (mid_1[3487:3480] < btm_1[3479:3472]) ? 1 : 0;
assign detect_min[434][21] = (mid_1[3487:3480] < btm_1[3487:3480]) ? 1 : 0;
assign detect_min[434][22] = (mid_1[3487:3480] < btm_1[3495:3488]) ? 1 : 0;
assign detect_min[434][23] = (mid_1[3487:3480] < btm_2[3479:3472]) ? 1 : 0;
assign detect_min[434][24] = (mid_1[3487:3480] < btm_2[3487:3480]) ? 1 : 0;
assign detect_min[434][25] = (mid_1[3487:3480] < btm_2[3495:3488]) ? 1 : 0;

assign detect_min[435][0] = (mid_1[3495:3488] < top_0[3487:3480]) ? 1 : 0;
assign detect_min[435][1] = (mid_1[3495:3488] < top_0[3495:3488]) ? 1 : 0;
assign detect_min[435][2] = (mid_1[3495:3488] < top_0[3503:3496]) ? 1 : 0;
assign detect_min[435][3] = (mid_1[3495:3488] < top_1[3487:3480]) ? 1 : 0;
assign detect_min[435][4] = (mid_1[3495:3488] < top_1[3495:3488]) ? 1 : 0;
assign detect_min[435][5] = (mid_1[3495:3488] < top_1[3503:3496]) ? 1 : 0;
assign detect_min[435][6] = (mid_1[3495:3488] < top_2[3487:3480]) ? 1 : 0;
assign detect_min[435][7] = (mid_1[3495:3488] < top_2[3495:3488]) ? 1 : 0;
assign detect_min[435][8] = (mid_1[3495:3488] < top_2[3503:3496]) ? 1 : 0;
assign detect_min[435][9] = (mid_1[3495:3488] < mid_0[3487:3480]) ? 1 : 0;
assign detect_min[435][10] = (mid_1[3495:3488] < mid_0[3495:3488]) ? 1 : 0;
assign detect_min[435][11] = (mid_1[3495:3488] < mid_0[3503:3496]) ? 1 : 0;
assign detect_min[435][12] = (mid_1[3495:3488] < mid_1[3487:3480]) ? 1 : 0;
assign detect_min[435][13] = (mid_1[3495:3488] < mid_1[3503:3496]) ? 1 : 0;
assign detect_min[435][14] = (mid_1[3495:3488] < mid_2[3487:3480]) ? 1 : 0;
assign detect_min[435][15] = (mid_1[3495:3488] < mid_2[3495:3488]) ? 1 : 0;
assign detect_min[435][16] = (mid_1[3495:3488] < mid_2[3503:3496]) ? 1 : 0;
assign detect_min[435][17] = (mid_1[3495:3488] < btm_0[3487:3480]) ? 1 : 0;
assign detect_min[435][18] = (mid_1[3495:3488] < btm_0[3495:3488]) ? 1 : 0;
assign detect_min[435][19] = (mid_1[3495:3488] < btm_0[3503:3496]) ? 1 : 0;
assign detect_min[435][20] = (mid_1[3495:3488] < btm_1[3487:3480]) ? 1 : 0;
assign detect_min[435][21] = (mid_1[3495:3488] < btm_1[3495:3488]) ? 1 : 0;
assign detect_min[435][22] = (mid_1[3495:3488] < btm_1[3503:3496]) ? 1 : 0;
assign detect_min[435][23] = (mid_1[3495:3488] < btm_2[3487:3480]) ? 1 : 0;
assign detect_min[435][24] = (mid_1[3495:3488] < btm_2[3495:3488]) ? 1 : 0;
assign detect_min[435][25] = (mid_1[3495:3488] < btm_2[3503:3496]) ? 1 : 0;

assign detect_min[436][0] = (mid_1[3503:3496] < top_0[3495:3488]) ? 1 : 0;
assign detect_min[436][1] = (mid_1[3503:3496] < top_0[3503:3496]) ? 1 : 0;
assign detect_min[436][2] = (mid_1[3503:3496] < top_0[3511:3504]) ? 1 : 0;
assign detect_min[436][3] = (mid_1[3503:3496] < top_1[3495:3488]) ? 1 : 0;
assign detect_min[436][4] = (mid_1[3503:3496] < top_1[3503:3496]) ? 1 : 0;
assign detect_min[436][5] = (mid_1[3503:3496] < top_1[3511:3504]) ? 1 : 0;
assign detect_min[436][6] = (mid_1[3503:3496] < top_2[3495:3488]) ? 1 : 0;
assign detect_min[436][7] = (mid_1[3503:3496] < top_2[3503:3496]) ? 1 : 0;
assign detect_min[436][8] = (mid_1[3503:3496] < top_2[3511:3504]) ? 1 : 0;
assign detect_min[436][9] = (mid_1[3503:3496] < mid_0[3495:3488]) ? 1 : 0;
assign detect_min[436][10] = (mid_1[3503:3496] < mid_0[3503:3496]) ? 1 : 0;
assign detect_min[436][11] = (mid_1[3503:3496] < mid_0[3511:3504]) ? 1 : 0;
assign detect_min[436][12] = (mid_1[3503:3496] < mid_1[3495:3488]) ? 1 : 0;
assign detect_min[436][13] = (mid_1[3503:3496] < mid_1[3511:3504]) ? 1 : 0;
assign detect_min[436][14] = (mid_1[3503:3496] < mid_2[3495:3488]) ? 1 : 0;
assign detect_min[436][15] = (mid_1[3503:3496] < mid_2[3503:3496]) ? 1 : 0;
assign detect_min[436][16] = (mid_1[3503:3496] < mid_2[3511:3504]) ? 1 : 0;
assign detect_min[436][17] = (mid_1[3503:3496] < btm_0[3495:3488]) ? 1 : 0;
assign detect_min[436][18] = (mid_1[3503:3496] < btm_0[3503:3496]) ? 1 : 0;
assign detect_min[436][19] = (mid_1[3503:3496] < btm_0[3511:3504]) ? 1 : 0;
assign detect_min[436][20] = (mid_1[3503:3496] < btm_1[3495:3488]) ? 1 : 0;
assign detect_min[436][21] = (mid_1[3503:3496] < btm_1[3503:3496]) ? 1 : 0;
assign detect_min[436][22] = (mid_1[3503:3496] < btm_1[3511:3504]) ? 1 : 0;
assign detect_min[436][23] = (mid_1[3503:3496] < btm_2[3495:3488]) ? 1 : 0;
assign detect_min[436][24] = (mid_1[3503:3496] < btm_2[3503:3496]) ? 1 : 0;
assign detect_min[436][25] = (mid_1[3503:3496] < btm_2[3511:3504]) ? 1 : 0;

assign detect_min[437][0] = (mid_1[3511:3504] < top_0[3503:3496]) ? 1 : 0;
assign detect_min[437][1] = (mid_1[3511:3504] < top_0[3511:3504]) ? 1 : 0;
assign detect_min[437][2] = (mid_1[3511:3504] < top_0[3519:3512]) ? 1 : 0;
assign detect_min[437][3] = (mid_1[3511:3504] < top_1[3503:3496]) ? 1 : 0;
assign detect_min[437][4] = (mid_1[3511:3504] < top_1[3511:3504]) ? 1 : 0;
assign detect_min[437][5] = (mid_1[3511:3504] < top_1[3519:3512]) ? 1 : 0;
assign detect_min[437][6] = (mid_1[3511:3504] < top_2[3503:3496]) ? 1 : 0;
assign detect_min[437][7] = (mid_1[3511:3504] < top_2[3511:3504]) ? 1 : 0;
assign detect_min[437][8] = (mid_1[3511:3504] < top_2[3519:3512]) ? 1 : 0;
assign detect_min[437][9] = (mid_1[3511:3504] < mid_0[3503:3496]) ? 1 : 0;
assign detect_min[437][10] = (mid_1[3511:3504] < mid_0[3511:3504]) ? 1 : 0;
assign detect_min[437][11] = (mid_1[3511:3504] < mid_0[3519:3512]) ? 1 : 0;
assign detect_min[437][12] = (mid_1[3511:3504] < mid_1[3503:3496]) ? 1 : 0;
assign detect_min[437][13] = (mid_1[3511:3504] < mid_1[3519:3512]) ? 1 : 0;
assign detect_min[437][14] = (mid_1[3511:3504] < mid_2[3503:3496]) ? 1 : 0;
assign detect_min[437][15] = (mid_1[3511:3504] < mid_2[3511:3504]) ? 1 : 0;
assign detect_min[437][16] = (mid_1[3511:3504] < mid_2[3519:3512]) ? 1 : 0;
assign detect_min[437][17] = (mid_1[3511:3504] < btm_0[3503:3496]) ? 1 : 0;
assign detect_min[437][18] = (mid_1[3511:3504] < btm_0[3511:3504]) ? 1 : 0;
assign detect_min[437][19] = (mid_1[3511:3504] < btm_0[3519:3512]) ? 1 : 0;
assign detect_min[437][20] = (mid_1[3511:3504] < btm_1[3503:3496]) ? 1 : 0;
assign detect_min[437][21] = (mid_1[3511:3504] < btm_1[3511:3504]) ? 1 : 0;
assign detect_min[437][22] = (mid_1[3511:3504] < btm_1[3519:3512]) ? 1 : 0;
assign detect_min[437][23] = (mid_1[3511:3504] < btm_2[3503:3496]) ? 1 : 0;
assign detect_min[437][24] = (mid_1[3511:3504] < btm_2[3511:3504]) ? 1 : 0;
assign detect_min[437][25] = (mid_1[3511:3504] < btm_2[3519:3512]) ? 1 : 0;

assign detect_min[438][0] = (mid_1[3519:3512] < top_0[3511:3504]) ? 1 : 0;
assign detect_min[438][1] = (mid_1[3519:3512] < top_0[3519:3512]) ? 1 : 0;
assign detect_min[438][2] = (mid_1[3519:3512] < top_0[3527:3520]) ? 1 : 0;
assign detect_min[438][3] = (mid_1[3519:3512] < top_1[3511:3504]) ? 1 : 0;
assign detect_min[438][4] = (mid_1[3519:3512] < top_1[3519:3512]) ? 1 : 0;
assign detect_min[438][5] = (mid_1[3519:3512] < top_1[3527:3520]) ? 1 : 0;
assign detect_min[438][6] = (mid_1[3519:3512] < top_2[3511:3504]) ? 1 : 0;
assign detect_min[438][7] = (mid_1[3519:3512] < top_2[3519:3512]) ? 1 : 0;
assign detect_min[438][8] = (mid_1[3519:3512] < top_2[3527:3520]) ? 1 : 0;
assign detect_min[438][9] = (mid_1[3519:3512] < mid_0[3511:3504]) ? 1 : 0;
assign detect_min[438][10] = (mid_1[3519:3512] < mid_0[3519:3512]) ? 1 : 0;
assign detect_min[438][11] = (mid_1[3519:3512] < mid_0[3527:3520]) ? 1 : 0;
assign detect_min[438][12] = (mid_1[3519:3512] < mid_1[3511:3504]) ? 1 : 0;
assign detect_min[438][13] = (mid_1[3519:3512] < mid_1[3527:3520]) ? 1 : 0;
assign detect_min[438][14] = (mid_1[3519:3512] < mid_2[3511:3504]) ? 1 : 0;
assign detect_min[438][15] = (mid_1[3519:3512] < mid_2[3519:3512]) ? 1 : 0;
assign detect_min[438][16] = (mid_1[3519:3512] < mid_2[3527:3520]) ? 1 : 0;
assign detect_min[438][17] = (mid_1[3519:3512] < btm_0[3511:3504]) ? 1 : 0;
assign detect_min[438][18] = (mid_1[3519:3512] < btm_0[3519:3512]) ? 1 : 0;
assign detect_min[438][19] = (mid_1[3519:3512] < btm_0[3527:3520]) ? 1 : 0;
assign detect_min[438][20] = (mid_1[3519:3512] < btm_1[3511:3504]) ? 1 : 0;
assign detect_min[438][21] = (mid_1[3519:3512] < btm_1[3519:3512]) ? 1 : 0;
assign detect_min[438][22] = (mid_1[3519:3512] < btm_1[3527:3520]) ? 1 : 0;
assign detect_min[438][23] = (mid_1[3519:3512] < btm_2[3511:3504]) ? 1 : 0;
assign detect_min[438][24] = (mid_1[3519:3512] < btm_2[3519:3512]) ? 1 : 0;
assign detect_min[438][25] = (mid_1[3519:3512] < btm_2[3527:3520]) ? 1 : 0;

assign detect_min[439][0] = (mid_1[3527:3520] < top_0[3519:3512]) ? 1 : 0;
assign detect_min[439][1] = (mid_1[3527:3520] < top_0[3527:3520]) ? 1 : 0;
assign detect_min[439][2] = (mid_1[3527:3520] < top_0[3535:3528]) ? 1 : 0;
assign detect_min[439][3] = (mid_1[3527:3520] < top_1[3519:3512]) ? 1 : 0;
assign detect_min[439][4] = (mid_1[3527:3520] < top_1[3527:3520]) ? 1 : 0;
assign detect_min[439][5] = (mid_1[3527:3520] < top_1[3535:3528]) ? 1 : 0;
assign detect_min[439][6] = (mid_1[3527:3520] < top_2[3519:3512]) ? 1 : 0;
assign detect_min[439][7] = (mid_1[3527:3520] < top_2[3527:3520]) ? 1 : 0;
assign detect_min[439][8] = (mid_1[3527:3520] < top_2[3535:3528]) ? 1 : 0;
assign detect_min[439][9] = (mid_1[3527:3520] < mid_0[3519:3512]) ? 1 : 0;
assign detect_min[439][10] = (mid_1[3527:3520] < mid_0[3527:3520]) ? 1 : 0;
assign detect_min[439][11] = (mid_1[3527:3520] < mid_0[3535:3528]) ? 1 : 0;
assign detect_min[439][12] = (mid_1[3527:3520] < mid_1[3519:3512]) ? 1 : 0;
assign detect_min[439][13] = (mid_1[3527:3520] < mid_1[3535:3528]) ? 1 : 0;
assign detect_min[439][14] = (mid_1[3527:3520] < mid_2[3519:3512]) ? 1 : 0;
assign detect_min[439][15] = (mid_1[3527:3520] < mid_2[3527:3520]) ? 1 : 0;
assign detect_min[439][16] = (mid_1[3527:3520] < mid_2[3535:3528]) ? 1 : 0;
assign detect_min[439][17] = (mid_1[3527:3520] < btm_0[3519:3512]) ? 1 : 0;
assign detect_min[439][18] = (mid_1[3527:3520] < btm_0[3527:3520]) ? 1 : 0;
assign detect_min[439][19] = (mid_1[3527:3520] < btm_0[3535:3528]) ? 1 : 0;
assign detect_min[439][20] = (mid_1[3527:3520] < btm_1[3519:3512]) ? 1 : 0;
assign detect_min[439][21] = (mid_1[3527:3520] < btm_1[3527:3520]) ? 1 : 0;
assign detect_min[439][22] = (mid_1[3527:3520] < btm_1[3535:3528]) ? 1 : 0;
assign detect_min[439][23] = (mid_1[3527:3520] < btm_2[3519:3512]) ? 1 : 0;
assign detect_min[439][24] = (mid_1[3527:3520] < btm_2[3527:3520]) ? 1 : 0;
assign detect_min[439][25] = (mid_1[3527:3520] < btm_2[3535:3528]) ? 1 : 0;

assign detect_min[440][0] = (mid_1[3535:3528] < top_0[3527:3520]) ? 1 : 0;
assign detect_min[440][1] = (mid_1[3535:3528] < top_0[3535:3528]) ? 1 : 0;
assign detect_min[440][2] = (mid_1[3535:3528] < top_0[3543:3536]) ? 1 : 0;
assign detect_min[440][3] = (mid_1[3535:3528] < top_1[3527:3520]) ? 1 : 0;
assign detect_min[440][4] = (mid_1[3535:3528] < top_1[3535:3528]) ? 1 : 0;
assign detect_min[440][5] = (mid_1[3535:3528] < top_1[3543:3536]) ? 1 : 0;
assign detect_min[440][6] = (mid_1[3535:3528] < top_2[3527:3520]) ? 1 : 0;
assign detect_min[440][7] = (mid_1[3535:3528] < top_2[3535:3528]) ? 1 : 0;
assign detect_min[440][8] = (mid_1[3535:3528] < top_2[3543:3536]) ? 1 : 0;
assign detect_min[440][9] = (mid_1[3535:3528] < mid_0[3527:3520]) ? 1 : 0;
assign detect_min[440][10] = (mid_1[3535:3528] < mid_0[3535:3528]) ? 1 : 0;
assign detect_min[440][11] = (mid_1[3535:3528] < mid_0[3543:3536]) ? 1 : 0;
assign detect_min[440][12] = (mid_1[3535:3528] < mid_1[3527:3520]) ? 1 : 0;
assign detect_min[440][13] = (mid_1[3535:3528] < mid_1[3543:3536]) ? 1 : 0;
assign detect_min[440][14] = (mid_1[3535:3528] < mid_2[3527:3520]) ? 1 : 0;
assign detect_min[440][15] = (mid_1[3535:3528] < mid_2[3535:3528]) ? 1 : 0;
assign detect_min[440][16] = (mid_1[3535:3528] < mid_2[3543:3536]) ? 1 : 0;
assign detect_min[440][17] = (mid_1[3535:3528] < btm_0[3527:3520]) ? 1 : 0;
assign detect_min[440][18] = (mid_1[3535:3528] < btm_0[3535:3528]) ? 1 : 0;
assign detect_min[440][19] = (mid_1[3535:3528] < btm_0[3543:3536]) ? 1 : 0;
assign detect_min[440][20] = (mid_1[3535:3528] < btm_1[3527:3520]) ? 1 : 0;
assign detect_min[440][21] = (mid_1[3535:3528] < btm_1[3535:3528]) ? 1 : 0;
assign detect_min[440][22] = (mid_1[3535:3528] < btm_1[3543:3536]) ? 1 : 0;
assign detect_min[440][23] = (mid_1[3535:3528] < btm_2[3527:3520]) ? 1 : 0;
assign detect_min[440][24] = (mid_1[3535:3528] < btm_2[3535:3528]) ? 1 : 0;
assign detect_min[440][25] = (mid_1[3535:3528] < btm_2[3543:3536]) ? 1 : 0;

assign detect_min[441][0] = (mid_1[3543:3536] < top_0[3535:3528]) ? 1 : 0;
assign detect_min[441][1] = (mid_1[3543:3536] < top_0[3543:3536]) ? 1 : 0;
assign detect_min[441][2] = (mid_1[3543:3536] < top_0[3551:3544]) ? 1 : 0;
assign detect_min[441][3] = (mid_1[3543:3536] < top_1[3535:3528]) ? 1 : 0;
assign detect_min[441][4] = (mid_1[3543:3536] < top_1[3543:3536]) ? 1 : 0;
assign detect_min[441][5] = (mid_1[3543:3536] < top_1[3551:3544]) ? 1 : 0;
assign detect_min[441][6] = (mid_1[3543:3536] < top_2[3535:3528]) ? 1 : 0;
assign detect_min[441][7] = (mid_1[3543:3536] < top_2[3543:3536]) ? 1 : 0;
assign detect_min[441][8] = (mid_1[3543:3536] < top_2[3551:3544]) ? 1 : 0;
assign detect_min[441][9] = (mid_1[3543:3536] < mid_0[3535:3528]) ? 1 : 0;
assign detect_min[441][10] = (mid_1[3543:3536] < mid_0[3543:3536]) ? 1 : 0;
assign detect_min[441][11] = (mid_1[3543:3536] < mid_0[3551:3544]) ? 1 : 0;
assign detect_min[441][12] = (mid_1[3543:3536] < mid_1[3535:3528]) ? 1 : 0;
assign detect_min[441][13] = (mid_1[3543:3536] < mid_1[3551:3544]) ? 1 : 0;
assign detect_min[441][14] = (mid_1[3543:3536] < mid_2[3535:3528]) ? 1 : 0;
assign detect_min[441][15] = (mid_1[3543:3536] < mid_2[3543:3536]) ? 1 : 0;
assign detect_min[441][16] = (mid_1[3543:3536] < mid_2[3551:3544]) ? 1 : 0;
assign detect_min[441][17] = (mid_1[3543:3536] < btm_0[3535:3528]) ? 1 : 0;
assign detect_min[441][18] = (mid_1[3543:3536] < btm_0[3543:3536]) ? 1 : 0;
assign detect_min[441][19] = (mid_1[3543:3536] < btm_0[3551:3544]) ? 1 : 0;
assign detect_min[441][20] = (mid_1[3543:3536] < btm_1[3535:3528]) ? 1 : 0;
assign detect_min[441][21] = (mid_1[3543:3536] < btm_1[3543:3536]) ? 1 : 0;
assign detect_min[441][22] = (mid_1[3543:3536] < btm_1[3551:3544]) ? 1 : 0;
assign detect_min[441][23] = (mid_1[3543:3536] < btm_2[3535:3528]) ? 1 : 0;
assign detect_min[441][24] = (mid_1[3543:3536] < btm_2[3543:3536]) ? 1 : 0;
assign detect_min[441][25] = (mid_1[3543:3536] < btm_2[3551:3544]) ? 1 : 0;

assign detect_min[442][0] = (mid_1[3551:3544] < top_0[3543:3536]) ? 1 : 0;
assign detect_min[442][1] = (mid_1[3551:3544] < top_0[3551:3544]) ? 1 : 0;
assign detect_min[442][2] = (mid_1[3551:3544] < top_0[3559:3552]) ? 1 : 0;
assign detect_min[442][3] = (mid_1[3551:3544] < top_1[3543:3536]) ? 1 : 0;
assign detect_min[442][4] = (mid_1[3551:3544] < top_1[3551:3544]) ? 1 : 0;
assign detect_min[442][5] = (mid_1[3551:3544] < top_1[3559:3552]) ? 1 : 0;
assign detect_min[442][6] = (mid_1[3551:3544] < top_2[3543:3536]) ? 1 : 0;
assign detect_min[442][7] = (mid_1[3551:3544] < top_2[3551:3544]) ? 1 : 0;
assign detect_min[442][8] = (mid_1[3551:3544] < top_2[3559:3552]) ? 1 : 0;
assign detect_min[442][9] = (mid_1[3551:3544] < mid_0[3543:3536]) ? 1 : 0;
assign detect_min[442][10] = (mid_1[3551:3544] < mid_0[3551:3544]) ? 1 : 0;
assign detect_min[442][11] = (mid_1[3551:3544] < mid_0[3559:3552]) ? 1 : 0;
assign detect_min[442][12] = (mid_1[3551:3544] < mid_1[3543:3536]) ? 1 : 0;
assign detect_min[442][13] = (mid_1[3551:3544] < mid_1[3559:3552]) ? 1 : 0;
assign detect_min[442][14] = (mid_1[3551:3544] < mid_2[3543:3536]) ? 1 : 0;
assign detect_min[442][15] = (mid_1[3551:3544] < mid_2[3551:3544]) ? 1 : 0;
assign detect_min[442][16] = (mid_1[3551:3544] < mid_2[3559:3552]) ? 1 : 0;
assign detect_min[442][17] = (mid_1[3551:3544] < btm_0[3543:3536]) ? 1 : 0;
assign detect_min[442][18] = (mid_1[3551:3544] < btm_0[3551:3544]) ? 1 : 0;
assign detect_min[442][19] = (mid_1[3551:3544] < btm_0[3559:3552]) ? 1 : 0;
assign detect_min[442][20] = (mid_1[3551:3544] < btm_1[3543:3536]) ? 1 : 0;
assign detect_min[442][21] = (mid_1[3551:3544] < btm_1[3551:3544]) ? 1 : 0;
assign detect_min[442][22] = (mid_1[3551:3544] < btm_1[3559:3552]) ? 1 : 0;
assign detect_min[442][23] = (mid_1[3551:3544] < btm_2[3543:3536]) ? 1 : 0;
assign detect_min[442][24] = (mid_1[3551:3544] < btm_2[3551:3544]) ? 1 : 0;
assign detect_min[442][25] = (mid_1[3551:3544] < btm_2[3559:3552]) ? 1 : 0;

assign detect_min[443][0] = (mid_1[3559:3552] < top_0[3551:3544]) ? 1 : 0;
assign detect_min[443][1] = (mid_1[3559:3552] < top_0[3559:3552]) ? 1 : 0;
assign detect_min[443][2] = (mid_1[3559:3552] < top_0[3567:3560]) ? 1 : 0;
assign detect_min[443][3] = (mid_1[3559:3552] < top_1[3551:3544]) ? 1 : 0;
assign detect_min[443][4] = (mid_1[3559:3552] < top_1[3559:3552]) ? 1 : 0;
assign detect_min[443][5] = (mid_1[3559:3552] < top_1[3567:3560]) ? 1 : 0;
assign detect_min[443][6] = (mid_1[3559:3552] < top_2[3551:3544]) ? 1 : 0;
assign detect_min[443][7] = (mid_1[3559:3552] < top_2[3559:3552]) ? 1 : 0;
assign detect_min[443][8] = (mid_1[3559:3552] < top_2[3567:3560]) ? 1 : 0;
assign detect_min[443][9] = (mid_1[3559:3552] < mid_0[3551:3544]) ? 1 : 0;
assign detect_min[443][10] = (mid_1[3559:3552] < mid_0[3559:3552]) ? 1 : 0;
assign detect_min[443][11] = (mid_1[3559:3552] < mid_0[3567:3560]) ? 1 : 0;
assign detect_min[443][12] = (mid_1[3559:3552] < mid_1[3551:3544]) ? 1 : 0;
assign detect_min[443][13] = (mid_1[3559:3552] < mid_1[3567:3560]) ? 1 : 0;
assign detect_min[443][14] = (mid_1[3559:3552] < mid_2[3551:3544]) ? 1 : 0;
assign detect_min[443][15] = (mid_1[3559:3552] < mid_2[3559:3552]) ? 1 : 0;
assign detect_min[443][16] = (mid_1[3559:3552] < mid_2[3567:3560]) ? 1 : 0;
assign detect_min[443][17] = (mid_1[3559:3552] < btm_0[3551:3544]) ? 1 : 0;
assign detect_min[443][18] = (mid_1[3559:3552] < btm_0[3559:3552]) ? 1 : 0;
assign detect_min[443][19] = (mid_1[3559:3552] < btm_0[3567:3560]) ? 1 : 0;
assign detect_min[443][20] = (mid_1[3559:3552] < btm_1[3551:3544]) ? 1 : 0;
assign detect_min[443][21] = (mid_1[3559:3552] < btm_1[3559:3552]) ? 1 : 0;
assign detect_min[443][22] = (mid_1[3559:3552] < btm_1[3567:3560]) ? 1 : 0;
assign detect_min[443][23] = (mid_1[3559:3552] < btm_2[3551:3544]) ? 1 : 0;
assign detect_min[443][24] = (mid_1[3559:3552] < btm_2[3559:3552]) ? 1 : 0;
assign detect_min[443][25] = (mid_1[3559:3552] < btm_2[3567:3560]) ? 1 : 0;

assign detect_min[444][0] = (mid_1[3567:3560] < top_0[3559:3552]) ? 1 : 0;
assign detect_min[444][1] = (mid_1[3567:3560] < top_0[3567:3560]) ? 1 : 0;
assign detect_min[444][2] = (mid_1[3567:3560] < top_0[3575:3568]) ? 1 : 0;
assign detect_min[444][3] = (mid_1[3567:3560] < top_1[3559:3552]) ? 1 : 0;
assign detect_min[444][4] = (mid_1[3567:3560] < top_1[3567:3560]) ? 1 : 0;
assign detect_min[444][5] = (mid_1[3567:3560] < top_1[3575:3568]) ? 1 : 0;
assign detect_min[444][6] = (mid_1[3567:3560] < top_2[3559:3552]) ? 1 : 0;
assign detect_min[444][7] = (mid_1[3567:3560] < top_2[3567:3560]) ? 1 : 0;
assign detect_min[444][8] = (mid_1[3567:3560] < top_2[3575:3568]) ? 1 : 0;
assign detect_min[444][9] = (mid_1[3567:3560] < mid_0[3559:3552]) ? 1 : 0;
assign detect_min[444][10] = (mid_1[3567:3560] < mid_0[3567:3560]) ? 1 : 0;
assign detect_min[444][11] = (mid_1[3567:3560] < mid_0[3575:3568]) ? 1 : 0;
assign detect_min[444][12] = (mid_1[3567:3560] < mid_1[3559:3552]) ? 1 : 0;
assign detect_min[444][13] = (mid_1[3567:3560] < mid_1[3575:3568]) ? 1 : 0;
assign detect_min[444][14] = (mid_1[3567:3560] < mid_2[3559:3552]) ? 1 : 0;
assign detect_min[444][15] = (mid_1[3567:3560] < mid_2[3567:3560]) ? 1 : 0;
assign detect_min[444][16] = (mid_1[3567:3560] < mid_2[3575:3568]) ? 1 : 0;
assign detect_min[444][17] = (mid_1[3567:3560] < btm_0[3559:3552]) ? 1 : 0;
assign detect_min[444][18] = (mid_1[3567:3560] < btm_0[3567:3560]) ? 1 : 0;
assign detect_min[444][19] = (mid_1[3567:3560] < btm_0[3575:3568]) ? 1 : 0;
assign detect_min[444][20] = (mid_1[3567:3560] < btm_1[3559:3552]) ? 1 : 0;
assign detect_min[444][21] = (mid_1[3567:3560] < btm_1[3567:3560]) ? 1 : 0;
assign detect_min[444][22] = (mid_1[3567:3560] < btm_1[3575:3568]) ? 1 : 0;
assign detect_min[444][23] = (mid_1[3567:3560] < btm_2[3559:3552]) ? 1 : 0;
assign detect_min[444][24] = (mid_1[3567:3560] < btm_2[3567:3560]) ? 1 : 0;
assign detect_min[444][25] = (mid_1[3567:3560] < btm_2[3575:3568]) ? 1 : 0;

assign detect_min[445][0] = (mid_1[3575:3568] < top_0[3567:3560]) ? 1 : 0;
assign detect_min[445][1] = (mid_1[3575:3568] < top_0[3575:3568]) ? 1 : 0;
assign detect_min[445][2] = (mid_1[3575:3568] < top_0[3583:3576]) ? 1 : 0;
assign detect_min[445][3] = (mid_1[3575:3568] < top_1[3567:3560]) ? 1 : 0;
assign detect_min[445][4] = (mid_1[3575:3568] < top_1[3575:3568]) ? 1 : 0;
assign detect_min[445][5] = (mid_1[3575:3568] < top_1[3583:3576]) ? 1 : 0;
assign detect_min[445][6] = (mid_1[3575:3568] < top_2[3567:3560]) ? 1 : 0;
assign detect_min[445][7] = (mid_1[3575:3568] < top_2[3575:3568]) ? 1 : 0;
assign detect_min[445][8] = (mid_1[3575:3568] < top_2[3583:3576]) ? 1 : 0;
assign detect_min[445][9] = (mid_1[3575:3568] < mid_0[3567:3560]) ? 1 : 0;
assign detect_min[445][10] = (mid_1[3575:3568] < mid_0[3575:3568]) ? 1 : 0;
assign detect_min[445][11] = (mid_1[3575:3568] < mid_0[3583:3576]) ? 1 : 0;
assign detect_min[445][12] = (mid_1[3575:3568] < mid_1[3567:3560]) ? 1 : 0;
assign detect_min[445][13] = (mid_1[3575:3568] < mid_1[3583:3576]) ? 1 : 0;
assign detect_min[445][14] = (mid_1[3575:3568] < mid_2[3567:3560]) ? 1 : 0;
assign detect_min[445][15] = (mid_1[3575:3568] < mid_2[3575:3568]) ? 1 : 0;
assign detect_min[445][16] = (mid_1[3575:3568] < mid_2[3583:3576]) ? 1 : 0;
assign detect_min[445][17] = (mid_1[3575:3568] < btm_0[3567:3560]) ? 1 : 0;
assign detect_min[445][18] = (mid_1[3575:3568] < btm_0[3575:3568]) ? 1 : 0;
assign detect_min[445][19] = (mid_1[3575:3568] < btm_0[3583:3576]) ? 1 : 0;
assign detect_min[445][20] = (mid_1[3575:3568] < btm_1[3567:3560]) ? 1 : 0;
assign detect_min[445][21] = (mid_1[3575:3568] < btm_1[3575:3568]) ? 1 : 0;
assign detect_min[445][22] = (mid_1[3575:3568] < btm_1[3583:3576]) ? 1 : 0;
assign detect_min[445][23] = (mid_1[3575:3568] < btm_2[3567:3560]) ? 1 : 0;
assign detect_min[445][24] = (mid_1[3575:3568] < btm_2[3575:3568]) ? 1 : 0;
assign detect_min[445][25] = (mid_1[3575:3568] < btm_2[3583:3576]) ? 1 : 0;

assign detect_min[446][0] = (mid_1[3583:3576] < top_0[3575:3568]) ? 1 : 0;
assign detect_min[446][1] = (mid_1[3583:3576] < top_0[3583:3576]) ? 1 : 0;
assign detect_min[446][2] = (mid_1[3583:3576] < top_0[3591:3584]) ? 1 : 0;
assign detect_min[446][3] = (mid_1[3583:3576] < top_1[3575:3568]) ? 1 : 0;
assign detect_min[446][4] = (mid_1[3583:3576] < top_1[3583:3576]) ? 1 : 0;
assign detect_min[446][5] = (mid_1[3583:3576] < top_1[3591:3584]) ? 1 : 0;
assign detect_min[446][6] = (mid_1[3583:3576] < top_2[3575:3568]) ? 1 : 0;
assign detect_min[446][7] = (mid_1[3583:3576] < top_2[3583:3576]) ? 1 : 0;
assign detect_min[446][8] = (mid_1[3583:3576] < top_2[3591:3584]) ? 1 : 0;
assign detect_min[446][9] = (mid_1[3583:3576] < mid_0[3575:3568]) ? 1 : 0;
assign detect_min[446][10] = (mid_1[3583:3576] < mid_0[3583:3576]) ? 1 : 0;
assign detect_min[446][11] = (mid_1[3583:3576] < mid_0[3591:3584]) ? 1 : 0;
assign detect_min[446][12] = (mid_1[3583:3576] < mid_1[3575:3568]) ? 1 : 0;
assign detect_min[446][13] = (mid_1[3583:3576] < mid_1[3591:3584]) ? 1 : 0;
assign detect_min[446][14] = (mid_1[3583:3576] < mid_2[3575:3568]) ? 1 : 0;
assign detect_min[446][15] = (mid_1[3583:3576] < mid_2[3583:3576]) ? 1 : 0;
assign detect_min[446][16] = (mid_1[3583:3576] < mid_2[3591:3584]) ? 1 : 0;
assign detect_min[446][17] = (mid_1[3583:3576] < btm_0[3575:3568]) ? 1 : 0;
assign detect_min[446][18] = (mid_1[3583:3576] < btm_0[3583:3576]) ? 1 : 0;
assign detect_min[446][19] = (mid_1[3583:3576] < btm_0[3591:3584]) ? 1 : 0;
assign detect_min[446][20] = (mid_1[3583:3576] < btm_1[3575:3568]) ? 1 : 0;
assign detect_min[446][21] = (mid_1[3583:3576] < btm_1[3583:3576]) ? 1 : 0;
assign detect_min[446][22] = (mid_1[3583:3576] < btm_1[3591:3584]) ? 1 : 0;
assign detect_min[446][23] = (mid_1[3583:3576] < btm_2[3575:3568]) ? 1 : 0;
assign detect_min[446][24] = (mid_1[3583:3576] < btm_2[3583:3576]) ? 1 : 0;
assign detect_min[446][25] = (mid_1[3583:3576] < btm_2[3591:3584]) ? 1 : 0;

assign detect_min[447][0] = (mid_1[3591:3584] < top_0[3583:3576]) ? 1 : 0;
assign detect_min[447][1] = (mid_1[3591:3584] < top_0[3591:3584]) ? 1 : 0;
assign detect_min[447][2] = (mid_1[3591:3584] < top_0[3599:3592]) ? 1 : 0;
assign detect_min[447][3] = (mid_1[3591:3584] < top_1[3583:3576]) ? 1 : 0;
assign detect_min[447][4] = (mid_1[3591:3584] < top_1[3591:3584]) ? 1 : 0;
assign detect_min[447][5] = (mid_1[3591:3584] < top_1[3599:3592]) ? 1 : 0;
assign detect_min[447][6] = (mid_1[3591:3584] < top_2[3583:3576]) ? 1 : 0;
assign detect_min[447][7] = (mid_1[3591:3584] < top_2[3591:3584]) ? 1 : 0;
assign detect_min[447][8] = (mid_1[3591:3584] < top_2[3599:3592]) ? 1 : 0;
assign detect_min[447][9] = (mid_1[3591:3584] < mid_0[3583:3576]) ? 1 : 0;
assign detect_min[447][10] = (mid_1[3591:3584] < mid_0[3591:3584]) ? 1 : 0;
assign detect_min[447][11] = (mid_1[3591:3584] < mid_0[3599:3592]) ? 1 : 0;
assign detect_min[447][12] = (mid_1[3591:3584] < mid_1[3583:3576]) ? 1 : 0;
assign detect_min[447][13] = (mid_1[3591:3584] < mid_1[3599:3592]) ? 1 : 0;
assign detect_min[447][14] = (mid_1[3591:3584] < mid_2[3583:3576]) ? 1 : 0;
assign detect_min[447][15] = (mid_1[3591:3584] < mid_2[3591:3584]) ? 1 : 0;
assign detect_min[447][16] = (mid_1[3591:3584] < mid_2[3599:3592]) ? 1 : 0;
assign detect_min[447][17] = (mid_1[3591:3584] < btm_0[3583:3576]) ? 1 : 0;
assign detect_min[447][18] = (mid_1[3591:3584] < btm_0[3591:3584]) ? 1 : 0;
assign detect_min[447][19] = (mid_1[3591:3584] < btm_0[3599:3592]) ? 1 : 0;
assign detect_min[447][20] = (mid_1[3591:3584] < btm_1[3583:3576]) ? 1 : 0;
assign detect_min[447][21] = (mid_1[3591:3584] < btm_1[3591:3584]) ? 1 : 0;
assign detect_min[447][22] = (mid_1[3591:3584] < btm_1[3599:3592]) ? 1 : 0;
assign detect_min[447][23] = (mid_1[3591:3584] < btm_2[3583:3576]) ? 1 : 0;
assign detect_min[447][24] = (mid_1[3591:3584] < btm_2[3591:3584]) ? 1 : 0;
assign detect_min[447][25] = (mid_1[3591:3584] < btm_2[3599:3592]) ? 1 : 0;

assign detect_min[448][0] = (mid_1[3599:3592] < top_0[3591:3584]) ? 1 : 0;
assign detect_min[448][1] = (mid_1[3599:3592] < top_0[3599:3592]) ? 1 : 0;
assign detect_min[448][2] = (mid_1[3599:3592] < top_0[3607:3600]) ? 1 : 0;
assign detect_min[448][3] = (mid_1[3599:3592] < top_1[3591:3584]) ? 1 : 0;
assign detect_min[448][4] = (mid_1[3599:3592] < top_1[3599:3592]) ? 1 : 0;
assign detect_min[448][5] = (mid_1[3599:3592] < top_1[3607:3600]) ? 1 : 0;
assign detect_min[448][6] = (mid_1[3599:3592] < top_2[3591:3584]) ? 1 : 0;
assign detect_min[448][7] = (mid_1[3599:3592] < top_2[3599:3592]) ? 1 : 0;
assign detect_min[448][8] = (mid_1[3599:3592] < top_2[3607:3600]) ? 1 : 0;
assign detect_min[448][9] = (mid_1[3599:3592] < mid_0[3591:3584]) ? 1 : 0;
assign detect_min[448][10] = (mid_1[3599:3592] < mid_0[3599:3592]) ? 1 : 0;
assign detect_min[448][11] = (mid_1[3599:3592] < mid_0[3607:3600]) ? 1 : 0;
assign detect_min[448][12] = (mid_1[3599:3592] < mid_1[3591:3584]) ? 1 : 0;
assign detect_min[448][13] = (mid_1[3599:3592] < mid_1[3607:3600]) ? 1 : 0;
assign detect_min[448][14] = (mid_1[3599:3592] < mid_2[3591:3584]) ? 1 : 0;
assign detect_min[448][15] = (mid_1[3599:3592] < mid_2[3599:3592]) ? 1 : 0;
assign detect_min[448][16] = (mid_1[3599:3592] < mid_2[3607:3600]) ? 1 : 0;
assign detect_min[448][17] = (mid_1[3599:3592] < btm_0[3591:3584]) ? 1 : 0;
assign detect_min[448][18] = (mid_1[3599:3592] < btm_0[3599:3592]) ? 1 : 0;
assign detect_min[448][19] = (mid_1[3599:3592] < btm_0[3607:3600]) ? 1 : 0;
assign detect_min[448][20] = (mid_1[3599:3592] < btm_1[3591:3584]) ? 1 : 0;
assign detect_min[448][21] = (mid_1[3599:3592] < btm_1[3599:3592]) ? 1 : 0;
assign detect_min[448][22] = (mid_1[3599:3592] < btm_1[3607:3600]) ? 1 : 0;
assign detect_min[448][23] = (mid_1[3599:3592] < btm_2[3591:3584]) ? 1 : 0;
assign detect_min[448][24] = (mid_1[3599:3592] < btm_2[3599:3592]) ? 1 : 0;
assign detect_min[448][25] = (mid_1[3599:3592] < btm_2[3607:3600]) ? 1 : 0;

assign detect_min[449][0] = (mid_1[3607:3600] < top_0[3599:3592]) ? 1 : 0;
assign detect_min[449][1] = (mid_1[3607:3600] < top_0[3607:3600]) ? 1 : 0;
assign detect_min[449][2] = (mid_1[3607:3600] < top_0[3615:3608]) ? 1 : 0;
assign detect_min[449][3] = (mid_1[3607:3600] < top_1[3599:3592]) ? 1 : 0;
assign detect_min[449][4] = (mid_1[3607:3600] < top_1[3607:3600]) ? 1 : 0;
assign detect_min[449][5] = (mid_1[3607:3600] < top_1[3615:3608]) ? 1 : 0;
assign detect_min[449][6] = (mid_1[3607:3600] < top_2[3599:3592]) ? 1 : 0;
assign detect_min[449][7] = (mid_1[3607:3600] < top_2[3607:3600]) ? 1 : 0;
assign detect_min[449][8] = (mid_1[3607:3600] < top_2[3615:3608]) ? 1 : 0;
assign detect_min[449][9] = (mid_1[3607:3600] < mid_0[3599:3592]) ? 1 : 0;
assign detect_min[449][10] = (mid_1[3607:3600] < mid_0[3607:3600]) ? 1 : 0;
assign detect_min[449][11] = (mid_1[3607:3600] < mid_0[3615:3608]) ? 1 : 0;
assign detect_min[449][12] = (mid_1[3607:3600] < mid_1[3599:3592]) ? 1 : 0;
assign detect_min[449][13] = (mid_1[3607:3600] < mid_1[3615:3608]) ? 1 : 0;
assign detect_min[449][14] = (mid_1[3607:3600] < mid_2[3599:3592]) ? 1 : 0;
assign detect_min[449][15] = (mid_1[3607:3600] < mid_2[3607:3600]) ? 1 : 0;
assign detect_min[449][16] = (mid_1[3607:3600] < mid_2[3615:3608]) ? 1 : 0;
assign detect_min[449][17] = (mid_1[3607:3600] < btm_0[3599:3592]) ? 1 : 0;
assign detect_min[449][18] = (mid_1[3607:3600] < btm_0[3607:3600]) ? 1 : 0;
assign detect_min[449][19] = (mid_1[3607:3600] < btm_0[3615:3608]) ? 1 : 0;
assign detect_min[449][20] = (mid_1[3607:3600] < btm_1[3599:3592]) ? 1 : 0;
assign detect_min[449][21] = (mid_1[3607:3600] < btm_1[3607:3600]) ? 1 : 0;
assign detect_min[449][22] = (mid_1[3607:3600] < btm_1[3615:3608]) ? 1 : 0;
assign detect_min[449][23] = (mid_1[3607:3600] < btm_2[3599:3592]) ? 1 : 0;
assign detect_min[449][24] = (mid_1[3607:3600] < btm_2[3607:3600]) ? 1 : 0;
assign detect_min[449][25] = (mid_1[3607:3600] < btm_2[3615:3608]) ? 1 : 0;

assign detect_min[450][0] = (mid_1[3615:3608] < top_0[3607:3600]) ? 1 : 0;
assign detect_min[450][1] = (mid_1[3615:3608] < top_0[3615:3608]) ? 1 : 0;
assign detect_min[450][2] = (mid_1[3615:3608] < top_0[3623:3616]) ? 1 : 0;
assign detect_min[450][3] = (mid_1[3615:3608] < top_1[3607:3600]) ? 1 : 0;
assign detect_min[450][4] = (mid_1[3615:3608] < top_1[3615:3608]) ? 1 : 0;
assign detect_min[450][5] = (mid_1[3615:3608] < top_1[3623:3616]) ? 1 : 0;
assign detect_min[450][6] = (mid_1[3615:3608] < top_2[3607:3600]) ? 1 : 0;
assign detect_min[450][7] = (mid_1[3615:3608] < top_2[3615:3608]) ? 1 : 0;
assign detect_min[450][8] = (mid_1[3615:3608] < top_2[3623:3616]) ? 1 : 0;
assign detect_min[450][9] = (mid_1[3615:3608] < mid_0[3607:3600]) ? 1 : 0;
assign detect_min[450][10] = (mid_1[3615:3608] < mid_0[3615:3608]) ? 1 : 0;
assign detect_min[450][11] = (mid_1[3615:3608] < mid_0[3623:3616]) ? 1 : 0;
assign detect_min[450][12] = (mid_1[3615:3608] < mid_1[3607:3600]) ? 1 : 0;
assign detect_min[450][13] = (mid_1[3615:3608] < mid_1[3623:3616]) ? 1 : 0;
assign detect_min[450][14] = (mid_1[3615:3608] < mid_2[3607:3600]) ? 1 : 0;
assign detect_min[450][15] = (mid_1[3615:3608] < mid_2[3615:3608]) ? 1 : 0;
assign detect_min[450][16] = (mid_1[3615:3608] < mid_2[3623:3616]) ? 1 : 0;
assign detect_min[450][17] = (mid_1[3615:3608] < btm_0[3607:3600]) ? 1 : 0;
assign detect_min[450][18] = (mid_1[3615:3608] < btm_0[3615:3608]) ? 1 : 0;
assign detect_min[450][19] = (mid_1[3615:3608] < btm_0[3623:3616]) ? 1 : 0;
assign detect_min[450][20] = (mid_1[3615:3608] < btm_1[3607:3600]) ? 1 : 0;
assign detect_min[450][21] = (mid_1[3615:3608] < btm_1[3615:3608]) ? 1 : 0;
assign detect_min[450][22] = (mid_1[3615:3608] < btm_1[3623:3616]) ? 1 : 0;
assign detect_min[450][23] = (mid_1[3615:3608] < btm_2[3607:3600]) ? 1 : 0;
assign detect_min[450][24] = (mid_1[3615:3608] < btm_2[3615:3608]) ? 1 : 0;
assign detect_min[450][25] = (mid_1[3615:3608] < btm_2[3623:3616]) ? 1 : 0;

assign detect_min[451][0] = (mid_1[3623:3616] < top_0[3615:3608]) ? 1 : 0;
assign detect_min[451][1] = (mid_1[3623:3616] < top_0[3623:3616]) ? 1 : 0;
assign detect_min[451][2] = (mid_1[3623:3616] < top_0[3631:3624]) ? 1 : 0;
assign detect_min[451][3] = (mid_1[3623:3616] < top_1[3615:3608]) ? 1 : 0;
assign detect_min[451][4] = (mid_1[3623:3616] < top_1[3623:3616]) ? 1 : 0;
assign detect_min[451][5] = (mid_1[3623:3616] < top_1[3631:3624]) ? 1 : 0;
assign detect_min[451][6] = (mid_1[3623:3616] < top_2[3615:3608]) ? 1 : 0;
assign detect_min[451][7] = (mid_1[3623:3616] < top_2[3623:3616]) ? 1 : 0;
assign detect_min[451][8] = (mid_1[3623:3616] < top_2[3631:3624]) ? 1 : 0;
assign detect_min[451][9] = (mid_1[3623:3616] < mid_0[3615:3608]) ? 1 : 0;
assign detect_min[451][10] = (mid_1[3623:3616] < mid_0[3623:3616]) ? 1 : 0;
assign detect_min[451][11] = (mid_1[3623:3616] < mid_0[3631:3624]) ? 1 : 0;
assign detect_min[451][12] = (mid_1[3623:3616] < mid_1[3615:3608]) ? 1 : 0;
assign detect_min[451][13] = (mid_1[3623:3616] < mid_1[3631:3624]) ? 1 : 0;
assign detect_min[451][14] = (mid_1[3623:3616] < mid_2[3615:3608]) ? 1 : 0;
assign detect_min[451][15] = (mid_1[3623:3616] < mid_2[3623:3616]) ? 1 : 0;
assign detect_min[451][16] = (mid_1[3623:3616] < mid_2[3631:3624]) ? 1 : 0;
assign detect_min[451][17] = (mid_1[3623:3616] < btm_0[3615:3608]) ? 1 : 0;
assign detect_min[451][18] = (mid_1[3623:3616] < btm_0[3623:3616]) ? 1 : 0;
assign detect_min[451][19] = (mid_1[3623:3616] < btm_0[3631:3624]) ? 1 : 0;
assign detect_min[451][20] = (mid_1[3623:3616] < btm_1[3615:3608]) ? 1 : 0;
assign detect_min[451][21] = (mid_1[3623:3616] < btm_1[3623:3616]) ? 1 : 0;
assign detect_min[451][22] = (mid_1[3623:3616] < btm_1[3631:3624]) ? 1 : 0;
assign detect_min[451][23] = (mid_1[3623:3616] < btm_2[3615:3608]) ? 1 : 0;
assign detect_min[451][24] = (mid_1[3623:3616] < btm_2[3623:3616]) ? 1 : 0;
assign detect_min[451][25] = (mid_1[3623:3616] < btm_2[3631:3624]) ? 1 : 0;

assign detect_min[452][0] = (mid_1[3631:3624] < top_0[3623:3616]) ? 1 : 0;
assign detect_min[452][1] = (mid_1[3631:3624] < top_0[3631:3624]) ? 1 : 0;
assign detect_min[452][2] = (mid_1[3631:3624] < top_0[3639:3632]) ? 1 : 0;
assign detect_min[452][3] = (mid_1[3631:3624] < top_1[3623:3616]) ? 1 : 0;
assign detect_min[452][4] = (mid_1[3631:3624] < top_1[3631:3624]) ? 1 : 0;
assign detect_min[452][5] = (mid_1[3631:3624] < top_1[3639:3632]) ? 1 : 0;
assign detect_min[452][6] = (mid_1[3631:3624] < top_2[3623:3616]) ? 1 : 0;
assign detect_min[452][7] = (mid_1[3631:3624] < top_2[3631:3624]) ? 1 : 0;
assign detect_min[452][8] = (mid_1[3631:3624] < top_2[3639:3632]) ? 1 : 0;
assign detect_min[452][9] = (mid_1[3631:3624] < mid_0[3623:3616]) ? 1 : 0;
assign detect_min[452][10] = (mid_1[3631:3624] < mid_0[3631:3624]) ? 1 : 0;
assign detect_min[452][11] = (mid_1[3631:3624] < mid_0[3639:3632]) ? 1 : 0;
assign detect_min[452][12] = (mid_1[3631:3624] < mid_1[3623:3616]) ? 1 : 0;
assign detect_min[452][13] = (mid_1[3631:3624] < mid_1[3639:3632]) ? 1 : 0;
assign detect_min[452][14] = (mid_1[3631:3624] < mid_2[3623:3616]) ? 1 : 0;
assign detect_min[452][15] = (mid_1[3631:3624] < mid_2[3631:3624]) ? 1 : 0;
assign detect_min[452][16] = (mid_1[3631:3624] < mid_2[3639:3632]) ? 1 : 0;
assign detect_min[452][17] = (mid_1[3631:3624] < btm_0[3623:3616]) ? 1 : 0;
assign detect_min[452][18] = (mid_1[3631:3624] < btm_0[3631:3624]) ? 1 : 0;
assign detect_min[452][19] = (mid_1[3631:3624] < btm_0[3639:3632]) ? 1 : 0;
assign detect_min[452][20] = (mid_1[3631:3624] < btm_1[3623:3616]) ? 1 : 0;
assign detect_min[452][21] = (mid_1[3631:3624] < btm_1[3631:3624]) ? 1 : 0;
assign detect_min[452][22] = (mid_1[3631:3624] < btm_1[3639:3632]) ? 1 : 0;
assign detect_min[452][23] = (mid_1[3631:3624] < btm_2[3623:3616]) ? 1 : 0;
assign detect_min[452][24] = (mid_1[3631:3624] < btm_2[3631:3624]) ? 1 : 0;
assign detect_min[452][25] = (mid_1[3631:3624] < btm_2[3639:3632]) ? 1 : 0;

assign detect_min[453][0] = (mid_1[3639:3632] < top_0[3631:3624]) ? 1 : 0;
assign detect_min[453][1] = (mid_1[3639:3632] < top_0[3639:3632]) ? 1 : 0;
assign detect_min[453][2] = (mid_1[3639:3632] < top_0[3647:3640]) ? 1 : 0;
assign detect_min[453][3] = (mid_1[3639:3632] < top_1[3631:3624]) ? 1 : 0;
assign detect_min[453][4] = (mid_1[3639:3632] < top_1[3639:3632]) ? 1 : 0;
assign detect_min[453][5] = (mid_1[3639:3632] < top_1[3647:3640]) ? 1 : 0;
assign detect_min[453][6] = (mid_1[3639:3632] < top_2[3631:3624]) ? 1 : 0;
assign detect_min[453][7] = (mid_1[3639:3632] < top_2[3639:3632]) ? 1 : 0;
assign detect_min[453][8] = (mid_1[3639:3632] < top_2[3647:3640]) ? 1 : 0;
assign detect_min[453][9] = (mid_1[3639:3632] < mid_0[3631:3624]) ? 1 : 0;
assign detect_min[453][10] = (mid_1[3639:3632] < mid_0[3639:3632]) ? 1 : 0;
assign detect_min[453][11] = (mid_1[3639:3632] < mid_0[3647:3640]) ? 1 : 0;
assign detect_min[453][12] = (mid_1[3639:3632] < mid_1[3631:3624]) ? 1 : 0;
assign detect_min[453][13] = (mid_1[3639:3632] < mid_1[3647:3640]) ? 1 : 0;
assign detect_min[453][14] = (mid_1[3639:3632] < mid_2[3631:3624]) ? 1 : 0;
assign detect_min[453][15] = (mid_1[3639:3632] < mid_2[3639:3632]) ? 1 : 0;
assign detect_min[453][16] = (mid_1[3639:3632] < mid_2[3647:3640]) ? 1 : 0;
assign detect_min[453][17] = (mid_1[3639:3632] < btm_0[3631:3624]) ? 1 : 0;
assign detect_min[453][18] = (mid_1[3639:3632] < btm_0[3639:3632]) ? 1 : 0;
assign detect_min[453][19] = (mid_1[3639:3632] < btm_0[3647:3640]) ? 1 : 0;
assign detect_min[453][20] = (mid_1[3639:3632] < btm_1[3631:3624]) ? 1 : 0;
assign detect_min[453][21] = (mid_1[3639:3632] < btm_1[3639:3632]) ? 1 : 0;
assign detect_min[453][22] = (mid_1[3639:3632] < btm_1[3647:3640]) ? 1 : 0;
assign detect_min[453][23] = (mid_1[3639:3632] < btm_2[3631:3624]) ? 1 : 0;
assign detect_min[453][24] = (mid_1[3639:3632] < btm_2[3639:3632]) ? 1 : 0;
assign detect_min[453][25] = (mid_1[3639:3632] < btm_2[3647:3640]) ? 1 : 0;

assign detect_min[454][0] = (mid_1[3647:3640] < top_0[3639:3632]) ? 1 : 0;
assign detect_min[454][1] = (mid_1[3647:3640] < top_0[3647:3640]) ? 1 : 0;
assign detect_min[454][2] = (mid_1[3647:3640] < top_0[3655:3648]) ? 1 : 0;
assign detect_min[454][3] = (mid_1[3647:3640] < top_1[3639:3632]) ? 1 : 0;
assign detect_min[454][4] = (mid_1[3647:3640] < top_1[3647:3640]) ? 1 : 0;
assign detect_min[454][5] = (mid_1[3647:3640] < top_1[3655:3648]) ? 1 : 0;
assign detect_min[454][6] = (mid_1[3647:3640] < top_2[3639:3632]) ? 1 : 0;
assign detect_min[454][7] = (mid_1[3647:3640] < top_2[3647:3640]) ? 1 : 0;
assign detect_min[454][8] = (mid_1[3647:3640] < top_2[3655:3648]) ? 1 : 0;
assign detect_min[454][9] = (mid_1[3647:3640] < mid_0[3639:3632]) ? 1 : 0;
assign detect_min[454][10] = (mid_1[3647:3640] < mid_0[3647:3640]) ? 1 : 0;
assign detect_min[454][11] = (mid_1[3647:3640] < mid_0[3655:3648]) ? 1 : 0;
assign detect_min[454][12] = (mid_1[3647:3640] < mid_1[3639:3632]) ? 1 : 0;
assign detect_min[454][13] = (mid_1[3647:3640] < mid_1[3655:3648]) ? 1 : 0;
assign detect_min[454][14] = (mid_1[3647:3640] < mid_2[3639:3632]) ? 1 : 0;
assign detect_min[454][15] = (mid_1[3647:3640] < mid_2[3647:3640]) ? 1 : 0;
assign detect_min[454][16] = (mid_1[3647:3640] < mid_2[3655:3648]) ? 1 : 0;
assign detect_min[454][17] = (mid_1[3647:3640] < btm_0[3639:3632]) ? 1 : 0;
assign detect_min[454][18] = (mid_1[3647:3640] < btm_0[3647:3640]) ? 1 : 0;
assign detect_min[454][19] = (mid_1[3647:3640] < btm_0[3655:3648]) ? 1 : 0;
assign detect_min[454][20] = (mid_1[3647:3640] < btm_1[3639:3632]) ? 1 : 0;
assign detect_min[454][21] = (mid_1[3647:3640] < btm_1[3647:3640]) ? 1 : 0;
assign detect_min[454][22] = (mid_1[3647:3640] < btm_1[3655:3648]) ? 1 : 0;
assign detect_min[454][23] = (mid_1[3647:3640] < btm_2[3639:3632]) ? 1 : 0;
assign detect_min[454][24] = (mid_1[3647:3640] < btm_2[3647:3640]) ? 1 : 0;
assign detect_min[454][25] = (mid_1[3647:3640] < btm_2[3655:3648]) ? 1 : 0;

assign detect_min[455][0] = (mid_1[3655:3648] < top_0[3647:3640]) ? 1 : 0;
assign detect_min[455][1] = (mid_1[3655:3648] < top_0[3655:3648]) ? 1 : 0;
assign detect_min[455][2] = (mid_1[3655:3648] < top_0[3663:3656]) ? 1 : 0;
assign detect_min[455][3] = (mid_1[3655:3648] < top_1[3647:3640]) ? 1 : 0;
assign detect_min[455][4] = (mid_1[3655:3648] < top_1[3655:3648]) ? 1 : 0;
assign detect_min[455][5] = (mid_1[3655:3648] < top_1[3663:3656]) ? 1 : 0;
assign detect_min[455][6] = (mid_1[3655:3648] < top_2[3647:3640]) ? 1 : 0;
assign detect_min[455][7] = (mid_1[3655:3648] < top_2[3655:3648]) ? 1 : 0;
assign detect_min[455][8] = (mid_1[3655:3648] < top_2[3663:3656]) ? 1 : 0;
assign detect_min[455][9] = (mid_1[3655:3648] < mid_0[3647:3640]) ? 1 : 0;
assign detect_min[455][10] = (mid_1[3655:3648] < mid_0[3655:3648]) ? 1 : 0;
assign detect_min[455][11] = (mid_1[3655:3648] < mid_0[3663:3656]) ? 1 : 0;
assign detect_min[455][12] = (mid_1[3655:3648] < mid_1[3647:3640]) ? 1 : 0;
assign detect_min[455][13] = (mid_1[3655:3648] < mid_1[3663:3656]) ? 1 : 0;
assign detect_min[455][14] = (mid_1[3655:3648] < mid_2[3647:3640]) ? 1 : 0;
assign detect_min[455][15] = (mid_1[3655:3648] < mid_2[3655:3648]) ? 1 : 0;
assign detect_min[455][16] = (mid_1[3655:3648] < mid_2[3663:3656]) ? 1 : 0;
assign detect_min[455][17] = (mid_1[3655:3648] < btm_0[3647:3640]) ? 1 : 0;
assign detect_min[455][18] = (mid_1[3655:3648] < btm_0[3655:3648]) ? 1 : 0;
assign detect_min[455][19] = (mid_1[3655:3648] < btm_0[3663:3656]) ? 1 : 0;
assign detect_min[455][20] = (mid_1[3655:3648] < btm_1[3647:3640]) ? 1 : 0;
assign detect_min[455][21] = (mid_1[3655:3648] < btm_1[3655:3648]) ? 1 : 0;
assign detect_min[455][22] = (mid_1[3655:3648] < btm_1[3663:3656]) ? 1 : 0;
assign detect_min[455][23] = (mid_1[3655:3648] < btm_2[3647:3640]) ? 1 : 0;
assign detect_min[455][24] = (mid_1[3655:3648] < btm_2[3655:3648]) ? 1 : 0;
assign detect_min[455][25] = (mid_1[3655:3648] < btm_2[3663:3656]) ? 1 : 0;

assign detect_min[456][0] = (mid_1[3663:3656] < top_0[3655:3648]) ? 1 : 0;
assign detect_min[456][1] = (mid_1[3663:3656] < top_0[3663:3656]) ? 1 : 0;
assign detect_min[456][2] = (mid_1[3663:3656] < top_0[3671:3664]) ? 1 : 0;
assign detect_min[456][3] = (mid_1[3663:3656] < top_1[3655:3648]) ? 1 : 0;
assign detect_min[456][4] = (mid_1[3663:3656] < top_1[3663:3656]) ? 1 : 0;
assign detect_min[456][5] = (mid_1[3663:3656] < top_1[3671:3664]) ? 1 : 0;
assign detect_min[456][6] = (mid_1[3663:3656] < top_2[3655:3648]) ? 1 : 0;
assign detect_min[456][7] = (mid_1[3663:3656] < top_2[3663:3656]) ? 1 : 0;
assign detect_min[456][8] = (mid_1[3663:3656] < top_2[3671:3664]) ? 1 : 0;
assign detect_min[456][9] = (mid_1[3663:3656] < mid_0[3655:3648]) ? 1 : 0;
assign detect_min[456][10] = (mid_1[3663:3656] < mid_0[3663:3656]) ? 1 : 0;
assign detect_min[456][11] = (mid_1[3663:3656] < mid_0[3671:3664]) ? 1 : 0;
assign detect_min[456][12] = (mid_1[3663:3656] < mid_1[3655:3648]) ? 1 : 0;
assign detect_min[456][13] = (mid_1[3663:3656] < mid_1[3671:3664]) ? 1 : 0;
assign detect_min[456][14] = (mid_1[3663:3656] < mid_2[3655:3648]) ? 1 : 0;
assign detect_min[456][15] = (mid_1[3663:3656] < mid_2[3663:3656]) ? 1 : 0;
assign detect_min[456][16] = (mid_1[3663:3656] < mid_2[3671:3664]) ? 1 : 0;
assign detect_min[456][17] = (mid_1[3663:3656] < btm_0[3655:3648]) ? 1 : 0;
assign detect_min[456][18] = (mid_1[3663:3656] < btm_0[3663:3656]) ? 1 : 0;
assign detect_min[456][19] = (mid_1[3663:3656] < btm_0[3671:3664]) ? 1 : 0;
assign detect_min[456][20] = (mid_1[3663:3656] < btm_1[3655:3648]) ? 1 : 0;
assign detect_min[456][21] = (mid_1[3663:3656] < btm_1[3663:3656]) ? 1 : 0;
assign detect_min[456][22] = (mid_1[3663:3656] < btm_1[3671:3664]) ? 1 : 0;
assign detect_min[456][23] = (mid_1[3663:3656] < btm_2[3655:3648]) ? 1 : 0;
assign detect_min[456][24] = (mid_1[3663:3656] < btm_2[3663:3656]) ? 1 : 0;
assign detect_min[456][25] = (mid_1[3663:3656] < btm_2[3671:3664]) ? 1 : 0;

assign detect_min[457][0] = (mid_1[3671:3664] < top_0[3663:3656]) ? 1 : 0;
assign detect_min[457][1] = (mid_1[3671:3664] < top_0[3671:3664]) ? 1 : 0;
assign detect_min[457][2] = (mid_1[3671:3664] < top_0[3679:3672]) ? 1 : 0;
assign detect_min[457][3] = (mid_1[3671:3664] < top_1[3663:3656]) ? 1 : 0;
assign detect_min[457][4] = (mid_1[3671:3664] < top_1[3671:3664]) ? 1 : 0;
assign detect_min[457][5] = (mid_1[3671:3664] < top_1[3679:3672]) ? 1 : 0;
assign detect_min[457][6] = (mid_1[3671:3664] < top_2[3663:3656]) ? 1 : 0;
assign detect_min[457][7] = (mid_1[3671:3664] < top_2[3671:3664]) ? 1 : 0;
assign detect_min[457][8] = (mid_1[3671:3664] < top_2[3679:3672]) ? 1 : 0;
assign detect_min[457][9] = (mid_1[3671:3664] < mid_0[3663:3656]) ? 1 : 0;
assign detect_min[457][10] = (mid_1[3671:3664] < mid_0[3671:3664]) ? 1 : 0;
assign detect_min[457][11] = (mid_1[3671:3664] < mid_0[3679:3672]) ? 1 : 0;
assign detect_min[457][12] = (mid_1[3671:3664] < mid_1[3663:3656]) ? 1 : 0;
assign detect_min[457][13] = (mid_1[3671:3664] < mid_1[3679:3672]) ? 1 : 0;
assign detect_min[457][14] = (mid_1[3671:3664] < mid_2[3663:3656]) ? 1 : 0;
assign detect_min[457][15] = (mid_1[3671:3664] < mid_2[3671:3664]) ? 1 : 0;
assign detect_min[457][16] = (mid_1[3671:3664] < mid_2[3679:3672]) ? 1 : 0;
assign detect_min[457][17] = (mid_1[3671:3664] < btm_0[3663:3656]) ? 1 : 0;
assign detect_min[457][18] = (mid_1[3671:3664] < btm_0[3671:3664]) ? 1 : 0;
assign detect_min[457][19] = (mid_1[3671:3664] < btm_0[3679:3672]) ? 1 : 0;
assign detect_min[457][20] = (mid_1[3671:3664] < btm_1[3663:3656]) ? 1 : 0;
assign detect_min[457][21] = (mid_1[3671:3664] < btm_1[3671:3664]) ? 1 : 0;
assign detect_min[457][22] = (mid_1[3671:3664] < btm_1[3679:3672]) ? 1 : 0;
assign detect_min[457][23] = (mid_1[3671:3664] < btm_2[3663:3656]) ? 1 : 0;
assign detect_min[457][24] = (mid_1[3671:3664] < btm_2[3671:3664]) ? 1 : 0;
assign detect_min[457][25] = (mid_1[3671:3664] < btm_2[3679:3672]) ? 1 : 0;

assign detect_min[458][0] = (mid_1[3679:3672] < top_0[3671:3664]) ? 1 : 0;
assign detect_min[458][1] = (mid_1[3679:3672] < top_0[3679:3672]) ? 1 : 0;
assign detect_min[458][2] = (mid_1[3679:3672] < top_0[3687:3680]) ? 1 : 0;
assign detect_min[458][3] = (mid_1[3679:3672] < top_1[3671:3664]) ? 1 : 0;
assign detect_min[458][4] = (mid_1[3679:3672] < top_1[3679:3672]) ? 1 : 0;
assign detect_min[458][5] = (mid_1[3679:3672] < top_1[3687:3680]) ? 1 : 0;
assign detect_min[458][6] = (mid_1[3679:3672] < top_2[3671:3664]) ? 1 : 0;
assign detect_min[458][7] = (mid_1[3679:3672] < top_2[3679:3672]) ? 1 : 0;
assign detect_min[458][8] = (mid_1[3679:3672] < top_2[3687:3680]) ? 1 : 0;
assign detect_min[458][9] = (mid_1[3679:3672] < mid_0[3671:3664]) ? 1 : 0;
assign detect_min[458][10] = (mid_1[3679:3672] < mid_0[3679:3672]) ? 1 : 0;
assign detect_min[458][11] = (mid_1[3679:3672] < mid_0[3687:3680]) ? 1 : 0;
assign detect_min[458][12] = (mid_1[3679:3672] < mid_1[3671:3664]) ? 1 : 0;
assign detect_min[458][13] = (mid_1[3679:3672] < mid_1[3687:3680]) ? 1 : 0;
assign detect_min[458][14] = (mid_1[3679:3672] < mid_2[3671:3664]) ? 1 : 0;
assign detect_min[458][15] = (mid_1[3679:3672] < mid_2[3679:3672]) ? 1 : 0;
assign detect_min[458][16] = (mid_1[3679:3672] < mid_2[3687:3680]) ? 1 : 0;
assign detect_min[458][17] = (mid_1[3679:3672] < btm_0[3671:3664]) ? 1 : 0;
assign detect_min[458][18] = (mid_1[3679:3672] < btm_0[3679:3672]) ? 1 : 0;
assign detect_min[458][19] = (mid_1[3679:3672] < btm_0[3687:3680]) ? 1 : 0;
assign detect_min[458][20] = (mid_1[3679:3672] < btm_1[3671:3664]) ? 1 : 0;
assign detect_min[458][21] = (mid_1[3679:3672] < btm_1[3679:3672]) ? 1 : 0;
assign detect_min[458][22] = (mid_1[3679:3672] < btm_1[3687:3680]) ? 1 : 0;
assign detect_min[458][23] = (mid_1[3679:3672] < btm_2[3671:3664]) ? 1 : 0;
assign detect_min[458][24] = (mid_1[3679:3672] < btm_2[3679:3672]) ? 1 : 0;
assign detect_min[458][25] = (mid_1[3679:3672] < btm_2[3687:3680]) ? 1 : 0;

assign detect_min[459][0] = (mid_1[3687:3680] < top_0[3679:3672]) ? 1 : 0;
assign detect_min[459][1] = (mid_1[3687:3680] < top_0[3687:3680]) ? 1 : 0;
assign detect_min[459][2] = (mid_1[3687:3680] < top_0[3695:3688]) ? 1 : 0;
assign detect_min[459][3] = (mid_1[3687:3680] < top_1[3679:3672]) ? 1 : 0;
assign detect_min[459][4] = (mid_1[3687:3680] < top_1[3687:3680]) ? 1 : 0;
assign detect_min[459][5] = (mid_1[3687:3680] < top_1[3695:3688]) ? 1 : 0;
assign detect_min[459][6] = (mid_1[3687:3680] < top_2[3679:3672]) ? 1 : 0;
assign detect_min[459][7] = (mid_1[3687:3680] < top_2[3687:3680]) ? 1 : 0;
assign detect_min[459][8] = (mid_1[3687:3680] < top_2[3695:3688]) ? 1 : 0;
assign detect_min[459][9] = (mid_1[3687:3680] < mid_0[3679:3672]) ? 1 : 0;
assign detect_min[459][10] = (mid_1[3687:3680] < mid_0[3687:3680]) ? 1 : 0;
assign detect_min[459][11] = (mid_1[3687:3680] < mid_0[3695:3688]) ? 1 : 0;
assign detect_min[459][12] = (mid_1[3687:3680] < mid_1[3679:3672]) ? 1 : 0;
assign detect_min[459][13] = (mid_1[3687:3680] < mid_1[3695:3688]) ? 1 : 0;
assign detect_min[459][14] = (mid_1[3687:3680] < mid_2[3679:3672]) ? 1 : 0;
assign detect_min[459][15] = (mid_1[3687:3680] < mid_2[3687:3680]) ? 1 : 0;
assign detect_min[459][16] = (mid_1[3687:3680] < mid_2[3695:3688]) ? 1 : 0;
assign detect_min[459][17] = (mid_1[3687:3680] < btm_0[3679:3672]) ? 1 : 0;
assign detect_min[459][18] = (mid_1[3687:3680] < btm_0[3687:3680]) ? 1 : 0;
assign detect_min[459][19] = (mid_1[3687:3680] < btm_0[3695:3688]) ? 1 : 0;
assign detect_min[459][20] = (mid_1[3687:3680] < btm_1[3679:3672]) ? 1 : 0;
assign detect_min[459][21] = (mid_1[3687:3680] < btm_1[3687:3680]) ? 1 : 0;
assign detect_min[459][22] = (mid_1[3687:3680] < btm_1[3695:3688]) ? 1 : 0;
assign detect_min[459][23] = (mid_1[3687:3680] < btm_2[3679:3672]) ? 1 : 0;
assign detect_min[459][24] = (mid_1[3687:3680] < btm_2[3687:3680]) ? 1 : 0;
assign detect_min[459][25] = (mid_1[3687:3680] < btm_2[3695:3688]) ? 1 : 0;

assign detect_min[460][0] = (mid_1[3695:3688] < top_0[3687:3680]) ? 1 : 0;
assign detect_min[460][1] = (mid_1[3695:3688] < top_0[3695:3688]) ? 1 : 0;
assign detect_min[460][2] = (mid_1[3695:3688] < top_0[3703:3696]) ? 1 : 0;
assign detect_min[460][3] = (mid_1[3695:3688] < top_1[3687:3680]) ? 1 : 0;
assign detect_min[460][4] = (mid_1[3695:3688] < top_1[3695:3688]) ? 1 : 0;
assign detect_min[460][5] = (mid_1[3695:3688] < top_1[3703:3696]) ? 1 : 0;
assign detect_min[460][6] = (mid_1[3695:3688] < top_2[3687:3680]) ? 1 : 0;
assign detect_min[460][7] = (mid_1[3695:3688] < top_2[3695:3688]) ? 1 : 0;
assign detect_min[460][8] = (mid_1[3695:3688] < top_2[3703:3696]) ? 1 : 0;
assign detect_min[460][9] = (mid_1[3695:3688] < mid_0[3687:3680]) ? 1 : 0;
assign detect_min[460][10] = (mid_1[3695:3688] < mid_0[3695:3688]) ? 1 : 0;
assign detect_min[460][11] = (mid_1[3695:3688] < mid_0[3703:3696]) ? 1 : 0;
assign detect_min[460][12] = (mid_1[3695:3688] < mid_1[3687:3680]) ? 1 : 0;
assign detect_min[460][13] = (mid_1[3695:3688] < mid_1[3703:3696]) ? 1 : 0;
assign detect_min[460][14] = (mid_1[3695:3688] < mid_2[3687:3680]) ? 1 : 0;
assign detect_min[460][15] = (mid_1[3695:3688] < mid_2[3695:3688]) ? 1 : 0;
assign detect_min[460][16] = (mid_1[3695:3688] < mid_2[3703:3696]) ? 1 : 0;
assign detect_min[460][17] = (mid_1[3695:3688] < btm_0[3687:3680]) ? 1 : 0;
assign detect_min[460][18] = (mid_1[3695:3688] < btm_0[3695:3688]) ? 1 : 0;
assign detect_min[460][19] = (mid_1[3695:3688] < btm_0[3703:3696]) ? 1 : 0;
assign detect_min[460][20] = (mid_1[3695:3688] < btm_1[3687:3680]) ? 1 : 0;
assign detect_min[460][21] = (mid_1[3695:3688] < btm_1[3695:3688]) ? 1 : 0;
assign detect_min[460][22] = (mid_1[3695:3688] < btm_1[3703:3696]) ? 1 : 0;
assign detect_min[460][23] = (mid_1[3695:3688] < btm_2[3687:3680]) ? 1 : 0;
assign detect_min[460][24] = (mid_1[3695:3688] < btm_2[3695:3688]) ? 1 : 0;
assign detect_min[460][25] = (mid_1[3695:3688] < btm_2[3703:3696]) ? 1 : 0;

assign detect_min[461][0] = (mid_1[3703:3696] < top_0[3695:3688]) ? 1 : 0;
assign detect_min[461][1] = (mid_1[3703:3696] < top_0[3703:3696]) ? 1 : 0;
assign detect_min[461][2] = (mid_1[3703:3696] < top_0[3711:3704]) ? 1 : 0;
assign detect_min[461][3] = (mid_1[3703:3696] < top_1[3695:3688]) ? 1 : 0;
assign detect_min[461][4] = (mid_1[3703:3696] < top_1[3703:3696]) ? 1 : 0;
assign detect_min[461][5] = (mid_1[3703:3696] < top_1[3711:3704]) ? 1 : 0;
assign detect_min[461][6] = (mid_1[3703:3696] < top_2[3695:3688]) ? 1 : 0;
assign detect_min[461][7] = (mid_1[3703:3696] < top_2[3703:3696]) ? 1 : 0;
assign detect_min[461][8] = (mid_1[3703:3696] < top_2[3711:3704]) ? 1 : 0;
assign detect_min[461][9] = (mid_1[3703:3696] < mid_0[3695:3688]) ? 1 : 0;
assign detect_min[461][10] = (mid_1[3703:3696] < mid_0[3703:3696]) ? 1 : 0;
assign detect_min[461][11] = (mid_1[3703:3696] < mid_0[3711:3704]) ? 1 : 0;
assign detect_min[461][12] = (mid_1[3703:3696] < mid_1[3695:3688]) ? 1 : 0;
assign detect_min[461][13] = (mid_1[3703:3696] < mid_1[3711:3704]) ? 1 : 0;
assign detect_min[461][14] = (mid_1[3703:3696] < mid_2[3695:3688]) ? 1 : 0;
assign detect_min[461][15] = (mid_1[3703:3696] < mid_2[3703:3696]) ? 1 : 0;
assign detect_min[461][16] = (mid_1[3703:3696] < mid_2[3711:3704]) ? 1 : 0;
assign detect_min[461][17] = (mid_1[3703:3696] < btm_0[3695:3688]) ? 1 : 0;
assign detect_min[461][18] = (mid_1[3703:3696] < btm_0[3703:3696]) ? 1 : 0;
assign detect_min[461][19] = (mid_1[3703:3696] < btm_0[3711:3704]) ? 1 : 0;
assign detect_min[461][20] = (mid_1[3703:3696] < btm_1[3695:3688]) ? 1 : 0;
assign detect_min[461][21] = (mid_1[3703:3696] < btm_1[3703:3696]) ? 1 : 0;
assign detect_min[461][22] = (mid_1[3703:3696] < btm_1[3711:3704]) ? 1 : 0;
assign detect_min[461][23] = (mid_1[3703:3696] < btm_2[3695:3688]) ? 1 : 0;
assign detect_min[461][24] = (mid_1[3703:3696] < btm_2[3703:3696]) ? 1 : 0;
assign detect_min[461][25] = (mid_1[3703:3696] < btm_2[3711:3704]) ? 1 : 0;

assign detect_min[462][0] = (mid_1[3711:3704] < top_0[3703:3696]) ? 1 : 0;
assign detect_min[462][1] = (mid_1[3711:3704] < top_0[3711:3704]) ? 1 : 0;
assign detect_min[462][2] = (mid_1[3711:3704] < top_0[3719:3712]) ? 1 : 0;
assign detect_min[462][3] = (mid_1[3711:3704] < top_1[3703:3696]) ? 1 : 0;
assign detect_min[462][4] = (mid_1[3711:3704] < top_1[3711:3704]) ? 1 : 0;
assign detect_min[462][5] = (mid_1[3711:3704] < top_1[3719:3712]) ? 1 : 0;
assign detect_min[462][6] = (mid_1[3711:3704] < top_2[3703:3696]) ? 1 : 0;
assign detect_min[462][7] = (mid_1[3711:3704] < top_2[3711:3704]) ? 1 : 0;
assign detect_min[462][8] = (mid_1[3711:3704] < top_2[3719:3712]) ? 1 : 0;
assign detect_min[462][9] = (mid_1[3711:3704] < mid_0[3703:3696]) ? 1 : 0;
assign detect_min[462][10] = (mid_1[3711:3704] < mid_0[3711:3704]) ? 1 : 0;
assign detect_min[462][11] = (mid_1[3711:3704] < mid_0[3719:3712]) ? 1 : 0;
assign detect_min[462][12] = (mid_1[3711:3704] < mid_1[3703:3696]) ? 1 : 0;
assign detect_min[462][13] = (mid_1[3711:3704] < mid_1[3719:3712]) ? 1 : 0;
assign detect_min[462][14] = (mid_1[3711:3704] < mid_2[3703:3696]) ? 1 : 0;
assign detect_min[462][15] = (mid_1[3711:3704] < mid_2[3711:3704]) ? 1 : 0;
assign detect_min[462][16] = (mid_1[3711:3704] < mid_2[3719:3712]) ? 1 : 0;
assign detect_min[462][17] = (mid_1[3711:3704] < btm_0[3703:3696]) ? 1 : 0;
assign detect_min[462][18] = (mid_1[3711:3704] < btm_0[3711:3704]) ? 1 : 0;
assign detect_min[462][19] = (mid_1[3711:3704] < btm_0[3719:3712]) ? 1 : 0;
assign detect_min[462][20] = (mid_1[3711:3704] < btm_1[3703:3696]) ? 1 : 0;
assign detect_min[462][21] = (mid_1[3711:3704] < btm_1[3711:3704]) ? 1 : 0;
assign detect_min[462][22] = (mid_1[3711:3704] < btm_1[3719:3712]) ? 1 : 0;
assign detect_min[462][23] = (mid_1[3711:3704] < btm_2[3703:3696]) ? 1 : 0;
assign detect_min[462][24] = (mid_1[3711:3704] < btm_2[3711:3704]) ? 1 : 0;
assign detect_min[462][25] = (mid_1[3711:3704] < btm_2[3719:3712]) ? 1 : 0;

assign detect_min[463][0] = (mid_1[3719:3712] < top_0[3711:3704]) ? 1 : 0;
assign detect_min[463][1] = (mid_1[3719:3712] < top_0[3719:3712]) ? 1 : 0;
assign detect_min[463][2] = (mid_1[3719:3712] < top_0[3727:3720]) ? 1 : 0;
assign detect_min[463][3] = (mid_1[3719:3712] < top_1[3711:3704]) ? 1 : 0;
assign detect_min[463][4] = (mid_1[3719:3712] < top_1[3719:3712]) ? 1 : 0;
assign detect_min[463][5] = (mid_1[3719:3712] < top_1[3727:3720]) ? 1 : 0;
assign detect_min[463][6] = (mid_1[3719:3712] < top_2[3711:3704]) ? 1 : 0;
assign detect_min[463][7] = (mid_1[3719:3712] < top_2[3719:3712]) ? 1 : 0;
assign detect_min[463][8] = (mid_1[3719:3712] < top_2[3727:3720]) ? 1 : 0;
assign detect_min[463][9] = (mid_1[3719:3712] < mid_0[3711:3704]) ? 1 : 0;
assign detect_min[463][10] = (mid_1[3719:3712] < mid_0[3719:3712]) ? 1 : 0;
assign detect_min[463][11] = (mid_1[3719:3712] < mid_0[3727:3720]) ? 1 : 0;
assign detect_min[463][12] = (mid_1[3719:3712] < mid_1[3711:3704]) ? 1 : 0;
assign detect_min[463][13] = (mid_1[3719:3712] < mid_1[3727:3720]) ? 1 : 0;
assign detect_min[463][14] = (mid_1[3719:3712] < mid_2[3711:3704]) ? 1 : 0;
assign detect_min[463][15] = (mid_1[3719:3712] < mid_2[3719:3712]) ? 1 : 0;
assign detect_min[463][16] = (mid_1[3719:3712] < mid_2[3727:3720]) ? 1 : 0;
assign detect_min[463][17] = (mid_1[3719:3712] < btm_0[3711:3704]) ? 1 : 0;
assign detect_min[463][18] = (mid_1[3719:3712] < btm_0[3719:3712]) ? 1 : 0;
assign detect_min[463][19] = (mid_1[3719:3712] < btm_0[3727:3720]) ? 1 : 0;
assign detect_min[463][20] = (mid_1[3719:3712] < btm_1[3711:3704]) ? 1 : 0;
assign detect_min[463][21] = (mid_1[3719:3712] < btm_1[3719:3712]) ? 1 : 0;
assign detect_min[463][22] = (mid_1[3719:3712] < btm_1[3727:3720]) ? 1 : 0;
assign detect_min[463][23] = (mid_1[3719:3712] < btm_2[3711:3704]) ? 1 : 0;
assign detect_min[463][24] = (mid_1[3719:3712] < btm_2[3719:3712]) ? 1 : 0;
assign detect_min[463][25] = (mid_1[3719:3712] < btm_2[3727:3720]) ? 1 : 0;

assign detect_min[464][0] = (mid_1[3727:3720] < top_0[3719:3712]) ? 1 : 0;
assign detect_min[464][1] = (mid_1[3727:3720] < top_0[3727:3720]) ? 1 : 0;
assign detect_min[464][2] = (mid_1[3727:3720] < top_0[3735:3728]) ? 1 : 0;
assign detect_min[464][3] = (mid_1[3727:3720] < top_1[3719:3712]) ? 1 : 0;
assign detect_min[464][4] = (mid_1[3727:3720] < top_1[3727:3720]) ? 1 : 0;
assign detect_min[464][5] = (mid_1[3727:3720] < top_1[3735:3728]) ? 1 : 0;
assign detect_min[464][6] = (mid_1[3727:3720] < top_2[3719:3712]) ? 1 : 0;
assign detect_min[464][7] = (mid_1[3727:3720] < top_2[3727:3720]) ? 1 : 0;
assign detect_min[464][8] = (mid_1[3727:3720] < top_2[3735:3728]) ? 1 : 0;
assign detect_min[464][9] = (mid_1[3727:3720] < mid_0[3719:3712]) ? 1 : 0;
assign detect_min[464][10] = (mid_1[3727:3720] < mid_0[3727:3720]) ? 1 : 0;
assign detect_min[464][11] = (mid_1[3727:3720] < mid_0[3735:3728]) ? 1 : 0;
assign detect_min[464][12] = (mid_1[3727:3720] < mid_1[3719:3712]) ? 1 : 0;
assign detect_min[464][13] = (mid_1[3727:3720] < mid_1[3735:3728]) ? 1 : 0;
assign detect_min[464][14] = (mid_1[3727:3720] < mid_2[3719:3712]) ? 1 : 0;
assign detect_min[464][15] = (mid_1[3727:3720] < mid_2[3727:3720]) ? 1 : 0;
assign detect_min[464][16] = (mid_1[3727:3720] < mid_2[3735:3728]) ? 1 : 0;
assign detect_min[464][17] = (mid_1[3727:3720] < btm_0[3719:3712]) ? 1 : 0;
assign detect_min[464][18] = (mid_1[3727:3720] < btm_0[3727:3720]) ? 1 : 0;
assign detect_min[464][19] = (mid_1[3727:3720] < btm_0[3735:3728]) ? 1 : 0;
assign detect_min[464][20] = (mid_1[3727:3720] < btm_1[3719:3712]) ? 1 : 0;
assign detect_min[464][21] = (mid_1[3727:3720] < btm_1[3727:3720]) ? 1 : 0;
assign detect_min[464][22] = (mid_1[3727:3720] < btm_1[3735:3728]) ? 1 : 0;
assign detect_min[464][23] = (mid_1[3727:3720] < btm_2[3719:3712]) ? 1 : 0;
assign detect_min[464][24] = (mid_1[3727:3720] < btm_2[3727:3720]) ? 1 : 0;
assign detect_min[464][25] = (mid_1[3727:3720] < btm_2[3735:3728]) ? 1 : 0;

assign detect_min[465][0] = (mid_1[3735:3728] < top_0[3727:3720]) ? 1 : 0;
assign detect_min[465][1] = (mid_1[3735:3728] < top_0[3735:3728]) ? 1 : 0;
assign detect_min[465][2] = (mid_1[3735:3728] < top_0[3743:3736]) ? 1 : 0;
assign detect_min[465][3] = (mid_1[3735:3728] < top_1[3727:3720]) ? 1 : 0;
assign detect_min[465][4] = (mid_1[3735:3728] < top_1[3735:3728]) ? 1 : 0;
assign detect_min[465][5] = (mid_1[3735:3728] < top_1[3743:3736]) ? 1 : 0;
assign detect_min[465][6] = (mid_1[3735:3728] < top_2[3727:3720]) ? 1 : 0;
assign detect_min[465][7] = (mid_1[3735:3728] < top_2[3735:3728]) ? 1 : 0;
assign detect_min[465][8] = (mid_1[3735:3728] < top_2[3743:3736]) ? 1 : 0;
assign detect_min[465][9] = (mid_1[3735:3728] < mid_0[3727:3720]) ? 1 : 0;
assign detect_min[465][10] = (mid_1[3735:3728] < mid_0[3735:3728]) ? 1 : 0;
assign detect_min[465][11] = (mid_1[3735:3728] < mid_0[3743:3736]) ? 1 : 0;
assign detect_min[465][12] = (mid_1[3735:3728] < mid_1[3727:3720]) ? 1 : 0;
assign detect_min[465][13] = (mid_1[3735:3728] < mid_1[3743:3736]) ? 1 : 0;
assign detect_min[465][14] = (mid_1[3735:3728] < mid_2[3727:3720]) ? 1 : 0;
assign detect_min[465][15] = (mid_1[3735:3728] < mid_2[3735:3728]) ? 1 : 0;
assign detect_min[465][16] = (mid_1[3735:3728] < mid_2[3743:3736]) ? 1 : 0;
assign detect_min[465][17] = (mid_1[3735:3728] < btm_0[3727:3720]) ? 1 : 0;
assign detect_min[465][18] = (mid_1[3735:3728] < btm_0[3735:3728]) ? 1 : 0;
assign detect_min[465][19] = (mid_1[3735:3728] < btm_0[3743:3736]) ? 1 : 0;
assign detect_min[465][20] = (mid_1[3735:3728] < btm_1[3727:3720]) ? 1 : 0;
assign detect_min[465][21] = (mid_1[3735:3728] < btm_1[3735:3728]) ? 1 : 0;
assign detect_min[465][22] = (mid_1[3735:3728] < btm_1[3743:3736]) ? 1 : 0;
assign detect_min[465][23] = (mid_1[3735:3728] < btm_2[3727:3720]) ? 1 : 0;
assign detect_min[465][24] = (mid_1[3735:3728] < btm_2[3735:3728]) ? 1 : 0;
assign detect_min[465][25] = (mid_1[3735:3728] < btm_2[3743:3736]) ? 1 : 0;

assign detect_min[466][0] = (mid_1[3743:3736] < top_0[3735:3728]) ? 1 : 0;
assign detect_min[466][1] = (mid_1[3743:3736] < top_0[3743:3736]) ? 1 : 0;
assign detect_min[466][2] = (mid_1[3743:3736] < top_0[3751:3744]) ? 1 : 0;
assign detect_min[466][3] = (mid_1[3743:3736] < top_1[3735:3728]) ? 1 : 0;
assign detect_min[466][4] = (mid_1[3743:3736] < top_1[3743:3736]) ? 1 : 0;
assign detect_min[466][5] = (mid_1[3743:3736] < top_1[3751:3744]) ? 1 : 0;
assign detect_min[466][6] = (mid_1[3743:3736] < top_2[3735:3728]) ? 1 : 0;
assign detect_min[466][7] = (mid_1[3743:3736] < top_2[3743:3736]) ? 1 : 0;
assign detect_min[466][8] = (mid_1[3743:3736] < top_2[3751:3744]) ? 1 : 0;
assign detect_min[466][9] = (mid_1[3743:3736] < mid_0[3735:3728]) ? 1 : 0;
assign detect_min[466][10] = (mid_1[3743:3736] < mid_0[3743:3736]) ? 1 : 0;
assign detect_min[466][11] = (mid_1[3743:3736] < mid_0[3751:3744]) ? 1 : 0;
assign detect_min[466][12] = (mid_1[3743:3736] < mid_1[3735:3728]) ? 1 : 0;
assign detect_min[466][13] = (mid_1[3743:3736] < mid_1[3751:3744]) ? 1 : 0;
assign detect_min[466][14] = (mid_1[3743:3736] < mid_2[3735:3728]) ? 1 : 0;
assign detect_min[466][15] = (mid_1[3743:3736] < mid_2[3743:3736]) ? 1 : 0;
assign detect_min[466][16] = (mid_1[3743:3736] < mid_2[3751:3744]) ? 1 : 0;
assign detect_min[466][17] = (mid_1[3743:3736] < btm_0[3735:3728]) ? 1 : 0;
assign detect_min[466][18] = (mid_1[3743:3736] < btm_0[3743:3736]) ? 1 : 0;
assign detect_min[466][19] = (mid_1[3743:3736] < btm_0[3751:3744]) ? 1 : 0;
assign detect_min[466][20] = (mid_1[3743:3736] < btm_1[3735:3728]) ? 1 : 0;
assign detect_min[466][21] = (mid_1[3743:3736] < btm_1[3743:3736]) ? 1 : 0;
assign detect_min[466][22] = (mid_1[3743:3736] < btm_1[3751:3744]) ? 1 : 0;
assign detect_min[466][23] = (mid_1[3743:3736] < btm_2[3735:3728]) ? 1 : 0;
assign detect_min[466][24] = (mid_1[3743:3736] < btm_2[3743:3736]) ? 1 : 0;
assign detect_min[466][25] = (mid_1[3743:3736] < btm_2[3751:3744]) ? 1 : 0;

assign detect_min[467][0] = (mid_1[3751:3744] < top_0[3743:3736]) ? 1 : 0;
assign detect_min[467][1] = (mid_1[3751:3744] < top_0[3751:3744]) ? 1 : 0;
assign detect_min[467][2] = (mid_1[3751:3744] < top_0[3759:3752]) ? 1 : 0;
assign detect_min[467][3] = (mid_1[3751:3744] < top_1[3743:3736]) ? 1 : 0;
assign detect_min[467][4] = (mid_1[3751:3744] < top_1[3751:3744]) ? 1 : 0;
assign detect_min[467][5] = (mid_1[3751:3744] < top_1[3759:3752]) ? 1 : 0;
assign detect_min[467][6] = (mid_1[3751:3744] < top_2[3743:3736]) ? 1 : 0;
assign detect_min[467][7] = (mid_1[3751:3744] < top_2[3751:3744]) ? 1 : 0;
assign detect_min[467][8] = (mid_1[3751:3744] < top_2[3759:3752]) ? 1 : 0;
assign detect_min[467][9] = (mid_1[3751:3744] < mid_0[3743:3736]) ? 1 : 0;
assign detect_min[467][10] = (mid_1[3751:3744] < mid_0[3751:3744]) ? 1 : 0;
assign detect_min[467][11] = (mid_1[3751:3744] < mid_0[3759:3752]) ? 1 : 0;
assign detect_min[467][12] = (mid_1[3751:3744] < mid_1[3743:3736]) ? 1 : 0;
assign detect_min[467][13] = (mid_1[3751:3744] < mid_1[3759:3752]) ? 1 : 0;
assign detect_min[467][14] = (mid_1[3751:3744] < mid_2[3743:3736]) ? 1 : 0;
assign detect_min[467][15] = (mid_1[3751:3744] < mid_2[3751:3744]) ? 1 : 0;
assign detect_min[467][16] = (mid_1[3751:3744] < mid_2[3759:3752]) ? 1 : 0;
assign detect_min[467][17] = (mid_1[3751:3744] < btm_0[3743:3736]) ? 1 : 0;
assign detect_min[467][18] = (mid_1[3751:3744] < btm_0[3751:3744]) ? 1 : 0;
assign detect_min[467][19] = (mid_1[3751:3744] < btm_0[3759:3752]) ? 1 : 0;
assign detect_min[467][20] = (mid_1[3751:3744] < btm_1[3743:3736]) ? 1 : 0;
assign detect_min[467][21] = (mid_1[3751:3744] < btm_1[3751:3744]) ? 1 : 0;
assign detect_min[467][22] = (mid_1[3751:3744] < btm_1[3759:3752]) ? 1 : 0;
assign detect_min[467][23] = (mid_1[3751:3744] < btm_2[3743:3736]) ? 1 : 0;
assign detect_min[467][24] = (mid_1[3751:3744] < btm_2[3751:3744]) ? 1 : 0;
assign detect_min[467][25] = (mid_1[3751:3744] < btm_2[3759:3752]) ? 1 : 0;

assign detect_min[468][0] = (mid_1[3759:3752] < top_0[3751:3744]) ? 1 : 0;
assign detect_min[468][1] = (mid_1[3759:3752] < top_0[3759:3752]) ? 1 : 0;
assign detect_min[468][2] = (mid_1[3759:3752] < top_0[3767:3760]) ? 1 : 0;
assign detect_min[468][3] = (mid_1[3759:3752] < top_1[3751:3744]) ? 1 : 0;
assign detect_min[468][4] = (mid_1[3759:3752] < top_1[3759:3752]) ? 1 : 0;
assign detect_min[468][5] = (mid_1[3759:3752] < top_1[3767:3760]) ? 1 : 0;
assign detect_min[468][6] = (mid_1[3759:3752] < top_2[3751:3744]) ? 1 : 0;
assign detect_min[468][7] = (mid_1[3759:3752] < top_2[3759:3752]) ? 1 : 0;
assign detect_min[468][8] = (mid_1[3759:3752] < top_2[3767:3760]) ? 1 : 0;
assign detect_min[468][9] = (mid_1[3759:3752] < mid_0[3751:3744]) ? 1 : 0;
assign detect_min[468][10] = (mid_1[3759:3752] < mid_0[3759:3752]) ? 1 : 0;
assign detect_min[468][11] = (mid_1[3759:3752] < mid_0[3767:3760]) ? 1 : 0;
assign detect_min[468][12] = (mid_1[3759:3752] < mid_1[3751:3744]) ? 1 : 0;
assign detect_min[468][13] = (mid_1[3759:3752] < mid_1[3767:3760]) ? 1 : 0;
assign detect_min[468][14] = (mid_1[3759:3752] < mid_2[3751:3744]) ? 1 : 0;
assign detect_min[468][15] = (mid_1[3759:3752] < mid_2[3759:3752]) ? 1 : 0;
assign detect_min[468][16] = (mid_1[3759:3752] < mid_2[3767:3760]) ? 1 : 0;
assign detect_min[468][17] = (mid_1[3759:3752] < btm_0[3751:3744]) ? 1 : 0;
assign detect_min[468][18] = (mid_1[3759:3752] < btm_0[3759:3752]) ? 1 : 0;
assign detect_min[468][19] = (mid_1[3759:3752] < btm_0[3767:3760]) ? 1 : 0;
assign detect_min[468][20] = (mid_1[3759:3752] < btm_1[3751:3744]) ? 1 : 0;
assign detect_min[468][21] = (mid_1[3759:3752] < btm_1[3759:3752]) ? 1 : 0;
assign detect_min[468][22] = (mid_1[3759:3752] < btm_1[3767:3760]) ? 1 : 0;
assign detect_min[468][23] = (mid_1[3759:3752] < btm_2[3751:3744]) ? 1 : 0;
assign detect_min[468][24] = (mid_1[3759:3752] < btm_2[3759:3752]) ? 1 : 0;
assign detect_min[468][25] = (mid_1[3759:3752] < btm_2[3767:3760]) ? 1 : 0;

assign detect_min[469][0] = (mid_1[3767:3760] < top_0[3759:3752]) ? 1 : 0;
assign detect_min[469][1] = (mid_1[3767:3760] < top_0[3767:3760]) ? 1 : 0;
assign detect_min[469][2] = (mid_1[3767:3760] < top_0[3775:3768]) ? 1 : 0;
assign detect_min[469][3] = (mid_1[3767:3760] < top_1[3759:3752]) ? 1 : 0;
assign detect_min[469][4] = (mid_1[3767:3760] < top_1[3767:3760]) ? 1 : 0;
assign detect_min[469][5] = (mid_1[3767:3760] < top_1[3775:3768]) ? 1 : 0;
assign detect_min[469][6] = (mid_1[3767:3760] < top_2[3759:3752]) ? 1 : 0;
assign detect_min[469][7] = (mid_1[3767:3760] < top_2[3767:3760]) ? 1 : 0;
assign detect_min[469][8] = (mid_1[3767:3760] < top_2[3775:3768]) ? 1 : 0;
assign detect_min[469][9] = (mid_1[3767:3760] < mid_0[3759:3752]) ? 1 : 0;
assign detect_min[469][10] = (mid_1[3767:3760] < mid_0[3767:3760]) ? 1 : 0;
assign detect_min[469][11] = (mid_1[3767:3760] < mid_0[3775:3768]) ? 1 : 0;
assign detect_min[469][12] = (mid_1[3767:3760] < mid_1[3759:3752]) ? 1 : 0;
assign detect_min[469][13] = (mid_1[3767:3760] < mid_1[3775:3768]) ? 1 : 0;
assign detect_min[469][14] = (mid_1[3767:3760] < mid_2[3759:3752]) ? 1 : 0;
assign detect_min[469][15] = (mid_1[3767:3760] < mid_2[3767:3760]) ? 1 : 0;
assign detect_min[469][16] = (mid_1[3767:3760] < mid_2[3775:3768]) ? 1 : 0;
assign detect_min[469][17] = (mid_1[3767:3760] < btm_0[3759:3752]) ? 1 : 0;
assign detect_min[469][18] = (mid_1[3767:3760] < btm_0[3767:3760]) ? 1 : 0;
assign detect_min[469][19] = (mid_1[3767:3760] < btm_0[3775:3768]) ? 1 : 0;
assign detect_min[469][20] = (mid_1[3767:3760] < btm_1[3759:3752]) ? 1 : 0;
assign detect_min[469][21] = (mid_1[3767:3760] < btm_1[3767:3760]) ? 1 : 0;
assign detect_min[469][22] = (mid_1[3767:3760] < btm_1[3775:3768]) ? 1 : 0;
assign detect_min[469][23] = (mid_1[3767:3760] < btm_2[3759:3752]) ? 1 : 0;
assign detect_min[469][24] = (mid_1[3767:3760] < btm_2[3767:3760]) ? 1 : 0;
assign detect_min[469][25] = (mid_1[3767:3760] < btm_2[3775:3768]) ? 1 : 0;

assign detect_min[470][0] = (mid_1[3775:3768] < top_0[3767:3760]) ? 1 : 0;
assign detect_min[470][1] = (mid_1[3775:3768] < top_0[3775:3768]) ? 1 : 0;
assign detect_min[470][2] = (mid_1[3775:3768] < top_0[3783:3776]) ? 1 : 0;
assign detect_min[470][3] = (mid_1[3775:3768] < top_1[3767:3760]) ? 1 : 0;
assign detect_min[470][4] = (mid_1[3775:3768] < top_1[3775:3768]) ? 1 : 0;
assign detect_min[470][5] = (mid_1[3775:3768] < top_1[3783:3776]) ? 1 : 0;
assign detect_min[470][6] = (mid_1[3775:3768] < top_2[3767:3760]) ? 1 : 0;
assign detect_min[470][7] = (mid_1[3775:3768] < top_2[3775:3768]) ? 1 : 0;
assign detect_min[470][8] = (mid_1[3775:3768] < top_2[3783:3776]) ? 1 : 0;
assign detect_min[470][9] = (mid_1[3775:3768] < mid_0[3767:3760]) ? 1 : 0;
assign detect_min[470][10] = (mid_1[3775:3768] < mid_0[3775:3768]) ? 1 : 0;
assign detect_min[470][11] = (mid_1[3775:3768] < mid_0[3783:3776]) ? 1 : 0;
assign detect_min[470][12] = (mid_1[3775:3768] < mid_1[3767:3760]) ? 1 : 0;
assign detect_min[470][13] = (mid_1[3775:3768] < mid_1[3783:3776]) ? 1 : 0;
assign detect_min[470][14] = (mid_1[3775:3768] < mid_2[3767:3760]) ? 1 : 0;
assign detect_min[470][15] = (mid_1[3775:3768] < mid_2[3775:3768]) ? 1 : 0;
assign detect_min[470][16] = (mid_1[3775:3768] < mid_2[3783:3776]) ? 1 : 0;
assign detect_min[470][17] = (mid_1[3775:3768] < btm_0[3767:3760]) ? 1 : 0;
assign detect_min[470][18] = (mid_1[3775:3768] < btm_0[3775:3768]) ? 1 : 0;
assign detect_min[470][19] = (mid_1[3775:3768] < btm_0[3783:3776]) ? 1 : 0;
assign detect_min[470][20] = (mid_1[3775:3768] < btm_1[3767:3760]) ? 1 : 0;
assign detect_min[470][21] = (mid_1[3775:3768] < btm_1[3775:3768]) ? 1 : 0;
assign detect_min[470][22] = (mid_1[3775:3768] < btm_1[3783:3776]) ? 1 : 0;
assign detect_min[470][23] = (mid_1[3775:3768] < btm_2[3767:3760]) ? 1 : 0;
assign detect_min[470][24] = (mid_1[3775:3768] < btm_2[3775:3768]) ? 1 : 0;
assign detect_min[470][25] = (mid_1[3775:3768] < btm_2[3783:3776]) ? 1 : 0;

assign detect_min[471][0] = (mid_1[3783:3776] < top_0[3775:3768]) ? 1 : 0;
assign detect_min[471][1] = (mid_1[3783:3776] < top_0[3783:3776]) ? 1 : 0;
assign detect_min[471][2] = (mid_1[3783:3776] < top_0[3791:3784]) ? 1 : 0;
assign detect_min[471][3] = (mid_1[3783:3776] < top_1[3775:3768]) ? 1 : 0;
assign detect_min[471][4] = (mid_1[3783:3776] < top_1[3783:3776]) ? 1 : 0;
assign detect_min[471][5] = (mid_1[3783:3776] < top_1[3791:3784]) ? 1 : 0;
assign detect_min[471][6] = (mid_1[3783:3776] < top_2[3775:3768]) ? 1 : 0;
assign detect_min[471][7] = (mid_1[3783:3776] < top_2[3783:3776]) ? 1 : 0;
assign detect_min[471][8] = (mid_1[3783:3776] < top_2[3791:3784]) ? 1 : 0;
assign detect_min[471][9] = (mid_1[3783:3776] < mid_0[3775:3768]) ? 1 : 0;
assign detect_min[471][10] = (mid_1[3783:3776] < mid_0[3783:3776]) ? 1 : 0;
assign detect_min[471][11] = (mid_1[3783:3776] < mid_0[3791:3784]) ? 1 : 0;
assign detect_min[471][12] = (mid_1[3783:3776] < mid_1[3775:3768]) ? 1 : 0;
assign detect_min[471][13] = (mid_1[3783:3776] < mid_1[3791:3784]) ? 1 : 0;
assign detect_min[471][14] = (mid_1[3783:3776] < mid_2[3775:3768]) ? 1 : 0;
assign detect_min[471][15] = (mid_1[3783:3776] < mid_2[3783:3776]) ? 1 : 0;
assign detect_min[471][16] = (mid_1[3783:3776] < mid_2[3791:3784]) ? 1 : 0;
assign detect_min[471][17] = (mid_1[3783:3776] < btm_0[3775:3768]) ? 1 : 0;
assign detect_min[471][18] = (mid_1[3783:3776] < btm_0[3783:3776]) ? 1 : 0;
assign detect_min[471][19] = (mid_1[3783:3776] < btm_0[3791:3784]) ? 1 : 0;
assign detect_min[471][20] = (mid_1[3783:3776] < btm_1[3775:3768]) ? 1 : 0;
assign detect_min[471][21] = (mid_1[3783:3776] < btm_1[3783:3776]) ? 1 : 0;
assign detect_min[471][22] = (mid_1[3783:3776] < btm_1[3791:3784]) ? 1 : 0;
assign detect_min[471][23] = (mid_1[3783:3776] < btm_2[3775:3768]) ? 1 : 0;
assign detect_min[471][24] = (mid_1[3783:3776] < btm_2[3783:3776]) ? 1 : 0;
assign detect_min[471][25] = (mid_1[3783:3776] < btm_2[3791:3784]) ? 1 : 0;

assign detect_min[472][0] = (mid_1[3791:3784] < top_0[3783:3776]) ? 1 : 0;
assign detect_min[472][1] = (mid_1[3791:3784] < top_0[3791:3784]) ? 1 : 0;
assign detect_min[472][2] = (mid_1[3791:3784] < top_0[3799:3792]) ? 1 : 0;
assign detect_min[472][3] = (mid_1[3791:3784] < top_1[3783:3776]) ? 1 : 0;
assign detect_min[472][4] = (mid_1[3791:3784] < top_1[3791:3784]) ? 1 : 0;
assign detect_min[472][5] = (mid_1[3791:3784] < top_1[3799:3792]) ? 1 : 0;
assign detect_min[472][6] = (mid_1[3791:3784] < top_2[3783:3776]) ? 1 : 0;
assign detect_min[472][7] = (mid_1[3791:3784] < top_2[3791:3784]) ? 1 : 0;
assign detect_min[472][8] = (mid_1[3791:3784] < top_2[3799:3792]) ? 1 : 0;
assign detect_min[472][9] = (mid_1[3791:3784] < mid_0[3783:3776]) ? 1 : 0;
assign detect_min[472][10] = (mid_1[3791:3784] < mid_0[3791:3784]) ? 1 : 0;
assign detect_min[472][11] = (mid_1[3791:3784] < mid_0[3799:3792]) ? 1 : 0;
assign detect_min[472][12] = (mid_1[3791:3784] < mid_1[3783:3776]) ? 1 : 0;
assign detect_min[472][13] = (mid_1[3791:3784] < mid_1[3799:3792]) ? 1 : 0;
assign detect_min[472][14] = (mid_1[3791:3784] < mid_2[3783:3776]) ? 1 : 0;
assign detect_min[472][15] = (mid_1[3791:3784] < mid_2[3791:3784]) ? 1 : 0;
assign detect_min[472][16] = (mid_1[3791:3784] < mid_2[3799:3792]) ? 1 : 0;
assign detect_min[472][17] = (mid_1[3791:3784] < btm_0[3783:3776]) ? 1 : 0;
assign detect_min[472][18] = (mid_1[3791:3784] < btm_0[3791:3784]) ? 1 : 0;
assign detect_min[472][19] = (mid_1[3791:3784] < btm_0[3799:3792]) ? 1 : 0;
assign detect_min[472][20] = (mid_1[3791:3784] < btm_1[3783:3776]) ? 1 : 0;
assign detect_min[472][21] = (mid_1[3791:3784] < btm_1[3791:3784]) ? 1 : 0;
assign detect_min[472][22] = (mid_1[3791:3784] < btm_1[3799:3792]) ? 1 : 0;
assign detect_min[472][23] = (mid_1[3791:3784] < btm_2[3783:3776]) ? 1 : 0;
assign detect_min[472][24] = (mid_1[3791:3784] < btm_2[3791:3784]) ? 1 : 0;
assign detect_min[472][25] = (mid_1[3791:3784] < btm_2[3799:3792]) ? 1 : 0;

assign detect_min[473][0] = (mid_1[3799:3792] < top_0[3791:3784]) ? 1 : 0;
assign detect_min[473][1] = (mid_1[3799:3792] < top_0[3799:3792]) ? 1 : 0;
assign detect_min[473][2] = (mid_1[3799:3792] < top_0[3807:3800]) ? 1 : 0;
assign detect_min[473][3] = (mid_1[3799:3792] < top_1[3791:3784]) ? 1 : 0;
assign detect_min[473][4] = (mid_1[3799:3792] < top_1[3799:3792]) ? 1 : 0;
assign detect_min[473][5] = (mid_1[3799:3792] < top_1[3807:3800]) ? 1 : 0;
assign detect_min[473][6] = (mid_1[3799:3792] < top_2[3791:3784]) ? 1 : 0;
assign detect_min[473][7] = (mid_1[3799:3792] < top_2[3799:3792]) ? 1 : 0;
assign detect_min[473][8] = (mid_1[3799:3792] < top_2[3807:3800]) ? 1 : 0;
assign detect_min[473][9] = (mid_1[3799:3792] < mid_0[3791:3784]) ? 1 : 0;
assign detect_min[473][10] = (mid_1[3799:3792] < mid_0[3799:3792]) ? 1 : 0;
assign detect_min[473][11] = (mid_1[3799:3792] < mid_0[3807:3800]) ? 1 : 0;
assign detect_min[473][12] = (mid_1[3799:3792] < mid_1[3791:3784]) ? 1 : 0;
assign detect_min[473][13] = (mid_1[3799:3792] < mid_1[3807:3800]) ? 1 : 0;
assign detect_min[473][14] = (mid_1[3799:3792] < mid_2[3791:3784]) ? 1 : 0;
assign detect_min[473][15] = (mid_1[3799:3792] < mid_2[3799:3792]) ? 1 : 0;
assign detect_min[473][16] = (mid_1[3799:3792] < mid_2[3807:3800]) ? 1 : 0;
assign detect_min[473][17] = (mid_1[3799:3792] < btm_0[3791:3784]) ? 1 : 0;
assign detect_min[473][18] = (mid_1[3799:3792] < btm_0[3799:3792]) ? 1 : 0;
assign detect_min[473][19] = (mid_1[3799:3792] < btm_0[3807:3800]) ? 1 : 0;
assign detect_min[473][20] = (mid_1[3799:3792] < btm_1[3791:3784]) ? 1 : 0;
assign detect_min[473][21] = (mid_1[3799:3792] < btm_1[3799:3792]) ? 1 : 0;
assign detect_min[473][22] = (mid_1[3799:3792] < btm_1[3807:3800]) ? 1 : 0;
assign detect_min[473][23] = (mid_1[3799:3792] < btm_2[3791:3784]) ? 1 : 0;
assign detect_min[473][24] = (mid_1[3799:3792] < btm_2[3799:3792]) ? 1 : 0;
assign detect_min[473][25] = (mid_1[3799:3792] < btm_2[3807:3800]) ? 1 : 0;

assign detect_min[474][0] = (mid_1[3807:3800] < top_0[3799:3792]) ? 1 : 0;
assign detect_min[474][1] = (mid_1[3807:3800] < top_0[3807:3800]) ? 1 : 0;
assign detect_min[474][2] = (mid_1[3807:3800] < top_0[3815:3808]) ? 1 : 0;
assign detect_min[474][3] = (mid_1[3807:3800] < top_1[3799:3792]) ? 1 : 0;
assign detect_min[474][4] = (mid_1[3807:3800] < top_1[3807:3800]) ? 1 : 0;
assign detect_min[474][5] = (mid_1[3807:3800] < top_1[3815:3808]) ? 1 : 0;
assign detect_min[474][6] = (mid_1[3807:3800] < top_2[3799:3792]) ? 1 : 0;
assign detect_min[474][7] = (mid_1[3807:3800] < top_2[3807:3800]) ? 1 : 0;
assign detect_min[474][8] = (mid_1[3807:3800] < top_2[3815:3808]) ? 1 : 0;
assign detect_min[474][9] = (mid_1[3807:3800] < mid_0[3799:3792]) ? 1 : 0;
assign detect_min[474][10] = (mid_1[3807:3800] < mid_0[3807:3800]) ? 1 : 0;
assign detect_min[474][11] = (mid_1[3807:3800] < mid_0[3815:3808]) ? 1 : 0;
assign detect_min[474][12] = (mid_1[3807:3800] < mid_1[3799:3792]) ? 1 : 0;
assign detect_min[474][13] = (mid_1[3807:3800] < mid_1[3815:3808]) ? 1 : 0;
assign detect_min[474][14] = (mid_1[3807:3800] < mid_2[3799:3792]) ? 1 : 0;
assign detect_min[474][15] = (mid_1[3807:3800] < mid_2[3807:3800]) ? 1 : 0;
assign detect_min[474][16] = (mid_1[3807:3800] < mid_2[3815:3808]) ? 1 : 0;
assign detect_min[474][17] = (mid_1[3807:3800] < btm_0[3799:3792]) ? 1 : 0;
assign detect_min[474][18] = (mid_1[3807:3800] < btm_0[3807:3800]) ? 1 : 0;
assign detect_min[474][19] = (mid_1[3807:3800] < btm_0[3815:3808]) ? 1 : 0;
assign detect_min[474][20] = (mid_1[3807:3800] < btm_1[3799:3792]) ? 1 : 0;
assign detect_min[474][21] = (mid_1[3807:3800] < btm_1[3807:3800]) ? 1 : 0;
assign detect_min[474][22] = (mid_1[3807:3800] < btm_1[3815:3808]) ? 1 : 0;
assign detect_min[474][23] = (mid_1[3807:3800] < btm_2[3799:3792]) ? 1 : 0;
assign detect_min[474][24] = (mid_1[3807:3800] < btm_2[3807:3800]) ? 1 : 0;
assign detect_min[474][25] = (mid_1[3807:3800] < btm_2[3815:3808]) ? 1 : 0;

assign detect_min[475][0] = (mid_1[3815:3808] < top_0[3807:3800]) ? 1 : 0;
assign detect_min[475][1] = (mid_1[3815:3808] < top_0[3815:3808]) ? 1 : 0;
assign detect_min[475][2] = (mid_1[3815:3808] < top_0[3823:3816]) ? 1 : 0;
assign detect_min[475][3] = (mid_1[3815:3808] < top_1[3807:3800]) ? 1 : 0;
assign detect_min[475][4] = (mid_1[3815:3808] < top_1[3815:3808]) ? 1 : 0;
assign detect_min[475][5] = (mid_1[3815:3808] < top_1[3823:3816]) ? 1 : 0;
assign detect_min[475][6] = (mid_1[3815:3808] < top_2[3807:3800]) ? 1 : 0;
assign detect_min[475][7] = (mid_1[3815:3808] < top_2[3815:3808]) ? 1 : 0;
assign detect_min[475][8] = (mid_1[3815:3808] < top_2[3823:3816]) ? 1 : 0;
assign detect_min[475][9] = (mid_1[3815:3808] < mid_0[3807:3800]) ? 1 : 0;
assign detect_min[475][10] = (mid_1[3815:3808] < mid_0[3815:3808]) ? 1 : 0;
assign detect_min[475][11] = (mid_1[3815:3808] < mid_0[3823:3816]) ? 1 : 0;
assign detect_min[475][12] = (mid_1[3815:3808] < mid_1[3807:3800]) ? 1 : 0;
assign detect_min[475][13] = (mid_1[3815:3808] < mid_1[3823:3816]) ? 1 : 0;
assign detect_min[475][14] = (mid_1[3815:3808] < mid_2[3807:3800]) ? 1 : 0;
assign detect_min[475][15] = (mid_1[3815:3808] < mid_2[3815:3808]) ? 1 : 0;
assign detect_min[475][16] = (mid_1[3815:3808] < mid_2[3823:3816]) ? 1 : 0;
assign detect_min[475][17] = (mid_1[3815:3808] < btm_0[3807:3800]) ? 1 : 0;
assign detect_min[475][18] = (mid_1[3815:3808] < btm_0[3815:3808]) ? 1 : 0;
assign detect_min[475][19] = (mid_1[3815:3808] < btm_0[3823:3816]) ? 1 : 0;
assign detect_min[475][20] = (mid_1[3815:3808] < btm_1[3807:3800]) ? 1 : 0;
assign detect_min[475][21] = (mid_1[3815:3808] < btm_1[3815:3808]) ? 1 : 0;
assign detect_min[475][22] = (mid_1[3815:3808] < btm_1[3823:3816]) ? 1 : 0;
assign detect_min[475][23] = (mid_1[3815:3808] < btm_2[3807:3800]) ? 1 : 0;
assign detect_min[475][24] = (mid_1[3815:3808] < btm_2[3815:3808]) ? 1 : 0;
assign detect_min[475][25] = (mid_1[3815:3808] < btm_2[3823:3816]) ? 1 : 0;

assign detect_min[476][0] = (mid_1[3823:3816] < top_0[3815:3808]) ? 1 : 0;
assign detect_min[476][1] = (mid_1[3823:3816] < top_0[3823:3816]) ? 1 : 0;
assign detect_min[476][2] = (mid_1[3823:3816] < top_0[3831:3824]) ? 1 : 0;
assign detect_min[476][3] = (mid_1[3823:3816] < top_1[3815:3808]) ? 1 : 0;
assign detect_min[476][4] = (mid_1[3823:3816] < top_1[3823:3816]) ? 1 : 0;
assign detect_min[476][5] = (mid_1[3823:3816] < top_1[3831:3824]) ? 1 : 0;
assign detect_min[476][6] = (mid_1[3823:3816] < top_2[3815:3808]) ? 1 : 0;
assign detect_min[476][7] = (mid_1[3823:3816] < top_2[3823:3816]) ? 1 : 0;
assign detect_min[476][8] = (mid_1[3823:3816] < top_2[3831:3824]) ? 1 : 0;
assign detect_min[476][9] = (mid_1[3823:3816] < mid_0[3815:3808]) ? 1 : 0;
assign detect_min[476][10] = (mid_1[3823:3816] < mid_0[3823:3816]) ? 1 : 0;
assign detect_min[476][11] = (mid_1[3823:3816] < mid_0[3831:3824]) ? 1 : 0;
assign detect_min[476][12] = (mid_1[3823:3816] < mid_1[3815:3808]) ? 1 : 0;
assign detect_min[476][13] = (mid_1[3823:3816] < mid_1[3831:3824]) ? 1 : 0;
assign detect_min[476][14] = (mid_1[3823:3816] < mid_2[3815:3808]) ? 1 : 0;
assign detect_min[476][15] = (mid_1[3823:3816] < mid_2[3823:3816]) ? 1 : 0;
assign detect_min[476][16] = (mid_1[3823:3816] < mid_2[3831:3824]) ? 1 : 0;
assign detect_min[476][17] = (mid_1[3823:3816] < btm_0[3815:3808]) ? 1 : 0;
assign detect_min[476][18] = (mid_1[3823:3816] < btm_0[3823:3816]) ? 1 : 0;
assign detect_min[476][19] = (mid_1[3823:3816] < btm_0[3831:3824]) ? 1 : 0;
assign detect_min[476][20] = (mid_1[3823:3816] < btm_1[3815:3808]) ? 1 : 0;
assign detect_min[476][21] = (mid_1[3823:3816] < btm_1[3823:3816]) ? 1 : 0;
assign detect_min[476][22] = (mid_1[3823:3816] < btm_1[3831:3824]) ? 1 : 0;
assign detect_min[476][23] = (mid_1[3823:3816] < btm_2[3815:3808]) ? 1 : 0;
assign detect_min[476][24] = (mid_1[3823:3816] < btm_2[3823:3816]) ? 1 : 0;
assign detect_min[476][25] = (mid_1[3823:3816] < btm_2[3831:3824]) ? 1 : 0;

assign detect_min[477][0] = (mid_1[3831:3824] < top_0[3823:3816]) ? 1 : 0;
assign detect_min[477][1] = (mid_1[3831:3824] < top_0[3831:3824]) ? 1 : 0;
assign detect_min[477][2] = (mid_1[3831:3824] < top_0[3839:3832]) ? 1 : 0;
assign detect_min[477][3] = (mid_1[3831:3824] < top_1[3823:3816]) ? 1 : 0;
assign detect_min[477][4] = (mid_1[3831:3824] < top_1[3831:3824]) ? 1 : 0;
assign detect_min[477][5] = (mid_1[3831:3824] < top_1[3839:3832]) ? 1 : 0;
assign detect_min[477][6] = (mid_1[3831:3824] < top_2[3823:3816]) ? 1 : 0;
assign detect_min[477][7] = (mid_1[3831:3824] < top_2[3831:3824]) ? 1 : 0;
assign detect_min[477][8] = (mid_1[3831:3824] < top_2[3839:3832]) ? 1 : 0;
assign detect_min[477][9] = (mid_1[3831:3824] < mid_0[3823:3816]) ? 1 : 0;
assign detect_min[477][10] = (mid_1[3831:3824] < mid_0[3831:3824]) ? 1 : 0;
assign detect_min[477][11] = (mid_1[3831:3824] < mid_0[3839:3832]) ? 1 : 0;
assign detect_min[477][12] = (mid_1[3831:3824] < mid_1[3823:3816]) ? 1 : 0;
assign detect_min[477][13] = (mid_1[3831:3824] < mid_1[3839:3832]) ? 1 : 0;
assign detect_min[477][14] = (mid_1[3831:3824] < mid_2[3823:3816]) ? 1 : 0;
assign detect_min[477][15] = (mid_1[3831:3824] < mid_2[3831:3824]) ? 1 : 0;
assign detect_min[477][16] = (mid_1[3831:3824] < mid_2[3839:3832]) ? 1 : 0;
assign detect_min[477][17] = (mid_1[3831:3824] < btm_0[3823:3816]) ? 1 : 0;
assign detect_min[477][18] = (mid_1[3831:3824] < btm_0[3831:3824]) ? 1 : 0;
assign detect_min[477][19] = (mid_1[3831:3824] < btm_0[3839:3832]) ? 1 : 0;
assign detect_min[477][20] = (mid_1[3831:3824] < btm_1[3823:3816]) ? 1 : 0;
assign detect_min[477][21] = (mid_1[3831:3824] < btm_1[3831:3824]) ? 1 : 0;
assign detect_min[477][22] = (mid_1[3831:3824] < btm_1[3839:3832]) ? 1 : 0;
assign detect_min[477][23] = (mid_1[3831:3824] < btm_2[3823:3816]) ? 1 : 0;
assign detect_min[477][24] = (mid_1[3831:3824] < btm_2[3831:3824]) ? 1 : 0;
assign detect_min[477][25] = (mid_1[3831:3824] < btm_2[3839:3832]) ? 1 : 0;

assign detect_min[478][0] = (mid_1[3839:3832] < top_0[3831:3824]) ? 1 : 0;
assign detect_min[478][1] = (mid_1[3839:3832] < top_0[3839:3832]) ? 1 : 0;
assign detect_min[478][2] = (mid_1[3839:3832] < top_0[3847:3840]) ? 1 : 0;
assign detect_min[478][3] = (mid_1[3839:3832] < top_1[3831:3824]) ? 1 : 0;
assign detect_min[478][4] = (mid_1[3839:3832] < top_1[3839:3832]) ? 1 : 0;
assign detect_min[478][5] = (mid_1[3839:3832] < top_1[3847:3840]) ? 1 : 0;
assign detect_min[478][6] = (mid_1[3839:3832] < top_2[3831:3824]) ? 1 : 0;
assign detect_min[478][7] = (mid_1[3839:3832] < top_2[3839:3832]) ? 1 : 0;
assign detect_min[478][8] = (mid_1[3839:3832] < top_2[3847:3840]) ? 1 : 0;
assign detect_min[478][9] = (mid_1[3839:3832] < mid_0[3831:3824]) ? 1 : 0;
assign detect_min[478][10] = (mid_1[3839:3832] < mid_0[3839:3832]) ? 1 : 0;
assign detect_min[478][11] = (mid_1[3839:3832] < mid_0[3847:3840]) ? 1 : 0;
assign detect_min[478][12] = (mid_1[3839:3832] < mid_1[3831:3824]) ? 1 : 0;
assign detect_min[478][13] = (mid_1[3839:3832] < mid_1[3847:3840]) ? 1 : 0;
assign detect_min[478][14] = (mid_1[3839:3832] < mid_2[3831:3824]) ? 1 : 0;
assign detect_min[478][15] = (mid_1[3839:3832] < mid_2[3839:3832]) ? 1 : 0;
assign detect_min[478][16] = (mid_1[3839:3832] < mid_2[3847:3840]) ? 1 : 0;
assign detect_min[478][17] = (mid_1[3839:3832] < btm_0[3831:3824]) ? 1 : 0;
assign detect_min[478][18] = (mid_1[3839:3832] < btm_0[3839:3832]) ? 1 : 0;
assign detect_min[478][19] = (mid_1[3839:3832] < btm_0[3847:3840]) ? 1 : 0;
assign detect_min[478][20] = (mid_1[3839:3832] < btm_1[3831:3824]) ? 1 : 0;
assign detect_min[478][21] = (mid_1[3839:3832] < btm_1[3839:3832]) ? 1 : 0;
assign detect_min[478][22] = (mid_1[3839:3832] < btm_1[3847:3840]) ? 1 : 0;
assign detect_min[478][23] = (mid_1[3839:3832] < btm_2[3831:3824]) ? 1 : 0;
assign detect_min[478][24] = (mid_1[3839:3832] < btm_2[3839:3832]) ? 1 : 0;
assign detect_min[478][25] = (mid_1[3839:3832] < btm_2[3847:3840]) ? 1 : 0;

assign detect_min[479][0] = (mid_1[3847:3840] < top_0[3839:3832]) ? 1 : 0;
assign detect_min[479][1] = (mid_1[3847:3840] < top_0[3847:3840]) ? 1 : 0;
assign detect_min[479][2] = (mid_1[3847:3840] < top_0[3855:3848]) ? 1 : 0;
assign detect_min[479][3] = (mid_1[3847:3840] < top_1[3839:3832]) ? 1 : 0;
assign detect_min[479][4] = (mid_1[3847:3840] < top_1[3847:3840]) ? 1 : 0;
assign detect_min[479][5] = (mid_1[3847:3840] < top_1[3855:3848]) ? 1 : 0;
assign detect_min[479][6] = (mid_1[3847:3840] < top_2[3839:3832]) ? 1 : 0;
assign detect_min[479][7] = (mid_1[3847:3840] < top_2[3847:3840]) ? 1 : 0;
assign detect_min[479][8] = (mid_1[3847:3840] < top_2[3855:3848]) ? 1 : 0;
assign detect_min[479][9] = (mid_1[3847:3840] < mid_0[3839:3832]) ? 1 : 0;
assign detect_min[479][10] = (mid_1[3847:3840] < mid_0[3847:3840]) ? 1 : 0;
assign detect_min[479][11] = (mid_1[3847:3840] < mid_0[3855:3848]) ? 1 : 0;
assign detect_min[479][12] = (mid_1[3847:3840] < mid_1[3839:3832]) ? 1 : 0;
assign detect_min[479][13] = (mid_1[3847:3840] < mid_1[3855:3848]) ? 1 : 0;
assign detect_min[479][14] = (mid_1[3847:3840] < mid_2[3839:3832]) ? 1 : 0;
assign detect_min[479][15] = (mid_1[3847:3840] < mid_2[3847:3840]) ? 1 : 0;
assign detect_min[479][16] = (mid_1[3847:3840] < mid_2[3855:3848]) ? 1 : 0;
assign detect_min[479][17] = (mid_1[3847:3840] < btm_0[3839:3832]) ? 1 : 0;
assign detect_min[479][18] = (mid_1[3847:3840] < btm_0[3847:3840]) ? 1 : 0;
assign detect_min[479][19] = (mid_1[3847:3840] < btm_0[3855:3848]) ? 1 : 0;
assign detect_min[479][20] = (mid_1[3847:3840] < btm_1[3839:3832]) ? 1 : 0;
assign detect_min[479][21] = (mid_1[3847:3840] < btm_1[3847:3840]) ? 1 : 0;
assign detect_min[479][22] = (mid_1[3847:3840] < btm_1[3855:3848]) ? 1 : 0;
assign detect_min[479][23] = (mid_1[3847:3840] < btm_2[3839:3832]) ? 1 : 0;
assign detect_min[479][24] = (mid_1[3847:3840] < btm_2[3847:3840]) ? 1 : 0;
assign detect_min[479][25] = (mid_1[3847:3840] < btm_2[3855:3848]) ? 1 : 0;

assign detect_min[480][0] = (mid_1[3855:3848] < top_0[3847:3840]) ? 1 : 0;
assign detect_min[480][1] = (mid_1[3855:3848] < top_0[3855:3848]) ? 1 : 0;
assign detect_min[480][2] = (mid_1[3855:3848] < top_0[3863:3856]) ? 1 : 0;
assign detect_min[480][3] = (mid_1[3855:3848] < top_1[3847:3840]) ? 1 : 0;
assign detect_min[480][4] = (mid_1[3855:3848] < top_1[3855:3848]) ? 1 : 0;
assign detect_min[480][5] = (mid_1[3855:3848] < top_1[3863:3856]) ? 1 : 0;
assign detect_min[480][6] = (mid_1[3855:3848] < top_2[3847:3840]) ? 1 : 0;
assign detect_min[480][7] = (mid_1[3855:3848] < top_2[3855:3848]) ? 1 : 0;
assign detect_min[480][8] = (mid_1[3855:3848] < top_2[3863:3856]) ? 1 : 0;
assign detect_min[480][9] = (mid_1[3855:3848] < mid_0[3847:3840]) ? 1 : 0;
assign detect_min[480][10] = (mid_1[3855:3848] < mid_0[3855:3848]) ? 1 : 0;
assign detect_min[480][11] = (mid_1[3855:3848] < mid_0[3863:3856]) ? 1 : 0;
assign detect_min[480][12] = (mid_1[3855:3848] < mid_1[3847:3840]) ? 1 : 0;
assign detect_min[480][13] = (mid_1[3855:3848] < mid_1[3863:3856]) ? 1 : 0;
assign detect_min[480][14] = (mid_1[3855:3848] < mid_2[3847:3840]) ? 1 : 0;
assign detect_min[480][15] = (mid_1[3855:3848] < mid_2[3855:3848]) ? 1 : 0;
assign detect_min[480][16] = (mid_1[3855:3848] < mid_2[3863:3856]) ? 1 : 0;
assign detect_min[480][17] = (mid_1[3855:3848] < btm_0[3847:3840]) ? 1 : 0;
assign detect_min[480][18] = (mid_1[3855:3848] < btm_0[3855:3848]) ? 1 : 0;
assign detect_min[480][19] = (mid_1[3855:3848] < btm_0[3863:3856]) ? 1 : 0;
assign detect_min[480][20] = (mid_1[3855:3848] < btm_1[3847:3840]) ? 1 : 0;
assign detect_min[480][21] = (mid_1[3855:3848] < btm_1[3855:3848]) ? 1 : 0;
assign detect_min[480][22] = (mid_1[3855:3848] < btm_1[3863:3856]) ? 1 : 0;
assign detect_min[480][23] = (mid_1[3855:3848] < btm_2[3847:3840]) ? 1 : 0;
assign detect_min[480][24] = (mid_1[3855:3848] < btm_2[3855:3848]) ? 1 : 0;
assign detect_min[480][25] = (mid_1[3855:3848] < btm_2[3863:3856]) ? 1 : 0;

assign detect_min[481][0] = (mid_1[3863:3856] < top_0[3855:3848]) ? 1 : 0;
assign detect_min[481][1] = (mid_1[3863:3856] < top_0[3863:3856]) ? 1 : 0;
assign detect_min[481][2] = (mid_1[3863:3856] < top_0[3871:3864]) ? 1 : 0;
assign detect_min[481][3] = (mid_1[3863:3856] < top_1[3855:3848]) ? 1 : 0;
assign detect_min[481][4] = (mid_1[3863:3856] < top_1[3863:3856]) ? 1 : 0;
assign detect_min[481][5] = (mid_1[3863:3856] < top_1[3871:3864]) ? 1 : 0;
assign detect_min[481][6] = (mid_1[3863:3856] < top_2[3855:3848]) ? 1 : 0;
assign detect_min[481][7] = (mid_1[3863:3856] < top_2[3863:3856]) ? 1 : 0;
assign detect_min[481][8] = (mid_1[3863:3856] < top_2[3871:3864]) ? 1 : 0;
assign detect_min[481][9] = (mid_1[3863:3856] < mid_0[3855:3848]) ? 1 : 0;
assign detect_min[481][10] = (mid_1[3863:3856] < mid_0[3863:3856]) ? 1 : 0;
assign detect_min[481][11] = (mid_1[3863:3856] < mid_0[3871:3864]) ? 1 : 0;
assign detect_min[481][12] = (mid_1[3863:3856] < mid_1[3855:3848]) ? 1 : 0;
assign detect_min[481][13] = (mid_1[3863:3856] < mid_1[3871:3864]) ? 1 : 0;
assign detect_min[481][14] = (mid_1[3863:3856] < mid_2[3855:3848]) ? 1 : 0;
assign detect_min[481][15] = (mid_1[3863:3856] < mid_2[3863:3856]) ? 1 : 0;
assign detect_min[481][16] = (mid_1[3863:3856] < mid_2[3871:3864]) ? 1 : 0;
assign detect_min[481][17] = (mid_1[3863:3856] < btm_0[3855:3848]) ? 1 : 0;
assign detect_min[481][18] = (mid_1[3863:3856] < btm_0[3863:3856]) ? 1 : 0;
assign detect_min[481][19] = (mid_1[3863:3856] < btm_0[3871:3864]) ? 1 : 0;
assign detect_min[481][20] = (mid_1[3863:3856] < btm_1[3855:3848]) ? 1 : 0;
assign detect_min[481][21] = (mid_1[3863:3856] < btm_1[3863:3856]) ? 1 : 0;
assign detect_min[481][22] = (mid_1[3863:3856] < btm_1[3871:3864]) ? 1 : 0;
assign detect_min[481][23] = (mid_1[3863:3856] < btm_2[3855:3848]) ? 1 : 0;
assign detect_min[481][24] = (mid_1[3863:3856] < btm_2[3863:3856]) ? 1 : 0;
assign detect_min[481][25] = (mid_1[3863:3856] < btm_2[3871:3864]) ? 1 : 0;

assign detect_min[482][0] = (mid_1[3871:3864] < top_0[3863:3856]) ? 1 : 0;
assign detect_min[482][1] = (mid_1[3871:3864] < top_0[3871:3864]) ? 1 : 0;
assign detect_min[482][2] = (mid_1[3871:3864] < top_0[3879:3872]) ? 1 : 0;
assign detect_min[482][3] = (mid_1[3871:3864] < top_1[3863:3856]) ? 1 : 0;
assign detect_min[482][4] = (mid_1[3871:3864] < top_1[3871:3864]) ? 1 : 0;
assign detect_min[482][5] = (mid_1[3871:3864] < top_1[3879:3872]) ? 1 : 0;
assign detect_min[482][6] = (mid_1[3871:3864] < top_2[3863:3856]) ? 1 : 0;
assign detect_min[482][7] = (mid_1[3871:3864] < top_2[3871:3864]) ? 1 : 0;
assign detect_min[482][8] = (mid_1[3871:3864] < top_2[3879:3872]) ? 1 : 0;
assign detect_min[482][9] = (mid_1[3871:3864] < mid_0[3863:3856]) ? 1 : 0;
assign detect_min[482][10] = (mid_1[3871:3864] < mid_0[3871:3864]) ? 1 : 0;
assign detect_min[482][11] = (mid_1[3871:3864] < mid_0[3879:3872]) ? 1 : 0;
assign detect_min[482][12] = (mid_1[3871:3864] < mid_1[3863:3856]) ? 1 : 0;
assign detect_min[482][13] = (mid_1[3871:3864] < mid_1[3879:3872]) ? 1 : 0;
assign detect_min[482][14] = (mid_1[3871:3864] < mid_2[3863:3856]) ? 1 : 0;
assign detect_min[482][15] = (mid_1[3871:3864] < mid_2[3871:3864]) ? 1 : 0;
assign detect_min[482][16] = (mid_1[3871:3864] < mid_2[3879:3872]) ? 1 : 0;
assign detect_min[482][17] = (mid_1[3871:3864] < btm_0[3863:3856]) ? 1 : 0;
assign detect_min[482][18] = (mid_1[3871:3864] < btm_0[3871:3864]) ? 1 : 0;
assign detect_min[482][19] = (mid_1[3871:3864] < btm_0[3879:3872]) ? 1 : 0;
assign detect_min[482][20] = (mid_1[3871:3864] < btm_1[3863:3856]) ? 1 : 0;
assign detect_min[482][21] = (mid_1[3871:3864] < btm_1[3871:3864]) ? 1 : 0;
assign detect_min[482][22] = (mid_1[3871:3864] < btm_1[3879:3872]) ? 1 : 0;
assign detect_min[482][23] = (mid_1[3871:3864] < btm_2[3863:3856]) ? 1 : 0;
assign detect_min[482][24] = (mid_1[3871:3864] < btm_2[3871:3864]) ? 1 : 0;
assign detect_min[482][25] = (mid_1[3871:3864] < btm_2[3879:3872]) ? 1 : 0;

assign detect_min[483][0] = (mid_1[3879:3872] < top_0[3871:3864]) ? 1 : 0;
assign detect_min[483][1] = (mid_1[3879:3872] < top_0[3879:3872]) ? 1 : 0;
assign detect_min[483][2] = (mid_1[3879:3872] < top_0[3887:3880]) ? 1 : 0;
assign detect_min[483][3] = (mid_1[3879:3872] < top_1[3871:3864]) ? 1 : 0;
assign detect_min[483][4] = (mid_1[3879:3872] < top_1[3879:3872]) ? 1 : 0;
assign detect_min[483][5] = (mid_1[3879:3872] < top_1[3887:3880]) ? 1 : 0;
assign detect_min[483][6] = (mid_1[3879:3872] < top_2[3871:3864]) ? 1 : 0;
assign detect_min[483][7] = (mid_1[3879:3872] < top_2[3879:3872]) ? 1 : 0;
assign detect_min[483][8] = (mid_1[3879:3872] < top_2[3887:3880]) ? 1 : 0;
assign detect_min[483][9] = (mid_1[3879:3872] < mid_0[3871:3864]) ? 1 : 0;
assign detect_min[483][10] = (mid_1[3879:3872] < mid_0[3879:3872]) ? 1 : 0;
assign detect_min[483][11] = (mid_1[3879:3872] < mid_0[3887:3880]) ? 1 : 0;
assign detect_min[483][12] = (mid_1[3879:3872] < mid_1[3871:3864]) ? 1 : 0;
assign detect_min[483][13] = (mid_1[3879:3872] < mid_1[3887:3880]) ? 1 : 0;
assign detect_min[483][14] = (mid_1[3879:3872] < mid_2[3871:3864]) ? 1 : 0;
assign detect_min[483][15] = (mid_1[3879:3872] < mid_2[3879:3872]) ? 1 : 0;
assign detect_min[483][16] = (mid_1[3879:3872] < mid_2[3887:3880]) ? 1 : 0;
assign detect_min[483][17] = (mid_1[3879:3872] < btm_0[3871:3864]) ? 1 : 0;
assign detect_min[483][18] = (mid_1[3879:3872] < btm_0[3879:3872]) ? 1 : 0;
assign detect_min[483][19] = (mid_1[3879:3872] < btm_0[3887:3880]) ? 1 : 0;
assign detect_min[483][20] = (mid_1[3879:3872] < btm_1[3871:3864]) ? 1 : 0;
assign detect_min[483][21] = (mid_1[3879:3872] < btm_1[3879:3872]) ? 1 : 0;
assign detect_min[483][22] = (mid_1[3879:3872] < btm_1[3887:3880]) ? 1 : 0;
assign detect_min[483][23] = (mid_1[3879:3872] < btm_2[3871:3864]) ? 1 : 0;
assign detect_min[483][24] = (mid_1[3879:3872] < btm_2[3879:3872]) ? 1 : 0;
assign detect_min[483][25] = (mid_1[3879:3872] < btm_2[3887:3880]) ? 1 : 0;

assign detect_min[484][0] = (mid_1[3887:3880] < top_0[3879:3872]) ? 1 : 0;
assign detect_min[484][1] = (mid_1[3887:3880] < top_0[3887:3880]) ? 1 : 0;
assign detect_min[484][2] = (mid_1[3887:3880] < top_0[3895:3888]) ? 1 : 0;
assign detect_min[484][3] = (mid_1[3887:3880] < top_1[3879:3872]) ? 1 : 0;
assign detect_min[484][4] = (mid_1[3887:3880] < top_1[3887:3880]) ? 1 : 0;
assign detect_min[484][5] = (mid_1[3887:3880] < top_1[3895:3888]) ? 1 : 0;
assign detect_min[484][6] = (mid_1[3887:3880] < top_2[3879:3872]) ? 1 : 0;
assign detect_min[484][7] = (mid_1[3887:3880] < top_2[3887:3880]) ? 1 : 0;
assign detect_min[484][8] = (mid_1[3887:3880] < top_2[3895:3888]) ? 1 : 0;
assign detect_min[484][9] = (mid_1[3887:3880] < mid_0[3879:3872]) ? 1 : 0;
assign detect_min[484][10] = (mid_1[3887:3880] < mid_0[3887:3880]) ? 1 : 0;
assign detect_min[484][11] = (mid_1[3887:3880] < mid_0[3895:3888]) ? 1 : 0;
assign detect_min[484][12] = (mid_1[3887:3880] < mid_1[3879:3872]) ? 1 : 0;
assign detect_min[484][13] = (mid_1[3887:3880] < mid_1[3895:3888]) ? 1 : 0;
assign detect_min[484][14] = (mid_1[3887:3880] < mid_2[3879:3872]) ? 1 : 0;
assign detect_min[484][15] = (mid_1[3887:3880] < mid_2[3887:3880]) ? 1 : 0;
assign detect_min[484][16] = (mid_1[3887:3880] < mid_2[3895:3888]) ? 1 : 0;
assign detect_min[484][17] = (mid_1[3887:3880] < btm_0[3879:3872]) ? 1 : 0;
assign detect_min[484][18] = (mid_1[3887:3880] < btm_0[3887:3880]) ? 1 : 0;
assign detect_min[484][19] = (mid_1[3887:3880] < btm_0[3895:3888]) ? 1 : 0;
assign detect_min[484][20] = (mid_1[3887:3880] < btm_1[3879:3872]) ? 1 : 0;
assign detect_min[484][21] = (mid_1[3887:3880] < btm_1[3887:3880]) ? 1 : 0;
assign detect_min[484][22] = (mid_1[3887:3880] < btm_1[3895:3888]) ? 1 : 0;
assign detect_min[484][23] = (mid_1[3887:3880] < btm_2[3879:3872]) ? 1 : 0;
assign detect_min[484][24] = (mid_1[3887:3880] < btm_2[3887:3880]) ? 1 : 0;
assign detect_min[484][25] = (mid_1[3887:3880] < btm_2[3895:3888]) ? 1 : 0;

assign detect_min[485][0] = (mid_1[3895:3888] < top_0[3887:3880]) ? 1 : 0;
assign detect_min[485][1] = (mid_1[3895:3888] < top_0[3895:3888]) ? 1 : 0;
assign detect_min[485][2] = (mid_1[3895:3888] < top_0[3903:3896]) ? 1 : 0;
assign detect_min[485][3] = (mid_1[3895:3888] < top_1[3887:3880]) ? 1 : 0;
assign detect_min[485][4] = (mid_1[3895:3888] < top_1[3895:3888]) ? 1 : 0;
assign detect_min[485][5] = (mid_1[3895:3888] < top_1[3903:3896]) ? 1 : 0;
assign detect_min[485][6] = (mid_1[3895:3888] < top_2[3887:3880]) ? 1 : 0;
assign detect_min[485][7] = (mid_1[3895:3888] < top_2[3895:3888]) ? 1 : 0;
assign detect_min[485][8] = (mid_1[3895:3888] < top_2[3903:3896]) ? 1 : 0;
assign detect_min[485][9] = (mid_1[3895:3888] < mid_0[3887:3880]) ? 1 : 0;
assign detect_min[485][10] = (mid_1[3895:3888] < mid_0[3895:3888]) ? 1 : 0;
assign detect_min[485][11] = (mid_1[3895:3888] < mid_0[3903:3896]) ? 1 : 0;
assign detect_min[485][12] = (mid_1[3895:3888] < mid_1[3887:3880]) ? 1 : 0;
assign detect_min[485][13] = (mid_1[3895:3888] < mid_1[3903:3896]) ? 1 : 0;
assign detect_min[485][14] = (mid_1[3895:3888] < mid_2[3887:3880]) ? 1 : 0;
assign detect_min[485][15] = (mid_1[3895:3888] < mid_2[3895:3888]) ? 1 : 0;
assign detect_min[485][16] = (mid_1[3895:3888] < mid_2[3903:3896]) ? 1 : 0;
assign detect_min[485][17] = (mid_1[3895:3888] < btm_0[3887:3880]) ? 1 : 0;
assign detect_min[485][18] = (mid_1[3895:3888] < btm_0[3895:3888]) ? 1 : 0;
assign detect_min[485][19] = (mid_1[3895:3888] < btm_0[3903:3896]) ? 1 : 0;
assign detect_min[485][20] = (mid_1[3895:3888] < btm_1[3887:3880]) ? 1 : 0;
assign detect_min[485][21] = (mid_1[3895:3888] < btm_1[3895:3888]) ? 1 : 0;
assign detect_min[485][22] = (mid_1[3895:3888] < btm_1[3903:3896]) ? 1 : 0;
assign detect_min[485][23] = (mid_1[3895:3888] < btm_2[3887:3880]) ? 1 : 0;
assign detect_min[485][24] = (mid_1[3895:3888] < btm_2[3895:3888]) ? 1 : 0;
assign detect_min[485][25] = (mid_1[3895:3888] < btm_2[3903:3896]) ? 1 : 0;

assign detect_min[486][0] = (mid_1[3903:3896] < top_0[3895:3888]) ? 1 : 0;
assign detect_min[486][1] = (mid_1[3903:3896] < top_0[3903:3896]) ? 1 : 0;
assign detect_min[486][2] = (mid_1[3903:3896] < top_0[3911:3904]) ? 1 : 0;
assign detect_min[486][3] = (mid_1[3903:3896] < top_1[3895:3888]) ? 1 : 0;
assign detect_min[486][4] = (mid_1[3903:3896] < top_1[3903:3896]) ? 1 : 0;
assign detect_min[486][5] = (mid_1[3903:3896] < top_1[3911:3904]) ? 1 : 0;
assign detect_min[486][6] = (mid_1[3903:3896] < top_2[3895:3888]) ? 1 : 0;
assign detect_min[486][7] = (mid_1[3903:3896] < top_2[3903:3896]) ? 1 : 0;
assign detect_min[486][8] = (mid_1[3903:3896] < top_2[3911:3904]) ? 1 : 0;
assign detect_min[486][9] = (mid_1[3903:3896] < mid_0[3895:3888]) ? 1 : 0;
assign detect_min[486][10] = (mid_1[3903:3896] < mid_0[3903:3896]) ? 1 : 0;
assign detect_min[486][11] = (mid_1[3903:3896] < mid_0[3911:3904]) ? 1 : 0;
assign detect_min[486][12] = (mid_1[3903:3896] < mid_1[3895:3888]) ? 1 : 0;
assign detect_min[486][13] = (mid_1[3903:3896] < mid_1[3911:3904]) ? 1 : 0;
assign detect_min[486][14] = (mid_1[3903:3896] < mid_2[3895:3888]) ? 1 : 0;
assign detect_min[486][15] = (mid_1[3903:3896] < mid_2[3903:3896]) ? 1 : 0;
assign detect_min[486][16] = (mid_1[3903:3896] < mid_2[3911:3904]) ? 1 : 0;
assign detect_min[486][17] = (mid_1[3903:3896] < btm_0[3895:3888]) ? 1 : 0;
assign detect_min[486][18] = (mid_1[3903:3896] < btm_0[3903:3896]) ? 1 : 0;
assign detect_min[486][19] = (mid_1[3903:3896] < btm_0[3911:3904]) ? 1 : 0;
assign detect_min[486][20] = (mid_1[3903:3896] < btm_1[3895:3888]) ? 1 : 0;
assign detect_min[486][21] = (mid_1[3903:3896] < btm_1[3903:3896]) ? 1 : 0;
assign detect_min[486][22] = (mid_1[3903:3896] < btm_1[3911:3904]) ? 1 : 0;
assign detect_min[486][23] = (mid_1[3903:3896] < btm_2[3895:3888]) ? 1 : 0;
assign detect_min[486][24] = (mid_1[3903:3896] < btm_2[3903:3896]) ? 1 : 0;
assign detect_min[486][25] = (mid_1[3903:3896] < btm_2[3911:3904]) ? 1 : 0;

assign detect_min[487][0] = (mid_1[3911:3904] < top_0[3903:3896]) ? 1 : 0;
assign detect_min[487][1] = (mid_1[3911:3904] < top_0[3911:3904]) ? 1 : 0;
assign detect_min[487][2] = (mid_1[3911:3904] < top_0[3919:3912]) ? 1 : 0;
assign detect_min[487][3] = (mid_1[3911:3904] < top_1[3903:3896]) ? 1 : 0;
assign detect_min[487][4] = (mid_1[3911:3904] < top_1[3911:3904]) ? 1 : 0;
assign detect_min[487][5] = (mid_1[3911:3904] < top_1[3919:3912]) ? 1 : 0;
assign detect_min[487][6] = (mid_1[3911:3904] < top_2[3903:3896]) ? 1 : 0;
assign detect_min[487][7] = (mid_1[3911:3904] < top_2[3911:3904]) ? 1 : 0;
assign detect_min[487][8] = (mid_1[3911:3904] < top_2[3919:3912]) ? 1 : 0;
assign detect_min[487][9] = (mid_1[3911:3904] < mid_0[3903:3896]) ? 1 : 0;
assign detect_min[487][10] = (mid_1[3911:3904] < mid_0[3911:3904]) ? 1 : 0;
assign detect_min[487][11] = (mid_1[3911:3904] < mid_0[3919:3912]) ? 1 : 0;
assign detect_min[487][12] = (mid_1[3911:3904] < mid_1[3903:3896]) ? 1 : 0;
assign detect_min[487][13] = (mid_1[3911:3904] < mid_1[3919:3912]) ? 1 : 0;
assign detect_min[487][14] = (mid_1[3911:3904] < mid_2[3903:3896]) ? 1 : 0;
assign detect_min[487][15] = (mid_1[3911:3904] < mid_2[3911:3904]) ? 1 : 0;
assign detect_min[487][16] = (mid_1[3911:3904] < mid_2[3919:3912]) ? 1 : 0;
assign detect_min[487][17] = (mid_1[3911:3904] < btm_0[3903:3896]) ? 1 : 0;
assign detect_min[487][18] = (mid_1[3911:3904] < btm_0[3911:3904]) ? 1 : 0;
assign detect_min[487][19] = (mid_1[3911:3904] < btm_0[3919:3912]) ? 1 : 0;
assign detect_min[487][20] = (mid_1[3911:3904] < btm_1[3903:3896]) ? 1 : 0;
assign detect_min[487][21] = (mid_1[3911:3904] < btm_1[3911:3904]) ? 1 : 0;
assign detect_min[487][22] = (mid_1[3911:3904] < btm_1[3919:3912]) ? 1 : 0;
assign detect_min[487][23] = (mid_1[3911:3904] < btm_2[3903:3896]) ? 1 : 0;
assign detect_min[487][24] = (mid_1[3911:3904] < btm_2[3911:3904]) ? 1 : 0;
assign detect_min[487][25] = (mid_1[3911:3904] < btm_2[3919:3912]) ? 1 : 0;

assign detect_min[488][0] = (mid_1[3919:3912] < top_0[3911:3904]) ? 1 : 0;
assign detect_min[488][1] = (mid_1[3919:3912] < top_0[3919:3912]) ? 1 : 0;
assign detect_min[488][2] = (mid_1[3919:3912] < top_0[3927:3920]) ? 1 : 0;
assign detect_min[488][3] = (mid_1[3919:3912] < top_1[3911:3904]) ? 1 : 0;
assign detect_min[488][4] = (mid_1[3919:3912] < top_1[3919:3912]) ? 1 : 0;
assign detect_min[488][5] = (mid_1[3919:3912] < top_1[3927:3920]) ? 1 : 0;
assign detect_min[488][6] = (mid_1[3919:3912] < top_2[3911:3904]) ? 1 : 0;
assign detect_min[488][7] = (mid_1[3919:3912] < top_2[3919:3912]) ? 1 : 0;
assign detect_min[488][8] = (mid_1[3919:3912] < top_2[3927:3920]) ? 1 : 0;
assign detect_min[488][9] = (mid_1[3919:3912] < mid_0[3911:3904]) ? 1 : 0;
assign detect_min[488][10] = (mid_1[3919:3912] < mid_0[3919:3912]) ? 1 : 0;
assign detect_min[488][11] = (mid_1[3919:3912] < mid_0[3927:3920]) ? 1 : 0;
assign detect_min[488][12] = (mid_1[3919:3912] < mid_1[3911:3904]) ? 1 : 0;
assign detect_min[488][13] = (mid_1[3919:3912] < mid_1[3927:3920]) ? 1 : 0;
assign detect_min[488][14] = (mid_1[3919:3912] < mid_2[3911:3904]) ? 1 : 0;
assign detect_min[488][15] = (mid_1[3919:3912] < mid_2[3919:3912]) ? 1 : 0;
assign detect_min[488][16] = (mid_1[3919:3912] < mid_2[3927:3920]) ? 1 : 0;
assign detect_min[488][17] = (mid_1[3919:3912] < btm_0[3911:3904]) ? 1 : 0;
assign detect_min[488][18] = (mid_1[3919:3912] < btm_0[3919:3912]) ? 1 : 0;
assign detect_min[488][19] = (mid_1[3919:3912] < btm_0[3927:3920]) ? 1 : 0;
assign detect_min[488][20] = (mid_1[3919:3912] < btm_1[3911:3904]) ? 1 : 0;
assign detect_min[488][21] = (mid_1[3919:3912] < btm_1[3919:3912]) ? 1 : 0;
assign detect_min[488][22] = (mid_1[3919:3912] < btm_1[3927:3920]) ? 1 : 0;
assign detect_min[488][23] = (mid_1[3919:3912] < btm_2[3911:3904]) ? 1 : 0;
assign detect_min[488][24] = (mid_1[3919:3912] < btm_2[3919:3912]) ? 1 : 0;
assign detect_min[488][25] = (mid_1[3919:3912] < btm_2[3927:3920]) ? 1 : 0;

assign detect_min[489][0] = (mid_1[3927:3920] < top_0[3919:3912]) ? 1 : 0;
assign detect_min[489][1] = (mid_1[3927:3920] < top_0[3927:3920]) ? 1 : 0;
assign detect_min[489][2] = (mid_1[3927:3920] < top_0[3935:3928]) ? 1 : 0;
assign detect_min[489][3] = (mid_1[3927:3920] < top_1[3919:3912]) ? 1 : 0;
assign detect_min[489][4] = (mid_1[3927:3920] < top_1[3927:3920]) ? 1 : 0;
assign detect_min[489][5] = (mid_1[3927:3920] < top_1[3935:3928]) ? 1 : 0;
assign detect_min[489][6] = (mid_1[3927:3920] < top_2[3919:3912]) ? 1 : 0;
assign detect_min[489][7] = (mid_1[3927:3920] < top_2[3927:3920]) ? 1 : 0;
assign detect_min[489][8] = (mid_1[3927:3920] < top_2[3935:3928]) ? 1 : 0;
assign detect_min[489][9] = (mid_1[3927:3920] < mid_0[3919:3912]) ? 1 : 0;
assign detect_min[489][10] = (mid_1[3927:3920] < mid_0[3927:3920]) ? 1 : 0;
assign detect_min[489][11] = (mid_1[3927:3920] < mid_0[3935:3928]) ? 1 : 0;
assign detect_min[489][12] = (mid_1[3927:3920] < mid_1[3919:3912]) ? 1 : 0;
assign detect_min[489][13] = (mid_1[3927:3920] < mid_1[3935:3928]) ? 1 : 0;
assign detect_min[489][14] = (mid_1[3927:3920] < mid_2[3919:3912]) ? 1 : 0;
assign detect_min[489][15] = (mid_1[3927:3920] < mid_2[3927:3920]) ? 1 : 0;
assign detect_min[489][16] = (mid_1[3927:3920] < mid_2[3935:3928]) ? 1 : 0;
assign detect_min[489][17] = (mid_1[3927:3920] < btm_0[3919:3912]) ? 1 : 0;
assign detect_min[489][18] = (mid_1[3927:3920] < btm_0[3927:3920]) ? 1 : 0;
assign detect_min[489][19] = (mid_1[3927:3920] < btm_0[3935:3928]) ? 1 : 0;
assign detect_min[489][20] = (mid_1[3927:3920] < btm_1[3919:3912]) ? 1 : 0;
assign detect_min[489][21] = (mid_1[3927:3920] < btm_1[3927:3920]) ? 1 : 0;
assign detect_min[489][22] = (mid_1[3927:3920] < btm_1[3935:3928]) ? 1 : 0;
assign detect_min[489][23] = (mid_1[3927:3920] < btm_2[3919:3912]) ? 1 : 0;
assign detect_min[489][24] = (mid_1[3927:3920] < btm_2[3927:3920]) ? 1 : 0;
assign detect_min[489][25] = (mid_1[3927:3920] < btm_2[3935:3928]) ? 1 : 0;

assign detect_min[490][0] = (mid_1[3935:3928] < top_0[3927:3920]) ? 1 : 0;
assign detect_min[490][1] = (mid_1[3935:3928] < top_0[3935:3928]) ? 1 : 0;
assign detect_min[490][2] = (mid_1[3935:3928] < top_0[3943:3936]) ? 1 : 0;
assign detect_min[490][3] = (mid_1[3935:3928] < top_1[3927:3920]) ? 1 : 0;
assign detect_min[490][4] = (mid_1[3935:3928] < top_1[3935:3928]) ? 1 : 0;
assign detect_min[490][5] = (mid_1[3935:3928] < top_1[3943:3936]) ? 1 : 0;
assign detect_min[490][6] = (mid_1[3935:3928] < top_2[3927:3920]) ? 1 : 0;
assign detect_min[490][7] = (mid_1[3935:3928] < top_2[3935:3928]) ? 1 : 0;
assign detect_min[490][8] = (mid_1[3935:3928] < top_2[3943:3936]) ? 1 : 0;
assign detect_min[490][9] = (mid_1[3935:3928] < mid_0[3927:3920]) ? 1 : 0;
assign detect_min[490][10] = (mid_1[3935:3928] < mid_0[3935:3928]) ? 1 : 0;
assign detect_min[490][11] = (mid_1[3935:3928] < mid_0[3943:3936]) ? 1 : 0;
assign detect_min[490][12] = (mid_1[3935:3928] < mid_1[3927:3920]) ? 1 : 0;
assign detect_min[490][13] = (mid_1[3935:3928] < mid_1[3943:3936]) ? 1 : 0;
assign detect_min[490][14] = (mid_1[3935:3928] < mid_2[3927:3920]) ? 1 : 0;
assign detect_min[490][15] = (mid_1[3935:3928] < mid_2[3935:3928]) ? 1 : 0;
assign detect_min[490][16] = (mid_1[3935:3928] < mid_2[3943:3936]) ? 1 : 0;
assign detect_min[490][17] = (mid_1[3935:3928] < btm_0[3927:3920]) ? 1 : 0;
assign detect_min[490][18] = (mid_1[3935:3928] < btm_0[3935:3928]) ? 1 : 0;
assign detect_min[490][19] = (mid_1[3935:3928] < btm_0[3943:3936]) ? 1 : 0;
assign detect_min[490][20] = (mid_1[3935:3928] < btm_1[3927:3920]) ? 1 : 0;
assign detect_min[490][21] = (mid_1[3935:3928] < btm_1[3935:3928]) ? 1 : 0;
assign detect_min[490][22] = (mid_1[3935:3928] < btm_1[3943:3936]) ? 1 : 0;
assign detect_min[490][23] = (mid_1[3935:3928] < btm_2[3927:3920]) ? 1 : 0;
assign detect_min[490][24] = (mid_1[3935:3928] < btm_2[3935:3928]) ? 1 : 0;
assign detect_min[490][25] = (mid_1[3935:3928] < btm_2[3943:3936]) ? 1 : 0;

assign detect_min[491][0] = (mid_1[3943:3936] < top_0[3935:3928]) ? 1 : 0;
assign detect_min[491][1] = (mid_1[3943:3936] < top_0[3943:3936]) ? 1 : 0;
assign detect_min[491][2] = (mid_1[3943:3936] < top_0[3951:3944]) ? 1 : 0;
assign detect_min[491][3] = (mid_1[3943:3936] < top_1[3935:3928]) ? 1 : 0;
assign detect_min[491][4] = (mid_1[3943:3936] < top_1[3943:3936]) ? 1 : 0;
assign detect_min[491][5] = (mid_1[3943:3936] < top_1[3951:3944]) ? 1 : 0;
assign detect_min[491][6] = (mid_1[3943:3936] < top_2[3935:3928]) ? 1 : 0;
assign detect_min[491][7] = (mid_1[3943:3936] < top_2[3943:3936]) ? 1 : 0;
assign detect_min[491][8] = (mid_1[3943:3936] < top_2[3951:3944]) ? 1 : 0;
assign detect_min[491][9] = (mid_1[3943:3936] < mid_0[3935:3928]) ? 1 : 0;
assign detect_min[491][10] = (mid_1[3943:3936] < mid_0[3943:3936]) ? 1 : 0;
assign detect_min[491][11] = (mid_1[3943:3936] < mid_0[3951:3944]) ? 1 : 0;
assign detect_min[491][12] = (mid_1[3943:3936] < mid_1[3935:3928]) ? 1 : 0;
assign detect_min[491][13] = (mid_1[3943:3936] < mid_1[3951:3944]) ? 1 : 0;
assign detect_min[491][14] = (mid_1[3943:3936] < mid_2[3935:3928]) ? 1 : 0;
assign detect_min[491][15] = (mid_1[3943:3936] < mid_2[3943:3936]) ? 1 : 0;
assign detect_min[491][16] = (mid_1[3943:3936] < mid_2[3951:3944]) ? 1 : 0;
assign detect_min[491][17] = (mid_1[3943:3936] < btm_0[3935:3928]) ? 1 : 0;
assign detect_min[491][18] = (mid_1[3943:3936] < btm_0[3943:3936]) ? 1 : 0;
assign detect_min[491][19] = (mid_1[3943:3936] < btm_0[3951:3944]) ? 1 : 0;
assign detect_min[491][20] = (mid_1[3943:3936] < btm_1[3935:3928]) ? 1 : 0;
assign detect_min[491][21] = (mid_1[3943:3936] < btm_1[3943:3936]) ? 1 : 0;
assign detect_min[491][22] = (mid_1[3943:3936] < btm_1[3951:3944]) ? 1 : 0;
assign detect_min[491][23] = (mid_1[3943:3936] < btm_2[3935:3928]) ? 1 : 0;
assign detect_min[491][24] = (mid_1[3943:3936] < btm_2[3943:3936]) ? 1 : 0;
assign detect_min[491][25] = (mid_1[3943:3936] < btm_2[3951:3944]) ? 1 : 0;

assign detect_min[492][0] = (mid_1[3951:3944] < top_0[3943:3936]) ? 1 : 0;
assign detect_min[492][1] = (mid_1[3951:3944] < top_0[3951:3944]) ? 1 : 0;
assign detect_min[492][2] = (mid_1[3951:3944] < top_0[3959:3952]) ? 1 : 0;
assign detect_min[492][3] = (mid_1[3951:3944] < top_1[3943:3936]) ? 1 : 0;
assign detect_min[492][4] = (mid_1[3951:3944] < top_1[3951:3944]) ? 1 : 0;
assign detect_min[492][5] = (mid_1[3951:3944] < top_1[3959:3952]) ? 1 : 0;
assign detect_min[492][6] = (mid_1[3951:3944] < top_2[3943:3936]) ? 1 : 0;
assign detect_min[492][7] = (mid_1[3951:3944] < top_2[3951:3944]) ? 1 : 0;
assign detect_min[492][8] = (mid_1[3951:3944] < top_2[3959:3952]) ? 1 : 0;
assign detect_min[492][9] = (mid_1[3951:3944] < mid_0[3943:3936]) ? 1 : 0;
assign detect_min[492][10] = (mid_1[3951:3944] < mid_0[3951:3944]) ? 1 : 0;
assign detect_min[492][11] = (mid_1[3951:3944] < mid_0[3959:3952]) ? 1 : 0;
assign detect_min[492][12] = (mid_1[3951:3944] < mid_1[3943:3936]) ? 1 : 0;
assign detect_min[492][13] = (mid_1[3951:3944] < mid_1[3959:3952]) ? 1 : 0;
assign detect_min[492][14] = (mid_1[3951:3944] < mid_2[3943:3936]) ? 1 : 0;
assign detect_min[492][15] = (mid_1[3951:3944] < mid_2[3951:3944]) ? 1 : 0;
assign detect_min[492][16] = (mid_1[3951:3944] < mid_2[3959:3952]) ? 1 : 0;
assign detect_min[492][17] = (mid_1[3951:3944] < btm_0[3943:3936]) ? 1 : 0;
assign detect_min[492][18] = (mid_1[3951:3944] < btm_0[3951:3944]) ? 1 : 0;
assign detect_min[492][19] = (mid_1[3951:3944] < btm_0[3959:3952]) ? 1 : 0;
assign detect_min[492][20] = (mid_1[3951:3944] < btm_1[3943:3936]) ? 1 : 0;
assign detect_min[492][21] = (mid_1[3951:3944] < btm_1[3951:3944]) ? 1 : 0;
assign detect_min[492][22] = (mid_1[3951:3944] < btm_1[3959:3952]) ? 1 : 0;
assign detect_min[492][23] = (mid_1[3951:3944] < btm_2[3943:3936]) ? 1 : 0;
assign detect_min[492][24] = (mid_1[3951:3944] < btm_2[3951:3944]) ? 1 : 0;
assign detect_min[492][25] = (mid_1[3951:3944] < btm_2[3959:3952]) ? 1 : 0;

assign detect_min[493][0] = (mid_1[3959:3952] < top_0[3951:3944]) ? 1 : 0;
assign detect_min[493][1] = (mid_1[3959:3952] < top_0[3959:3952]) ? 1 : 0;
assign detect_min[493][2] = (mid_1[3959:3952] < top_0[3967:3960]) ? 1 : 0;
assign detect_min[493][3] = (mid_1[3959:3952] < top_1[3951:3944]) ? 1 : 0;
assign detect_min[493][4] = (mid_1[3959:3952] < top_1[3959:3952]) ? 1 : 0;
assign detect_min[493][5] = (mid_1[3959:3952] < top_1[3967:3960]) ? 1 : 0;
assign detect_min[493][6] = (mid_1[3959:3952] < top_2[3951:3944]) ? 1 : 0;
assign detect_min[493][7] = (mid_1[3959:3952] < top_2[3959:3952]) ? 1 : 0;
assign detect_min[493][8] = (mid_1[3959:3952] < top_2[3967:3960]) ? 1 : 0;
assign detect_min[493][9] = (mid_1[3959:3952] < mid_0[3951:3944]) ? 1 : 0;
assign detect_min[493][10] = (mid_1[3959:3952] < mid_0[3959:3952]) ? 1 : 0;
assign detect_min[493][11] = (mid_1[3959:3952] < mid_0[3967:3960]) ? 1 : 0;
assign detect_min[493][12] = (mid_1[3959:3952] < mid_1[3951:3944]) ? 1 : 0;
assign detect_min[493][13] = (mid_1[3959:3952] < mid_1[3967:3960]) ? 1 : 0;
assign detect_min[493][14] = (mid_1[3959:3952] < mid_2[3951:3944]) ? 1 : 0;
assign detect_min[493][15] = (mid_1[3959:3952] < mid_2[3959:3952]) ? 1 : 0;
assign detect_min[493][16] = (mid_1[3959:3952] < mid_2[3967:3960]) ? 1 : 0;
assign detect_min[493][17] = (mid_1[3959:3952] < btm_0[3951:3944]) ? 1 : 0;
assign detect_min[493][18] = (mid_1[3959:3952] < btm_0[3959:3952]) ? 1 : 0;
assign detect_min[493][19] = (mid_1[3959:3952] < btm_0[3967:3960]) ? 1 : 0;
assign detect_min[493][20] = (mid_1[3959:3952] < btm_1[3951:3944]) ? 1 : 0;
assign detect_min[493][21] = (mid_1[3959:3952] < btm_1[3959:3952]) ? 1 : 0;
assign detect_min[493][22] = (mid_1[3959:3952] < btm_1[3967:3960]) ? 1 : 0;
assign detect_min[493][23] = (mid_1[3959:3952] < btm_2[3951:3944]) ? 1 : 0;
assign detect_min[493][24] = (mid_1[3959:3952] < btm_2[3959:3952]) ? 1 : 0;
assign detect_min[493][25] = (mid_1[3959:3952] < btm_2[3967:3960]) ? 1 : 0;

assign detect_min[494][0] = (mid_1[3967:3960] < top_0[3959:3952]) ? 1 : 0;
assign detect_min[494][1] = (mid_1[3967:3960] < top_0[3967:3960]) ? 1 : 0;
assign detect_min[494][2] = (mid_1[3967:3960] < top_0[3975:3968]) ? 1 : 0;
assign detect_min[494][3] = (mid_1[3967:3960] < top_1[3959:3952]) ? 1 : 0;
assign detect_min[494][4] = (mid_1[3967:3960] < top_1[3967:3960]) ? 1 : 0;
assign detect_min[494][5] = (mid_1[3967:3960] < top_1[3975:3968]) ? 1 : 0;
assign detect_min[494][6] = (mid_1[3967:3960] < top_2[3959:3952]) ? 1 : 0;
assign detect_min[494][7] = (mid_1[3967:3960] < top_2[3967:3960]) ? 1 : 0;
assign detect_min[494][8] = (mid_1[3967:3960] < top_2[3975:3968]) ? 1 : 0;
assign detect_min[494][9] = (mid_1[3967:3960] < mid_0[3959:3952]) ? 1 : 0;
assign detect_min[494][10] = (mid_1[3967:3960] < mid_0[3967:3960]) ? 1 : 0;
assign detect_min[494][11] = (mid_1[3967:3960] < mid_0[3975:3968]) ? 1 : 0;
assign detect_min[494][12] = (mid_1[3967:3960] < mid_1[3959:3952]) ? 1 : 0;
assign detect_min[494][13] = (mid_1[3967:3960] < mid_1[3975:3968]) ? 1 : 0;
assign detect_min[494][14] = (mid_1[3967:3960] < mid_2[3959:3952]) ? 1 : 0;
assign detect_min[494][15] = (mid_1[3967:3960] < mid_2[3967:3960]) ? 1 : 0;
assign detect_min[494][16] = (mid_1[3967:3960] < mid_2[3975:3968]) ? 1 : 0;
assign detect_min[494][17] = (mid_1[3967:3960] < btm_0[3959:3952]) ? 1 : 0;
assign detect_min[494][18] = (mid_1[3967:3960] < btm_0[3967:3960]) ? 1 : 0;
assign detect_min[494][19] = (mid_1[3967:3960] < btm_0[3975:3968]) ? 1 : 0;
assign detect_min[494][20] = (mid_1[3967:3960] < btm_1[3959:3952]) ? 1 : 0;
assign detect_min[494][21] = (mid_1[3967:3960] < btm_1[3967:3960]) ? 1 : 0;
assign detect_min[494][22] = (mid_1[3967:3960] < btm_1[3975:3968]) ? 1 : 0;
assign detect_min[494][23] = (mid_1[3967:3960] < btm_2[3959:3952]) ? 1 : 0;
assign detect_min[494][24] = (mid_1[3967:3960] < btm_2[3967:3960]) ? 1 : 0;
assign detect_min[494][25] = (mid_1[3967:3960] < btm_2[3975:3968]) ? 1 : 0;

assign detect_min[495][0] = (mid_1[3975:3968] < top_0[3967:3960]) ? 1 : 0;
assign detect_min[495][1] = (mid_1[3975:3968] < top_0[3975:3968]) ? 1 : 0;
assign detect_min[495][2] = (mid_1[3975:3968] < top_0[3983:3976]) ? 1 : 0;
assign detect_min[495][3] = (mid_1[3975:3968] < top_1[3967:3960]) ? 1 : 0;
assign detect_min[495][4] = (mid_1[3975:3968] < top_1[3975:3968]) ? 1 : 0;
assign detect_min[495][5] = (mid_1[3975:3968] < top_1[3983:3976]) ? 1 : 0;
assign detect_min[495][6] = (mid_1[3975:3968] < top_2[3967:3960]) ? 1 : 0;
assign detect_min[495][7] = (mid_1[3975:3968] < top_2[3975:3968]) ? 1 : 0;
assign detect_min[495][8] = (mid_1[3975:3968] < top_2[3983:3976]) ? 1 : 0;
assign detect_min[495][9] = (mid_1[3975:3968] < mid_0[3967:3960]) ? 1 : 0;
assign detect_min[495][10] = (mid_1[3975:3968] < mid_0[3975:3968]) ? 1 : 0;
assign detect_min[495][11] = (mid_1[3975:3968] < mid_0[3983:3976]) ? 1 : 0;
assign detect_min[495][12] = (mid_1[3975:3968] < mid_1[3967:3960]) ? 1 : 0;
assign detect_min[495][13] = (mid_1[3975:3968] < mid_1[3983:3976]) ? 1 : 0;
assign detect_min[495][14] = (mid_1[3975:3968] < mid_2[3967:3960]) ? 1 : 0;
assign detect_min[495][15] = (mid_1[3975:3968] < mid_2[3975:3968]) ? 1 : 0;
assign detect_min[495][16] = (mid_1[3975:3968] < mid_2[3983:3976]) ? 1 : 0;
assign detect_min[495][17] = (mid_1[3975:3968] < btm_0[3967:3960]) ? 1 : 0;
assign detect_min[495][18] = (mid_1[3975:3968] < btm_0[3975:3968]) ? 1 : 0;
assign detect_min[495][19] = (mid_1[3975:3968] < btm_0[3983:3976]) ? 1 : 0;
assign detect_min[495][20] = (mid_1[3975:3968] < btm_1[3967:3960]) ? 1 : 0;
assign detect_min[495][21] = (mid_1[3975:3968] < btm_1[3975:3968]) ? 1 : 0;
assign detect_min[495][22] = (mid_1[3975:3968] < btm_1[3983:3976]) ? 1 : 0;
assign detect_min[495][23] = (mid_1[3975:3968] < btm_2[3967:3960]) ? 1 : 0;
assign detect_min[495][24] = (mid_1[3975:3968] < btm_2[3975:3968]) ? 1 : 0;
assign detect_min[495][25] = (mid_1[3975:3968] < btm_2[3983:3976]) ? 1 : 0;

assign detect_min[496][0] = (mid_1[3983:3976] < top_0[3975:3968]) ? 1 : 0;
assign detect_min[496][1] = (mid_1[3983:3976] < top_0[3983:3976]) ? 1 : 0;
assign detect_min[496][2] = (mid_1[3983:3976] < top_0[3991:3984]) ? 1 : 0;
assign detect_min[496][3] = (mid_1[3983:3976] < top_1[3975:3968]) ? 1 : 0;
assign detect_min[496][4] = (mid_1[3983:3976] < top_1[3983:3976]) ? 1 : 0;
assign detect_min[496][5] = (mid_1[3983:3976] < top_1[3991:3984]) ? 1 : 0;
assign detect_min[496][6] = (mid_1[3983:3976] < top_2[3975:3968]) ? 1 : 0;
assign detect_min[496][7] = (mid_1[3983:3976] < top_2[3983:3976]) ? 1 : 0;
assign detect_min[496][8] = (mid_1[3983:3976] < top_2[3991:3984]) ? 1 : 0;
assign detect_min[496][9] = (mid_1[3983:3976] < mid_0[3975:3968]) ? 1 : 0;
assign detect_min[496][10] = (mid_1[3983:3976] < mid_0[3983:3976]) ? 1 : 0;
assign detect_min[496][11] = (mid_1[3983:3976] < mid_0[3991:3984]) ? 1 : 0;
assign detect_min[496][12] = (mid_1[3983:3976] < mid_1[3975:3968]) ? 1 : 0;
assign detect_min[496][13] = (mid_1[3983:3976] < mid_1[3991:3984]) ? 1 : 0;
assign detect_min[496][14] = (mid_1[3983:3976] < mid_2[3975:3968]) ? 1 : 0;
assign detect_min[496][15] = (mid_1[3983:3976] < mid_2[3983:3976]) ? 1 : 0;
assign detect_min[496][16] = (mid_1[3983:3976] < mid_2[3991:3984]) ? 1 : 0;
assign detect_min[496][17] = (mid_1[3983:3976] < btm_0[3975:3968]) ? 1 : 0;
assign detect_min[496][18] = (mid_1[3983:3976] < btm_0[3983:3976]) ? 1 : 0;
assign detect_min[496][19] = (mid_1[3983:3976] < btm_0[3991:3984]) ? 1 : 0;
assign detect_min[496][20] = (mid_1[3983:3976] < btm_1[3975:3968]) ? 1 : 0;
assign detect_min[496][21] = (mid_1[3983:3976] < btm_1[3983:3976]) ? 1 : 0;
assign detect_min[496][22] = (mid_1[3983:3976] < btm_1[3991:3984]) ? 1 : 0;
assign detect_min[496][23] = (mid_1[3983:3976] < btm_2[3975:3968]) ? 1 : 0;
assign detect_min[496][24] = (mid_1[3983:3976] < btm_2[3983:3976]) ? 1 : 0;
assign detect_min[496][25] = (mid_1[3983:3976] < btm_2[3991:3984]) ? 1 : 0;

assign detect_min[497][0] = (mid_1[3991:3984] < top_0[3983:3976]) ? 1 : 0;
assign detect_min[497][1] = (mid_1[3991:3984] < top_0[3991:3984]) ? 1 : 0;
assign detect_min[497][2] = (mid_1[3991:3984] < top_0[3999:3992]) ? 1 : 0;
assign detect_min[497][3] = (mid_1[3991:3984] < top_1[3983:3976]) ? 1 : 0;
assign detect_min[497][4] = (mid_1[3991:3984] < top_1[3991:3984]) ? 1 : 0;
assign detect_min[497][5] = (mid_1[3991:3984] < top_1[3999:3992]) ? 1 : 0;
assign detect_min[497][6] = (mid_1[3991:3984] < top_2[3983:3976]) ? 1 : 0;
assign detect_min[497][7] = (mid_1[3991:3984] < top_2[3991:3984]) ? 1 : 0;
assign detect_min[497][8] = (mid_1[3991:3984] < top_2[3999:3992]) ? 1 : 0;
assign detect_min[497][9] = (mid_1[3991:3984] < mid_0[3983:3976]) ? 1 : 0;
assign detect_min[497][10] = (mid_1[3991:3984] < mid_0[3991:3984]) ? 1 : 0;
assign detect_min[497][11] = (mid_1[3991:3984] < mid_0[3999:3992]) ? 1 : 0;
assign detect_min[497][12] = (mid_1[3991:3984] < mid_1[3983:3976]) ? 1 : 0;
assign detect_min[497][13] = (mid_1[3991:3984] < mid_1[3999:3992]) ? 1 : 0;
assign detect_min[497][14] = (mid_1[3991:3984] < mid_2[3983:3976]) ? 1 : 0;
assign detect_min[497][15] = (mid_1[3991:3984] < mid_2[3991:3984]) ? 1 : 0;
assign detect_min[497][16] = (mid_1[3991:3984] < mid_2[3999:3992]) ? 1 : 0;
assign detect_min[497][17] = (mid_1[3991:3984] < btm_0[3983:3976]) ? 1 : 0;
assign detect_min[497][18] = (mid_1[3991:3984] < btm_0[3991:3984]) ? 1 : 0;
assign detect_min[497][19] = (mid_1[3991:3984] < btm_0[3999:3992]) ? 1 : 0;
assign detect_min[497][20] = (mid_1[3991:3984] < btm_1[3983:3976]) ? 1 : 0;
assign detect_min[497][21] = (mid_1[3991:3984] < btm_1[3991:3984]) ? 1 : 0;
assign detect_min[497][22] = (mid_1[3991:3984] < btm_1[3999:3992]) ? 1 : 0;
assign detect_min[497][23] = (mid_1[3991:3984] < btm_2[3983:3976]) ? 1 : 0;
assign detect_min[497][24] = (mid_1[3991:3984] < btm_2[3991:3984]) ? 1 : 0;
assign detect_min[497][25] = (mid_1[3991:3984] < btm_2[3999:3992]) ? 1 : 0;

assign detect_min[498][0] = (mid_1[3999:3992] < top_0[3991:3984]) ? 1 : 0;
assign detect_min[498][1] = (mid_1[3999:3992] < top_0[3999:3992]) ? 1 : 0;
assign detect_min[498][2] = (mid_1[3999:3992] < top_0[4007:4000]) ? 1 : 0;
assign detect_min[498][3] = (mid_1[3999:3992] < top_1[3991:3984]) ? 1 : 0;
assign detect_min[498][4] = (mid_1[3999:3992] < top_1[3999:3992]) ? 1 : 0;
assign detect_min[498][5] = (mid_1[3999:3992] < top_1[4007:4000]) ? 1 : 0;
assign detect_min[498][6] = (mid_1[3999:3992] < top_2[3991:3984]) ? 1 : 0;
assign detect_min[498][7] = (mid_1[3999:3992] < top_2[3999:3992]) ? 1 : 0;
assign detect_min[498][8] = (mid_1[3999:3992] < top_2[4007:4000]) ? 1 : 0;
assign detect_min[498][9] = (mid_1[3999:3992] < mid_0[3991:3984]) ? 1 : 0;
assign detect_min[498][10] = (mid_1[3999:3992] < mid_0[3999:3992]) ? 1 : 0;
assign detect_min[498][11] = (mid_1[3999:3992] < mid_0[4007:4000]) ? 1 : 0;
assign detect_min[498][12] = (mid_1[3999:3992] < mid_1[3991:3984]) ? 1 : 0;
assign detect_min[498][13] = (mid_1[3999:3992] < mid_1[4007:4000]) ? 1 : 0;
assign detect_min[498][14] = (mid_1[3999:3992] < mid_2[3991:3984]) ? 1 : 0;
assign detect_min[498][15] = (mid_1[3999:3992] < mid_2[3999:3992]) ? 1 : 0;
assign detect_min[498][16] = (mid_1[3999:3992] < mid_2[4007:4000]) ? 1 : 0;
assign detect_min[498][17] = (mid_1[3999:3992] < btm_0[3991:3984]) ? 1 : 0;
assign detect_min[498][18] = (mid_1[3999:3992] < btm_0[3999:3992]) ? 1 : 0;
assign detect_min[498][19] = (mid_1[3999:3992] < btm_0[4007:4000]) ? 1 : 0;
assign detect_min[498][20] = (mid_1[3999:3992] < btm_1[3991:3984]) ? 1 : 0;
assign detect_min[498][21] = (mid_1[3999:3992] < btm_1[3999:3992]) ? 1 : 0;
assign detect_min[498][22] = (mid_1[3999:3992] < btm_1[4007:4000]) ? 1 : 0;
assign detect_min[498][23] = (mid_1[3999:3992] < btm_2[3991:3984]) ? 1 : 0;
assign detect_min[498][24] = (mid_1[3999:3992] < btm_2[3999:3992]) ? 1 : 0;
assign detect_min[498][25] = (mid_1[3999:3992] < btm_2[4007:4000]) ? 1 : 0;

assign detect_min[499][0] = (mid_1[4007:4000] < top_0[3999:3992]) ? 1 : 0;
assign detect_min[499][1] = (mid_1[4007:4000] < top_0[4007:4000]) ? 1 : 0;
assign detect_min[499][2] = (mid_1[4007:4000] < top_0[4015:4008]) ? 1 : 0;
assign detect_min[499][3] = (mid_1[4007:4000] < top_1[3999:3992]) ? 1 : 0;
assign detect_min[499][4] = (mid_1[4007:4000] < top_1[4007:4000]) ? 1 : 0;
assign detect_min[499][5] = (mid_1[4007:4000] < top_1[4015:4008]) ? 1 : 0;
assign detect_min[499][6] = (mid_1[4007:4000] < top_2[3999:3992]) ? 1 : 0;
assign detect_min[499][7] = (mid_1[4007:4000] < top_2[4007:4000]) ? 1 : 0;
assign detect_min[499][8] = (mid_1[4007:4000] < top_2[4015:4008]) ? 1 : 0;
assign detect_min[499][9] = (mid_1[4007:4000] < mid_0[3999:3992]) ? 1 : 0;
assign detect_min[499][10] = (mid_1[4007:4000] < mid_0[4007:4000]) ? 1 : 0;
assign detect_min[499][11] = (mid_1[4007:4000] < mid_0[4015:4008]) ? 1 : 0;
assign detect_min[499][12] = (mid_1[4007:4000] < mid_1[3999:3992]) ? 1 : 0;
assign detect_min[499][13] = (mid_1[4007:4000] < mid_1[4015:4008]) ? 1 : 0;
assign detect_min[499][14] = (mid_1[4007:4000] < mid_2[3999:3992]) ? 1 : 0;
assign detect_min[499][15] = (mid_1[4007:4000] < mid_2[4007:4000]) ? 1 : 0;
assign detect_min[499][16] = (mid_1[4007:4000] < mid_2[4015:4008]) ? 1 : 0;
assign detect_min[499][17] = (mid_1[4007:4000] < btm_0[3999:3992]) ? 1 : 0;
assign detect_min[499][18] = (mid_1[4007:4000] < btm_0[4007:4000]) ? 1 : 0;
assign detect_min[499][19] = (mid_1[4007:4000] < btm_0[4015:4008]) ? 1 : 0;
assign detect_min[499][20] = (mid_1[4007:4000] < btm_1[3999:3992]) ? 1 : 0;
assign detect_min[499][21] = (mid_1[4007:4000] < btm_1[4007:4000]) ? 1 : 0;
assign detect_min[499][22] = (mid_1[4007:4000] < btm_1[4015:4008]) ? 1 : 0;
assign detect_min[499][23] = (mid_1[4007:4000] < btm_2[3999:3992]) ? 1 : 0;
assign detect_min[499][24] = (mid_1[4007:4000] < btm_2[4007:4000]) ? 1 : 0;
assign detect_min[499][25] = (mid_1[4007:4000] < btm_2[4015:4008]) ? 1 : 0;

assign detect_min[500][0] = (mid_1[4015:4008] < top_0[4007:4000]) ? 1 : 0;
assign detect_min[500][1] = (mid_1[4015:4008] < top_0[4015:4008]) ? 1 : 0;
assign detect_min[500][2] = (mid_1[4015:4008] < top_0[4023:4016]) ? 1 : 0;
assign detect_min[500][3] = (mid_1[4015:4008] < top_1[4007:4000]) ? 1 : 0;
assign detect_min[500][4] = (mid_1[4015:4008] < top_1[4015:4008]) ? 1 : 0;
assign detect_min[500][5] = (mid_1[4015:4008] < top_1[4023:4016]) ? 1 : 0;
assign detect_min[500][6] = (mid_1[4015:4008] < top_2[4007:4000]) ? 1 : 0;
assign detect_min[500][7] = (mid_1[4015:4008] < top_2[4015:4008]) ? 1 : 0;
assign detect_min[500][8] = (mid_1[4015:4008] < top_2[4023:4016]) ? 1 : 0;
assign detect_min[500][9] = (mid_1[4015:4008] < mid_0[4007:4000]) ? 1 : 0;
assign detect_min[500][10] = (mid_1[4015:4008] < mid_0[4015:4008]) ? 1 : 0;
assign detect_min[500][11] = (mid_1[4015:4008] < mid_0[4023:4016]) ? 1 : 0;
assign detect_min[500][12] = (mid_1[4015:4008] < mid_1[4007:4000]) ? 1 : 0;
assign detect_min[500][13] = (mid_1[4015:4008] < mid_1[4023:4016]) ? 1 : 0;
assign detect_min[500][14] = (mid_1[4015:4008] < mid_2[4007:4000]) ? 1 : 0;
assign detect_min[500][15] = (mid_1[4015:4008] < mid_2[4015:4008]) ? 1 : 0;
assign detect_min[500][16] = (mid_1[4015:4008] < mid_2[4023:4016]) ? 1 : 0;
assign detect_min[500][17] = (mid_1[4015:4008] < btm_0[4007:4000]) ? 1 : 0;
assign detect_min[500][18] = (mid_1[4015:4008] < btm_0[4015:4008]) ? 1 : 0;
assign detect_min[500][19] = (mid_1[4015:4008] < btm_0[4023:4016]) ? 1 : 0;
assign detect_min[500][20] = (mid_1[4015:4008] < btm_1[4007:4000]) ? 1 : 0;
assign detect_min[500][21] = (mid_1[4015:4008] < btm_1[4015:4008]) ? 1 : 0;
assign detect_min[500][22] = (mid_1[4015:4008] < btm_1[4023:4016]) ? 1 : 0;
assign detect_min[500][23] = (mid_1[4015:4008] < btm_2[4007:4000]) ? 1 : 0;
assign detect_min[500][24] = (mid_1[4015:4008] < btm_2[4015:4008]) ? 1 : 0;
assign detect_min[500][25] = (mid_1[4015:4008] < btm_2[4023:4016]) ? 1 : 0;

assign detect_min[501][0] = (mid_1[4023:4016] < top_0[4015:4008]) ? 1 : 0;
assign detect_min[501][1] = (mid_1[4023:4016] < top_0[4023:4016]) ? 1 : 0;
assign detect_min[501][2] = (mid_1[4023:4016] < top_0[4031:4024]) ? 1 : 0;
assign detect_min[501][3] = (mid_1[4023:4016] < top_1[4015:4008]) ? 1 : 0;
assign detect_min[501][4] = (mid_1[4023:4016] < top_1[4023:4016]) ? 1 : 0;
assign detect_min[501][5] = (mid_1[4023:4016] < top_1[4031:4024]) ? 1 : 0;
assign detect_min[501][6] = (mid_1[4023:4016] < top_2[4015:4008]) ? 1 : 0;
assign detect_min[501][7] = (mid_1[4023:4016] < top_2[4023:4016]) ? 1 : 0;
assign detect_min[501][8] = (mid_1[4023:4016] < top_2[4031:4024]) ? 1 : 0;
assign detect_min[501][9] = (mid_1[4023:4016] < mid_0[4015:4008]) ? 1 : 0;
assign detect_min[501][10] = (mid_1[4023:4016] < mid_0[4023:4016]) ? 1 : 0;
assign detect_min[501][11] = (mid_1[4023:4016] < mid_0[4031:4024]) ? 1 : 0;
assign detect_min[501][12] = (mid_1[4023:4016] < mid_1[4015:4008]) ? 1 : 0;
assign detect_min[501][13] = (mid_1[4023:4016] < mid_1[4031:4024]) ? 1 : 0;
assign detect_min[501][14] = (mid_1[4023:4016] < mid_2[4015:4008]) ? 1 : 0;
assign detect_min[501][15] = (mid_1[4023:4016] < mid_2[4023:4016]) ? 1 : 0;
assign detect_min[501][16] = (mid_1[4023:4016] < mid_2[4031:4024]) ? 1 : 0;
assign detect_min[501][17] = (mid_1[4023:4016] < btm_0[4015:4008]) ? 1 : 0;
assign detect_min[501][18] = (mid_1[4023:4016] < btm_0[4023:4016]) ? 1 : 0;
assign detect_min[501][19] = (mid_1[4023:4016] < btm_0[4031:4024]) ? 1 : 0;
assign detect_min[501][20] = (mid_1[4023:4016] < btm_1[4015:4008]) ? 1 : 0;
assign detect_min[501][21] = (mid_1[4023:4016] < btm_1[4023:4016]) ? 1 : 0;
assign detect_min[501][22] = (mid_1[4023:4016] < btm_1[4031:4024]) ? 1 : 0;
assign detect_min[501][23] = (mid_1[4023:4016] < btm_2[4015:4008]) ? 1 : 0;
assign detect_min[501][24] = (mid_1[4023:4016] < btm_2[4023:4016]) ? 1 : 0;
assign detect_min[501][25] = (mid_1[4023:4016] < btm_2[4031:4024]) ? 1 : 0;

assign detect_min[502][0] = (mid_1[4031:4024] < top_0[4023:4016]) ? 1 : 0;
assign detect_min[502][1] = (mid_1[4031:4024] < top_0[4031:4024]) ? 1 : 0;
assign detect_min[502][2] = (mid_1[4031:4024] < top_0[4039:4032]) ? 1 : 0;
assign detect_min[502][3] = (mid_1[4031:4024] < top_1[4023:4016]) ? 1 : 0;
assign detect_min[502][4] = (mid_1[4031:4024] < top_1[4031:4024]) ? 1 : 0;
assign detect_min[502][5] = (mid_1[4031:4024] < top_1[4039:4032]) ? 1 : 0;
assign detect_min[502][6] = (mid_1[4031:4024] < top_2[4023:4016]) ? 1 : 0;
assign detect_min[502][7] = (mid_1[4031:4024] < top_2[4031:4024]) ? 1 : 0;
assign detect_min[502][8] = (mid_1[4031:4024] < top_2[4039:4032]) ? 1 : 0;
assign detect_min[502][9] = (mid_1[4031:4024] < mid_0[4023:4016]) ? 1 : 0;
assign detect_min[502][10] = (mid_1[4031:4024] < mid_0[4031:4024]) ? 1 : 0;
assign detect_min[502][11] = (mid_1[4031:4024] < mid_0[4039:4032]) ? 1 : 0;
assign detect_min[502][12] = (mid_1[4031:4024] < mid_1[4023:4016]) ? 1 : 0;
assign detect_min[502][13] = (mid_1[4031:4024] < mid_1[4039:4032]) ? 1 : 0;
assign detect_min[502][14] = (mid_1[4031:4024] < mid_2[4023:4016]) ? 1 : 0;
assign detect_min[502][15] = (mid_1[4031:4024] < mid_2[4031:4024]) ? 1 : 0;
assign detect_min[502][16] = (mid_1[4031:4024] < mid_2[4039:4032]) ? 1 : 0;
assign detect_min[502][17] = (mid_1[4031:4024] < btm_0[4023:4016]) ? 1 : 0;
assign detect_min[502][18] = (mid_1[4031:4024] < btm_0[4031:4024]) ? 1 : 0;
assign detect_min[502][19] = (mid_1[4031:4024] < btm_0[4039:4032]) ? 1 : 0;
assign detect_min[502][20] = (mid_1[4031:4024] < btm_1[4023:4016]) ? 1 : 0;
assign detect_min[502][21] = (mid_1[4031:4024] < btm_1[4031:4024]) ? 1 : 0;
assign detect_min[502][22] = (mid_1[4031:4024] < btm_1[4039:4032]) ? 1 : 0;
assign detect_min[502][23] = (mid_1[4031:4024] < btm_2[4023:4016]) ? 1 : 0;
assign detect_min[502][24] = (mid_1[4031:4024] < btm_2[4031:4024]) ? 1 : 0;
assign detect_min[502][25] = (mid_1[4031:4024] < btm_2[4039:4032]) ? 1 : 0;

assign detect_min[503][0] = (mid_1[4039:4032] < top_0[4031:4024]) ? 1 : 0;
assign detect_min[503][1] = (mid_1[4039:4032] < top_0[4039:4032]) ? 1 : 0;
assign detect_min[503][2] = (mid_1[4039:4032] < top_0[4047:4040]) ? 1 : 0;
assign detect_min[503][3] = (mid_1[4039:4032] < top_1[4031:4024]) ? 1 : 0;
assign detect_min[503][4] = (mid_1[4039:4032] < top_1[4039:4032]) ? 1 : 0;
assign detect_min[503][5] = (mid_1[4039:4032] < top_1[4047:4040]) ? 1 : 0;
assign detect_min[503][6] = (mid_1[4039:4032] < top_2[4031:4024]) ? 1 : 0;
assign detect_min[503][7] = (mid_1[4039:4032] < top_2[4039:4032]) ? 1 : 0;
assign detect_min[503][8] = (mid_1[4039:4032] < top_2[4047:4040]) ? 1 : 0;
assign detect_min[503][9] = (mid_1[4039:4032] < mid_0[4031:4024]) ? 1 : 0;
assign detect_min[503][10] = (mid_1[4039:4032] < mid_0[4039:4032]) ? 1 : 0;
assign detect_min[503][11] = (mid_1[4039:4032] < mid_0[4047:4040]) ? 1 : 0;
assign detect_min[503][12] = (mid_1[4039:4032] < mid_1[4031:4024]) ? 1 : 0;
assign detect_min[503][13] = (mid_1[4039:4032] < mid_1[4047:4040]) ? 1 : 0;
assign detect_min[503][14] = (mid_1[4039:4032] < mid_2[4031:4024]) ? 1 : 0;
assign detect_min[503][15] = (mid_1[4039:4032] < mid_2[4039:4032]) ? 1 : 0;
assign detect_min[503][16] = (mid_1[4039:4032] < mid_2[4047:4040]) ? 1 : 0;
assign detect_min[503][17] = (mid_1[4039:4032] < btm_0[4031:4024]) ? 1 : 0;
assign detect_min[503][18] = (mid_1[4039:4032] < btm_0[4039:4032]) ? 1 : 0;
assign detect_min[503][19] = (mid_1[4039:4032] < btm_0[4047:4040]) ? 1 : 0;
assign detect_min[503][20] = (mid_1[4039:4032] < btm_1[4031:4024]) ? 1 : 0;
assign detect_min[503][21] = (mid_1[4039:4032] < btm_1[4039:4032]) ? 1 : 0;
assign detect_min[503][22] = (mid_1[4039:4032] < btm_1[4047:4040]) ? 1 : 0;
assign detect_min[503][23] = (mid_1[4039:4032] < btm_2[4031:4024]) ? 1 : 0;
assign detect_min[503][24] = (mid_1[4039:4032] < btm_2[4039:4032]) ? 1 : 0;
assign detect_min[503][25] = (mid_1[4039:4032] < btm_2[4047:4040]) ? 1 : 0;

assign detect_min[504][0] = (mid_1[4047:4040] < top_0[4039:4032]) ? 1 : 0;
assign detect_min[504][1] = (mid_1[4047:4040] < top_0[4047:4040]) ? 1 : 0;
assign detect_min[504][2] = (mid_1[4047:4040] < top_0[4055:4048]) ? 1 : 0;
assign detect_min[504][3] = (mid_1[4047:4040] < top_1[4039:4032]) ? 1 : 0;
assign detect_min[504][4] = (mid_1[4047:4040] < top_1[4047:4040]) ? 1 : 0;
assign detect_min[504][5] = (mid_1[4047:4040] < top_1[4055:4048]) ? 1 : 0;
assign detect_min[504][6] = (mid_1[4047:4040] < top_2[4039:4032]) ? 1 : 0;
assign detect_min[504][7] = (mid_1[4047:4040] < top_2[4047:4040]) ? 1 : 0;
assign detect_min[504][8] = (mid_1[4047:4040] < top_2[4055:4048]) ? 1 : 0;
assign detect_min[504][9] = (mid_1[4047:4040] < mid_0[4039:4032]) ? 1 : 0;
assign detect_min[504][10] = (mid_1[4047:4040] < mid_0[4047:4040]) ? 1 : 0;
assign detect_min[504][11] = (mid_1[4047:4040] < mid_0[4055:4048]) ? 1 : 0;
assign detect_min[504][12] = (mid_1[4047:4040] < mid_1[4039:4032]) ? 1 : 0;
assign detect_min[504][13] = (mid_1[4047:4040] < mid_1[4055:4048]) ? 1 : 0;
assign detect_min[504][14] = (mid_1[4047:4040] < mid_2[4039:4032]) ? 1 : 0;
assign detect_min[504][15] = (mid_1[4047:4040] < mid_2[4047:4040]) ? 1 : 0;
assign detect_min[504][16] = (mid_1[4047:4040] < mid_2[4055:4048]) ? 1 : 0;
assign detect_min[504][17] = (mid_1[4047:4040] < btm_0[4039:4032]) ? 1 : 0;
assign detect_min[504][18] = (mid_1[4047:4040] < btm_0[4047:4040]) ? 1 : 0;
assign detect_min[504][19] = (mid_1[4047:4040] < btm_0[4055:4048]) ? 1 : 0;
assign detect_min[504][20] = (mid_1[4047:4040] < btm_1[4039:4032]) ? 1 : 0;
assign detect_min[504][21] = (mid_1[4047:4040] < btm_1[4047:4040]) ? 1 : 0;
assign detect_min[504][22] = (mid_1[4047:4040] < btm_1[4055:4048]) ? 1 : 0;
assign detect_min[504][23] = (mid_1[4047:4040] < btm_2[4039:4032]) ? 1 : 0;
assign detect_min[504][24] = (mid_1[4047:4040] < btm_2[4047:4040]) ? 1 : 0;
assign detect_min[504][25] = (mid_1[4047:4040] < btm_2[4055:4048]) ? 1 : 0;

assign detect_min[505][0] = (mid_1[4055:4048] < top_0[4047:4040]) ? 1 : 0;
assign detect_min[505][1] = (mid_1[4055:4048] < top_0[4055:4048]) ? 1 : 0;
assign detect_min[505][2] = (mid_1[4055:4048] < top_0[4063:4056]) ? 1 : 0;
assign detect_min[505][3] = (mid_1[4055:4048] < top_1[4047:4040]) ? 1 : 0;
assign detect_min[505][4] = (mid_1[4055:4048] < top_1[4055:4048]) ? 1 : 0;
assign detect_min[505][5] = (mid_1[4055:4048] < top_1[4063:4056]) ? 1 : 0;
assign detect_min[505][6] = (mid_1[4055:4048] < top_2[4047:4040]) ? 1 : 0;
assign detect_min[505][7] = (mid_1[4055:4048] < top_2[4055:4048]) ? 1 : 0;
assign detect_min[505][8] = (mid_1[4055:4048] < top_2[4063:4056]) ? 1 : 0;
assign detect_min[505][9] = (mid_1[4055:4048] < mid_0[4047:4040]) ? 1 : 0;
assign detect_min[505][10] = (mid_1[4055:4048] < mid_0[4055:4048]) ? 1 : 0;
assign detect_min[505][11] = (mid_1[4055:4048] < mid_0[4063:4056]) ? 1 : 0;
assign detect_min[505][12] = (mid_1[4055:4048] < mid_1[4047:4040]) ? 1 : 0;
assign detect_min[505][13] = (mid_1[4055:4048] < mid_1[4063:4056]) ? 1 : 0;
assign detect_min[505][14] = (mid_1[4055:4048] < mid_2[4047:4040]) ? 1 : 0;
assign detect_min[505][15] = (mid_1[4055:4048] < mid_2[4055:4048]) ? 1 : 0;
assign detect_min[505][16] = (mid_1[4055:4048] < mid_2[4063:4056]) ? 1 : 0;
assign detect_min[505][17] = (mid_1[4055:4048] < btm_0[4047:4040]) ? 1 : 0;
assign detect_min[505][18] = (mid_1[4055:4048] < btm_0[4055:4048]) ? 1 : 0;
assign detect_min[505][19] = (mid_1[4055:4048] < btm_0[4063:4056]) ? 1 : 0;
assign detect_min[505][20] = (mid_1[4055:4048] < btm_1[4047:4040]) ? 1 : 0;
assign detect_min[505][21] = (mid_1[4055:4048] < btm_1[4055:4048]) ? 1 : 0;
assign detect_min[505][22] = (mid_1[4055:4048] < btm_1[4063:4056]) ? 1 : 0;
assign detect_min[505][23] = (mid_1[4055:4048] < btm_2[4047:4040]) ? 1 : 0;
assign detect_min[505][24] = (mid_1[4055:4048] < btm_2[4055:4048]) ? 1 : 0;
assign detect_min[505][25] = (mid_1[4055:4048] < btm_2[4063:4056]) ? 1 : 0;

assign detect_min[506][0] = (mid_1[4063:4056] < top_0[4055:4048]) ? 1 : 0;
assign detect_min[506][1] = (mid_1[4063:4056] < top_0[4063:4056]) ? 1 : 0;
assign detect_min[506][2] = (mid_1[4063:4056] < top_0[4071:4064]) ? 1 : 0;
assign detect_min[506][3] = (mid_1[4063:4056] < top_1[4055:4048]) ? 1 : 0;
assign detect_min[506][4] = (mid_1[4063:4056] < top_1[4063:4056]) ? 1 : 0;
assign detect_min[506][5] = (mid_1[4063:4056] < top_1[4071:4064]) ? 1 : 0;
assign detect_min[506][6] = (mid_1[4063:4056] < top_2[4055:4048]) ? 1 : 0;
assign detect_min[506][7] = (mid_1[4063:4056] < top_2[4063:4056]) ? 1 : 0;
assign detect_min[506][8] = (mid_1[4063:4056] < top_2[4071:4064]) ? 1 : 0;
assign detect_min[506][9] = (mid_1[4063:4056] < mid_0[4055:4048]) ? 1 : 0;
assign detect_min[506][10] = (mid_1[4063:4056] < mid_0[4063:4056]) ? 1 : 0;
assign detect_min[506][11] = (mid_1[4063:4056] < mid_0[4071:4064]) ? 1 : 0;
assign detect_min[506][12] = (mid_1[4063:4056] < mid_1[4055:4048]) ? 1 : 0;
assign detect_min[506][13] = (mid_1[4063:4056] < mid_1[4071:4064]) ? 1 : 0;
assign detect_min[506][14] = (mid_1[4063:4056] < mid_2[4055:4048]) ? 1 : 0;
assign detect_min[506][15] = (mid_1[4063:4056] < mid_2[4063:4056]) ? 1 : 0;
assign detect_min[506][16] = (mid_1[4063:4056] < mid_2[4071:4064]) ? 1 : 0;
assign detect_min[506][17] = (mid_1[4063:4056] < btm_0[4055:4048]) ? 1 : 0;
assign detect_min[506][18] = (mid_1[4063:4056] < btm_0[4063:4056]) ? 1 : 0;
assign detect_min[506][19] = (mid_1[4063:4056] < btm_0[4071:4064]) ? 1 : 0;
assign detect_min[506][20] = (mid_1[4063:4056] < btm_1[4055:4048]) ? 1 : 0;
assign detect_min[506][21] = (mid_1[4063:4056] < btm_1[4063:4056]) ? 1 : 0;
assign detect_min[506][22] = (mid_1[4063:4056] < btm_1[4071:4064]) ? 1 : 0;
assign detect_min[506][23] = (mid_1[4063:4056] < btm_2[4055:4048]) ? 1 : 0;
assign detect_min[506][24] = (mid_1[4063:4056] < btm_2[4063:4056]) ? 1 : 0;
assign detect_min[506][25] = (mid_1[4063:4056] < btm_2[4071:4064]) ? 1 : 0;

assign detect_min[507][0] = (mid_1[4071:4064] < top_0[4063:4056]) ? 1 : 0;
assign detect_min[507][1] = (mid_1[4071:4064] < top_0[4071:4064]) ? 1 : 0;
assign detect_min[507][2] = (mid_1[4071:4064] < top_0[4079:4072]) ? 1 : 0;
assign detect_min[507][3] = (mid_1[4071:4064] < top_1[4063:4056]) ? 1 : 0;
assign detect_min[507][4] = (mid_1[4071:4064] < top_1[4071:4064]) ? 1 : 0;
assign detect_min[507][5] = (mid_1[4071:4064] < top_1[4079:4072]) ? 1 : 0;
assign detect_min[507][6] = (mid_1[4071:4064] < top_2[4063:4056]) ? 1 : 0;
assign detect_min[507][7] = (mid_1[4071:4064] < top_2[4071:4064]) ? 1 : 0;
assign detect_min[507][8] = (mid_1[4071:4064] < top_2[4079:4072]) ? 1 : 0;
assign detect_min[507][9] = (mid_1[4071:4064] < mid_0[4063:4056]) ? 1 : 0;
assign detect_min[507][10] = (mid_1[4071:4064] < mid_0[4071:4064]) ? 1 : 0;
assign detect_min[507][11] = (mid_1[4071:4064] < mid_0[4079:4072]) ? 1 : 0;
assign detect_min[507][12] = (mid_1[4071:4064] < mid_1[4063:4056]) ? 1 : 0;
assign detect_min[507][13] = (mid_1[4071:4064] < mid_1[4079:4072]) ? 1 : 0;
assign detect_min[507][14] = (mid_1[4071:4064] < mid_2[4063:4056]) ? 1 : 0;
assign detect_min[507][15] = (mid_1[4071:4064] < mid_2[4071:4064]) ? 1 : 0;
assign detect_min[507][16] = (mid_1[4071:4064] < mid_2[4079:4072]) ? 1 : 0;
assign detect_min[507][17] = (mid_1[4071:4064] < btm_0[4063:4056]) ? 1 : 0;
assign detect_min[507][18] = (mid_1[4071:4064] < btm_0[4071:4064]) ? 1 : 0;
assign detect_min[507][19] = (mid_1[4071:4064] < btm_0[4079:4072]) ? 1 : 0;
assign detect_min[507][20] = (mid_1[4071:4064] < btm_1[4063:4056]) ? 1 : 0;
assign detect_min[507][21] = (mid_1[4071:4064] < btm_1[4071:4064]) ? 1 : 0;
assign detect_min[507][22] = (mid_1[4071:4064] < btm_1[4079:4072]) ? 1 : 0;
assign detect_min[507][23] = (mid_1[4071:4064] < btm_2[4063:4056]) ? 1 : 0;
assign detect_min[507][24] = (mid_1[4071:4064] < btm_2[4071:4064]) ? 1 : 0;
assign detect_min[507][25] = (mid_1[4071:4064] < btm_2[4079:4072]) ? 1 : 0;

assign detect_min[508][0] = (mid_1[4079:4072] < top_0[4071:4064]) ? 1 : 0;
assign detect_min[508][1] = (mid_1[4079:4072] < top_0[4079:4072]) ? 1 : 0;
assign detect_min[508][2] = (mid_1[4079:4072] < top_0[4087:4080]) ? 1 : 0;
assign detect_min[508][3] = (mid_1[4079:4072] < top_1[4071:4064]) ? 1 : 0;
assign detect_min[508][4] = (mid_1[4079:4072] < top_1[4079:4072]) ? 1 : 0;
assign detect_min[508][5] = (mid_1[4079:4072] < top_1[4087:4080]) ? 1 : 0;
assign detect_min[508][6] = (mid_1[4079:4072] < top_2[4071:4064]) ? 1 : 0;
assign detect_min[508][7] = (mid_1[4079:4072] < top_2[4079:4072]) ? 1 : 0;
assign detect_min[508][8] = (mid_1[4079:4072] < top_2[4087:4080]) ? 1 : 0;
assign detect_min[508][9] = (mid_1[4079:4072] < mid_0[4071:4064]) ? 1 : 0;
assign detect_min[508][10] = (mid_1[4079:4072] < mid_0[4079:4072]) ? 1 : 0;
assign detect_min[508][11] = (mid_1[4079:4072] < mid_0[4087:4080]) ? 1 : 0;
assign detect_min[508][12] = (mid_1[4079:4072] < mid_1[4071:4064]) ? 1 : 0;
assign detect_min[508][13] = (mid_1[4079:4072] < mid_1[4087:4080]) ? 1 : 0;
assign detect_min[508][14] = (mid_1[4079:4072] < mid_2[4071:4064]) ? 1 : 0;
assign detect_min[508][15] = (mid_1[4079:4072] < mid_2[4079:4072]) ? 1 : 0;
assign detect_min[508][16] = (mid_1[4079:4072] < mid_2[4087:4080]) ? 1 : 0;
assign detect_min[508][17] = (mid_1[4079:4072] < btm_0[4071:4064]) ? 1 : 0;
assign detect_min[508][18] = (mid_1[4079:4072] < btm_0[4079:4072]) ? 1 : 0;
assign detect_min[508][19] = (mid_1[4079:4072] < btm_0[4087:4080]) ? 1 : 0;
assign detect_min[508][20] = (mid_1[4079:4072] < btm_1[4071:4064]) ? 1 : 0;
assign detect_min[508][21] = (mid_1[4079:4072] < btm_1[4079:4072]) ? 1 : 0;
assign detect_min[508][22] = (mid_1[4079:4072] < btm_1[4087:4080]) ? 1 : 0;
assign detect_min[508][23] = (mid_1[4079:4072] < btm_2[4071:4064]) ? 1 : 0;
assign detect_min[508][24] = (mid_1[4079:4072] < btm_2[4079:4072]) ? 1 : 0;
assign detect_min[508][25] = (mid_1[4079:4072] < btm_2[4087:4080]) ? 1 : 0;

assign detect_min[509][0] = (mid_1[4087:4080] < top_0[4079:4072]) ? 1 : 0;
assign detect_min[509][1] = (mid_1[4087:4080] < top_0[4087:4080]) ? 1 : 0;
assign detect_min[509][2] = (mid_1[4087:4080] < top_0[4095:4088]) ? 1 : 0;
assign detect_min[509][3] = (mid_1[4087:4080] < top_1[4079:4072]) ? 1 : 0;
assign detect_min[509][4] = (mid_1[4087:4080] < top_1[4087:4080]) ? 1 : 0;
assign detect_min[509][5] = (mid_1[4087:4080] < top_1[4095:4088]) ? 1 : 0;
assign detect_min[509][6] = (mid_1[4087:4080] < top_2[4079:4072]) ? 1 : 0;
assign detect_min[509][7] = (mid_1[4087:4080] < top_2[4087:4080]) ? 1 : 0;
assign detect_min[509][8] = (mid_1[4087:4080] < top_2[4095:4088]) ? 1 : 0;
assign detect_min[509][9] = (mid_1[4087:4080] < mid_0[4079:4072]) ? 1 : 0;
assign detect_min[509][10] = (mid_1[4087:4080] < mid_0[4087:4080]) ? 1 : 0;
assign detect_min[509][11] = (mid_1[4087:4080] < mid_0[4095:4088]) ? 1 : 0;
assign detect_min[509][12] = (mid_1[4087:4080] < mid_1[4079:4072]) ? 1 : 0;
assign detect_min[509][13] = (mid_1[4087:4080] < mid_1[4095:4088]) ? 1 : 0;
assign detect_min[509][14] = (mid_1[4087:4080] < mid_2[4079:4072]) ? 1 : 0;
assign detect_min[509][15] = (mid_1[4087:4080] < mid_2[4087:4080]) ? 1 : 0;
assign detect_min[509][16] = (mid_1[4087:4080] < mid_2[4095:4088]) ? 1 : 0;
assign detect_min[509][17] = (mid_1[4087:4080] < btm_0[4079:4072]) ? 1 : 0;
assign detect_min[509][18] = (mid_1[4087:4080] < btm_0[4087:4080]) ? 1 : 0;
assign detect_min[509][19] = (mid_1[4087:4080] < btm_0[4095:4088]) ? 1 : 0;
assign detect_min[509][20] = (mid_1[4087:4080] < btm_1[4079:4072]) ? 1 : 0;
assign detect_min[509][21] = (mid_1[4087:4080] < btm_1[4087:4080]) ? 1 : 0;
assign detect_min[509][22] = (mid_1[4087:4080] < btm_1[4095:4088]) ? 1 : 0;
assign detect_min[509][23] = (mid_1[4087:4080] < btm_2[4079:4072]) ? 1 : 0;
assign detect_min[509][24] = (mid_1[4087:4080] < btm_2[4087:4080]) ? 1 : 0;
assign detect_min[509][25] = (mid_1[4087:4080] < btm_2[4095:4088]) ? 1 : 0;

assign detect_min[510][0] = (mid_1[4095:4088] < top_0[4087:4080]) ? 1 : 0;
assign detect_min[510][1] = (mid_1[4095:4088] < top_0[4095:4088]) ? 1 : 0;
assign detect_min[510][2] = (mid_1[4095:4088] < top_0[4103:4096]) ? 1 : 0;
assign detect_min[510][3] = (mid_1[4095:4088] < top_1[4087:4080]) ? 1 : 0;
assign detect_min[510][4] = (mid_1[4095:4088] < top_1[4095:4088]) ? 1 : 0;
assign detect_min[510][5] = (mid_1[4095:4088] < top_1[4103:4096]) ? 1 : 0;
assign detect_min[510][6] = (mid_1[4095:4088] < top_2[4087:4080]) ? 1 : 0;
assign detect_min[510][7] = (mid_1[4095:4088] < top_2[4095:4088]) ? 1 : 0;
assign detect_min[510][8] = (mid_1[4095:4088] < top_2[4103:4096]) ? 1 : 0;
assign detect_min[510][9] = (mid_1[4095:4088] < mid_0[4087:4080]) ? 1 : 0;
assign detect_min[510][10] = (mid_1[4095:4088] < mid_0[4095:4088]) ? 1 : 0;
assign detect_min[510][11] = (mid_1[4095:4088] < mid_0[4103:4096]) ? 1 : 0;
assign detect_min[510][12] = (mid_1[4095:4088] < mid_1[4087:4080]) ? 1 : 0;
assign detect_min[510][13] = (mid_1[4095:4088] < mid_1[4103:4096]) ? 1 : 0;
assign detect_min[510][14] = (mid_1[4095:4088] < mid_2[4087:4080]) ? 1 : 0;
assign detect_min[510][15] = (mid_1[4095:4088] < mid_2[4095:4088]) ? 1 : 0;
assign detect_min[510][16] = (mid_1[4095:4088] < mid_2[4103:4096]) ? 1 : 0;
assign detect_min[510][17] = (mid_1[4095:4088] < btm_0[4087:4080]) ? 1 : 0;
assign detect_min[510][18] = (mid_1[4095:4088] < btm_0[4095:4088]) ? 1 : 0;
assign detect_min[510][19] = (mid_1[4095:4088] < btm_0[4103:4096]) ? 1 : 0;
assign detect_min[510][20] = (mid_1[4095:4088] < btm_1[4087:4080]) ? 1 : 0;
assign detect_min[510][21] = (mid_1[4095:4088] < btm_1[4095:4088]) ? 1 : 0;
assign detect_min[510][22] = (mid_1[4095:4088] < btm_1[4103:4096]) ? 1 : 0;
assign detect_min[510][23] = (mid_1[4095:4088] < btm_2[4087:4080]) ? 1 : 0;
assign detect_min[510][24] = (mid_1[4095:4088] < btm_2[4095:4088]) ? 1 : 0;
assign detect_min[510][25] = (mid_1[4095:4088] < btm_2[4103:4096]) ? 1 : 0;

assign detect_min[511][0] = (mid_1[4103:4096] < top_0[4095:4088]) ? 1 : 0;
assign detect_min[511][1] = (mid_1[4103:4096] < top_0[4103:4096]) ? 1 : 0;
assign detect_min[511][2] = (mid_1[4103:4096] < top_0[4111:4104]) ? 1 : 0;
assign detect_min[511][3] = (mid_1[4103:4096] < top_1[4095:4088]) ? 1 : 0;
assign detect_min[511][4] = (mid_1[4103:4096] < top_1[4103:4096]) ? 1 : 0;
assign detect_min[511][5] = (mid_1[4103:4096] < top_1[4111:4104]) ? 1 : 0;
assign detect_min[511][6] = (mid_1[4103:4096] < top_2[4095:4088]) ? 1 : 0;
assign detect_min[511][7] = (mid_1[4103:4096] < top_2[4103:4096]) ? 1 : 0;
assign detect_min[511][8] = (mid_1[4103:4096] < top_2[4111:4104]) ? 1 : 0;
assign detect_min[511][9] = (mid_1[4103:4096] < mid_0[4095:4088]) ? 1 : 0;
assign detect_min[511][10] = (mid_1[4103:4096] < mid_0[4103:4096]) ? 1 : 0;
assign detect_min[511][11] = (mid_1[4103:4096] < mid_0[4111:4104]) ? 1 : 0;
assign detect_min[511][12] = (mid_1[4103:4096] < mid_1[4095:4088]) ? 1 : 0;
assign detect_min[511][13] = (mid_1[4103:4096] < mid_1[4111:4104]) ? 1 : 0;
assign detect_min[511][14] = (mid_1[4103:4096] < mid_2[4095:4088]) ? 1 : 0;
assign detect_min[511][15] = (mid_1[4103:4096] < mid_2[4103:4096]) ? 1 : 0;
assign detect_min[511][16] = (mid_1[4103:4096] < mid_2[4111:4104]) ? 1 : 0;
assign detect_min[511][17] = (mid_1[4103:4096] < btm_0[4095:4088]) ? 1 : 0;
assign detect_min[511][18] = (mid_1[4103:4096] < btm_0[4103:4096]) ? 1 : 0;
assign detect_min[511][19] = (mid_1[4103:4096] < btm_0[4111:4104]) ? 1 : 0;
assign detect_min[511][20] = (mid_1[4103:4096] < btm_1[4095:4088]) ? 1 : 0;
assign detect_min[511][21] = (mid_1[4103:4096] < btm_1[4103:4096]) ? 1 : 0;
assign detect_min[511][22] = (mid_1[4103:4096] < btm_1[4111:4104]) ? 1 : 0;
assign detect_min[511][23] = (mid_1[4103:4096] < btm_2[4095:4088]) ? 1 : 0;
assign detect_min[511][24] = (mid_1[4103:4096] < btm_2[4103:4096]) ? 1 : 0;
assign detect_min[511][25] = (mid_1[4103:4096] < btm_2[4111:4104]) ? 1 : 0;

assign detect_min[512][0] = (mid_1[4111:4104] < top_0[4103:4096]) ? 1 : 0;
assign detect_min[512][1] = (mid_1[4111:4104] < top_0[4111:4104]) ? 1 : 0;
assign detect_min[512][2] = (mid_1[4111:4104] < top_0[4119:4112]) ? 1 : 0;
assign detect_min[512][3] = (mid_1[4111:4104] < top_1[4103:4096]) ? 1 : 0;
assign detect_min[512][4] = (mid_1[4111:4104] < top_1[4111:4104]) ? 1 : 0;
assign detect_min[512][5] = (mid_1[4111:4104] < top_1[4119:4112]) ? 1 : 0;
assign detect_min[512][6] = (mid_1[4111:4104] < top_2[4103:4096]) ? 1 : 0;
assign detect_min[512][7] = (mid_1[4111:4104] < top_2[4111:4104]) ? 1 : 0;
assign detect_min[512][8] = (mid_1[4111:4104] < top_2[4119:4112]) ? 1 : 0;
assign detect_min[512][9] = (mid_1[4111:4104] < mid_0[4103:4096]) ? 1 : 0;
assign detect_min[512][10] = (mid_1[4111:4104] < mid_0[4111:4104]) ? 1 : 0;
assign detect_min[512][11] = (mid_1[4111:4104] < mid_0[4119:4112]) ? 1 : 0;
assign detect_min[512][12] = (mid_1[4111:4104] < mid_1[4103:4096]) ? 1 : 0;
assign detect_min[512][13] = (mid_1[4111:4104] < mid_1[4119:4112]) ? 1 : 0;
assign detect_min[512][14] = (mid_1[4111:4104] < mid_2[4103:4096]) ? 1 : 0;
assign detect_min[512][15] = (mid_1[4111:4104] < mid_2[4111:4104]) ? 1 : 0;
assign detect_min[512][16] = (mid_1[4111:4104] < mid_2[4119:4112]) ? 1 : 0;
assign detect_min[512][17] = (mid_1[4111:4104] < btm_0[4103:4096]) ? 1 : 0;
assign detect_min[512][18] = (mid_1[4111:4104] < btm_0[4111:4104]) ? 1 : 0;
assign detect_min[512][19] = (mid_1[4111:4104] < btm_0[4119:4112]) ? 1 : 0;
assign detect_min[512][20] = (mid_1[4111:4104] < btm_1[4103:4096]) ? 1 : 0;
assign detect_min[512][21] = (mid_1[4111:4104] < btm_1[4111:4104]) ? 1 : 0;
assign detect_min[512][22] = (mid_1[4111:4104] < btm_1[4119:4112]) ? 1 : 0;
assign detect_min[512][23] = (mid_1[4111:4104] < btm_2[4103:4096]) ? 1 : 0;
assign detect_min[512][24] = (mid_1[4111:4104] < btm_2[4111:4104]) ? 1 : 0;
assign detect_min[512][25] = (mid_1[4111:4104] < btm_2[4119:4112]) ? 1 : 0;

assign detect_min[513][0] = (mid_1[4119:4112] < top_0[4111:4104]) ? 1 : 0;
assign detect_min[513][1] = (mid_1[4119:4112] < top_0[4119:4112]) ? 1 : 0;
assign detect_min[513][2] = (mid_1[4119:4112] < top_0[4127:4120]) ? 1 : 0;
assign detect_min[513][3] = (mid_1[4119:4112] < top_1[4111:4104]) ? 1 : 0;
assign detect_min[513][4] = (mid_1[4119:4112] < top_1[4119:4112]) ? 1 : 0;
assign detect_min[513][5] = (mid_1[4119:4112] < top_1[4127:4120]) ? 1 : 0;
assign detect_min[513][6] = (mid_1[4119:4112] < top_2[4111:4104]) ? 1 : 0;
assign detect_min[513][7] = (mid_1[4119:4112] < top_2[4119:4112]) ? 1 : 0;
assign detect_min[513][8] = (mid_1[4119:4112] < top_2[4127:4120]) ? 1 : 0;
assign detect_min[513][9] = (mid_1[4119:4112] < mid_0[4111:4104]) ? 1 : 0;
assign detect_min[513][10] = (mid_1[4119:4112] < mid_0[4119:4112]) ? 1 : 0;
assign detect_min[513][11] = (mid_1[4119:4112] < mid_0[4127:4120]) ? 1 : 0;
assign detect_min[513][12] = (mid_1[4119:4112] < mid_1[4111:4104]) ? 1 : 0;
assign detect_min[513][13] = (mid_1[4119:4112] < mid_1[4127:4120]) ? 1 : 0;
assign detect_min[513][14] = (mid_1[4119:4112] < mid_2[4111:4104]) ? 1 : 0;
assign detect_min[513][15] = (mid_1[4119:4112] < mid_2[4119:4112]) ? 1 : 0;
assign detect_min[513][16] = (mid_1[4119:4112] < mid_2[4127:4120]) ? 1 : 0;
assign detect_min[513][17] = (mid_1[4119:4112] < btm_0[4111:4104]) ? 1 : 0;
assign detect_min[513][18] = (mid_1[4119:4112] < btm_0[4119:4112]) ? 1 : 0;
assign detect_min[513][19] = (mid_1[4119:4112] < btm_0[4127:4120]) ? 1 : 0;
assign detect_min[513][20] = (mid_1[4119:4112] < btm_1[4111:4104]) ? 1 : 0;
assign detect_min[513][21] = (mid_1[4119:4112] < btm_1[4119:4112]) ? 1 : 0;
assign detect_min[513][22] = (mid_1[4119:4112] < btm_1[4127:4120]) ? 1 : 0;
assign detect_min[513][23] = (mid_1[4119:4112] < btm_2[4111:4104]) ? 1 : 0;
assign detect_min[513][24] = (mid_1[4119:4112] < btm_2[4119:4112]) ? 1 : 0;
assign detect_min[513][25] = (mid_1[4119:4112] < btm_2[4127:4120]) ? 1 : 0;

assign detect_min[514][0] = (mid_1[4127:4120] < top_0[4119:4112]) ? 1 : 0;
assign detect_min[514][1] = (mid_1[4127:4120] < top_0[4127:4120]) ? 1 : 0;
assign detect_min[514][2] = (mid_1[4127:4120] < top_0[4135:4128]) ? 1 : 0;
assign detect_min[514][3] = (mid_1[4127:4120] < top_1[4119:4112]) ? 1 : 0;
assign detect_min[514][4] = (mid_1[4127:4120] < top_1[4127:4120]) ? 1 : 0;
assign detect_min[514][5] = (mid_1[4127:4120] < top_1[4135:4128]) ? 1 : 0;
assign detect_min[514][6] = (mid_1[4127:4120] < top_2[4119:4112]) ? 1 : 0;
assign detect_min[514][7] = (mid_1[4127:4120] < top_2[4127:4120]) ? 1 : 0;
assign detect_min[514][8] = (mid_1[4127:4120] < top_2[4135:4128]) ? 1 : 0;
assign detect_min[514][9] = (mid_1[4127:4120] < mid_0[4119:4112]) ? 1 : 0;
assign detect_min[514][10] = (mid_1[4127:4120] < mid_0[4127:4120]) ? 1 : 0;
assign detect_min[514][11] = (mid_1[4127:4120] < mid_0[4135:4128]) ? 1 : 0;
assign detect_min[514][12] = (mid_1[4127:4120] < mid_1[4119:4112]) ? 1 : 0;
assign detect_min[514][13] = (mid_1[4127:4120] < mid_1[4135:4128]) ? 1 : 0;
assign detect_min[514][14] = (mid_1[4127:4120] < mid_2[4119:4112]) ? 1 : 0;
assign detect_min[514][15] = (mid_1[4127:4120] < mid_2[4127:4120]) ? 1 : 0;
assign detect_min[514][16] = (mid_1[4127:4120] < mid_2[4135:4128]) ? 1 : 0;
assign detect_min[514][17] = (mid_1[4127:4120] < btm_0[4119:4112]) ? 1 : 0;
assign detect_min[514][18] = (mid_1[4127:4120] < btm_0[4127:4120]) ? 1 : 0;
assign detect_min[514][19] = (mid_1[4127:4120] < btm_0[4135:4128]) ? 1 : 0;
assign detect_min[514][20] = (mid_1[4127:4120] < btm_1[4119:4112]) ? 1 : 0;
assign detect_min[514][21] = (mid_1[4127:4120] < btm_1[4127:4120]) ? 1 : 0;
assign detect_min[514][22] = (mid_1[4127:4120] < btm_1[4135:4128]) ? 1 : 0;
assign detect_min[514][23] = (mid_1[4127:4120] < btm_2[4119:4112]) ? 1 : 0;
assign detect_min[514][24] = (mid_1[4127:4120] < btm_2[4127:4120]) ? 1 : 0;
assign detect_min[514][25] = (mid_1[4127:4120] < btm_2[4135:4128]) ? 1 : 0;

assign detect_min[515][0] = (mid_1[4135:4128] < top_0[4127:4120]) ? 1 : 0;
assign detect_min[515][1] = (mid_1[4135:4128] < top_0[4135:4128]) ? 1 : 0;
assign detect_min[515][2] = (mid_1[4135:4128] < top_0[4143:4136]) ? 1 : 0;
assign detect_min[515][3] = (mid_1[4135:4128] < top_1[4127:4120]) ? 1 : 0;
assign detect_min[515][4] = (mid_1[4135:4128] < top_1[4135:4128]) ? 1 : 0;
assign detect_min[515][5] = (mid_1[4135:4128] < top_1[4143:4136]) ? 1 : 0;
assign detect_min[515][6] = (mid_1[4135:4128] < top_2[4127:4120]) ? 1 : 0;
assign detect_min[515][7] = (mid_1[4135:4128] < top_2[4135:4128]) ? 1 : 0;
assign detect_min[515][8] = (mid_1[4135:4128] < top_2[4143:4136]) ? 1 : 0;
assign detect_min[515][9] = (mid_1[4135:4128] < mid_0[4127:4120]) ? 1 : 0;
assign detect_min[515][10] = (mid_1[4135:4128] < mid_0[4135:4128]) ? 1 : 0;
assign detect_min[515][11] = (mid_1[4135:4128] < mid_0[4143:4136]) ? 1 : 0;
assign detect_min[515][12] = (mid_1[4135:4128] < mid_1[4127:4120]) ? 1 : 0;
assign detect_min[515][13] = (mid_1[4135:4128] < mid_1[4143:4136]) ? 1 : 0;
assign detect_min[515][14] = (mid_1[4135:4128] < mid_2[4127:4120]) ? 1 : 0;
assign detect_min[515][15] = (mid_1[4135:4128] < mid_2[4135:4128]) ? 1 : 0;
assign detect_min[515][16] = (mid_1[4135:4128] < mid_2[4143:4136]) ? 1 : 0;
assign detect_min[515][17] = (mid_1[4135:4128] < btm_0[4127:4120]) ? 1 : 0;
assign detect_min[515][18] = (mid_1[4135:4128] < btm_0[4135:4128]) ? 1 : 0;
assign detect_min[515][19] = (mid_1[4135:4128] < btm_0[4143:4136]) ? 1 : 0;
assign detect_min[515][20] = (mid_1[4135:4128] < btm_1[4127:4120]) ? 1 : 0;
assign detect_min[515][21] = (mid_1[4135:4128] < btm_1[4135:4128]) ? 1 : 0;
assign detect_min[515][22] = (mid_1[4135:4128] < btm_1[4143:4136]) ? 1 : 0;
assign detect_min[515][23] = (mid_1[4135:4128] < btm_2[4127:4120]) ? 1 : 0;
assign detect_min[515][24] = (mid_1[4135:4128] < btm_2[4135:4128]) ? 1 : 0;
assign detect_min[515][25] = (mid_1[4135:4128] < btm_2[4143:4136]) ? 1 : 0;

assign detect_min[516][0] = (mid_1[4143:4136] < top_0[4135:4128]) ? 1 : 0;
assign detect_min[516][1] = (mid_1[4143:4136] < top_0[4143:4136]) ? 1 : 0;
assign detect_min[516][2] = (mid_1[4143:4136] < top_0[4151:4144]) ? 1 : 0;
assign detect_min[516][3] = (mid_1[4143:4136] < top_1[4135:4128]) ? 1 : 0;
assign detect_min[516][4] = (mid_1[4143:4136] < top_1[4143:4136]) ? 1 : 0;
assign detect_min[516][5] = (mid_1[4143:4136] < top_1[4151:4144]) ? 1 : 0;
assign detect_min[516][6] = (mid_1[4143:4136] < top_2[4135:4128]) ? 1 : 0;
assign detect_min[516][7] = (mid_1[4143:4136] < top_2[4143:4136]) ? 1 : 0;
assign detect_min[516][8] = (mid_1[4143:4136] < top_2[4151:4144]) ? 1 : 0;
assign detect_min[516][9] = (mid_1[4143:4136] < mid_0[4135:4128]) ? 1 : 0;
assign detect_min[516][10] = (mid_1[4143:4136] < mid_0[4143:4136]) ? 1 : 0;
assign detect_min[516][11] = (mid_1[4143:4136] < mid_0[4151:4144]) ? 1 : 0;
assign detect_min[516][12] = (mid_1[4143:4136] < mid_1[4135:4128]) ? 1 : 0;
assign detect_min[516][13] = (mid_1[4143:4136] < mid_1[4151:4144]) ? 1 : 0;
assign detect_min[516][14] = (mid_1[4143:4136] < mid_2[4135:4128]) ? 1 : 0;
assign detect_min[516][15] = (mid_1[4143:4136] < mid_2[4143:4136]) ? 1 : 0;
assign detect_min[516][16] = (mid_1[4143:4136] < mid_2[4151:4144]) ? 1 : 0;
assign detect_min[516][17] = (mid_1[4143:4136] < btm_0[4135:4128]) ? 1 : 0;
assign detect_min[516][18] = (mid_1[4143:4136] < btm_0[4143:4136]) ? 1 : 0;
assign detect_min[516][19] = (mid_1[4143:4136] < btm_0[4151:4144]) ? 1 : 0;
assign detect_min[516][20] = (mid_1[4143:4136] < btm_1[4135:4128]) ? 1 : 0;
assign detect_min[516][21] = (mid_1[4143:4136] < btm_1[4143:4136]) ? 1 : 0;
assign detect_min[516][22] = (mid_1[4143:4136] < btm_1[4151:4144]) ? 1 : 0;
assign detect_min[516][23] = (mid_1[4143:4136] < btm_2[4135:4128]) ? 1 : 0;
assign detect_min[516][24] = (mid_1[4143:4136] < btm_2[4143:4136]) ? 1 : 0;
assign detect_min[516][25] = (mid_1[4143:4136] < btm_2[4151:4144]) ? 1 : 0;

assign detect_min[517][0] = (mid_1[4151:4144] < top_0[4143:4136]) ? 1 : 0;
assign detect_min[517][1] = (mid_1[4151:4144] < top_0[4151:4144]) ? 1 : 0;
assign detect_min[517][2] = (mid_1[4151:4144] < top_0[4159:4152]) ? 1 : 0;
assign detect_min[517][3] = (mid_1[4151:4144] < top_1[4143:4136]) ? 1 : 0;
assign detect_min[517][4] = (mid_1[4151:4144] < top_1[4151:4144]) ? 1 : 0;
assign detect_min[517][5] = (mid_1[4151:4144] < top_1[4159:4152]) ? 1 : 0;
assign detect_min[517][6] = (mid_1[4151:4144] < top_2[4143:4136]) ? 1 : 0;
assign detect_min[517][7] = (mid_1[4151:4144] < top_2[4151:4144]) ? 1 : 0;
assign detect_min[517][8] = (mid_1[4151:4144] < top_2[4159:4152]) ? 1 : 0;
assign detect_min[517][9] = (mid_1[4151:4144] < mid_0[4143:4136]) ? 1 : 0;
assign detect_min[517][10] = (mid_1[4151:4144] < mid_0[4151:4144]) ? 1 : 0;
assign detect_min[517][11] = (mid_1[4151:4144] < mid_0[4159:4152]) ? 1 : 0;
assign detect_min[517][12] = (mid_1[4151:4144] < mid_1[4143:4136]) ? 1 : 0;
assign detect_min[517][13] = (mid_1[4151:4144] < mid_1[4159:4152]) ? 1 : 0;
assign detect_min[517][14] = (mid_1[4151:4144] < mid_2[4143:4136]) ? 1 : 0;
assign detect_min[517][15] = (mid_1[4151:4144] < mid_2[4151:4144]) ? 1 : 0;
assign detect_min[517][16] = (mid_1[4151:4144] < mid_2[4159:4152]) ? 1 : 0;
assign detect_min[517][17] = (mid_1[4151:4144] < btm_0[4143:4136]) ? 1 : 0;
assign detect_min[517][18] = (mid_1[4151:4144] < btm_0[4151:4144]) ? 1 : 0;
assign detect_min[517][19] = (mid_1[4151:4144] < btm_0[4159:4152]) ? 1 : 0;
assign detect_min[517][20] = (mid_1[4151:4144] < btm_1[4143:4136]) ? 1 : 0;
assign detect_min[517][21] = (mid_1[4151:4144] < btm_1[4151:4144]) ? 1 : 0;
assign detect_min[517][22] = (mid_1[4151:4144] < btm_1[4159:4152]) ? 1 : 0;
assign detect_min[517][23] = (mid_1[4151:4144] < btm_2[4143:4136]) ? 1 : 0;
assign detect_min[517][24] = (mid_1[4151:4144] < btm_2[4151:4144]) ? 1 : 0;
assign detect_min[517][25] = (mid_1[4151:4144] < btm_2[4159:4152]) ? 1 : 0;

assign detect_min[518][0] = (mid_1[4159:4152] < top_0[4151:4144]) ? 1 : 0;
assign detect_min[518][1] = (mid_1[4159:4152] < top_0[4159:4152]) ? 1 : 0;
assign detect_min[518][2] = (mid_1[4159:4152] < top_0[4167:4160]) ? 1 : 0;
assign detect_min[518][3] = (mid_1[4159:4152] < top_1[4151:4144]) ? 1 : 0;
assign detect_min[518][4] = (mid_1[4159:4152] < top_1[4159:4152]) ? 1 : 0;
assign detect_min[518][5] = (mid_1[4159:4152] < top_1[4167:4160]) ? 1 : 0;
assign detect_min[518][6] = (mid_1[4159:4152] < top_2[4151:4144]) ? 1 : 0;
assign detect_min[518][7] = (mid_1[4159:4152] < top_2[4159:4152]) ? 1 : 0;
assign detect_min[518][8] = (mid_1[4159:4152] < top_2[4167:4160]) ? 1 : 0;
assign detect_min[518][9] = (mid_1[4159:4152] < mid_0[4151:4144]) ? 1 : 0;
assign detect_min[518][10] = (mid_1[4159:4152] < mid_0[4159:4152]) ? 1 : 0;
assign detect_min[518][11] = (mid_1[4159:4152] < mid_0[4167:4160]) ? 1 : 0;
assign detect_min[518][12] = (mid_1[4159:4152] < mid_1[4151:4144]) ? 1 : 0;
assign detect_min[518][13] = (mid_1[4159:4152] < mid_1[4167:4160]) ? 1 : 0;
assign detect_min[518][14] = (mid_1[4159:4152] < mid_2[4151:4144]) ? 1 : 0;
assign detect_min[518][15] = (mid_1[4159:4152] < mid_2[4159:4152]) ? 1 : 0;
assign detect_min[518][16] = (mid_1[4159:4152] < mid_2[4167:4160]) ? 1 : 0;
assign detect_min[518][17] = (mid_1[4159:4152] < btm_0[4151:4144]) ? 1 : 0;
assign detect_min[518][18] = (mid_1[4159:4152] < btm_0[4159:4152]) ? 1 : 0;
assign detect_min[518][19] = (mid_1[4159:4152] < btm_0[4167:4160]) ? 1 : 0;
assign detect_min[518][20] = (mid_1[4159:4152] < btm_1[4151:4144]) ? 1 : 0;
assign detect_min[518][21] = (mid_1[4159:4152] < btm_1[4159:4152]) ? 1 : 0;
assign detect_min[518][22] = (mid_1[4159:4152] < btm_1[4167:4160]) ? 1 : 0;
assign detect_min[518][23] = (mid_1[4159:4152] < btm_2[4151:4144]) ? 1 : 0;
assign detect_min[518][24] = (mid_1[4159:4152] < btm_2[4159:4152]) ? 1 : 0;
assign detect_min[518][25] = (mid_1[4159:4152] < btm_2[4167:4160]) ? 1 : 0;

assign detect_min[519][0] = (mid_1[4167:4160] < top_0[4159:4152]) ? 1 : 0;
assign detect_min[519][1] = (mid_1[4167:4160] < top_0[4167:4160]) ? 1 : 0;
assign detect_min[519][2] = (mid_1[4167:4160] < top_0[4175:4168]) ? 1 : 0;
assign detect_min[519][3] = (mid_1[4167:4160] < top_1[4159:4152]) ? 1 : 0;
assign detect_min[519][4] = (mid_1[4167:4160] < top_1[4167:4160]) ? 1 : 0;
assign detect_min[519][5] = (mid_1[4167:4160] < top_1[4175:4168]) ? 1 : 0;
assign detect_min[519][6] = (mid_1[4167:4160] < top_2[4159:4152]) ? 1 : 0;
assign detect_min[519][7] = (mid_1[4167:4160] < top_2[4167:4160]) ? 1 : 0;
assign detect_min[519][8] = (mid_1[4167:4160] < top_2[4175:4168]) ? 1 : 0;
assign detect_min[519][9] = (mid_1[4167:4160] < mid_0[4159:4152]) ? 1 : 0;
assign detect_min[519][10] = (mid_1[4167:4160] < mid_0[4167:4160]) ? 1 : 0;
assign detect_min[519][11] = (mid_1[4167:4160] < mid_0[4175:4168]) ? 1 : 0;
assign detect_min[519][12] = (mid_1[4167:4160] < mid_1[4159:4152]) ? 1 : 0;
assign detect_min[519][13] = (mid_1[4167:4160] < mid_1[4175:4168]) ? 1 : 0;
assign detect_min[519][14] = (mid_1[4167:4160] < mid_2[4159:4152]) ? 1 : 0;
assign detect_min[519][15] = (mid_1[4167:4160] < mid_2[4167:4160]) ? 1 : 0;
assign detect_min[519][16] = (mid_1[4167:4160] < mid_2[4175:4168]) ? 1 : 0;
assign detect_min[519][17] = (mid_1[4167:4160] < btm_0[4159:4152]) ? 1 : 0;
assign detect_min[519][18] = (mid_1[4167:4160] < btm_0[4167:4160]) ? 1 : 0;
assign detect_min[519][19] = (mid_1[4167:4160] < btm_0[4175:4168]) ? 1 : 0;
assign detect_min[519][20] = (mid_1[4167:4160] < btm_1[4159:4152]) ? 1 : 0;
assign detect_min[519][21] = (mid_1[4167:4160] < btm_1[4167:4160]) ? 1 : 0;
assign detect_min[519][22] = (mid_1[4167:4160] < btm_1[4175:4168]) ? 1 : 0;
assign detect_min[519][23] = (mid_1[4167:4160] < btm_2[4159:4152]) ? 1 : 0;
assign detect_min[519][24] = (mid_1[4167:4160] < btm_2[4167:4160]) ? 1 : 0;
assign detect_min[519][25] = (mid_1[4167:4160] < btm_2[4175:4168]) ? 1 : 0;

assign detect_min[520][0] = (mid_1[4175:4168] < top_0[4167:4160]) ? 1 : 0;
assign detect_min[520][1] = (mid_1[4175:4168] < top_0[4175:4168]) ? 1 : 0;
assign detect_min[520][2] = (mid_1[4175:4168] < top_0[4183:4176]) ? 1 : 0;
assign detect_min[520][3] = (mid_1[4175:4168] < top_1[4167:4160]) ? 1 : 0;
assign detect_min[520][4] = (mid_1[4175:4168] < top_1[4175:4168]) ? 1 : 0;
assign detect_min[520][5] = (mid_1[4175:4168] < top_1[4183:4176]) ? 1 : 0;
assign detect_min[520][6] = (mid_1[4175:4168] < top_2[4167:4160]) ? 1 : 0;
assign detect_min[520][7] = (mid_1[4175:4168] < top_2[4175:4168]) ? 1 : 0;
assign detect_min[520][8] = (mid_1[4175:4168] < top_2[4183:4176]) ? 1 : 0;
assign detect_min[520][9] = (mid_1[4175:4168] < mid_0[4167:4160]) ? 1 : 0;
assign detect_min[520][10] = (mid_1[4175:4168] < mid_0[4175:4168]) ? 1 : 0;
assign detect_min[520][11] = (mid_1[4175:4168] < mid_0[4183:4176]) ? 1 : 0;
assign detect_min[520][12] = (mid_1[4175:4168] < mid_1[4167:4160]) ? 1 : 0;
assign detect_min[520][13] = (mid_1[4175:4168] < mid_1[4183:4176]) ? 1 : 0;
assign detect_min[520][14] = (mid_1[4175:4168] < mid_2[4167:4160]) ? 1 : 0;
assign detect_min[520][15] = (mid_1[4175:4168] < mid_2[4175:4168]) ? 1 : 0;
assign detect_min[520][16] = (mid_1[4175:4168] < mid_2[4183:4176]) ? 1 : 0;
assign detect_min[520][17] = (mid_1[4175:4168] < btm_0[4167:4160]) ? 1 : 0;
assign detect_min[520][18] = (mid_1[4175:4168] < btm_0[4175:4168]) ? 1 : 0;
assign detect_min[520][19] = (mid_1[4175:4168] < btm_0[4183:4176]) ? 1 : 0;
assign detect_min[520][20] = (mid_1[4175:4168] < btm_1[4167:4160]) ? 1 : 0;
assign detect_min[520][21] = (mid_1[4175:4168] < btm_1[4175:4168]) ? 1 : 0;
assign detect_min[520][22] = (mid_1[4175:4168] < btm_1[4183:4176]) ? 1 : 0;
assign detect_min[520][23] = (mid_1[4175:4168] < btm_2[4167:4160]) ? 1 : 0;
assign detect_min[520][24] = (mid_1[4175:4168] < btm_2[4175:4168]) ? 1 : 0;
assign detect_min[520][25] = (mid_1[4175:4168] < btm_2[4183:4176]) ? 1 : 0;

assign detect_min[521][0] = (mid_1[4183:4176] < top_0[4175:4168]) ? 1 : 0;
assign detect_min[521][1] = (mid_1[4183:4176] < top_0[4183:4176]) ? 1 : 0;
assign detect_min[521][2] = (mid_1[4183:4176] < top_0[4191:4184]) ? 1 : 0;
assign detect_min[521][3] = (mid_1[4183:4176] < top_1[4175:4168]) ? 1 : 0;
assign detect_min[521][4] = (mid_1[4183:4176] < top_1[4183:4176]) ? 1 : 0;
assign detect_min[521][5] = (mid_1[4183:4176] < top_1[4191:4184]) ? 1 : 0;
assign detect_min[521][6] = (mid_1[4183:4176] < top_2[4175:4168]) ? 1 : 0;
assign detect_min[521][7] = (mid_1[4183:4176] < top_2[4183:4176]) ? 1 : 0;
assign detect_min[521][8] = (mid_1[4183:4176] < top_2[4191:4184]) ? 1 : 0;
assign detect_min[521][9] = (mid_1[4183:4176] < mid_0[4175:4168]) ? 1 : 0;
assign detect_min[521][10] = (mid_1[4183:4176] < mid_0[4183:4176]) ? 1 : 0;
assign detect_min[521][11] = (mid_1[4183:4176] < mid_0[4191:4184]) ? 1 : 0;
assign detect_min[521][12] = (mid_1[4183:4176] < mid_1[4175:4168]) ? 1 : 0;
assign detect_min[521][13] = (mid_1[4183:4176] < mid_1[4191:4184]) ? 1 : 0;
assign detect_min[521][14] = (mid_1[4183:4176] < mid_2[4175:4168]) ? 1 : 0;
assign detect_min[521][15] = (mid_1[4183:4176] < mid_2[4183:4176]) ? 1 : 0;
assign detect_min[521][16] = (mid_1[4183:4176] < mid_2[4191:4184]) ? 1 : 0;
assign detect_min[521][17] = (mid_1[4183:4176] < btm_0[4175:4168]) ? 1 : 0;
assign detect_min[521][18] = (mid_1[4183:4176] < btm_0[4183:4176]) ? 1 : 0;
assign detect_min[521][19] = (mid_1[4183:4176] < btm_0[4191:4184]) ? 1 : 0;
assign detect_min[521][20] = (mid_1[4183:4176] < btm_1[4175:4168]) ? 1 : 0;
assign detect_min[521][21] = (mid_1[4183:4176] < btm_1[4183:4176]) ? 1 : 0;
assign detect_min[521][22] = (mid_1[4183:4176] < btm_1[4191:4184]) ? 1 : 0;
assign detect_min[521][23] = (mid_1[4183:4176] < btm_2[4175:4168]) ? 1 : 0;
assign detect_min[521][24] = (mid_1[4183:4176] < btm_2[4183:4176]) ? 1 : 0;
assign detect_min[521][25] = (mid_1[4183:4176] < btm_2[4191:4184]) ? 1 : 0;

assign detect_min[522][0] = (mid_1[4191:4184] < top_0[4183:4176]) ? 1 : 0;
assign detect_min[522][1] = (mid_1[4191:4184] < top_0[4191:4184]) ? 1 : 0;
assign detect_min[522][2] = (mid_1[4191:4184] < top_0[4199:4192]) ? 1 : 0;
assign detect_min[522][3] = (mid_1[4191:4184] < top_1[4183:4176]) ? 1 : 0;
assign detect_min[522][4] = (mid_1[4191:4184] < top_1[4191:4184]) ? 1 : 0;
assign detect_min[522][5] = (mid_1[4191:4184] < top_1[4199:4192]) ? 1 : 0;
assign detect_min[522][6] = (mid_1[4191:4184] < top_2[4183:4176]) ? 1 : 0;
assign detect_min[522][7] = (mid_1[4191:4184] < top_2[4191:4184]) ? 1 : 0;
assign detect_min[522][8] = (mid_1[4191:4184] < top_2[4199:4192]) ? 1 : 0;
assign detect_min[522][9] = (mid_1[4191:4184] < mid_0[4183:4176]) ? 1 : 0;
assign detect_min[522][10] = (mid_1[4191:4184] < mid_0[4191:4184]) ? 1 : 0;
assign detect_min[522][11] = (mid_1[4191:4184] < mid_0[4199:4192]) ? 1 : 0;
assign detect_min[522][12] = (mid_1[4191:4184] < mid_1[4183:4176]) ? 1 : 0;
assign detect_min[522][13] = (mid_1[4191:4184] < mid_1[4199:4192]) ? 1 : 0;
assign detect_min[522][14] = (mid_1[4191:4184] < mid_2[4183:4176]) ? 1 : 0;
assign detect_min[522][15] = (mid_1[4191:4184] < mid_2[4191:4184]) ? 1 : 0;
assign detect_min[522][16] = (mid_1[4191:4184] < mid_2[4199:4192]) ? 1 : 0;
assign detect_min[522][17] = (mid_1[4191:4184] < btm_0[4183:4176]) ? 1 : 0;
assign detect_min[522][18] = (mid_1[4191:4184] < btm_0[4191:4184]) ? 1 : 0;
assign detect_min[522][19] = (mid_1[4191:4184] < btm_0[4199:4192]) ? 1 : 0;
assign detect_min[522][20] = (mid_1[4191:4184] < btm_1[4183:4176]) ? 1 : 0;
assign detect_min[522][21] = (mid_1[4191:4184] < btm_1[4191:4184]) ? 1 : 0;
assign detect_min[522][22] = (mid_1[4191:4184] < btm_1[4199:4192]) ? 1 : 0;
assign detect_min[522][23] = (mid_1[4191:4184] < btm_2[4183:4176]) ? 1 : 0;
assign detect_min[522][24] = (mid_1[4191:4184] < btm_2[4191:4184]) ? 1 : 0;
assign detect_min[522][25] = (mid_1[4191:4184] < btm_2[4199:4192]) ? 1 : 0;

assign detect_min[523][0] = (mid_1[4199:4192] < top_0[4191:4184]) ? 1 : 0;
assign detect_min[523][1] = (mid_1[4199:4192] < top_0[4199:4192]) ? 1 : 0;
assign detect_min[523][2] = (mid_1[4199:4192] < top_0[4207:4200]) ? 1 : 0;
assign detect_min[523][3] = (mid_1[4199:4192] < top_1[4191:4184]) ? 1 : 0;
assign detect_min[523][4] = (mid_1[4199:4192] < top_1[4199:4192]) ? 1 : 0;
assign detect_min[523][5] = (mid_1[4199:4192] < top_1[4207:4200]) ? 1 : 0;
assign detect_min[523][6] = (mid_1[4199:4192] < top_2[4191:4184]) ? 1 : 0;
assign detect_min[523][7] = (mid_1[4199:4192] < top_2[4199:4192]) ? 1 : 0;
assign detect_min[523][8] = (mid_1[4199:4192] < top_2[4207:4200]) ? 1 : 0;
assign detect_min[523][9] = (mid_1[4199:4192] < mid_0[4191:4184]) ? 1 : 0;
assign detect_min[523][10] = (mid_1[4199:4192] < mid_0[4199:4192]) ? 1 : 0;
assign detect_min[523][11] = (mid_1[4199:4192] < mid_0[4207:4200]) ? 1 : 0;
assign detect_min[523][12] = (mid_1[4199:4192] < mid_1[4191:4184]) ? 1 : 0;
assign detect_min[523][13] = (mid_1[4199:4192] < mid_1[4207:4200]) ? 1 : 0;
assign detect_min[523][14] = (mid_1[4199:4192] < mid_2[4191:4184]) ? 1 : 0;
assign detect_min[523][15] = (mid_1[4199:4192] < mid_2[4199:4192]) ? 1 : 0;
assign detect_min[523][16] = (mid_1[4199:4192] < mid_2[4207:4200]) ? 1 : 0;
assign detect_min[523][17] = (mid_1[4199:4192] < btm_0[4191:4184]) ? 1 : 0;
assign detect_min[523][18] = (mid_1[4199:4192] < btm_0[4199:4192]) ? 1 : 0;
assign detect_min[523][19] = (mid_1[4199:4192] < btm_0[4207:4200]) ? 1 : 0;
assign detect_min[523][20] = (mid_1[4199:4192] < btm_1[4191:4184]) ? 1 : 0;
assign detect_min[523][21] = (mid_1[4199:4192] < btm_1[4199:4192]) ? 1 : 0;
assign detect_min[523][22] = (mid_1[4199:4192] < btm_1[4207:4200]) ? 1 : 0;
assign detect_min[523][23] = (mid_1[4199:4192] < btm_2[4191:4184]) ? 1 : 0;
assign detect_min[523][24] = (mid_1[4199:4192] < btm_2[4199:4192]) ? 1 : 0;
assign detect_min[523][25] = (mid_1[4199:4192] < btm_2[4207:4200]) ? 1 : 0;

assign detect_min[524][0] = (mid_1[4207:4200] < top_0[4199:4192]) ? 1 : 0;
assign detect_min[524][1] = (mid_1[4207:4200] < top_0[4207:4200]) ? 1 : 0;
assign detect_min[524][2] = (mid_1[4207:4200] < top_0[4215:4208]) ? 1 : 0;
assign detect_min[524][3] = (mid_1[4207:4200] < top_1[4199:4192]) ? 1 : 0;
assign detect_min[524][4] = (mid_1[4207:4200] < top_1[4207:4200]) ? 1 : 0;
assign detect_min[524][5] = (mid_1[4207:4200] < top_1[4215:4208]) ? 1 : 0;
assign detect_min[524][6] = (mid_1[4207:4200] < top_2[4199:4192]) ? 1 : 0;
assign detect_min[524][7] = (mid_1[4207:4200] < top_2[4207:4200]) ? 1 : 0;
assign detect_min[524][8] = (mid_1[4207:4200] < top_2[4215:4208]) ? 1 : 0;
assign detect_min[524][9] = (mid_1[4207:4200] < mid_0[4199:4192]) ? 1 : 0;
assign detect_min[524][10] = (mid_1[4207:4200] < mid_0[4207:4200]) ? 1 : 0;
assign detect_min[524][11] = (mid_1[4207:4200] < mid_0[4215:4208]) ? 1 : 0;
assign detect_min[524][12] = (mid_1[4207:4200] < mid_1[4199:4192]) ? 1 : 0;
assign detect_min[524][13] = (mid_1[4207:4200] < mid_1[4215:4208]) ? 1 : 0;
assign detect_min[524][14] = (mid_1[4207:4200] < mid_2[4199:4192]) ? 1 : 0;
assign detect_min[524][15] = (mid_1[4207:4200] < mid_2[4207:4200]) ? 1 : 0;
assign detect_min[524][16] = (mid_1[4207:4200] < mid_2[4215:4208]) ? 1 : 0;
assign detect_min[524][17] = (mid_1[4207:4200] < btm_0[4199:4192]) ? 1 : 0;
assign detect_min[524][18] = (mid_1[4207:4200] < btm_0[4207:4200]) ? 1 : 0;
assign detect_min[524][19] = (mid_1[4207:4200] < btm_0[4215:4208]) ? 1 : 0;
assign detect_min[524][20] = (mid_1[4207:4200] < btm_1[4199:4192]) ? 1 : 0;
assign detect_min[524][21] = (mid_1[4207:4200] < btm_1[4207:4200]) ? 1 : 0;
assign detect_min[524][22] = (mid_1[4207:4200] < btm_1[4215:4208]) ? 1 : 0;
assign detect_min[524][23] = (mid_1[4207:4200] < btm_2[4199:4192]) ? 1 : 0;
assign detect_min[524][24] = (mid_1[4207:4200] < btm_2[4207:4200]) ? 1 : 0;
assign detect_min[524][25] = (mid_1[4207:4200] < btm_2[4215:4208]) ? 1 : 0;

assign detect_min[525][0] = (mid_1[4215:4208] < top_0[4207:4200]) ? 1 : 0;
assign detect_min[525][1] = (mid_1[4215:4208] < top_0[4215:4208]) ? 1 : 0;
assign detect_min[525][2] = (mid_1[4215:4208] < top_0[4223:4216]) ? 1 : 0;
assign detect_min[525][3] = (mid_1[4215:4208] < top_1[4207:4200]) ? 1 : 0;
assign detect_min[525][4] = (mid_1[4215:4208] < top_1[4215:4208]) ? 1 : 0;
assign detect_min[525][5] = (mid_1[4215:4208] < top_1[4223:4216]) ? 1 : 0;
assign detect_min[525][6] = (mid_1[4215:4208] < top_2[4207:4200]) ? 1 : 0;
assign detect_min[525][7] = (mid_1[4215:4208] < top_2[4215:4208]) ? 1 : 0;
assign detect_min[525][8] = (mid_1[4215:4208] < top_2[4223:4216]) ? 1 : 0;
assign detect_min[525][9] = (mid_1[4215:4208] < mid_0[4207:4200]) ? 1 : 0;
assign detect_min[525][10] = (mid_1[4215:4208] < mid_0[4215:4208]) ? 1 : 0;
assign detect_min[525][11] = (mid_1[4215:4208] < mid_0[4223:4216]) ? 1 : 0;
assign detect_min[525][12] = (mid_1[4215:4208] < mid_1[4207:4200]) ? 1 : 0;
assign detect_min[525][13] = (mid_1[4215:4208] < mid_1[4223:4216]) ? 1 : 0;
assign detect_min[525][14] = (mid_1[4215:4208] < mid_2[4207:4200]) ? 1 : 0;
assign detect_min[525][15] = (mid_1[4215:4208] < mid_2[4215:4208]) ? 1 : 0;
assign detect_min[525][16] = (mid_1[4215:4208] < mid_2[4223:4216]) ? 1 : 0;
assign detect_min[525][17] = (mid_1[4215:4208] < btm_0[4207:4200]) ? 1 : 0;
assign detect_min[525][18] = (mid_1[4215:4208] < btm_0[4215:4208]) ? 1 : 0;
assign detect_min[525][19] = (mid_1[4215:4208] < btm_0[4223:4216]) ? 1 : 0;
assign detect_min[525][20] = (mid_1[4215:4208] < btm_1[4207:4200]) ? 1 : 0;
assign detect_min[525][21] = (mid_1[4215:4208] < btm_1[4215:4208]) ? 1 : 0;
assign detect_min[525][22] = (mid_1[4215:4208] < btm_1[4223:4216]) ? 1 : 0;
assign detect_min[525][23] = (mid_1[4215:4208] < btm_2[4207:4200]) ? 1 : 0;
assign detect_min[525][24] = (mid_1[4215:4208] < btm_2[4215:4208]) ? 1 : 0;
assign detect_min[525][25] = (mid_1[4215:4208] < btm_2[4223:4216]) ? 1 : 0;

assign detect_min[526][0] = (mid_1[4223:4216] < top_0[4215:4208]) ? 1 : 0;
assign detect_min[526][1] = (mid_1[4223:4216] < top_0[4223:4216]) ? 1 : 0;
assign detect_min[526][2] = (mid_1[4223:4216] < top_0[4231:4224]) ? 1 : 0;
assign detect_min[526][3] = (mid_1[4223:4216] < top_1[4215:4208]) ? 1 : 0;
assign detect_min[526][4] = (mid_1[4223:4216] < top_1[4223:4216]) ? 1 : 0;
assign detect_min[526][5] = (mid_1[4223:4216] < top_1[4231:4224]) ? 1 : 0;
assign detect_min[526][6] = (mid_1[4223:4216] < top_2[4215:4208]) ? 1 : 0;
assign detect_min[526][7] = (mid_1[4223:4216] < top_2[4223:4216]) ? 1 : 0;
assign detect_min[526][8] = (mid_1[4223:4216] < top_2[4231:4224]) ? 1 : 0;
assign detect_min[526][9] = (mid_1[4223:4216] < mid_0[4215:4208]) ? 1 : 0;
assign detect_min[526][10] = (mid_1[4223:4216] < mid_0[4223:4216]) ? 1 : 0;
assign detect_min[526][11] = (mid_1[4223:4216] < mid_0[4231:4224]) ? 1 : 0;
assign detect_min[526][12] = (mid_1[4223:4216] < mid_1[4215:4208]) ? 1 : 0;
assign detect_min[526][13] = (mid_1[4223:4216] < mid_1[4231:4224]) ? 1 : 0;
assign detect_min[526][14] = (mid_1[4223:4216] < mid_2[4215:4208]) ? 1 : 0;
assign detect_min[526][15] = (mid_1[4223:4216] < mid_2[4223:4216]) ? 1 : 0;
assign detect_min[526][16] = (mid_1[4223:4216] < mid_2[4231:4224]) ? 1 : 0;
assign detect_min[526][17] = (mid_1[4223:4216] < btm_0[4215:4208]) ? 1 : 0;
assign detect_min[526][18] = (mid_1[4223:4216] < btm_0[4223:4216]) ? 1 : 0;
assign detect_min[526][19] = (mid_1[4223:4216] < btm_0[4231:4224]) ? 1 : 0;
assign detect_min[526][20] = (mid_1[4223:4216] < btm_1[4215:4208]) ? 1 : 0;
assign detect_min[526][21] = (mid_1[4223:4216] < btm_1[4223:4216]) ? 1 : 0;
assign detect_min[526][22] = (mid_1[4223:4216] < btm_1[4231:4224]) ? 1 : 0;
assign detect_min[526][23] = (mid_1[4223:4216] < btm_2[4215:4208]) ? 1 : 0;
assign detect_min[526][24] = (mid_1[4223:4216] < btm_2[4223:4216]) ? 1 : 0;
assign detect_min[526][25] = (mid_1[4223:4216] < btm_2[4231:4224]) ? 1 : 0;

assign detect_min[527][0] = (mid_1[4231:4224] < top_0[4223:4216]) ? 1 : 0;
assign detect_min[527][1] = (mid_1[4231:4224] < top_0[4231:4224]) ? 1 : 0;
assign detect_min[527][2] = (mid_1[4231:4224] < top_0[4239:4232]) ? 1 : 0;
assign detect_min[527][3] = (mid_1[4231:4224] < top_1[4223:4216]) ? 1 : 0;
assign detect_min[527][4] = (mid_1[4231:4224] < top_1[4231:4224]) ? 1 : 0;
assign detect_min[527][5] = (mid_1[4231:4224] < top_1[4239:4232]) ? 1 : 0;
assign detect_min[527][6] = (mid_1[4231:4224] < top_2[4223:4216]) ? 1 : 0;
assign detect_min[527][7] = (mid_1[4231:4224] < top_2[4231:4224]) ? 1 : 0;
assign detect_min[527][8] = (mid_1[4231:4224] < top_2[4239:4232]) ? 1 : 0;
assign detect_min[527][9] = (mid_1[4231:4224] < mid_0[4223:4216]) ? 1 : 0;
assign detect_min[527][10] = (mid_1[4231:4224] < mid_0[4231:4224]) ? 1 : 0;
assign detect_min[527][11] = (mid_1[4231:4224] < mid_0[4239:4232]) ? 1 : 0;
assign detect_min[527][12] = (mid_1[4231:4224] < mid_1[4223:4216]) ? 1 : 0;
assign detect_min[527][13] = (mid_1[4231:4224] < mid_1[4239:4232]) ? 1 : 0;
assign detect_min[527][14] = (mid_1[4231:4224] < mid_2[4223:4216]) ? 1 : 0;
assign detect_min[527][15] = (mid_1[4231:4224] < mid_2[4231:4224]) ? 1 : 0;
assign detect_min[527][16] = (mid_1[4231:4224] < mid_2[4239:4232]) ? 1 : 0;
assign detect_min[527][17] = (mid_1[4231:4224] < btm_0[4223:4216]) ? 1 : 0;
assign detect_min[527][18] = (mid_1[4231:4224] < btm_0[4231:4224]) ? 1 : 0;
assign detect_min[527][19] = (mid_1[4231:4224] < btm_0[4239:4232]) ? 1 : 0;
assign detect_min[527][20] = (mid_1[4231:4224] < btm_1[4223:4216]) ? 1 : 0;
assign detect_min[527][21] = (mid_1[4231:4224] < btm_1[4231:4224]) ? 1 : 0;
assign detect_min[527][22] = (mid_1[4231:4224] < btm_1[4239:4232]) ? 1 : 0;
assign detect_min[527][23] = (mid_1[4231:4224] < btm_2[4223:4216]) ? 1 : 0;
assign detect_min[527][24] = (mid_1[4231:4224] < btm_2[4231:4224]) ? 1 : 0;
assign detect_min[527][25] = (mid_1[4231:4224] < btm_2[4239:4232]) ? 1 : 0;

assign detect_min[528][0] = (mid_1[4239:4232] < top_0[4231:4224]) ? 1 : 0;
assign detect_min[528][1] = (mid_1[4239:4232] < top_0[4239:4232]) ? 1 : 0;
assign detect_min[528][2] = (mid_1[4239:4232] < top_0[4247:4240]) ? 1 : 0;
assign detect_min[528][3] = (mid_1[4239:4232] < top_1[4231:4224]) ? 1 : 0;
assign detect_min[528][4] = (mid_1[4239:4232] < top_1[4239:4232]) ? 1 : 0;
assign detect_min[528][5] = (mid_1[4239:4232] < top_1[4247:4240]) ? 1 : 0;
assign detect_min[528][6] = (mid_1[4239:4232] < top_2[4231:4224]) ? 1 : 0;
assign detect_min[528][7] = (mid_1[4239:4232] < top_2[4239:4232]) ? 1 : 0;
assign detect_min[528][8] = (mid_1[4239:4232] < top_2[4247:4240]) ? 1 : 0;
assign detect_min[528][9] = (mid_1[4239:4232] < mid_0[4231:4224]) ? 1 : 0;
assign detect_min[528][10] = (mid_1[4239:4232] < mid_0[4239:4232]) ? 1 : 0;
assign detect_min[528][11] = (mid_1[4239:4232] < mid_0[4247:4240]) ? 1 : 0;
assign detect_min[528][12] = (mid_1[4239:4232] < mid_1[4231:4224]) ? 1 : 0;
assign detect_min[528][13] = (mid_1[4239:4232] < mid_1[4247:4240]) ? 1 : 0;
assign detect_min[528][14] = (mid_1[4239:4232] < mid_2[4231:4224]) ? 1 : 0;
assign detect_min[528][15] = (mid_1[4239:4232] < mid_2[4239:4232]) ? 1 : 0;
assign detect_min[528][16] = (mid_1[4239:4232] < mid_2[4247:4240]) ? 1 : 0;
assign detect_min[528][17] = (mid_1[4239:4232] < btm_0[4231:4224]) ? 1 : 0;
assign detect_min[528][18] = (mid_1[4239:4232] < btm_0[4239:4232]) ? 1 : 0;
assign detect_min[528][19] = (mid_1[4239:4232] < btm_0[4247:4240]) ? 1 : 0;
assign detect_min[528][20] = (mid_1[4239:4232] < btm_1[4231:4224]) ? 1 : 0;
assign detect_min[528][21] = (mid_1[4239:4232] < btm_1[4239:4232]) ? 1 : 0;
assign detect_min[528][22] = (mid_1[4239:4232] < btm_1[4247:4240]) ? 1 : 0;
assign detect_min[528][23] = (mid_1[4239:4232] < btm_2[4231:4224]) ? 1 : 0;
assign detect_min[528][24] = (mid_1[4239:4232] < btm_2[4239:4232]) ? 1 : 0;
assign detect_min[528][25] = (mid_1[4239:4232] < btm_2[4247:4240]) ? 1 : 0;

assign detect_min[529][0] = (mid_1[4247:4240] < top_0[4239:4232]) ? 1 : 0;
assign detect_min[529][1] = (mid_1[4247:4240] < top_0[4247:4240]) ? 1 : 0;
assign detect_min[529][2] = (mid_1[4247:4240] < top_0[4255:4248]) ? 1 : 0;
assign detect_min[529][3] = (mid_1[4247:4240] < top_1[4239:4232]) ? 1 : 0;
assign detect_min[529][4] = (mid_1[4247:4240] < top_1[4247:4240]) ? 1 : 0;
assign detect_min[529][5] = (mid_1[4247:4240] < top_1[4255:4248]) ? 1 : 0;
assign detect_min[529][6] = (mid_1[4247:4240] < top_2[4239:4232]) ? 1 : 0;
assign detect_min[529][7] = (mid_1[4247:4240] < top_2[4247:4240]) ? 1 : 0;
assign detect_min[529][8] = (mid_1[4247:4240] < top_2[4255:4248]) ? 1 : 0;
assign detect_min[529][9] = (mid_1[4247:4240] < mid_0[4239:4232]) ? 1 : 0;
assign detect_min[529][10] = (mid_1[4247:4240] < mid_0[4247:4240]) ? 1 : 0;
assign detect_min[529][11] = (mid_1[4247:4240] < mid_0[4255:4248]) ? 1 : 0;
assign detect_min[529][12] = (mid_1[4247:4240] < mid_1[4239:4232]) ? 1 : 0;
assign detect_min[529][13] = (mid_1[4247:4240] < mid_1[4255:4248]) ? 1 : 0;
assign detect_min[529][14] = (mid_1[4247:4240] < mid_2[4239:4232]) ? 1 : 0;
assign detect_min[529][15] = (mid_1[4247:4240] < mid_2[4247:4240]) ? 1 : 0;
assign detect_min[529][16] = (mid_1[4247:4240] < mid_2[4255:4248]) ? 1 : 0;
assign detect_min[529][17] = (mid_1[4247:4240] < btm_0[4239:4232]) ? 1 : 0;
assign detect_min[529][18] = (mid_1[4247:4240] < btm_0[4247:4240]) ? 1 : 0;
assign detect_min[529][19] = (mid_1[4247:4240] < btm_0[4255:4248]) ? 1 : 0;
assign detect_min[529][20] = (mid_1[4247:4240] < btm_1[4239:4232]) ? 1 : 0;
assign detect_min[529][21] = (mid_1[4247:4240] < btm_1[4247:4240]) ? 1 : 0;
assign detect_min[529][22] = (mid_1[4247:4240] < btm_1[4255:4248]) ? 1 : 0;
assign detect_min[529][23] = (mid_1[4247:4240] < btm_2[4239:4232]) ? 1 : 0;
assign detect_min[529][24] = (mid_1[4247:4240] < btm_2[4247:4240]) ? 1 : 0;
assign detect_min[529][25] = (mid_1[4247:4240] < btm_2[4255:4248]) ? 1 : 0;

assign detect_min[530][0] = (mid_1[4255:4248] < top_0[4247:4240]) ? 1 : 0;
assign detect_min[530][1] = (mid_1[4255:4248] < top_0[4255:4248]) ? 1 : 0;
assign detect_min[530][2] = (mid_1[4255:4248] < top_0[4263:4256]) ? 1 : 0;
assign detect_min[530][3] = (mid_1[4255:4248] < top_1[4247:4240]) ? 1 : 0;
assign detect_min[530][4] = (mid_1[4255:4248] < top_1[4255:4248]) ? 1 : 0;
assign detect_min[530][5] = (mid_1[4255:4248] < top_1[4263:4256]) ? 1 : 0;
assign detect_min[530][6] = (mid_1[4255:4248] < top_2[4247:4240]) ? 1 : 0;
assign detect_min[530][7] = (mid_1[4255:4248] < top_2[4255:4248]) ? 1 : 0;
assign detect_min[530][8] = (mid_1[4255:4248] < top_2[4263:4256]) ? 1 : 0;
assign detect_min[530][9] = (mid_1[4255:4248] < mid_0[4247:4240]) ? 1 : 0;
assign detect_min[530][10] = (mid_1[4255:4248] < mid_0[4255:4248]) ? 1 : 0;
assign detect_min[530][11] = (mid_1[4255:4248] < mid_0[4263:4256]) ? 1 : 0;
assign detect_min[530][12] = (mid_1[4255:4248] < mid_1[4247:4240]) ? 1 : 0;
assign detect_min[530][13] = (mid_1[4255:4248] < mid_1[4263:4256]) ? 1 : 0;
assign detect_min[530][14] = (mid_1[4255:4248] < mid_2[4247:4240]) ? 1 : 0;
assign detect_min[530][15] = (mid_1[4255:4248] < mid_2[4255:4248]) ? 1 : 0;
assign detect_min[530][16] = (mid_1[4255:4248] < mid_2[4263:4256]) ? 1 : 0;
assign detect_min[530][17] = (mid_1[4255:4248] < btm_0[4247:4240]) ? 1 : 0;
assign detect_min[530][18] = (mid_1[4255:4248] < btm_0[4255:4248]) ? 1 : 0;
assign detect_min[530][19] = (mid_1[4255:4248] < btm_0[4263:4256]) ? 1 : 0;
assign detect_min[530][20] = (mid_1[4255:4248] < btm_1[4247:4240]) ? 1 : 0;
assign detect_min[530][21] = (mid_1[4255:4248] < btm_1[4255:4248]) ? 1 : 0;
assign detect_min[530][22] = (mid_1[4255:4248] < btm_1[4263:4256]) ? 1 : 0;
assign detect_min[530][23] = (mid_1[4255:4248] < btm_2[4247:4240]) ? 1 : 0;
assign detect_min[530][24] = (mid_1[4255:4248] < btm_2[4255:4248]) ? 1 : 0;
assign detect_min[530][25] = (mid_1[4255:4248] < btm_2[4263:4256]) ? 1 : 0;

assign detect_min[531][0] = (mid_1[4263:4256] < top_0[4255:4248]) ? 1 : 0;
assign detect_min[531][1] = (mid_1[4263:4256] < top_0[4263:4256]) ? 1 : 0;
assign detect_min[531][2] = (mid_1[4263:4256] < top_0[4271:4264]) ? 1 : 0;
assign detect_min[531][3] = (mid_1[4263:4256] < top_1[4255:4248]) ? 1 : 0;
assign detect_min[531][4] = (mid_1[4263:4256] < top_1[4263:4256]) ? 1 : 0;
assign detect_min[531][5] = (mid_1[4263:4256] < top_1[4271:4264]) ? 1 : 0;
assign detect_min[531][6] = (mid_1[4263:4256] < top_2[4255:4248]) ? 1 : 0;
assign detect_min[531][7] = (mid_1[4263:4256] < top_2[4263:4256]) ? 1 : 0;
assign detect_min[531][8] = (mid_1[4263:4256] < top_2[4271:4264]) ? 1 : 0;
assign detect_min[531][9] = (mid_1[4263:4256] < mid_0[4255:4248]) ? 1 : 0;
assign detect_min[531][10] = (mid_1[4263:4256] < mid_0[4263:4256]) ? 1 : 0;
assign detect_min[531][11] = (mid_1[4263:4256] < mid_0[4271:4264]) ? 1 : 0;
assign detect_min[531][12] = (mid_1[4263:4256] < mid_1[4255:4248]) ? 1 : 0;
assign detect_min[531][13] = (mid_1[4263:4256] < mid_1[4271:4264]) ? 1 : 0;
assign detect_min[531][14] = (mid_1[4263:4256] < mid_2[4255:4248]) ? 1 : 0;
assign detect_min[531][15] = (mid_1[4263:4256] < mid_2[4263:4256]) ? 1 : 0;
assign detect_min[531][16] = (mid_1[4263:4256] < mid_2[4271:4264]) ? 1 : 0;
assign detect_min[531][17] = (mid_1[4263:4256] < btm_0[4255:4248]) ? 1 : 0;
assign detect_min[531][18] = (mid_1[4263:4256] < btm_0[4263:4256]) ? 1 : 0;
assign detect_min[531][19] = (mid_1[4263:4256] < btm_0[4271:4264]) ? 1 : 0;
assign detect_min[531][20] = (mid_1[4263:4256] < btm_1[4255:4248]) ? 1 : 0;
assign detect_min[531][21] = (mid_1[4263:4256] < btm_1[4263:4256]) ? 1 : 0;
assign detect_min[531][22] = (mid_1[4263:4256] < btm_1[4271:4264]) ? 1 : 0;
assign detect_min[531][23] = (mid_1[4263:4256] < btm_2[4255:4248]) ? 1 : 0;
assign detect_min[531][24] = (mid_1[4263:4256] < btm_2[4263:4256]) ? 1 : 0;
assign detect_min[531][25] = (mid_1[4263:4256] < btm_2[4271:4264]) ? 1 : 0;

assign detect_min[532][0] = (mid_1[4271:4264] < top_0[4263:4256]) ? 1 : 0;
assign detect_min[532][1] = (mid_1[4271:4264] < top_0[4271:4264]) ? 1 : 0;
assign detect_min[532][2] = (mid_1[4271:4264] < top_0[4279:4272]) ? 1 : 0;
assign detect_min[532][3] = (mid_1[4271:4264] < top_1[4263:4256]) ? 1 : 0;
assign detect_min[532][4] = (mid_1[4271:4264] < top_1[4271:4264]) ? 1 : 0;
assign detect_min[532][5] = (mid_1[4271:4264] < top_1[4279:4272]) ? 1 : 0;
assign detect_min[532][6] = (mid_1[4271:4264] < top_2[4263:4256]) ? 1 : 0;
assign detect_min[532][7] = (mid_1[4271:4264] < top_2[4271:4264]) ? 1 : 0;
assign detect_min[532][8] = (mid_1[4271:4264] < top_2[4279:4272]) ? 1 : 0;
assign detect_min[532][9] = (mid_1[4271:4264] < mid_0[4263:4256]) ? 1 : 0;
assign detect_min[532][10] = (mid_1[4271:4264] < mid_0[4271:4264]) ? 1 : 0;
assign detect_min[532][11] = (mid_1[4271:4264] < mid_0[4279:4272]) ? 1 : 0;
assign detect_min[532][12] = (mid_1[4271:4264] < mid_1[4263:4256]) ? 1 : 0;
assign detect_min[532][13] = (mid_1[4271:4264] < mid_1[4279:4272]) ? 1 : 0;
assign detect_min[532][14] = (mid_1[4271:4264] < mid_2[4263:4256]) ? 1 : 0;
assign detect_min[532][15] = (mid_1[4271:4264] < mid_2[4271:4264]) ? 1 : 0;
assign detect_min[532][16] = (mid_1[4271:4264] < mid_2[4279:4272]) ? 1 : 0;
assign detect_min[532][17] = (mid_1[4271:4264] < btm_0[4263:4256]) ? 1 : 0;
assign detect_min[532][18] = (mid_1[4271:4264] < btm_0[4271:4264]) ? 1 : 0;
assign detect_min[532][19] = (mid_1[4271:4264] < btm_0[4279:4272]) ? 1 : 0;
assign detect_min[532][20] = (mid_1[4271:4264] < btm_1[4263:4256]) ? 1 : 0;
assign detect_min[532][21] = (mid_1[4271:4264] < btm_1[4271:4264]) ? 1 : 0;
assign detect_min[532][22] = (mid_1[4271:4264] < btm_1[4279:4272]) ? 1 : 0;
assign detect_min[532][23] = (mid_1[4271:4264] < btm_2[4263:4256]) ? 1 : 0;
assign detect_min[532][24] = (mid_1[4271:4264] < btm_2[4271:4264]) ? 1 : 0;
assign detect_min[532][25] = (mid_1[4271:4264] < btm_2[4279:4272]) ? 1 : 0;

assign detect_min[533][0] = (mid_1[4279:4272] < top_0[4271:4264]) ? 1 : 0;
assign detect_min[533][1] = (mid_1[4279:4272] < top_0[4279:4272]) ? 1 : 0;
assign detect_min[533][2] = (mid_1[4279:4272] < top_0[4287:4280]) ? 1 : 0;
assign detect_min[533][3] = (mid_1[4279:4272] < top_1[4271:4264]) ? 1 : 0;
assign detect_min[533][4] = (mid_1[4279:4272] < top_1[4279:4272]) ? 1 : 0;
assign detect_min[533][5] = (mid_1[4279:4272] < top_1[4287:4280]) ? 1 : 0;
assign detect_min[533][6] = (mid_1[4279:4272] < top_2[4271:4264]) ? 1 : 0;
assign detect_min[533][7] = (mid_1[4279:4272] < top_2[4279:4272]) ? 1 : 0;
assign detect_min[533][8] = (mid_1[4279:4272] < top_2[4287:4280]) ? 1 : 0;
assign detect_min[533][9] = (mid_1[4279:4272] < mid_0[4271:4264]) ? 1 : 0;
assign detect_min[533][10] = (mid_1[4279:4272] < mid_0[4279:4272]) ? 1 : 0;
assign detect_min[533][11] = (mid_1[4279:4272] < mid_0[4287:4280]) ? 1 : 0;
assign detect_min[533][12] = (mid_1[4279:4272] < mid_1[4271:4264]) ? 1 : 0;
assign detect_min[533][13] = (mid_1[4279:4272] < mid_1[4287:4280]) ? 1 : 0;
assign detect_min[533][14] = (mid_1[4279:4272] < mid_2[4271:4264]) ? 1 : 0;
assign detect_min[533][15] = (mid_1[4279:4272] < mid_2[4279:4272]) ? 1 : 0;
assign detect_min[533][16] = (mid_1[4279:4272] < mid_2[4287:4280]) ? 1 : 0;
assign detect_min[533][17] = (mid_1[4279:4272] < btm_0[4271:4264]) ? 1 : 0;
assign detect_min[533][18] = (mid_1[4279:4272] < btm_0[4279:4272]) ? 1 : 0;
assign detect_min[533][19] = (mid_1[4279:4272] < btm_0[4287:4280]) ? 1 : 0;
assign detect_min[533][20] = (mid_1[4279:4272] < btm_1[4271:4264]) ? 1 : 0;
assign detect_min[533][21] = (mid_1[4279:4272] < btm_1[4279:4272]) ? 1 : 0;
assign detect_min[533][22] = (mid_1[4279:4272] < btm_1[4287:4280]) ? 1 : 0;
assign detect_min[533][23] = (mid_1[4279:4272] < btm_2[4271:4264]) ? 1 : 0;
assign detect_min[533][24] = (mid_1[4279:4272] < btm_2[4279:4272]) ? 1 : 0;
assign detect_min[533][25] = (mid_1[4279:4272] < btm_2[4287:4280]) ? 1 : 0;

assign detect_min[534][0] = (mid_1[4287:4280] < top_0[4279:4272]) ? 1 : 0;
assign detect_min[534][1] = (mid_1[4287:4280] < top_0[4287:4280]) ? 1 : 0;
assign detect_min[534][2] = (mid_1[4287:4280] < top_0[4295:4288]) ? 1 : 0;
assign detect_min[534][3] = (mid_1[4287:4280] < top_1[4279:4272]) ? 1 : 0;
assign detect_min[534][4] = (mid_1[4287:4280] < top_1[4287:4280]) ? 1 : 0;
assign detect_min[534][5] = (mid_1[4287:4280] < top_1[4295:4288]) ? 1 : 0;
assign detect_min[534][6] = (mid_1[4287:4280] < top_2[4279:4272]) ? 1 : 0;
assign detect_min[534][7] = (mid_1[4287:4280] < top_2[4287:4280]) ? 1 : 0;
assign detect_min[534][8] = (mid_1[4287:4280] < top_2[4295:4288]) ? 1 : 0;
assign detect_min[534][9] = (mid_1[4287:4280] < mid_0[4279:4272]) ? 1 : 0;
assign detect_min[534][10] = (mid_1[4287:4280] < mid_0[4287:4280]) ? 1 : 0;
assign detect_min[534][11] = (mid_1[4287:4280] < mid_0[4295:4288]) ? 1 : 0;
assign detect_min[534][12] = (mid_1[4287:4280] < mid_1[4279:4272]) ? 1 : 0;
assign detect_min[534][13] = (mid_1[4287:4280] < mid_1[4295:4288]) ? 1 : 0;
assign detect_min[534][14] = (mid_1[4287:4280] < mid_2[4279:4272]) ? 1 : 0;
assign detect_min[534][15] = (mid_1[4287:4280] < mid_2[4287:4280]) ? 1 : 0;
assign detect_min[534][16] = (mid_1[4287:4280] < mid_2[4295:4288]) ? 1 : 0;
assign detect_min[534][17] = (mid_1[4287:4280] < btm_0[4279:4272]) ? 1 : 0;
assign detect_min[534][18] = (mid_1[4287:4280] < btm_0[4287:4280]) ? 1 : 0;
assign detect_min[534][19] = (mid_1[4287:4280] < btm_0[4295:4288]) ? 1 : 0;
assign detect_min[534][20] = (mid_1[4287:4280] < btm_1[4279:4272]) ? 1 : 0;
assign detect_min[534][21] = (mid_1[4287:4280] < btm_1[4287:4280]) ? 1 : 0;
assign detect_min[534][22] = (mid_1[4287:4280] < btm_1[4295:4288]) ? 1 : 0;
assign detect_min[534][23] = (mid_1[4287:4280] < btm_2[4279:4272]) ? 1 : 0;
assign detect_min[534][24] = (mid_1[4287:4280] < btm_2[4287:4280]) ? 1 : 0;
assign detect_min[534][25] = (mid_1[4287:4280] < btm_2[4295:4288]) ? 1 : 0;

assign detect_min[535][0] = (mid_1[4295:4288] < top_0[4287:4280]) ? 1 : 0;
assign detect_min[535][1] = (mid_1[4295:4288] < top_0[4295:4288]) ? 1 : 0;
assign detect_min[535][2] = (mid_1[4295:4288] < top_0[4303:4296]) ? 1 : 0;
assign detect_min[535][3] = (mid_1[4295:4288] < top_1[4287:4280]) ? 1 : 0;
assign detect_min[535][4] = (mid_1[4295:4288] < top_1[4295:4288]) ? 1 : 0;
assign detect_min[535][5] = (mid_1[4295:4288] < top_1[4303:4296]) ? 1 : 0;
assign detect_min[535][6] = (mid_1[4295:4288] < top_2[4287:4280]) ? 1 : 0;
assign detect_min[535][7] = (mid_1[4295:4288] < top_2[4295:4288]) ? 1 : 0;
assign detect_min[535][8] = (mid_1[4295:4288] < top_2[4303:4296]) ? 1 : 0;
assign detect_min[535][9] = (mid_1[4295:4288] < mid_0[4287:4280]) ? 1 : 0;
assign detect_min[535][10] = (mid_1[4295:4288] < mid_0[4295:4288]) ? 1 : 0;
assign detect_min[535][11] = (mid_1[4295:4288] < mid_0[4303:4296]) ? 1 : 0;
assign detect_min[535][12] = (mid_1[4295:4288] < mid_1[4287:4280]) ? 1 : 0;
assign detect_min[535][13] = (mid_1[4295:4288] < mid_1[4303:4296]) ? 1 : 0;
assign detect_min[535][14] = (mid_1[4295:4288] < mid_2[4287:4280]) ? 1 : 0;
assign detect_min[535][15] = (mid_1[4295:4288] < mid_2[4295:4288]) ? 1 : 0;
assign detect_min[535][16] = (mid_1[4295:4288] < mid_2[4303:4296]) ? 1 : 0;
assign detect_min[535][17] = (mid_1[4295:4288] < btm_0[4287:4280]) ? 1 : 0;
assign detect_min[535][18] = (mid_1[4295:4288] < btm_0[4295:4288]) ? 1 : 0;
assign detect_min[535][19] = (mid_1[4295:4288] < btm_0[4303:4296]) ? 1 : 0;
assign detect_min[535][20] = (mid_1[4295:4288] < btm_1[4287:4280]) ? 1 : 0;
assign detect_min[535][21] = (mid_1[4295:4288] < btm_1[4295:4288]) ? 1 : 0;
assign detect_min[535][22] = (mid_1[4295:4288] < btm_1[4303:4296]) ? 1 : 0;
assign detect_min[535][23] = (mid_1[4295:4288] < btm_2[4287:4280]) ? 1 : 0;
assign detect_min[535][24] = (mid_1[4295:4288] < btm_2[4295:4288]) ? 1 : 0;
assign detect_min[535][25] = (mid_1[4295:4288] < btm_2[4303:4296]) ? 1 : 0;

assign detect_min[536][0] = (mid_1[4303:4296] < top_0[4295:4288]) ? 1 : 0;
assign detect_min[536][1] = (mid_1[4303:4296] < top_0[4303:4296]) ? 1 : 0;
assign detect_min[536][2] = (mid_1[4303:4296] < top_0[4311:4304]) ? 1 : 0;
assign detect_min[536][3] = (mid_1[4303:4296] < top_1[4295:4288]) ? 1 : 0;
assign detect_min[536][4] = (mid_1[4303:4296] < top_1[4303:4296]) ? 1 : 0;
assign detect_min[536][5] = (mid_1[4303:4296] < top_1[4311:4304]) ? 1 : 0;
assign detect_min[536][6] = (mid_1[4303:4296] < top_2[4295:4288]) ? 1 : 0;
assign detect_min[536][7] = (mid_1[4303:4296] < top_2[4303:4296]) ? 1 : 0;
assign detect_min[536][8] = (mid_1[4303:4296] < top_2[4311:4304]) ? 1 : 0;
assign detect_min[536][9] = (mid_1[4303:4296] < mid_0[4295:4288]) ? 1 : 0;
assign detect_min[536][10] = (mid_1[4303:4296] < mid_0[4303:4296]) ? 1 : 0;
assign detect_min[536][11] = (mid_1[4303:4296] < mid_0[4311:4304]) ? 1 : 0;
assign detect_min[536][12] = (mid_1[4303:4296] < mid_1[4295:4288]) ? 1 : 0;
assign detect_min[536][13] = (mid_1[4303:4296] < mid_1[4311:4304]) ? 1 : 0;
assign detect_min[536][14] = (mid_1[4303:4296] < mid_2[4295:4288]) ? 1 : 0;
assign detect_min[536][15] = (mid_1[4303:4296] < mid_2[4303:4296]) ? 1 : 0;
assign detect_min[536][16] = (mid_1[4303:4296] < mid_2[4311:4304]) ? 1 : 0;
assign detect_min[536][17] = (mid_1[4303:4296] < btm_0[4295:4288]) ? 1 : 0;
assign detect_min[536][18] = (mid_1[4303:4296] < btm_0[4303:4296]) ? 1 : 0;
assign detect_min[536][19] = (mid_1[4303:4296] < btm_0[4311:4304]) ? 1 : 0;
assign detect_min[536][20] = (mid_1[4303:4296] < btm_1[4295:4288]) ? 1 : 0;
assign detect_min[536][21] = (mid_1[4303:4296] < btm_1[4303:4296]) ? 1 : 0;
assign detect_min[536][22] = (mid_1[4303:4296] < btm_1[4311:4304]) ? 1 : 0;
assign detect_min[536][23] = (mid_1[4303:4296] < btm_2[4295:4288]) ? 1 : 0;
assign detect_min[536][24] = (mid_1[4303:4296] < btm_2[4303:4296]) ? 1 : 0;
assign detect_min[536][25] = (mid_1[4303:4296] < btm_2[4311:4304]) ? 1 : 0;

assign detect_min[537][0] = (mid_1[4311:4304] < top_0[4303:4296]) ? 1 : 0;
assign detect_min[537][1] = (mid_1[4311:4304] < top_0[4311:4304]) ? 1 : 0;
assign detect_min[537][2] = (mid_1[4311:4304] < top_0[4319:4312]) ? 1 : 0;
assign detect_min[537][3] = (mid_1[4311:4304] < top_1[4303:4296]) ? 1 : 0;
assign detect_min[537][4] = (mid_1[4311:4304] < top_1[4311:4304]) ? 1 : 0;
assign detect_min[537][5] = (mid_1[4311:4304] < top_1[4319:4312]) ? 1 : 0;
assign detect_min[537][6] = (mid_1[4311:4304] < top_2[4303:4296]) ? 1 : 0;
assign detect_min[537][7] = (mid_1[4311:4304] < top_2[4311:4304]) ? 1 : 0;
assign detect_min[537][8] = (mid_1[4311:4304] < top_2[4319:4312]) ? 1 : 0;
assign detect_min[537][9] = (mid_1[4311:4304] < mid_0[4303:4296]) ? 1 : 0;
assign detect_min[537][10] = (mid_1[4311:4304] < mid_0[4311:4304]) ? 1 : 0;
assign detect_min[537][11] = (mid_1[4311:4304] < mid_0[4319:4312]) ? 1 : 0;
assign detect_min[537][12] = (mid_1[4311:4304] < mid_1[4303:4296]) ? 1 : 0;
assign detect_min[537][13] = (mid_1[4311:4304] < mid_1[4319:4312]) ? 1 : 0;
assign detect_min[537][14] = (mid_1[4311:4304] < mid_2[4303:4296]) ? 1 : 0;
assign detect_min[537][15] = (mid_1[4311:4304] < mid_2[4311:4304]) ? 1 : 0;
assign detect_min[537][16] = (mid_1[4311:4304] < mid_2[4319:4312]) ? 1 : 0;
assign detect_min[537][17] = (mid_1[4311:4304] < btm_0[4303:4296]) ? 1 : 0;
assign detect_min[537][18] = (mid_1[4311:4304] < btm_0[4311:4304]) ? 1 : 0;
assign detect_min[537][19] = (mid_1[4311:4304] < btm_0[4319:4312]) ? 1 : 0;
assign detect_min[537][20] = (mid_1[4311:4304] < btm_1[4303:4296]) ? 1 : 0;
assign detect_min[537][21] = (mid_1[4311:4304] < btm_1[4311:4304]) ? 1 : 0;
assign detect_min[537][22] = (mid_1[4311:4304] < btm_1[4319:4312]) ? 1 : 0;
assign detect_min[537][23] = (mid_1[4311:4304] < btm_2[4303:4296]) ? 1 : 0;
assign detect_min[537][24] = (mid_1[4311:4304] < btm_2[4311:4304]) ? 1 : 0;
assign detect_min[537][25] = (mid_1[4311:4304] < btm_2[4319:4312]) ? 1 : 0;

assign detect_min[538][0] = (mid_1[4319:4312] < top_0[4311:4304]) ? 1 : 0;
assign detect_min[538][1] = (mid_1[4319:4312] < top_0[4319:4312]) ? 1 : 0;
assign detect_min[538][2] = (mid_1[4319:4312] < top_0[4327:4320]) ? 1 : 0;
assign detect_min[538][3] = (mid_1[4319:4312] < top_1[4311:4304]) ? 1 : 0;
assign detect_min[538][4] = (mid_1[4319:4312] < top_1[4319:4312]) ? 1 : 0;
assign detect_min[538][5] = (mid_1[4319:4312] < top_1[4327:4320]) ? 1 : 0;
assign detect_min[538][6] = (mid_1[4319:4312] < top_2[4311:4304]) ? 1 : 0;
assign detect_min[538][7] = (mid_1[4319:4312] < top_2[4319:4312]) ? 1 : 0;
assign detect_min[538][8] = (mid_1[4319:4312] < top_2[4327:4320]) ? 1 : 0;
assign detect_min[538][9] = (mid_1[4319:4312] < mid_0[4311:4304]) ? 1 : 0;
assign detect_min[538][10] = (mid_1[4319:4312] < mid_0[4319:4312]) ? 1 : 0;
assign detect_min[538][11] = (mid_1[4319:4312] < mid_0[4327:4320]) ? 1 : 0;
assign detect_min[538][12] = (mid_1[4319:4312] < mid_1[4311:4304]) ? 1 : 0;
assign detect_min[538][13] = (mid_1[4319:4312] < mid_1[4327:4320]) ? 1 : 0;
assign detect_min[538][14] = (mid_1[4319:4312] < mid_2[4311:4304]) ? 1 : 0;
assign detect_min[538][15] = (mid_1[4319:4312] < mid_2[4319:4312]) ? 1 : 0;
assign detect_min[538][16] = (mid_1[4319:4312] < mid_2[4327:4320]) ? 1 : 0;
assign detect_min[538][17] = (mid_1[4319:4312] < btm_0[4311:4304]) ? 1 : 0;
assign detect_min[538][18] = (mid_1[4319:4312] < btm_0[4319:4312]) ? 1 : 0;
assign detect_min[538][19] = (mid_1[4319:4312] < btm_0[4327:4320]) ? 1 : 0;
assign detect_min[538][20] = (mid_1[4319:4312] < btm_1[4311:4304]) ? 1 : 0;
assign detect_min[538][21] = (mid_1[4319:4312] < btm_1[4319:4312]) ? 1 : 0;
assign detect_min[538][22] = (mid_1[4319:4312] < btm_1[4327:4320]) ? 1 : 0;
assign detect_min[538][23] = (mid_1[4319:4312] < btm_2[4311:4304]) ? 1 : 0;
assign detect_min[538][24] = (mid_1[4319:4312] < btm_2[4319:4312]) ? 1 : 0;
assign detect_min[538][25] = (mid_1[4319:4312] < btm_2[4327:4320]) ? 1 : 0;

assign detect_min[539][0] = (mid_1[4327:4320] < top_0[4319:4312]) ? 1 : 0;
assign detect_min[539][1] = (mid_1[4327:4320] < top_0[4327:4320]) ? 1 : 0;
assign detect_min[539][2] = (mid_1[4327:4320] < top_0[4335:4328]) ? 1 : 0;
assign detect_min[539][3] = (mid_1[4327:4320] < top_1[4319:4312]) ? 1 : 0;
assign detect_min[539][4] = (mid_1[4327:4320] < top_1[4327:4320]) ? 1 : 0;
assign detect_min[539][5] = (mid_1[4327:4320] < top_1[4335:4328]) ? 1 : 0;
assign detect_min[539][6] = (mid_1[4327:4320] < top_2[4319:4312]) ? 1 : 0;
assign detect_min[539][7] = (mid_1[4327:4320] < top_2[4327:4320]) ? 1 : 0;
assign detect_min[539][8] = (mid_1[4327:4320] < top_2[4335:4328]) ? 1 : 0;
assign detect_min[539][9] = (mid_1[4327:4320] < mid_0[4319:4312]) ? 1 : 0;
assign detect_min[539][10] = (mid_1[4327:4320] < mid_0[4327:4320]) ? 1 : 0;
assign detect_min[539][11] = (mid_1[4327:4320] < mid_0[4335:4328]) ? 1 : 0;
assign detect_min[539][12] = (mid_1[4327:4320] < mid_1[4319:4312]) ? 1 : 0;
assign detect_min[539][13] = (mid_1[4327:4320] < mid_1[4335:4328]) ? 1 : 0;
assign detect_min[539][14] = (mid_1[4327:4320] < mid_2[4319:4312]) ? 1 : 0;
assign detect_min[539][15] = (mid_1[4327:4320] < mid_2[4327:4320]) ? 1 : 0;
assign detect_min[539][16] = (mid_1[4327:4320] < mid_2[4335:4328]) ? 1 : 0;
assign detect_min[539][17] = (mid_1[4327:4320] < btm_0[4319:4312]) ? 1 : 0;
assign detect_min[539][18] = (mid_1[4327:4320] < btm_0[4327:4320]) ? 1 : 0;
assign detect_min[539][19] = (mid_1[4327:4320] < btm_0[4335:4328]) ? 1 : 0;
assign detect_min[539][20] = (mid_1[4327:4320] < btm_1[4319:4312]) ? 1 : 0;
assign detect_min[539][21] = (mid_1[4327:4320] < btm_1[4327:4320]) ? 1 : 0;
assign detect_min[539][22] = (mid_1[4327:4320] < btm_1[4335:4328]) ? 1 : 0;
assign detect_min[539][23] = (mid_1[4327:4320] < btm_2[4319:4312]) ? 1 : 0;
assign detect_min[539][24] = (mid_1[4327:4320] < btm_2[4327:4320]) ? 1 : 0;
assign detect_min[539][25] = (mid_1[4327:4320] < btm_2[4335:4328]) ? 1 : 0;

assign detect_min[540][0] = (mid_1[4335:4328] < top_0[4327:4320]) ? 1 : 0;
assign detect_min[540][1] = (mid_1[4335:4328] < top_0[4335:4328]) ? 1 : 0;
assign detect_min[540][2] = (mid_1[4335:4328] < top_0[4343:4336]) ? 1 : 0;
assign detect_min[540][3] = (mid_1[4335:4328] < top_1[4327:4320]) ? 1 : 0;
assign detect_min[540][4] = (mid_1[4335:4328] < top_1[4335:4328]) ? 1 : 0;
assign detect_min[540][5] = (mid_1[4335:4328] < top_1[4343:4336]) ? 1 : 0;
assign detect_min[540][6] = (mid_1[4335:4328] < top_2[4327:4320]) ? 1 : 0;
assign detect_min[540][7] = (mid_1[4335:4328] < top_2[4335:4328]) ? 1 : 0;
assign detect_min[540][8] = (mid_1[4335:4328] < top_2[4343:4336]) ? 1 : 0;
assign detect_min[540][9] = (mid_1[4335:4328] < mid_0[4327:4320]) ? 1 : 0;
assign detect_min[540][10] = (mid_1[4335:4328] < mid_0[4335:4328]) ? 1 : 0;
assign detect_min[540][11] = (mid_1[4335:4328] < mid_0[4343:4336]) ? 1 : 0;
assign detect_min[540][12] = (mid_1[4335:4328] < mid_1[4327:4320]) ? 1 : 0;
assign detect_min[540][13] = (mid_1[4335:4328] < mid_1[4343:4336]) ? 1 : 0;
assign detect_min[540][14] = (mid_1[4335:4328] < mid_2[4327:4320]) ? 1 : 0;
assign detect_min[540][15] = (mid_1[4335:4328] < mid_2[4335:4328]) ? 1 : 0;
assign detect_min[540][16] = (mid_1[4335:4328] < mid_2[4343:4336]) ? 1 : 0;
assign detect_min[540][17] = (mid_1[4335:4328] < btm_0[4327:4320]) ? 1 : 0;
assign detect_min[540][18] = (mid_1[4335:4328] < btm_0[4335:4328]) ? 1 : 0;
assign detect_min[540][19] = (mid_1[4335:4328] < btm_0[4343:4336]) ? 1 : 0;
assign detect_min[540][20] = (mid_1[4335:4328] < btm_1[4327:4320]) ? 1 : 0;
assign detect_min[540][21] = (mid_1[4335:4328] < btm_1[4335:4328]) ? 1 : 0;
assign detect_min[540][22] = (mid_1[4335:4328] < btm_1[4343:4336]) ? 1 : 0;
assign detect_min[540][23] = (mid_1[4335:4328] < btm_2[4327:4320]) ? 1 : 0;
assign detect_min[540][24] = (mid_1[4335:4328] < btm_2[4335:4328]) ? 1 : 0;
assign detect_min[540][25] = (mid_1[4335:4328] < btm_2[4343:4336]) ? 1 : 0;

assign detect_min[541][0] = (mid_1[4343:4336] < top_0[4335:4328]) ? 1 : 0;
assign detect_min[541][1] = (mid_1[4343:4336] < top_0[4343:4336]) ? 1 : 0;
assign detect_min[541][2] = (mid_1[4343:4336] < top_0[4351:4344]) ? 1 : 0;
assign detect_min[541][3] = (mid_1[4343:4336] < top_1[4335:4328]) ? 1 : 0;
assign detect_min[541][4] = (mid_1[4343:4336] < top_1[4343:4336]) ? 1 : 0;
assign detect_min[541][5] = (mid_1[4343:4336] < top_1[4351:4344]) ? 1 : 0;
assign detect_min[541][6] = (mid_1[4343:4336] < top_2[4335:4328]) ? 1 : 0;
assign detect_min[541][7] = (mid_1[4343:4336] < top_2[4343:4336]) ? 1 : 0;
assign detect_min[541][8] = (mid_1[4343:4336] < top_2[4351:4344]) ? 1 : 0;
assign detect_min[541][9] = (mid_1[4343:4336] < mid_0[4335:4328]) ? 1 : 0;
assign detect_min[541][10] = (mid_1[4343:4336] < mid_0[4343:4336]) ? 1 : 0;
assign detect_min[541][11] = (mid_1[4343:4336] < mid_0[4351:4344]) ? 1 : 0;
assign detect_min[541][12] = (mid_1[4343:4336] < mid_1[4335:4328]) ? 1 : 0;
assign detect_min[541][13] = (mid_1[4343:4336] < mid_1[4351:4344]) ? 1 : 0;
assign detect_min[541][14] = (mid_1[4343:4336] < mid_2[4335:4328]) ? 1 : 0;
assign detect_min[541][15] = (mid_1[4343:4336] < mid_2[4343:4336]) ? 1 : 0;
assign detect_min[541][16] = (mid_1[4343:4336] < mid_2[4351:4344]) ? 1 : 0;
assign detect_min[541][17] = (mid_1[4343:4336] < btm_0[4335:4328]) ? 1 : 0;
assign detect_min[541][18] = (mid_1[4343:4336] < btm_0[4343:4336]) ? 1 : 0;
assign detect_min[541][19] = (mid_1[4343:4336] < btm_0[4351:4344]) ? 1 : 0;
assign detect_min[541][20] = (mid_1[4343:4336] < btm_1[4335:4328]) ? 1 : 0;
assign detect_min[541][21] = (mid_1[4343:4336] < btm_1[4343:4336]) ? 1 : 0;
assign detect_min[541][22] = (mid_1[4343:4336] < btm_1[4351:4344]) ? 1 : 0;
assign detect_min[541][23] = (mid_1[4343:4336] < btm_2[4335:4328]) ? 1 : 0;
assign detect_min[541][24] = (mid_1[4343:4336] < btm_2[4343:4336]) ? 1 : 0;
assign detect_min[541][25] = (mid_1[4343:4336] < btm_2[4351:4344]) ? 1 : 0;

assign detect_min[542][0] = (mid_1[4351:4344] < top_0[4343:4336]) ? 1 : 0;
assign detect_min[542][1] = (mid_1[4351:4344] < top_0[4351:4344]) ? 1 : 0;
assign detect_min[542][2] = (mid_1[4351:4344] < top_0[4359:4352]) ? 1 : 0;
assign detect_min[542][3] = (mid_1[4351:4344] < top_1[4343:4336]) ? 1 : 0;
assign detect_min[542][4] = (mid_1[4351:4344] < top_1[4351:4344]) ? 1 : 0;
assign detect_min[542][5] = (mid_1[4351:4344] < top_1[4359:4352]) ? 1 : 0;
assign detect_min[542][6] = (mid_1[4351:4344] < top_2[4343:4336]) ? 1 : 0;
assign detect_min[542][7] = (mid_1[4351:4344] < top_2[4351:4344]) ? 1 : 0;
assign detect_min[542][8] = (mid_1[4351:4344] < top_2[4359:4352]) ? 1 : 0;
assign detect_min[542][9] = (mid_1[4351:4344] < mid_0[4343:4336]) ? 1 : 0;
assign detect_min[542][10] = (mid_1[4351:4344] < mid_0[4351:4344]) ? 1 : 0;
assign detect_min[542][11] = (mid_1[4351:4344] < mid_0[4359:4352]) ? 1 : 0;
assign detect_min[542][12] = (mid_1[4351:4344] < mid_1[4343:4336]) ? 1 : 0;
assign detect_min[542][13] = (mid_1[4351:4344] < mid_1[4359:4352]) ? 1 : 0;
assign detect_min[542][14] = (mid_1[4351:4344] < mid_2[4343:4336]) ? 1 : 0;
assign detect_min[542][15] = (mid_1[4351:4344] < mid_2[4351:4344]) ? 1 : 0;
assign detect_min[542][16] = (mid_1[4351:4344] < mid_2[4359:4352]) ? 1 : 0;
assign detect_min[542][17] = (mid_1[4351:4344] < btm_0[4343:4336]) ? 1 : 0;
assign detect_min[542][18] = (mid_1[4351:4344] < btm_0[4351:4344]) ? 1 : 0;
assign detect_min[542][19] = (mid_1[4351:4344] < btm_0[4359:4352]) ? 1 : 0;
assign detect_min[542][20] = (mid_1[4351:4344] < btm_1[4343:4336]) ? 1 : 0;
assign detect_min[542][21] = (mid_1[4351:4344] < btm_1[4351:4344]) ? 1 : 0;
assign detect_min[542][22] = (mid_1[4351:4344] < btm_1[4359:4352]) ? 1 : 0;
assign detect_min[542][23] = (mid_1[4351:4344] < btm_2[4343:4336]) ? 1 : 0;
assign detect_min[542][24] = (mid_1[4351:4344] < btm_2[4351:4344]) ? 1 : 0;
assign detect_min[542][25] = (mid_1[4351:4344] < btm_2[4359:4352]) ? 1 : 0;

assign detect_min[543][0] = (mid_1[4359:4352] < top_0[4351:4344]) ? 1 : 0;
assign detect_min[543][1] = (mid_1[4359:4352] < top_0[4359:4352]) ? 1 : 0;
assign detect_min[543][2] = (mid_1[4359:4352] < top_0[4367:4360]) ? 1 : 0;
assign detect_min[543][3] = (mid_1[4359:4352] < top_1[4351:4344]) ? 1 : 0;
assign detect_min[543][4] = (mid_1[4359:4352] < top_1[4359:4352]) ? 1 : 0;
assign detect_min[543][5] = (mid_1[4359:4352] < top_1[4367:4360]) ? 1 : 0;
assign detect_min[543][6] = (mid_1[4359:4352] < top_2[4351:4344]) ? 1 : 0;
assign detect_min[543][7] = (mid_1[4359:4352] < top_2[4359:4352]) ? 1 : 0;
assign detect_min[543][8] = (mid_1[4359:4352] < top_2[4367:4360]) ? 1 : 0;
assign detect_min[543][9] = (mid_1[4359:4352] < mid_0[4351:4344]) ? 1 : 0;
assign detect_min[543][10] = (mid_1[4359:4352] < mid_0[4359:4352]) ? 1 : 0;
assign detect_min[543][11] = (mid_1[4359:4352] < mid_0[4367:4360]) ? 1 : 0;
assign detect_min[543][12] = (mid_1[4359:4352] < mid_1[4351:4344]) ? 1 : 0;
assign detect_min[543][13] = (mid_1[4359:4352] < mid_1[4367:4360]) ? 1 : 0;
assign detect_min[543][14] = (mid_1[4359:4352] < mid_2[4351:4344]) ? 1 : 0;
assign detect_min[543][15] = (mid_1[4359:4352] < mid_2[4359:4352]) ? 1 : 0;
assign detect_min[543][16] = (mid_1[4359:4352] < mid_2[4367:4360]) ? 1 : 0;
assign detect_min[543][17] = (mid_1[4359:4352] < btm_0[4351:4344]) ? 1 : 0;
assign detect_min[543][18] = (mid_1[4359:4352] < btm_0[4359:4352]) ? 1 : 0;
assign detect_min[543][19] = (mid_1[4359:4352] < btm_0[4367:4360]) ? 1 : 0;
assign detect_min[543][20] = (mid_1[4359:4352] < btm_1[4351:4344]) ? 1 : 0;
assign detect_min[543][21] = (mid_1[4359:4352] < btm_1[4359:4352]) ? 1 : 0;
assign detect_min[543][22] = (mid_1[4359:4352] < btm_1[4367:4360]) ? 1 : 0;
assign detect_min[543][23] = (mid_1[4359:4352] < btm_2[4351:4344]) ? 1 : 0;
assign detect_min[543][24] = (mid_1[4359:4352] < btm_2[4359:4352]) ? 1 : 0;
assign detect_min[543][25] = (mid_1[4359:4352] < btm_2[4367:4360]) ? 1 : 0;

assign detect_min[544][0] = (mid_1[4367:4360] < top_0[4359:4352]) ? 1 : 0;
assign detect_min[544][1] = (mid_1[4367:4360] < top_0[4367:4360]) ? 1 : 0;
assign detect_min[544][2] = (mid_1[4367:4360] < top_0[4375:4368]) ? 1 : 0;
assign detect_min[544][3] = (mid_1[4367:4360] < top_1[4359:4352]) ? 1 : 0;
assign detect_min[544][4] = (mid_1[4367:4360] < top_1[4367:4360]) ? 1 : 0;
assign detect_min[544][5] = (mid_1[4367:4360] < top_1[4375:4368]) ? 1 : 0;
assign detect_min[544][6] = (mid_1[4367:4360] < top_2[4359:4352]) ? 1 : 0;
assign detect_min[544][7] = (mid_1[4367:4360] < top_2[4367:4360]) ? 1 : 0;
assign detect_min[544][8] = (mid_1[4367:4360] < top_2[4375:4368]) ? 1 : 0;
assign detect_min[544][9] = (mid_1[4367:4360] < mid_0[4359:4352]) ? 1 : 0;
assign detect_min[544][10] = (mid_1[4367:4360] < mid_0[4367:4360]) ? 1 : 0;
assign detect_min[544][11] = (mid_1[4367:4360] < mid_0[4375:4368]) ? 1 : 0;
assign detect_min[544][12] = (mid_1[4367:4360] < mid_1[4359:4352]) ? 1 : 0;
assign detect_min[544][13] = (mid_1[4367:4360] < mid_1[4375:4368]) ? 1 : 0;
assign detect_min[544][14] = (mid_1[4367:4360] < mid_2[4359:4352]) ? 1 : 0;
assign detect_min[544][15] = (mid_1[4367:4360] < mid_2[4367:4360]) ? 1 : 0;
assign detect_min[544][16] = (mid_1[4367:4360] < mid_2[4375:4368]) ? 1 : 0;
assign detect_min[544][17] = (mid_1[4367:4360] < btm_0[4359:4352]) ? 1 : 0;
assign detect_min[544][18] = (mid_1[4367:4360] < btm_0[4367:4360]) ? 1 : 0;
assign detect_min[544][19] = (mid_1[4367:4360] < btm_0[4375:4368]) ? 1 : 0;
assign detect_min[544][20] = (mid_1[4367:4360] < btm_1[4359:4352]) ? 1 : 0;
assign detect_min[544][21] = (mid_1[4367:4360] < btm_1[4367:4360]) ? 1 : 0;
assign detect_min[544][22] = (mid_1[4367:4360] < btm_1[4375:4368]) ? 1 : 0;
assign detect_min[544][23] = (mid_1[4367:4360] < btm_2[4359:4352]) ? 1 : 0;
assign detect_min[544][24] = (mid_1[4367:4360] < btm_2[4367:4360]) ? 1 : 0;
assign detect_min[544][25] = (mid_1[4367:4360] < btm_2[4375:4368]) ? 1 : 0;

assign detect_min[545][0] = (mid_1[4375:4368] < top_0[4367:4360]) ? 1 : 0;
assign detect_min[545][1] = (mid_1[4375:4368] < top_0[4375:4368]) ? 1 : 0;
assign detect_min[545][2] = (mid_1[4375:4368] < top_0[4383:4376]) ? 1 : 0;
assign detect_min[545][3] = (mid_1[4375:4368] < top_1[4367:4360]) ? 1 : 0;
assign detect_min[545][4] = (mid_1[4375:4368] < top_1[4375:4368]) ? 1 : 0;
assign detect_min[545][5] = (mid_1[4375:4368] < top_1[4383:4376]) ? 1 : 0;
assign detect_min[545][6] = (mid_1[4375:4368] < top_2[4367:4360]) ? 1 : 0;
assign detect_min[545][7] = (mid_1[4375:4368] < top_2[4375:4368]) ? 1 : 0;
assign detect_min[545][8] = (mid_1[4375:4368] < top_2[4383:4376]) ? 1 : 0;
assign detect_min[545][9] = (mid_1[4375:4368] < mid_0[4367:4360]) ? 1 : 0;
assign detect_min[545][10] = (mid_1[4375:4368] < mid_0[4375:4368]) ? 1 : 0;
assign detect_min[545][11] = (mid_1[4375:4368] < mid_0[4383:4376]) ? 1 : 0;
assign detect_min[545][12] = (mid_1[4375:4368] < mid_1[4367:4360]) ? 1 : 0;
assign detect_min[545][13] = (mid_1[4375:4368] < mid_1[4383:4376]) ? 1 : 0;
assign detect_min[545][14] = (mid_1[4375:4368] < mid_2[4367:4360]) ? 1 : 0;
assign detect_min[545][15] = (mid_1[4375:4368] < mid_2[4375:4368]) ? 1 : 0;
assign detect_min[545][16] = (mid_1[4375:4368] < mid_2[4383:4376]) ? 1 : 0;
assign detect_min[545][17] = (mid_1[4375:4368] < btm_0[4367:4360]) ? 1 : 0;
assign detect_min[545][18] = (mid_1[4375:4368] < btm_0[4375:4368]) ? 1 : 0;
assign detect_min[545][19] = (mid_1[4375:4368] < btm_0[4383:4376]) ? 1 : 0;
assign detect_min[545][20] = (mid_1[4375:4368] < btm_1[4367:4360]) ? 1 : 0;
assign detect_min[545][21] = (mid_1[4375:4368] < btm_1[4375:4368]) ? 1 : 0;
assign detect_min[545][22] = (mid_1[4375:4368] < btm_1[4383:4376]) ? 1 : 0;
assign detect_min[545][23] = (mid_1[4375:4368] < btm_2[4367:4360]) ? 1 : 0;
assign detect_min[545][24] = (mid_1[4375:4368] < btm_2[4375:4368]) ? 1 : 0;
assign detect_min[545][25] = (mid_1[4375:4368] < btm_2[4383:4376]) ? 1 : 0;

assign detect_min[546][0] = (mid_1[4383:4376] < top_0[4375:4368]) ? 1 : 0;
assign detect_min[546][1] = (mid_1[4383:4376] < top_0[4383:4376]) ? 1 : 0;
assign detect_min[546][2] = (mid_1[4383:4376] < top_0[4391:4384]) ? 1 : 0;
assign detect_min[546][3] = (mid_1[4383:4376] < top_1[4375:4368]) ? 1 : 0;
assign detect_min[546][4] = (mid_1[4383:4376] < top_1[4383:4376]) ? 1 : 0;
assign detect_min[546][5] = (mid_1[4383:4376] < top_1[4391:4384]) ? 1 : 0;
assign detect_min[546][6] = (mid_1[4383:4376] < top_2[4375:4368]) ? 1 : 0;
assign detect_min[546][7] = (mid_1[4383:4376] < top_2[4383:4376]) ? 1 : 0;
assign detect_min[546][8] = (mid_1[4383:4376] < top_2[4391:4384]) ? 1 : 0;
assign detect_min[546][9] = (mid_1[4383:4376] < mid_0[4375:4368]) ? 1 : 0;
assign detect_min[546][10] = (mid_1[4383:4376] < mid_0[4383:4376]) ? 1 : 0;
assign detect_min[546][11] = (mid_1[4383:4376] < mid_0[4391:4384]) ? 1 : 0;
assign detect_min[546][12] = (mid_1[4383:4376] < mid_1[4375:4368]) ? 1 : 0;
assign detect_min[546][13] = (mid_1[4383:4376] < mid_1[4391:4384]) ? 1 : 0;
assign detect_min[546][14] = (mid_1[4383:4376] < mid_2[4375:4368]) ? 1 : 0;
assign detect_min[546][15] = (mid_1[4383:4376] < mid_2[4383:4376]) ? 1 : 0;
assign detect_min[546][16] = (mid_1[4383:4376] < mid_2[4391:4384]) ? 1 : 0;
assign detect_min[546][17] = (mid_1[4383:4376] < btm_0[4375:4368]) ? 1 : 0;
assign detect_min[546][18] = (mid_1[4383:4376] < btm_0[4383:4376]) ? 1 : 0;
assign detect_min[546][19] = (mid_1[4383:4376] < btm_0[4391:4384]) ? 1 : 0;
assign detect_min[546][20] = (mid_1[4383:4376] < btm_1[4375:4368]) ? 1 : 0;
assign detect_min[546][21] = (mid_1[4383:4376] < btm_1[4383:4376]) ? 1 : 0;
assign detect_min[546][22] = (mid_1[4383:4376] < btm_1[4391:4384]) ? 1 : 0;
assign detect_min[546][23] = (mid_1[4383:4376] < btm_2[4375:4368]) ? 1 : 0;
assign detect_min[546][24] = (mid_1[4383:4376] < btm_2[4383:4376]) ? 1 : 0;
assign detect_min[546][25] = (mid_1[4383:4376] < btm_2[4391:4384]) ? 1 : 0;

assign detect_min[547][0] = (mid_1[4391:4384] < top_0[4383:4376]) ? 1 : 0;
assign detect_min[547][1] = (mid_1[4391:4384] < top_0[4391:4384]) ? 1 : 0;
assign detect_min[547][2] = (mid_1[4391:4384] < top_0[4399:4392]) ? 1 : 0;
assign detect_min[547][3] = (mid_1[4391:4384] < top_1[4383:4376]) ? 1 : 0;
assign detect_min[547][4] = (mid_1[4391:4384] < top_1[4391:4384]) ? 1 : 0;
assign detect_min[547][5] = (mid_1[4391:4384] < top_1[4399:4392]) ? 1 : 0;
assign detect_min[547][6] = (mid_1[4391:4384] < top_2[4383:4376]) ? 1 : 0;
assign detect_min[547][7] = (mid_1[4391:4384] < top_2[4391:4384]) ? 1 : 0;
assign detect_min[547][8] = (mid_1[4391:4384] < top_2[4399:4392]) ? 1 : 0;
assign detect_min[547][9] = (mid_1[4391:4384] < mid_0[4383:4376]) ? 1 : 0;
assign detect_min[547][10] = (mid_1[4391:4384] < mid_0[4391:4384]) ? 1 : 0;
assign detect_min[547][11] = (mid_1[4391:4384] < mid_0[4399:4392]) ? 1 : 0;
assign detect_min[547][12] = (mid_1[4391:4384] < mid_1[4383:4376]) ? 1 : 0;
assign detect_min[547][13] = (mid_1[4391:4384] < mid_1[4399:4392]) ? 1 : 0;
assign detect_min[547][14] = (mid_1[4391:4384] < mid_2[4383:4376]) ? 1 : 0;
assign detect_min[547][15] = (mid_1[4391:4384] < mid_2[4391:4384]) ? 1 : 0;
assign detect_min[547][16] = (mid_1[4391:4384] < mid_2[4399:4392]) ? 1 : 0;
assign detect_min[547][17] = (mid_1[4391:4384] < btm_0[4383:4376]) ? 1 : 0;
assign detect_min[547][18] = (mid_1[4391:4384] < btm_0[4391:4384]) ? 1 : 0;
assign detect_min[547][19] = (mid_1[4391:4384] < btm_0[4399:4392]) ? 1 : 0;
assign detect_min[547][20] = (mid_1[4391:4384] < btm_1[4383:4376]) ? 1 : 0;
assign detect_min[547][21] = (mid_1[4391:4384] < btm_1[4391:4384]) ? 1 : 0;
assign detect_min[547][22] = (mid_1[4391:4384] < btm_1[4399:4392]) ? 1 : 0;
assign detect_min[547][23] = (mid_1[4391:4384] < btm_2[4383:4376]) ? 1 : 0;
assign detect_min[547][24] = (mid_1[4391:4384] < btm_2[4391:4384]) ? 1 : 0;
assign detect_min[547][25] = (mid_1[4391:4384] < btm_2[4399:4392]) ? 1 : 0;

assign detect_min[548][0] = (mid_1[4399:4392] < top_0[4391:4384]) ? 1 : 0;
assign detect_min[548][1] = (mid_1[4399:4392] < top_0[4399:4392]) ? 1 : 0;
assign detect_min[548][2] = (mid_1[4399:4392] < top_0[4407:4400]) ? 1 : 0;
assign detect_min[548][3] = (mid_1[4399:4392] < top_1[4391:4384]) ? 1 : 0;
assign detect_min[548][4] = (mid_1[4399:4392] < top_1[4399:4392]) ? 1 : 0;
assign detect_min[548][5] = (mid_1[4399:4392] < top_1[4407:4400]) ? 1 : 0;
assign detect_min[548][6] = (mid_1[4399:4392] < top_2[4391:4384]) ? 1 : 0;
assign detect_min[548][7] = (mid_1[4399:4392] < top_2[4399:4392]) ? 1 : 0;
assign detect_min[548][8] = (mid_1[4399:4392] < top_2[4407:4400]) ? 1 : 0;
assign detect_min[548][9] = (mid_1[4399:4392] < mid_0[4391:4384]) ? 1 : 0;
assign detect_min[548][10] = (mid_1[4399:4392] < mid_0[4399:4392]) ? 1 : 0;
assign detect_min[548][11] = (mid_1[4399:4392] < mid_0[4407:4400]) ? 1 : 0;
assign detect_min[548][12] = (mid_1[4399:4392] < mid_1[4391:4384]) ? 1 : 0;
assign detect_min[548][13] = (mid_1[4399:4392] < mid_1[4407:4400]) ? 1 : 0;
assign detect_min[548][14] = (mid_1[4399:4392] < mid_2[4391:4384]) ? 1 : 0;
assign detect_min[548][15] = (mid_1[4399:4392] < mid_2[4399:4392]) ? 1 : 0;
assign detect_min[548][16] = (mid_1[4399:4392] < mid_2[4407:4400]) ? 1 : 0;
assign detect_min[548][17] = (mid_1[4399:4392] < btm_0[4391:4384]) ? 1 : 0;
assign detect_min[548][18] = (mid_1[4399:4392] < btm_0[4399:4392]) ? 1 : 0;
assign detect_min[548][19] = (mid_1[4399:4392] < btm_0[4407:4400]) ? 1 : 0;
assign detect_min[548][20] = (mid_1[4399:4392] < btm_1[4391:4384]) ? 1 : 0;
assign detect_min[548][21] = (mid_1[4399:4392] < btm_1[4399:4392]) ? 1 : 0;
assign detect_min[548][22] = (mid_1[4399:4392] < btm_1[4407:4400]) ? 1 : 0;
assign detect_min[548][23] = (mid_1[4399:4392] < btm_2[4391:4384]) ? 1 : 0;
assign detect_min[548][24] = (mid_1[4399:4392] < btm_2[4399:4392]) ? 1 : 0;
assign detect_min[548][25] = (mid_1[4399:4392] < btm_2[4407:4400]) ? 1 : 0;

assign detect_min[549][0] = (mid_1[4407:4400] < top_0[4399:4392]) ? 1 : 0;
assign detect_min[549][1] = (mid_1[4407:4400] < top_0[4407:4400]) ? 1 : 0;
assign detect_min[549][2] = (mid_1[4407:4400] < top_0[4415:4408]) ? 1 : 0;
assign detect_min[549][3] = (mid_1[4407:4400] < top_1[4399:4392]) ? 1 : 0;
assign detect_min[549][4] = (mid_1[4407:4400] < top_1[4407:4400]) ? 1 : 0;
assign detect_min[549][5] = (mid_1[4407:4400] < top_1[4415:4408]) ? 1 : 0;
assign detect_min[549][6] = (mid_1[4407:4400] < top_2[4399:4392]) ? 1 : 0;
assign detect_min[549][7] = (mid_1[4407:4400] < top_2[4407:4400]) ? 1 : 0;
assign detect_min[549][8] = (mid_1[4407:4400] < top_2[4415:4408]) ? 1 : 0;
assign detect_min[549][9] = (mid_1[4407:4400] < mid_0[4399:4392]) ? 1 : 0;
assign detect_min[549][10] = (mid_1[4407:4400] < mid_0[4407:4400]) ? 1 : 0;
assign detect_min[549][11] = (mid_1[4407:4400] < mid_0[4415:4408]) ? 1 : 0;
assign detect_min[549][12] = (mid_1[4407:4400] < mid_1[4399:4392]) ? 1 : 0;
assign detect_min[549][13] = (mid_1[4407:4400] < mid_1[4415:4408]) ? 1 : 0;
assign detect_min[549][14] = (mid_1[4407:4400] < mid_2[4399:4392]) ? 1 : 0;
assign detect_min[549][15] = (mid_1[4407:4400] < mid_2[4407:4400]) ? 1 : 0;
assign detect_min[549][16] = (mid_1[4407:4400] < mid_2[4415:4408]) ? 1 : 0;
assign detect_min[549][17] = (mid_1[4407:4400] < btm_0[4399:4392]) ? 1 : 0;
assign detect_min[549][18] = (mid_1[4407:4400] < btm_0[4407:4400]) ? 1 : 0;
assign detect_min[549][19] = (mid_1[4407:4400] < btm_0[4415:4408]) ? 1 : 0;
assign detect_min[549][20] = (mid_1[4407:4400] < btm_1[4399:4392]) ? 1 : 0;
assign detect_min[549][21] = (mid_1[4407:4400] < btm_1[4407:4400]) ? 1 : 0;
assign detect_min[549][22] = (mid_1[4407:4400] < btm_1[4415:4408]) ? 1 : 0;
assign detect_min[549][23] = (mid_1[4407:4400] < btm_2[4399:4392]) ? 1 : 0;
assign detect_min[549][24] = (mid_1[4407:4400] < btm_2[4407:4400]) ? 1 : 0;
assign detect_min[549][25] = (mid_1[4407:4400] < btm_2[4415:4408]) ? 1 : 0;

assign detect_min[550][0] = (mid_1[4415:4408] < top_0[4407:4400]) ? 1 : 0;
assign detect_min[550][1] = (mid_1[4415:4408] < top_0[4415:4408]) ? 1 : 0;
assign detect_min[550][2] = (mid_1[4415:4408] < top_0[4423:4416]) ? 1 : 0;
assign detect_min[550][3] = (mid_1[4415:4408] < top_1[4407:4400]) ? 1 : 0;
assign detect_min[550][4] = (mid_1[4415:4408] < top_1[4415:4408]) ? 1 : 0;
assign detect_min[550][5] = (mid_1[4415:4408] < top_1[4423:4416]) ? 1 : 0;
assign detect_min[550][6] = (mid_1[4415:4408] < top_2[4407:4400]) ? 1 : 0;
assign detect_min[550][7] = (mid_1[4415:4408] < top_2[4415:4408]) ? 1 : 0;
assign detect_min[550][8] = (mid_1[4415:4408] < top_2[4423:4416]) ? 1 : 0;
assign detect_min[550][9] = (mid_1[4415:4408] < mid_0[4407:4400]) ? 1 : 0;
assign detect_min[550][10] = (mid_1[4415:4408] < mid_0[4415:4408]) ? 1 : 0;
assign detect_min[550][11] = (mid_1[4415:4408] < mid_0[4423:4416]) ? 1 : 0;
assign detect_min[550][12] = (mid_1[4415:4408] < mid_1[4407:4400]) ? 1 : 0;
assign detect_min[550][13] = (mid_1[4415:4408] < mid_1[4423:4416]) ? 1 : 0;
assign detect_min[550][14] = (mid_1[4415:4408] < mid_2[4407:4400]) ? 1 : 0;
assign detect_min[550][15] = (mid_1[4415:4408] < mid_2[4415:4408]) ? 1 : 0;
assign detect_min[550][16] = (mid_1[4415:4408] < mid_2[4423:4416]) ? 1 : 0;
assign detect_min[550][17] = (mid_1[4415:4408] < btm_0[4407:4400]) ? 1 : 0;
assign detect_min[550][18] = (mid_1[4415:4408] < btm_0[4415:4408]) ? 1 : 0;
assign detect_min[550][19] = (mid_1[4415:4408] < btm_0[4423:4416]) ? 1 : 0;
assign detect_min[550][20] = (mid_1[4415:4408] < btm_1[4407:4400]) ? 1 : 0;
assign detect_min[550][21] = (mid_1[4415:4408] < btm_1[4415:4408]) ? 1 : 0;
assign detect_min[550][22] = (mid_1[4415:4408] < btm_1[4423:4416]) ? 1 : 0;
assign detect_min[550][23] = (mid_1[4415:4408] < btm_2[4407:4400]) ? 1 : 0;
assign detect_min[550][24] = (mid_1[4415:4408] < btm_2[4415:4408]) ? 1 : 0;
assign detect_min[550][25] = (mid_1[4415:4408] < btm_2[4423:4416]) ? 1 : 0;

assign detect_min[551][0] = (mid_1[4423:4416] < top_0[4415:4408]) ? 1 : 0;
assign detect_min[551][1] = (mid_1[4423:4416] < top_0[4423:4416]) ? 1 : 0;
assign detect_min[551][2] = (mid_1[4423:4416] < top_0[4431:4424]) ? 1 : 0;
assign detect_min[551][3] = (mid_1[4423:4416] < top_1[4415:4408]) ? 1 : 0;
assign detect_min[551][4] = (mid_1[4423:4416] < top_1[4423:4416]) ? 1 : 0;
assign detect_min[551][5] = (mid_1[4423:4416] < top_1[4431:4424]) ? 1 : 0;
assign detect_min[551][6] = (mid_1[4423:4416] < top_2[4415:4408]) ? 1 : 0;
assign detect_min[551][7] = (mid_1[4423:4416] < top_2[4423:4416]) ? 1 : 0;
assign detect_min[551][8] = (mid_1[4423:4416] < top_2[4431:4424]) ? 1 : 0;
assign detect_min[551][9] = (mid_1[4423:4416] < mid_0[4415:4408]) ? 1 : 0;
assign detect_min[551][10] = (mid_1[4423:4416] < mid_0[4423:4416]) ? 1 : 0;
assign detect_min[551][11] = (mid_1[4423:4416] < mid_0[4431:4424]) ? 1 : 0;
assign detect_min[551][12] = (mid_1[4423:4416] < mid_1[4415:4408]) ? 1 : 0;
assign detect_min[551][13] = (mid_1[4423:4416] < mid_1[4431:4424]) ? 1 : 0;
assign detect_min[551][14] = (mid_1[4423:4416] < mid_2[4415:4408]) ? 1 : 0;
assign detect_min[551][15] = (mid_1[4423:4416] < mid_2[4423:4416]) ? 1 : 0;
assign detect_min[551][16] = (mid_1[4423:4416] < mid_2[4431:4424]) ? 1 : 0;
assign detect_min[551][17] = (mid_1[4423:4416] < btm_0[4415:4408]) ? 1 : 0;
assign detect_min[551][18] = (mid_1[4423:4416] < btm_0[4423:4416]) ? 1 : 0;
assign detect_min[551][19] = (mid_1[4423:4416] < btm_0[4431:4424]) ? 1 : 0;
assign detect_min[551][20] = (mid_1[4423:4416] < btm_1[4415:4408]) ? 1 : 0;
assign detect_min[551][21] = (mid_1[4423:4416] < btm_1[4423:4416]) ? 1 : 0;
assign detect_min[551][22] = (mid_1[4423:4416] < btm_1[4431:4424]) ? 1 : 0;
assign detect_min[551][23] = (mid_1[4423:4416] < btm_2[4415:4408]) ? 1 : 0;
assign detect_min[551][24] = (mid_1[4423:4416] < btm_2[4423:4416]) ? 1 : 0;
assign detect_min[551][25] = (mid_1[4423:4416] < btm_2[4431:4424]) ? 1 : 0;

assign detect_min[552][0] = (mid_1[4431:4424] < top_0[4423:4416]) ? 1 : 0;
assign detect_min[552][1] = (mid_1[4431:4424] < top_0[4431:4424]) ? 1 : 0;
assign detect_min[552][2] = (mid_1[4431:4424] < top_0[4439:4432]) ? 1 : 0;
assign detect_min[552][3] = (mid_1[4431:4424] < top_1[4423:4416]) ? 1 : 0;
assign detect_min[552][4] = (mid_1[4431:4424] < top_1[4431:4424]) ? 1 : 0;
assign detect_min[552][5] = (mid_1[4431:4424] < top_1[4439:4432]) ? 1 : 0;
assign detect_min[552][6] = (mid_1[4431:4424] < top_2[4423:4416]) ? 1 : 0;
assign detect_min[552][7] = (mid_1[4431:4424] < top_2[4431:4424]) ? 1 : 0;
assign detect_min[552][8] = (mid_1[4431:4424] < top_2[4439:4432]) ? 1 : 0;
assign detect_min[552][9] = (mid_1[4431:4424] < mid_0[4423:4416]) ? 1 : 0;
assign detect_min[552][10] = (mid_1[4431:4424] < mid_0[4431:4424]) ? 1 : 0;
assign detect_min[552][11] = (mid_1[4431:4424] < mid_0[4439:4432]) ? 1 : 0;
assign detect_min[552][12] = (mid_1[4431:4424] < mid_1[4423:4416]) ? 1 : 0;
assign detect_min[552][13] = (mid_1[4431:4424] < mid_1[4439:4432]) ? 1 : 0;
assign detect_min[552][14] = (mid_1[4431:4424] < mid_2[4423:4416]) ? 1 : 0;
assign detect_min[552][15] = (mid_1[4431:4424] < mid_2[4431:4424]) ? 1 : 0;
assign detect_min[552][16] = (mid_1[4431:4424] < mid_2[4439:4432]) ? 1 : 0;
assign detect_min[552][17] = (mid_1[4431:4424] < btm_0[4423:4416]) ? 1 : 0;
assign detect_min[552][18] = (mid_1[4431:4424] < btm_0[4431:4424]) ? 1 : 0;
assign detect_min[552][19] = (mid_1[4431:4424] < btm_0[4439:4432]) ? 1 : 0;
assign detect_min[552][20] = (mid_1[4431:4424] < btm_1[4423:4416]) ? 1 : 0;
assign detect_min[552][21] = (mid_1[4431:4424] < btm_1[4431:4424]) ? 1 : 0;
assign detect_min[552][22] = (mid_1[4431:4424] < btm_1[4439:4432]) ? 1 : 0;
assign detect_min[552][23] = (mid_1[4431:4424] < btm_2[4423:4416]) ? 1 : 0;
assign detect_min[552][24] = (mid_1[4431:4424] < btm_2[4431:4424]) ? 1 : 0;
assign detect_min[552][25] = (mid_1[4431:4424] < btm_2[4439:4432]) ? 1 : 0;

assign detect_min[553][0] = (mid_1[4439:4432] < top_0[4431:4424]) ? 1 : 0;
assign detect_min[553][1] = (mid_1[4439:4432] < top_0[4439:4432]) ? 1 : 0;
assign detect_min[553][2] = (mid_1[4439:4432] < top_0[4447:4440]) ? 1 : 0;
assign detect_min[553][3] = (mid_1[4439:4432] < top_1[4431:4424]) ? 1 : 0;
assign detect_min[553][4] = (mid_1[4439:4432] < top_1[4439:4432]) ? 1 : 0;
assign detect_min[553][5] = (mid_1[4439:4432] < top_1[4447:4440]) ? 1 : 0;
assign detect_min[553][6] = (mid_1[4439:4432] < top_2[4431:4424]) ? 1 : 0;
assign detect_min[553][7] = (mid_1[4439:4432] < top_2[4439:4432]) ? 1 : 0;
assign detect_min[553][8] = (mid_1[4439:4432] < top_2[4447:4440]) ? 1 : 0;
assign detect_min[553][9] = (mid_1[4439:4432] < mid_0[4431:4424]) ? 1 : 0;
assign detect_min[553][10] = (mid_1[4439:4432] < mid_0[4439:4432]) ? 1 : 0;
assign detect_min[553][11] = (mid_1[4439:4432] < mid_0[4447:4440]) ? 1 : 0;
assign detect_min[553][12] = (mid_1[4439:4432] < mid_1[4431:4424]) ? 1 : 0;
assign detect_min[553][13] = (mid_1[4439:4432] < mid_1[4447:4440]) ? 1 : 0;
assign detect_min[553][14] = (mid_1[4439:4432] < mid_2[4431:4424]) ? 1 : 0;
assign detect_min[553][15] = (mid_1[4439:4432] < mid_2[4439:4432]) ? 1 : 0;
assign detect_min[553][16] = (mid_1[4439:4432] < mid_2[4447:4440]) ? 1 : 0;
assign detect_min[553][17] = (mid_1[4439:4432] < btm_0[4431:4424]) ? 1 : 0;
assign detect_min[553][18] = (mid_1[4439:4432] < btm_0[4439:4432]) ? 1 : 0;
assign detect_min[553][19] = (mid_1[4439:4432] < btm_0[4447:4440]) ? 1 : 0;
assign detect_min[553][20] = (mid_1[4439:4432] < btm_1[4431:4424]) ? 1 : 0;
assign detect_min[553][21] = (mid_1[4439:4432] < btm_1[4439:4432]) ? 1 : 0;
assign detect_min[553][22] = (mid_1[4439:4432] < btm_1[4447:4440]) ? 1 : 0;
assign detect_min[553][23] = (mid_1[4439:4432] < btm_2[4431:4424]) ? 1 : 0;
assign detect_min[553][24] = (mid_1[4439:4432] < btm_2[4439:4432]) ? 1 : 0;
assign detect_min[553][25] = (mid_1[4439:4432] < btm_2[4447:4440]) ? 1 : 0;

assign detect_min[554][0] = (mid_1[4447:4440] < top_0[4439:4432]) ? 1 : 0;
assign detect_min[554][1] = (mid_1[4447:4440] < top_0[4447:4440]) ? 1 : 0;
assign detect_min[554][2] = (mid_1[4447:4440] < top_0[4455:4448]) ? 1 : 0;
assign detect_min[554][3] = (mid_1[4447:4440] < top_1[4439:4432]) ? 1 : 0;
assign detect_min[554][4] = (mid_1[4447:4440] < top_1[4447:4440]) ? 1 : 0;
assign detect_min[554][5] = (mid_1[4447:4440] < top_1[4455:4448]) ? 1 : 0;
assign detect_min[554][6] = (mid_1[4447:4440] < top_2[4439:4432]) ? 1 : 0;
assign detect_min[554][7] = (mid_1[4447:4440] < top_2[4447:4440]) ? 1 : 0;
assign detect_min[554][8] = (mid_1[4447:4440] < top_2[4455:4448]) ? 1 : 0;
assign detect_min[554][9] = (mid_1[4447:4440] < mid_0[4439:4432]) ? 1 : 0;
assign detect_min[554][10] = (mid_1[4447:4440] < mid_0[4447:4440]) ? 1 : 0;
assign detect_min[554][11] = (mid_1[4447:4440] < mid_0[4455:4448]) ? 1 : 0;
assign detect_min[554][12] = (mid_1[4447:4440] < mid_1[4439:4432]) ? 1 : 0;
assign detect_min[554][13] = (mid_1[4447:4440] < mid_1[4455:4448]) ? 1 : 0;
assign detect_min[554][14] = (mid_1[4447:4440] < mid_2[4439:4432]) ? 1 : 0;
assign detect_min[554][15] = (mid_1[4447:4440] < mid_2[4447:4440]) ? 1 : 0;
assign detect_min[554][16] = (mid_1[4447:4440] < mid_2[4455:4448]) ? 1 : 0;
assign detect_min[554][17] = (mid_1[4447:4440] < btm_0[4439:4432]) ? 1 : 0;
assign detect_min[554][18] = (mid_1[4447:4440] < btm_0[4447:4440]) ? 1 : 0;
assign detect_min[554][19] = (mid_1[4447:4440] < btm_0[4455:4448]) ? 1 : 0;
assign detect_min[554][20] = (mid_1[4447:4440] < btm_1[4439:4432]) ? 1 : 0;
assign detect_min[554][21] = (mid_1[4447:4440] < btm_1[4447:4440]) ? 1 : 0;
assign detect_min[554][22] = (mid_1[4447:4440] < btm_1[4455:4448]) ? 1 : 0;
assign detect_min[554][23] = (mid_1[4447:4440] < btm_2[4439:4432]) ? 1 : 0;
assign detect_min[554][24] = (mid_1[4447:4440] < btm_2[4447:4440]) ? 1 : 0;
assign detect_min[554][25] = (mid_1[4447:4440] < btm_2[4455:4448]) ? 1 : 0;

assign detect_min[555][0] = (mid_1[4455:4448] < top_0[4447:4440]) ? 1 : 0;
assign detect_min[555][1] = (mid_1[4455:4448] < top_0[4455:4448]) ? 1 : 0;
assign detect_min[555][2] = (mid_1[4455:4448] < top_0[4463:4456]) ? 1 : 0;
assign detect_min[555][3] = (mid_1[4455:4448] < top_1[4447:4440]) ? 1 : 0;
assign detect_min[555][4] = (mid_1[4455:4448] < top_1[4455:4448]) ? 1 : 0;
assign detect_min[555][5] = (mid_1[4455:4448] < top_1[4463:4456]) ? 1 : 0;
assign detect_min[555][6] = (mid_1[4455:4448] < top_2[4447:4440]) ? 1 : 0;
assign detect_min[555][7] = (mid_1[4455:4448] < top_2[4455:4448]) ? 1 : 0;
assign detect_min[555][8] = (mid_1[4455:4448] < top_2[4463:4456]) ? 1 : 0;
assign detect_min[555][9] = (mid_1[4455:4448] < mid_0[4447:4440]) ? 1 : 0;
assign detect_min[555][10] = (mid_1[4455:4448] < mid_0[4455:4448]) ? 1 : 0;
assign detect_min[555][11] = (mid_1[4455:4448] < mid_0[4463:4456]) ? 1 : 0;
assign detect_min[555][12] = (mid_1[4455:4448] < mid_1[4447:4440]) ? 1 : 0;
assign detect_min[555][13] = (mid_1[4455:4448] < mid_1[4463:4456]) ? 1 : 0;
assign detect_min[555][14] = (mid_1[4455:4448] < mid_2[4447:4440]) ? 1 : 0;
assign detect_min[555][15] = (mid_1[4455:4448] < mid_2[4455:4448]) ? 1 : 0;
assign detect_min[555][16] = (mid_1[4455:4448] < mid_2[4463:4456]) ? 1 : 0;
assign detect_min[555][17] = (mid_1[4455:4448] < btm_0[4447:4440]) ? 1 : 0;
assign detect_min[555][18] = (mid_1[4455:4448] < btm_0[4455:4448]) ? 1 : 0;
assign detect_min[555][19] = (mid_1[4455:4448] < btm_0[4463:4456]) ? 1 : 0;
assign detect_min[555][20] = (mid_1[4455:4448] < btm_1[4447:4440]) ? 1 : 0;
assign detect_min[555][21] = (mid_1[4455:4448] < btm_1[4455:4448]) ? 1 : 0;
assign detect_min[555][22] = (mid_1[4455:4448] < btm_1[4463:4456]) ? 1 : 0;
assign detect_min[555][23] = (mid_1[4455:4448] < btm_2[4447:4440]) ? 1 : 0;
assign detect_min[555][24] = (mid_1[4455:4448] < btm_2[4455:4448]) ? 1 : 0;
assign detect_min[555][25] = (mid_1[4455:4448] < btm_2[4463:4456]) ? 1 : 0;

assign detect_min[556][0] = (mid_1[4463:4456] < top_0[4455:4448]) ? 1 : 0;
assign detect_min[556][1] = (mid_1[4463:4456] < top_0[4463:4456]) ? 1 : 0;
assign detect_min[556][2] = (mid_1[4463:4456] < top_0[4471:4464]) ? 1 : 0;
assign detect_min[556][3] = (mid_1[4463:4456] < top_1[4455:4448]) ? 1 : 0;
assign detect_min[556][4] = (mid_1[4463:4456] < top_1[4463:4456]) ? 1 : 0;
assign detect_min[556][5] = (mid_1[4463:4456] < top_1[4471:4464]) ? 1 : 0;
assign detect_min[556][6] = (mid_1[4463:4456] < top_2[4455:4448]) ? 1 : 0;
assign detect_min[556][7] = (mid_1[4463:4456] < top_2[4463:4456]) ? 1 : 0;
assign detect_min[556][8] = (mid_1[4463:4456] < top_2[4471:4464]) ? 1 : 0;
assign detect_min[556][9] = (mid_1[4463:4456] < mid_0[4455:4448]) ? 1 : 0;
assign detect_min[556][10] = (mid_1[4463:4456] < mid_0[4463:4456]) ? 1 : 0;
assign detect_min[556][11] = (mid_1[4463:4456] < mid_0[4471:4464]) ? 1 : 0;
assign detect_min[556][12] = (mid_1[4463:4456] < mid_1[4455:4448]) ? 1 : 0;
assign detect_min[556][13] = (mid_1[4463:4456] < mid_1[4471:4464]) ? 1 : 0;
assign detect_min[556][14] = (mid_1[4463:4456] < mid_2[4455:4448]) ? 1 : 0;
assign detect_min[556][15] = (mid_1[4463:4456] < mid_2[4463:4456]) ? 1 : 0;
assign detect_min[556][16] = (mid_1[4463:4456] < mid_2[4471:4464]) ? 1 : 0;
assign detect_min[556][17] = (mid_1[4463:4456] < btm_0[4455:4448]) ? 1 : 0;
assign detect_min[556][18] = (mid_1[4463:4456] < btm_0[4463:4456]) ? 1 : 0;
assign detect_min[556][19] = (mid_1[4463:4456] < btm_0[4471:4464]) ? 1 : 0;
assign detect_min[556][20] = (mid_1[4463:4456] < btm_1[4455:4448]) ? 1 : 0;
assign detect_min[556][21] = (mid_1[4463:4456] < btm_1[4463:4456]) ? 1 : 0;
assign detect_min[556][22] = (mid_1[4463:4456] < btm_1[4471:4464]) ? 1 : 0;
assign detect_min[556][23] = (mid_1[4463:4456] < btm_2[4455:4448]) ? 1 : 0;
assign detect_min[556][24] = (mid_1[4463:4456] < btm_2[4463:4456]) ? 1 : 0;
assign detect_min[556][25] = (mid_1[4463:4456] < btm_2[4471:4464]) ? 1 : 0;

assign detect_min[557][0] = (mid_1[4471:4464] < top_0[4463:4456]) ? 1 : 0;
assign detect_min[557][1] = (mid_1[4471:4464] < top_0[4471:4464]) ? 1 : 0;
assign detect_min[557][2] = (mid_1[4471:4464] < top_0[4479:4472]) ? 1 : 0;
assign detect_min[557][3] = (mid_1[4471:4464] < top_1[4463:4456]) ? 1 : 0;
assign detect_min[557][4] = (mid_1[4471:4464] < top_1[4471:4464]) ? 1 : 0;
assign detect_min[557][5] = (mid_1[4471:4464] < top_1[4479:4472]) ? 1 : 0;
assign detect_min[557][6] = (mid_1[4471:4464] < top_2[4463:4456]) ? 1 : 0;
assign detect_min[557][7] = (mid_1[4471:4464] < top_2[4471:4464]) ? 1 : 0;
assign detect_min[557][8] = (mid_1[4471:4464] < top_2[4479:4472]) ? 1 : 0;
assign detect_min[557][9] = (mid_1[4471:4464] < mid_0[4463:4456]) ? 1 : 0;
assign detect_min[557][10] = (mid_1[4471:4464] < mid_0[4471:4464]) ? 1 : 0;
assign detect_min[557][11] = (mid_1[4471:4464] < mid_0[4479:4472]) ? 1 : 0;
assign detect_min[557][12] = (mid_1[4471:4464] < mid_1[4463:4456]) ? 1 : 0;
assign detect_min[557][13] = (mid_1[4471:4464] < mid_1[4479:4472]) ? 1 : 0;
assign detect_min[557][14] = (mid_1[4471:4464] < mid_2[4463:4456]) ? 1 : 0;
assign detect_min[557][15] = (mid_1[4471:4464] < mid_2[4471:4464]) ? 1 : 0;
assign detect_min[557][16] = (mid_1[4471:4464] < mid_2[4479:4472]) ? 1 : 0;
assign detect_min[557][17] = (mid_1[4471:4464] < btm_0[4463:4456]) ? 1 : 0;
assign detect_min[557][18] = (mid_1[4471:4464] < btm_0[4471:4464]) ? 1 : 0;
assign detect_min[557][19] = (mid_1[4471:4464] < btm_0[4479:4472]) ? 1 : 0;
assign detect_min[557][20] = (mid_1[4471:4464] < btm_1[4463:4456]) ? 1 : 0;
assign detect_min[557][21] = (mid_1[4471:4464] < btm_1[4471:4464]) ? 1 : 0;
assign detect_min[557][22] = (mid_1[4471:4464] < btm_1[4479:4472]) ? 1 : 0;
assign detect_min[557][23] = (mid_1[4471:4464] < btm_2[4463:4456]) ? 1 : 0;
assign detect_min[557][24] = (mid_1[4471:4464] < btm_2[4471:4464]) ? 1 : 0;
assign detect_min[557][25] = (mid_1[4471:4464] < btm_2[4479:4472]) ? 1 : 0;

assign detect_min[558][0] = (mid_1[4479:4472] < top_0[4471:4464]) ? 1 : 0;
assign detect_min[558][1] = (mid_1[4479:4472] < top_0[4479:4472]) ? 1 : 0;
assign detect_min[558][2] = (mid_1[4479:4472] < top_0[4487:4480]) ? 1 : 0;
assign detect_min[558][3] = (mid_1[4479:4472] < top_1[4471:4464]) ? 1 : 0;
assign detect_min[558][4] = (mid_1[4479:4472] < top_1[4479:4472]) ? 1 : 0;
assign detect_min[558][5] = (mid_1[4479:4472] < top_1[4487:4480]) ? 1 : 0;
assign detect_min[558][6] = (mid_1[4479:4472] < top_2[4471:4464]) ? 1 : 0;
assign detect_min[558][7] = (mid_1[4479:4472] < top_2[4479:4472]) ? 1 : 0;
assign detect_min[558][8] = (mid_1[4479:4472] < top_2[4487:4480]) ? 1 : 0;
assign detect_min[558][9] = (mid_1[4479:4472] < mid_0[4471:4464]) ? 1 : 0;
assign detect_min[558][10] = (mid_1[4479:4472] < mid_0[4479:4472]) ? 1 : 0;
assign detect_min[558][11] = (mid_1[4479:4472] < mid_0[4487:4480]) ? 1 : 0;
assign detect_min[558][12] = (mid_1[4479:4472] < mid_1[4471:4464]) ? 1 : 0;
assign detect_min[558][13] = (mid_1[4479:4472] < mid_1[4487:4480]) ? 1 : 0;
assign detect_min[558][14] = (mid_1[4479:4472] < mid_2[4471:4464]) ? 1 : 0;
assign detect_min[558][15] = (mid_1[4479:4472] < mid_2[4479:4472]) ? 1 : 0;
assign detect_min[558][16] = (mid_1[4479:4472] < mid_2[4487:4480]) ? 1 : 0;
assign detect_min[558][17] = (mid_1[4479:4472] < btm_0[4471:4464]) ? 1 : 0;
assign detect_min[558][18] = (mid_1[4479:4472] < btm_0[4479:4472]) ? 1 : 0;
assign detect_min[558][19] = (mid_1[4479:4472] < btm_0[4487:4480]) ? 1 : 0;
assign detect_min[558][20] = (mid_1[4479:4472] < btm_1[4471:4464]) ? 1 : 0;
assign detect_min[558][21] = (mid_1[4479:4472] < btm_1[4479:4472]) ? 1 : 0;
assign detect_min[558][22] = (mid_1[4479:4472] < btm_1[4487:4480]) ? 1 : 0;
assign detect_min[558][23] = (mid_1[4479:4472] < btm_2[4471:4464]) ? 1 : 0;
assign detect_min[558][24] = (mid_1[4479:4472] < btm_2[4479:4472]) ? 1 : 0;
assign detect_min[558][25] = (mid_1[4479:4472] < btm_2[4487:4480]) ? 1 : 0;

assign detect_min[559][0] = (mid_1[4487:4480] < top_0[4479:4472]) ? 1 : 0;
assign detect_min[559][1] = (mid_1[4487:4480] < top_0[4487:4480]) ? 1 : 0;
assign detect_min[559][2] = (mid_1[4487:4480] < top_0[4495:4488]) ? 1 : 0;
assign detect_min[559][3] = (mid_1[4487:4480] < top_1[4479:4472]) ? 1 : 0;
assign detect_min[559][4] = (mid_1[4487:4480] < top_1[4487:4480]) ? 1 : 0;
assign detect_min[559][5] = (mid_1[4487:4480] < top_1[4495:4488]) ? 1 : 0;
assign detect_min[559][6] = (mid_1[4487:4480] < top_2[4479:4472]) ? 1 : 0;
assign detect_min[559][7] = (mid_1[4487:4480] < top_2[4487:4480]) ? 1 : 0;
assign detect_min[559][8] = (mid_1[4487:4480] < top_2[4495:4488]) ? 1 : 0;
assign detect_min[559][9] = (mid_1[4487:4480] < mid_0[4479:4472]) ? 1 : 0;
assign detect_min[559][10] = (mid_1[4487:4480] < mid_0[4487:4480]) ? 1 : 0;
assign detect_min[559][11] = (mid_1[4487:4480] < mid_0[4495:4488]) ? 1 : 0;
assign detect_min[559][12] = (mid_1[4487:4480] < mid_1[4479:4472]) ? 1 : 0;
assign detect_min[559][13] = (mid_1[4487:4480] < mid_1[4495:4488]) ? 1 : 0;
assign detect_min[559][14] = (mid_1[4487:4480] < mid_2[4479:4472]) ? 1 : 0;
assign detect_min[559][15] = (mid_1[4487:4480] < mid_2[4487:4480]) ? 1 : 0;
assign detect_min[559][16] = (mid_1[4487:4480] < mid_2[4495:4488]) ? 1 : 0;
assign detect_min[559][17] = (mid_1[4487:4480] < btm_0[4479:4472]) ? 1 : 0;
assign detect_min[559][18] = (mid_1[4487:4480] < btm_0[4487:4480]) ? 1 : 0;
assign detect_min[559][19] = (mid_1[4487:4480] < btm_0[4495:4488]) ? 1 : 0;
assign detect_min[559][20] = (mid_1[4487:4480] < btm_1[4479:4472]) ? 1 : 0;
assign detect_min[559][21] = (mid_1[4487:4480] < btm_1[4487:4480]) ? 1 : 0;
assign detect_min[559][22] = (mid_1[4487:4480] < btm_1[4495:4488]) ? 1 : 0;
assign detect_min[559][23] = (mid_1[4487:4480] < btm_2[4479:4472]) ? 1 : 0;
assign detect_min[559][24] = (mid_1[4487:4480] < btm_2[4487:4480]) ? 1 : 0;
assign detect_min[559][25] = (mid_1[4487:4480] < btm_2[4495:4488]) ? 1 : 0;

assign detect_min[560][0] = (mid_1[4495:4488] < top_0[4487:4480]) ? 1 : 0;
assign detect_min[560][1] = (mid_1[4495:4488] < top_0[4495:4488]) ? 1 : 0;
assign detect_min[560][2] = (mid_1[4495:4488] < top_0[4503:4496]) ? 1 : 0;
assign detect_min[560][3] = (mid_1[4495:4488] < top_1[4487:4480]) ? 1 : 0;
assign detect_min[560][4] = (mid_1[4495:4488] < top_1[4495:4488]) ? 1 : 0;
assign detect_min[560][5] = (mid_1[4495:4488] < top_1[4503:4496]) ? 1 : 0;
assign detect_min[560][6] = (mid_1[4495:4488] < top_2[4487:4480]) ? 1 : 0;
assign detect_min[560][7] = (mid_1[4495:4488] < top_2[4495:4488]) ? 1 : 0;
assign detect_min[560][8] = (mid_1[4495:4488] < top_2[4503:4496]) ? 1 : 0;
assign detect_min[560][9] = (mid_1[4495:4488] < mid_0[4487:4480]) ? 1 : 0;
assign detect_min[560][10] = (mid_1[4495:4488] < mid_0[4495:4488]) ? 1 : 0;
assign detect_min[560][11] = (mid_1[4495:4488] < mid_0[4503:4496]) ? 1 : 0;
assign detect_min[560][12] = (mid_1[4495:4488] < mid_1[4487:4480]) ? 1 : 0;
assign detect_min[560][13] = (mid_1[4495:4488] < mid_1[4503:4496]) ? 1 : 0;
assign detect_min[560][14] = (mid_1[4495:4488] < mid_2[4487:4480]) ? 1 : 0;
assign detect_min[560][15] = (mid_1[4495:4488] < mid_2[4495:4488]) ? 1 : 0;
assign detect_min[560][16] = (mid_1[4495:4488] < mid_2[4503:4496]) ? 1 : 0;
assign detect_min[560][17] = (mid_1[4495:4488] < btm_0[4487:4480]) ? 1 : 0;
assign detect_min[560][18] = (mid_1[4495:4488] < btm_0[4495:4488]) ? 1 : 0;
assign detect_min[560][19] = (mid_1[4495:4488] < btm_0[4503:4496]) ? 1 : 0;
assign detect_min[560][20] = (mid_1[4495:4488] < btm_1[4487:4480]) ? 1 : 0;
assign detect_min[560][21] = (mid_1[4495:4488] < btm_1[4495:4488]) ? 1 : 0;
assign detect_min[560][22] = (mid_1[4495:4488] < btm_1[4503:4496]) ? 1 : 0;
assign detect_min[560][23] = (mid_1[4495:4488] < btm_2[4487:4480]) ? 1 : 0;
assign detect_min[560][24] = (mid_1[4495:4488] < btm_2[4495:4488]) ? 1 : 0;
assign detect_min[560][25] = (mid_1[4495:4488] < btm_2[4503:4496]) ? 1 : 0;

assign detect_min[561][0] = (mid_1[4503:4496] < top_0[4495:4488]) ? 1 : 0;
assign detect_min[561][1] = (mid_1[4503:4496] < top_0[4503:4496]) ? 1 : 0;
assign detect_min[561][2] = (mid_1[4503:4496] < top_0[4511:4504]) ? 1 : 0;
assign detect_min[561][3] = (mid_1[4503:4496] < top_1[4495:4488]) ? 1 : 0;
assign detect_min[561][4] = (mid_1[4503:4496] < top_1[4503:4496]) ? 1 : 0;
assign detect_min[561][5] = (mid_1[4503:4496] < top_1[4511:4504]) ? 1 : 0;
assign detect_min[561][6] = (mid_1[4503:4496] < top_2[4495:4488]) ? 1 : 0;
assign detect_min[561][7] = (mid_1[4503:4496] < top_2[4503:4496]) ? 1 : 0;
assign detect_min[561][8] = (mid_1[4503:4496] < top_2[4511:4504]) ? 1 : 0;
assign detect_min[561][9] = (mid_1[4503:4496] < mid_0[4495:4488]) ? 1 : 0;
assign detect_min[561][10] = (mid_1[4503:4496] < mid_0[4503:4496]) ? 1 : 0;
assign detect_min[561][11] = (mid_1[4503:4496] < mid_0[4511:4504]) ? 1 : 0;
assign detect_min[561][12] = (mid_1[4503:4496] < mid_1[4495:4488]) ? 1 : 0;
assign detect_min[561][13] = (mid_1[4503:4496] < mid_1[4511:4504]) ? 1 : 0;
assign detect_min[561][14] = (mid_1[4503:4496] < mid_2[4495:4488]) ? 1 : 0;
assign detect_min[561][15] = (mid_1[4503:4496] < mid_2[4503:4496]) ? 1 : 0;
assign detect_min[561][16] = (mid_1[4503:4496] < mid_2[4511:4504]) ? 1 : 0;
assign detect_min[561][17] = (mid_1[4503:4496] < btm_0[4495:4488]) ? 1 : 0;
assign detect_min[561][18] = (mid_1[4503:4496] < btm_0[4503:4496]) ? 1 : 0;
assign detect_min[561][19] = (mid_1[4503:4496] < btm_0[4511:4504]) ? 1 : 0;
assign detect_min[561][20] = (mid_1[4503:4496] < btm_1[4495:4488]) ? 1 : 0;
assign detect_min[561][21] = (mid_1[4503:4496] < btm_1[4503:4496]) ? 1 : 0;
assign detect_min[561][22] = (mid_1[4503:4496] < btm_1[4511:4504]) ? 1 : 0;
assign detect_min[561][23] = (mid_1[4503:4496] < btm_2[4495:4488]) ? 1 : 0;
assign detect_min[561][24] = (mid_1[4503:4496] < btm_2[4503:4496]) ? 1 : 0;
assign detect_min[561][25] = (mid_1[4503:4496] < btm_2[4511:4504]) ? 1 : 0;

assign detect_min[562][0] = (mid_1[4511:4504] < top_0[4503:4496]) ? 1 : 0;
assign detect_min[562][1] = (mid_1[4511:4504] < top_0[4511:4504]) ? 1 : 0;
assign detect_min[562][2] = (mid_1[4511:4504] < top_0[4519:4512]) ? 1 : 0;
assign detect_min[562][3] = (mid_1[4511:4504] < top_1[4503:4496]) ? 1 : 0;
assign detect_min[562][4] = (mid_1[4511:4504] < top_1[4511:4504]) ? 1 : 0;
assign detect_min[562][5] = (mid_1[4511:4504] < top_1[4519:4512]) ? 1 : 0;
assign detect_min[562][6] = (mid_1[4511:4504] < top_2[4503:4496]) ? 1 : 0;
assign detect_min[562][7] = (mid_1[4511:4504] < top_2[4511:4504]) ? 1 : 0;
assign detect_min[562][8] = (mid_1[4511:4504] < top_2[4519:4512]) ? 1 : 0;
assign detect_min[562][9] = (mid_1[4511:4504] < mid_0[4503:4496]) ? 1 : 0;
assign detect_min[562][10] = (mid_1[4511:4504] < mid_0[4511:4504]) ? 1 : 0;
assign detect_min[562][11] = (mid_1[4511:4504] < mid_0[4519:4512]) ? 1 : 0;
assign detect_min[562][12] = (mid_1[4511:4504] < mid_1[4503:4496]) ? 1 : 0;
assign detect_min[562][13] = (mid_1[4511:4504] < mid_1[4519:4512]) ? 1 : 0;
assign detect_min[562][14] = (mid_1[4511:4504] < mid_2[4503:4496]) ? 1 : 0;
assign detect_min[562][15] = (mid_1[4511:4504] < mid_2[4511:4504]) ? 1 : 0;
assign detect_min[562][16] = (mid_1[4511:4504] < mid_2[4519:4512]) ? 1 : 0;
assign detect_min[562][17] = (mid_1[4511:4504] < btm_0[4503:4496]) ? 1 : 0;
assign detect_min[562][18] = (mid_1[4511:4504] < btm_0[4511:4504]) ? 1 : 0;
assign detect_min[562][19] = (mid_1[4511:4504] < btm_0[4519:4512]) ? 1 : 0;
assign detect_min[562][20] = (mid_1[4511:4504] < btm_1[4503:4496]) ? 1 : 0;
assign detect_min[562][21] = (mid_1[4511:4504] < btm_1[4511:4504]) ? 1 : 0;
assign detect_min[562][22] = (mid_1[4511:4504] < btm_1[4519:4512]) ? 1 : 0;
assign detect_min[562][23] = (mid_1[4511:4504] < btm_2[4503:4496]) ? 1 : 0;
assign detect_min[562][24] = (mid_1[4511:4504] < btm_2[4511:4504]) ? 1 : 0;
assign detect_min[562][25] = (mid_1[4511:4504] < btm_2[4519:4512]) ? 1 : 0;

assign detect_min[563][0] = (mid_1[4519:4512] < top_0[4511:4504]) ? 1 : 0;
assign detect_min[563][1] = (mid_1[4519:4512] < top_0[4519:4512]) ? 1 : 0;
assign detect_min[563][2] = (mid_1[4519:4512] < top_0[4527:4520]) ? 1 : 0;
assign detect_min[563][3] = (mid_1[4519:4512] < top_1[4511:4504]) ? 1 : 0;
assign detect_min[563][4] = (mid_1[4519:4512] < top_1[4519:4512]) ? 1 : 0;
assign detect_min[563][5] = (mid_1[4519:4512] < top_1[4527:4520]) ? 1 : 0;
assign detect_min[563][6] = (mid_1[4519:4512] < top_2[4511:4504]) ? 1 : 0;
assign detect_min[563][7] = (mid_1[4519:4512] < top_2[4519:4512]) ? 1 : 0;
assign detect_min[563][8] = (mid_1[4519:4512] < top_2[4527:4520]) ? 1 : 0;
assign detect_min[563][9] = (mid_1[4519:4512] < mid_0[4511:4504]) ? 1 : 0;
assign detect_min[563][10] = (mid_1[4519:4512] < mid_0[4519:4512]) ? 1 : 0;
assign detect_min[563][11] = (mid_1[4519:4512] < mid_0[4527:4520]) ? 1 : 0;
assign detect_min[563][12] = (mid_1[4519:4512] < mid_1[4511:4504]) ? 1 : 0;
assign detect_min[563][13] = (mid_1[4519:4512] < mid_1[4527:4520]) ? 1 : 0;
assign detect_min[563][14] = (mid_1[4519:4512] < mid_2[4511:4504]) ? 1 : 0;
assign detect_min[563][15] = (mid_1[4519:4512] < mid_2[4519:4512]) ? 1 : 0;
assign detect_min[563][16] = (mid_1[4519:4512] < mid_2[4527:4520]) ? 1 : 0;
assign detect_min[563][17] = (mid_1[4519:4512] < btm_0[4511:4504]) ? 1 : 0;
assign detect_min[563][18] = (mid_1[4519:4512] < btm_0[4519:4512]) ? 1 : 0;
assign detect_min[563][19] = (mid_1[4519:4512] < btm_0[4527:4520]) ? 1 : 0;
assign detect_min[563][20] = (mid_1[4519:4512] < btm_1[4511:4504]) ? 1 : 0;
assign detect_min[563][21] = (mid_1[4519:4512] < btm_1[4519:4512]) ? 1 : 0;
assign detect_min[563][22] = (mid_1[4519:4512] < btm_1[4527:4520]) ? 1 : 0;
assign detect_min[563][23] = (mid_1[4519:4512] < btm_2[4511:4504]) ? 1 : 0;
assign detect_min[563][24] = (mid_1[4519:4512] < btm_2[4519:4512]) ? 1 : 0;
assign detect_min[563][25] = (mid_1[4519:4512] < btm_2[4527:4520]) ? 1 : 0;

assign detect_min[564][0] = (mid_1[4527:4520] < top_0[4519:4512]) ? 1 : 0;
assign detect_min[564][1] = (mid_1[4527:4520] < top_0[4527:4520]) ? 1 : 0;
assign detect_min[564][2] = (mid_1[4527:4520] < top_0[4535:4528]) ? 1 : 0;
assign detect_min[564][3] = (mid_1[4527:4520] < top_1[4519:4512]) ? 1 : 0;
assign detect_min[564][4] = (mid_1[4527:4520] < top_1[4527:4520]) ? 1 : 0;
assign detect_min[564][5] = (mid_1[4527:4520] < top_1[4535:4528]) ? 1 : 0;
assign detect_min[564][6] = (mid_1[4527:4520] < top_2[4519:4512]) ? 1 : 0;
assign detect_min[564][7] = (mid_1[4527:4520] < top_2[4527:4520]) ? 1 : 0;
assign detect_min[564][8] = (mid_1[4527:4520] < top_2[4535:4528]) ? 1 : 0;
assign detect_min[564][9] = (mid_1[4527:4520] < mid_0[4519:4512]) ? 1 : 0;
assign detect_min[564][10] = (mid_1[4527:4520] < mid_0[4527:4520]) ? 1 : 0;
assign detect_min[564][11] = (mid_1[4527:4520] < mid_0[4535:4528]) ? 1 : 0;
assign detect_min[564][12] = (mid_1[4527:4520] < mid_1[4519:4512]) ? 1 : 0;
assign detect_min[564][13] = (mid_1[4527:4520] < mid_1[4535:4528]) ? 1 : 0;
assign detect_min[564][14] = (mid_1[4527:4520] < mid_2[4519:4512]) ? 1 : 0;
assign detect_min[564][15] = (mid_1[4527:4520] < mid_2[4527:4520]) ? 1 : 0;
assign detect_min[564][16] = (mid_1[4527:4520] < mid_2[4535:4528]) ? 1 : 0;
assign detect_min[564][17] = (mid_1[4527:4520] < btm_0[4519:4512]) ? 1 : 0;
assign detect_min[564][18] = (mid_1[4527:4520] < btm_0[4527:4520]) ? 1 : 0;
assign detect_min[564][19] = (mid_1[4527:4520] < btm_0[4535:4528]) ? 1 : 0;
assign detect_min[564][20] = (mid_1[4527:4520] < btm_1[4519:4512]) ? 1 : 0;
assign detect_min[564][21] = (mid_1[4527:4520] < btm_1[4527:4520]) ? 1 : 0;
assign detect_min[564][22] = (mid_1[4527:4520] < btm_1[4535:4528]) ? 1 : 0;
assign detect_min[564][23] = (mid_1[4527:4520] < btm_2[4519:4512]) ? 1 : 0;
assign detect_min[564][24] = (mid_1[4527:4520] < btm_2[4527:4520]) ? 1 : 0;
assign detect_min[564][25] = (mid_1[4527:4520] < btm_2[4535:4528]) ? 1 : 0;

assign detect_min[565][0] = (mid_1[4535:4528] < top_0[4527:4520]) ? 1 : 0;
assign detect_min[565][1] = (mid_1[4535:4528] < top_0[4535:4528]) ? 1 : 0;
assign detect_min[565][2] = (mid_1[4535:4528] < top_0[4543:4536]) ? 1 : 0;
assign detect_min[565][3] = (mid_1[4535:4528] < top_1[4527:4520]) ? 1 : 0;
assign detect_min[565][4] = (mid_1[4535:4528] < top_1[4535:4528]) ? 1 : 0;
assign detect_min[565][5] = (mid_1[4535:4528] < top_1[4543:4536]) ? 1 : 0;
assign detect_min[565][6] = (mid_1[4535:4528] < top_2[4527:4520]) ? 1 : 0;
assign detect_min[565][7] = (mid_1[4535:4528] < top_2[4535:4528]) ? 1 : 0;
assign detect_min[565][8] = (mid_1[4535:4528] < top_2[4543:4536]) ? 1 : 0;
assign detect_min[565][9] = (mid_1[4535:4528] < mid_0[4527:4520]) ? 1 : 0;
assign detect_min[565][10] = (mid_1[4535:4528] < mid_0[4535:4528]) ? 1 : 0;
assign detect_min[565][11] = (mid_1[4535:4528] < mid_0[4543:4536]) ? 1 : 0;
assign detect_min[565][12] = (mid_1[4535:4528] < mid_1[4527:4520]) ? 1 : 0;
assign detect_min[565][13] = (mid_1[4535:4528] < mid_1[4543:4536]) ? 1 : 0;
assign detect_min[565][14] = (mid_1[4535:4528] < mid_2[4527:4520]) ? 1 : 0;
assign detect_min[565][15] = (mid_1[4535:4528] < mid_2[4535:4528]) ? 1 : 0;
assign detect_min[565][16] = (mid_1[4535:4528] < mid_2[4543:4536]) ? 1 : 0;
assign detect_min[565][17] = (mid_1[4535:4528] < btm_0[4527:4520]) ? 1 : 0;
assign detect_min[565][18] = (mid_1[4535:4528] < btm_0[4535:4528]) ? 1 : 0;
assign detect_min[565][19] = (mid_1[4535:4528] < btm_0[4543:4536]) ? 1 : 0;
assign detect_min[565][20] = (mid_1[4535:4528] < btm_1[4527:4520]) ? 1 : 0;
assign detect_min[565][21] = (mid_1[4535:4528] < btm_1[4535:4528]) ? 1 : 0;
assign detect_min[565][22] = (mid_1[4535:4528] < btm_1[4543:4536]) ? 1 : 0;
assign detect_min[565][23] = (mid_1[4535:4528] < btm_2[4527:4520]) ? 1 : 0;
assign detect_min[565][24] = (mid_1[4535:4528] < btm_2[4535:4528]) ? 1 : 0;
assign detect_min[565][25] = (mid_1[4535:4528] < btm_2[4543:4536]) ? 1 : 0;

assign detect_min[566][0] = (mid_1[4543:4536] < top_0[4535:4528]) ? 1 : 0;
assign detect_min[566][1] = (mid_1[4543:4536] < top_0[4543:4536]) ? 1 : 0;
assign detect_min[566][2] = (mid_1[4543:4536] < top_0[4551:4544]) ? 1 : 0;
assign detect_min[566][3] = (mid_1[4543:4536] < top_1[4535:4528]) ? 1 : 0;
assign detect_min[566][4] = (mid_1[4543:4536] < top_1[4543:4536]) ? 1 : 0;
assign detect_min[566][5] = (mid_1[4543:4536] < top_1[4551:4544]) ? 1 : 0;
assign detect_min[566][6] = (mid_1[4543:4536] < top_2[4535:4528]) ? 1 : 0;
assign detect_min[566][7] = (mid_1[4543:4536] < top_2[4543:4536]) ? 1 : 0;
assign detect_min[566][8] = (mid_1[4543:4536] < top_2[4551:4544]) ? 1 : 0;
assign detect_min[566][9] = (mid_1[4543:4536] < mid_0[4535:4528]) ? 1 : 0;
assign detect_min[566][10] = (mid_1[4543:4536] < mid_0[4543:4536]) ? 1 : 0;
assign detect_min[566][11] = (mid_1[4543:4536] < mid_0[4551:4544]) ? 1 : 0;
assign detect_min[566][12] = (mid_1[4543:4536] < mid_1[4535:4528]) ? 1 : 0;
assign detect_min[566][13] = (mid_1[4543:4536] < mid_1[4551:4544]) ? 1 : 0;
assign detect_min[566][14] = (mid_1[4543:4536] < mid_2[4535:4528]) ? 1 : 0;
assign detect_min[566][15] = (mid_1[4543:4536] < mid_2[4543:4536]) ? 1 : 0;
assign detect_min[566][16] = (mid_1[4543:4536] < mid_2[4551:4544]) ? 1 : 0;
assign detect_min[566][17] = (mid_1[4543:4536] < btm_0[4535:4528]) ? 1 : 0;
assign detect_min[566][18] = (mid_1[4543:4536] < btm_0[4543:4536]) ? 1 : 0;
assign detect_min[566][19] = (mid_1[4543:4536] < btm_0[4551:4544]) ? 1 : 0;
assign detect_min[566][20] = (mid_1[4543:4536] < btm_1[4535:4528]) ? 1 : 0;
assign detect_min[566][21] = (mid_1[4543:4536] < btm_1[4543:4536]) ? 1 : 0;
assign detect_min[566][22] = (mid_1[4543:4536] < btm_1[4551:4544]) ? 1 : 0;
assign detect_min[566][23] = (mid_1[4543:4536] < btm_2[4535:4528]) ? 1 : 0;
assign detect_min[566][24] = (mid_1[4543:4536] < btm_2[4543:4536]) ? 1 : 0;
assign detect_min[566][25] = (mid_1[4543:4536] < btm_2[4551:4544]) ? 1 : 0;

assign detect_min[567][0] = (mid_1[4551:4544] < top_0[4543:4536]) ? 1 : 0;
assign detect_min[567][1] = (mid_1[4551:4544] < top_0[4551:4544]) ? 1 : 0;
assign detect_min[567][2] = (mid_1[4551:4544] < top_0[4559:4552]) ? 1 : 0;
assign detect_min[567][3] = (mid_1[4551:4544] < top_1[4543:4536]) ? 1 : 0;
assign detect_min[567][4] = (mid_1[4551:4544] < top_1[4551:4544]) ? 1 : 0;
assign detect_min[567][5] = (mid_1[4551:4544] < top_1[4559:4552]) ? 1 : 0;
assign detect_min[567][6] = (mid_1[4551:4544] < top_2[4543:4536]) ? 1 : 0;
assign detect_min[567][7] = (mid_1[4551:4544] < top_2[4551:4544]) ? 1 : 0;
assign detect_min[567][8] = (mid_1[4551:4544] < top_2[4559:4552]) ? 1 : 0;
assign detect_min[567][9] = (mid_1[4551:4544] < mid_0[4543:4536]) ? 1 : 0;
assign detect_min[567][10] = (mid_1[4551:4544] < mid_0[4551:4544]) ? 1 : 0;
assign detect_min[567][11] = (mid_1[4551:4544] < mid_0[4559:4552]) ? 1 : 0;
assign detect_min[567][12] = (mid_1[4551:4544] < mid_1[4543:4536]) ? 1 : 0;
assign detect_min[567][13] = (mid_1[4551:4544] < mid_1[4559:4552]) ? 1 : 0;
assign detect_min[567][14] = (mid_1[4551:4544] < mid_2[4543:4536]) ? 1 : 0;
assign detect_min[567][15] = (mid_1[4551:4544] < mid_2[4551:4544]) ? 1 : 0;
assign detect_min[567][16] = (mid_1[4551:4544] < mid_2[4559:4552]) ? 1 : 0;
assign detect_min[567][17] = (mid_1[4551:4544] < btm_0[4543:4536]) ? 1 : 0;
assign detect_min[567][18] = (mid_1[4551:4544] < btm_0[4551:4544]) ? 1 : 0;
assign detect_min[567][19] = (mid_1[4551:4544] < btm_0[4559:4552]) ? 1 : 0;
assign detect_min[567][20] = (mid_1[4551:4544] < btm_1[4543:4536]) ? 1 : 0;
assign detect_min[567][21] = (mid_1[4551:4544] < btm_1[4551:4544]) ? 1 : 0;
assign detect_min[567][22] = (mid_1[4551:4544] < btm_1[4559:4552]) ? 1 : 0;
assign detect_min[567][23] = (mid_1[4551:4544] < btm_2[4543:4536]) ? 1 : 0;
assign detect_min[567][24] = (mid_1[4551:4544] < btm_2[4551:4544]) ? 1 : 0;
assign detect_min[567][25] = (mid_1[4551:4544] < btm_2[4559:4552]) ? 1 : 0;

assign detect_min[568][0] = (mid_1[4559:4552] < top_0[4551:4544]) ? 1 : 0;
assign detect_min[568][1] = (mid_1[4559:4552] < top_0[4559:4552]) ? 1 : 0;
assign detect_min[568][2] = (mid_1[4559:4552] < top_0[4567:4560]) ? 1 : 0;
assign detect_min[568][3] = (mid_1[4559:4552] < top_1[4551:4544]) ? 1 : 0;
assign detect_min[568][4] = (mid_1[4559:4552] < top_1[4559:4552]) ? 1 : 0;
assign detect_min[568][5] = (mid_1[4559:4552] < top_1[4567:4560]) ? 1 : 0;
assign detect_min[568][6] = (mid_1[4559:4552] < top_2[4551:4544]) ? 1 : 0;
assign detect_min[568][7] = (mid_1[4559:4552] < top_2[4559:4552]) ? 1 : 0;
assign detect_min[568][8] = (mid_1[4559:4552] < top_2[4567:4560]) ? 1 : 0;
assign detect_min[568][9] = (mid_1[4559:4552] < mid_0[4551:4544]) ? 1 : 0;
assign detect_min[568][10] = (mid_1[4559:4552] < mid_0[4559:4552]) ? 1 : 0;
assign detect_min[568][11] = (mid_1[4559:4552] < mid_0[4567:4560]) ? 1 : 0;
assign detect_min[568][12] = (mid_1[4559:4552] < mid_1[4551:4544]) ? 1 : 0;
assign detect_min[568][13] = (mid_1[4559:4552] < mid_1[4567:4560]) ? 1 : 0;
assign detect_min[568][14] = (mid_1[4559:4552] < mid_2[4551:4544]) ? 1 : 0;
assign detect_min[568][15] = (mid_1[4559:4552] < mid_2[4559:4552]) ? 1 : 0;
assign detect_min[568][16] = (mid_1[4559:4552] < mid_2[4567:4560]) ? 1 : 0;
assign detect_min[568][17] = (mid_1[4559:4552] < btm_0[4551:4544]) ? 1 : 0;
assign detect_min[568][18] = (mid_1[4559:4552] < btm_0[4559:4552]) ? 1 : 0;
assign detect_min[568][19] = (mid_1[4559:4552] < btm_0[4567:4560]) ? 1 : 0;
assign detect_min[568][20] = (mid_1[4559:4552] < btm_1[4551:4544]) ? 1 : 0;
assign detect_min[568][21] = (mid_1[4559:4552] < btm_1[4559:4552]) ? 1 : 0;
assign detect_min[568][22] = (mid_1[4559:4552] < btm_1[4567:4560]) ? 1 : 0;
assign detect_min[568][23] = (mid_1[4559:4552] < btm_2[4551:4544]) ? 1 : 0;
assign detect_min[568][24] = (mid_1[4559:4552] < btm_2[4559:4552]) ? 1 : 0;
assign detect_min[568][25] = (mid_1[4559:4552] < btm_2[4567:4560]) ? 1 : 0;

assign detect_min[569][0] = (mid_1[4567:4560] < top_0[4559:4552]) ? 1 : 0;
assign detect_min[569][1] = (mid_1[4567:4560] < top_0[4567:4560]) ? 1 : 0;
assign detect_min[569][2] = (mid_1[4567:4560] < top_0[4575:4568]) ? 1 : 0;
assign detect_min[569][3] = (mid_1[4567:4560] < top_1[4559:4552]) ? 1 : 0;
assign detect_min[569][4] = (mid_1[4567:4560] < top_1[4567:4560]) ? 1 : 0;
assign detect_min[569][5] = (mid_1[4567:4560] < top_1[4575:4568]) ? 1 : 0;
assign detect_min[569][6] = (mid_1[4567:4560] < top_2[4559:4552]) ? 1 : 0;
assign detect_min[569][7] = (mid_1[4567:4560] < top_2[4567:4560]) ? 1 : 0;
assign detect_min[569][8] = (mid_1[4567:4560] < top_2[4575:4568]) ? 1 : 0;
assign detect_min[569][9] = (mid_1[4567:4560] < mid_0[4559:4552]) ? 1 : 0;
assign detect_min[569][10] = (mid_1[4567:4560] < mid_0[4567:4560]) ? 1 : 0;
assign detect_min[569][11] = (mid_1[4567:4560] < mid_0[4575:4568]) ? 1 : 0;
assign detect_min[569][12] = (mid_1[4567:4560] < mid_1[4559:4552]) ? 1 : 0;
assign detect_min[569][13] = (mid_1[4567:4560] < mid_1[4575:4568]) ? 1 : 0;
assign detect_min[569][14] = (mid_1[4567:4560] < mid_2[4559:4552]) ? 1 : 0;
assign detect_min[569][15] = (mid_1[4567:4560] < mid_2[4567:4560]) ? 1 : 0;
assign detect_min[569][16] = (mid_1[4567:4560] < mid_2[4575:4568]) ? 1 : 0;
assign detect_min[569][17] = (mid_1[4567:4560] < btm_0[4559:4552]) ? 1 : 0;
assign detect_min[569][18] = (mid_1[4567:4560] < btm_0[4567:4560]) ? 1 : 0;
assign detect_min[569][19] = (mid_1[4567:4560] < btm_0[4575:4568]) ? 1 : 0;
assign detect_min[569][20] = (mid_1[4567:4560] < btm_1[4559:4552]) ? 1 : 0;
assign detect_min[569][21] = (mid_1[4567:4560] < btm_1[4567:4560]) ? 1 : 0;
assign detect_min[569][22] = (mid_1[4567:4560] < btm_1[4575:4568]) ? 1 : 0;
assign detect_min[569][23] = (mid_1[4567:4560] < btm_2[4559:4552]) ? 1 : 0;
assign detect_min[569][24] = (mid_1[4567:4560] < btm_2[4567:4560]) ? 1 : 0;
assign detect_min[569][25] = (mid_1[4567:4560] < btm_2[4575:4568]) ? 1 : 0;

assign detect_min[570][0] = (mid_1[4575:4568] < top_0[4567:4560]) ? 1 : 0;
assign detect_min[570][1] = (mid_1[4575:4568] < top_0[4575:4568]) ? 1 : 0;
assign detect_min[570][2] = (mid_1[4575:4568] < top_0[4583:4576]) ? 1 : 0;
assign detect_min[570][3] = (mid_1[4575:4568] < top_1[4567:4560]) ? 1 : 0;
assign detect_min[570][4] = (mid_1[4575:4568] < top_1[4575:4568]) ? 1 : 0;
assign detect_min[570][5] = (mid_1[4575:4568] < top_1[4583:4576]) ? 1 : 0;
assign detect_min[570][6] = (mid_1[4575:4568] < top_2[4567:4560]) ? 1 : 0;
assign detect_min[570][7] = (mid_1[4575:4568] < top_2[4575:4568]) ? 1 : 0;
assign detect_min[570][8] = (mid_1[4575:4568] < top_2[4583:4576]) ? 1 : 0;
assign detect_min[570][9] = (mid_1[4575:4568] < mid_0[4567:4560]) ? 1 : 0;
assign detect_min[570][10] = (mid_1[4575:4568] < mid_0[4575:4568]) ? 1 : 0;
assign detect_min[570][11] = (mid_1[4575:4568] < mid_0[4583:4576]) ? 1 : 0;
assign detect_min[570][12] = (mid_1[4575:4568] < mid_1[4567:4560]) ? 1 : 0;
assign detect_min[570][13] = (mid_1[4575:4568] < mid_1[4583:4576]) ? 1 : 0;
assign detect_min[570][14] = (mid_1[4575:4568] < mid_2[4567:4560]) ? 1 : 0;
assign detect_min[570][15] = (mid_1[4575:4568] < mid_2[4575:4568]) ? 1 : 0;
assign detect_min[570][16] = (mid_1[4575:4568] < mid_2[4583:4576]) ? 1 : 0;
assign detect_min[570][17] = (mid_1[4575:4568] < btm_0[4567:4560]) ? 1 : 0;
assign detect_min[570][18] = (mid_1[4575:4568] < btm_0[4575:4568]) ? 1 : 0;
assign detect_min[570][19] = (mid_1[4575:4568] < btm_0[4583:4576]) ? 1 : 0;
assign detect_min[570][20] = (mid_1[4575:4568] < btm_1[4567:4560]) ? 1 : 0;
assign detect_min[570][21] = (mid_1[4575:4568] < btm_1[4575:4568]) ? 1 : 0;
assign detect_min[570][22] = (mid_1[4575:4568] < btm_1[4583:4576]) ? 1 : 0;
assign detect_min[570][23] = (mid_1[4575:4568] < btm_2[4567:4560]) ? 1 : 0;
assign detect_min[570][24] = (mid_1[4575:4568] < btm_2[4575:4568]) ? 1 : 0;
assign detect_min[570][25] = (mid_1[4575:4568] < btm_2[4583:4576]) ? 1 : 0;

assign detect_min[571][0] = (mid_1[4583:4576] < top_0[4575:4568]) ? 1 : 0;
assign detect_min[571][1] = (mid_1[4583:4576] < top_0[4583:4576]) ? 1 : 0;
assign detect_min[571][2] = (mid_1[4583:4576] < top_0[4591:4584]) ? 1 : 0;
assign detect_min[571][3] = (mid_1[4583:4576] < top_1[4575:4568]) ? 1 : 0;
assign detect_min[571][4] = (mid_1[4583:4576] < top_1[4583:4576]) ? 1 : 0;
assign detect_min[571][5] = (mid_1[4583:4576] < top_1[4591:4584]) ? 1 : 0;
assign detect_min[571][6] = (mid_1[4583:4576] < top_2[4575:4568]) ? 1 : 0;
assign detect_min[571][7] = (mid_1[4583:4576] < top_2[4583:4576]) ? 1 : 0;
assign detect_min[571][8] = (mid_1[4583:4576] < top_2[4591:4584]) ? 1 : 0;
assign detect_min[571][9] = (mid_1[4583:4576] < mid_0[4575:4568]) ? 1 : 0;
assign detect_min[571][10] = (mid_1[4583:4576] < mid_0[4583:4576]) ? 1 : 0;
assign detect_min[571][11] = (mid_1[4583:4576] < mid_0[4591:4584]) ? 1 : 0;
assign detect_min[571][12] = (mid_1[4583:4576] < mid_1[4575:4568]) ? 1 : 0;
assign detect_min[571][13] = (mid_1[4583:4576] < mid_1[4591:4584]) ? 1 : 0;
assign detect_min[571][14] = (mid_1[4583:4576] < mid_2[4575:4568]) ? 1 : 0;
assign detect_min[571][15] = (mid_1[4583:4576] < mid_2[4583:4576]) ? 1 : 0;
assign detect_min[571][16] = (mid_1[4583:4576] < mid_2[4591:4584]) ? 1 : 0;
assign detect_min[571][17] = (mid_1[4583:4576] < btm_0[4575:4568]) ? 1 : 0;
assign detect_min[571][18] = (mid_1[4583:4576] < btm_0[4583:4576]) ? 1 : 0;
assign detect_min[571][19] = (mid_1[4583:4576] < btm_0[4591:4584]) ? 1 : 0;
assign detect_min[571][20] = (mid_1[4583:4576] < btm_1[4575:4568]) ? 1 : 0;
assign detect_min[571][21] = (mid_1[4583:4576] < btm_1[4583:4576]) ? 1 : 0;
assign detect_min[571][22] = (mid_1[4583:4576] < btm_1[4591:4584]) ? 1 : 0;
assign detect_min[571][23] = (mid_1[4583:4576] < btm_2[4575:4568]) ? 1 : 0;
assign detect_min[571][24] = (mid_1[4583:4576] < btm_2[4583:4576]) ? 1 : 0;
assign detect_min[571][25] = (mid_1[4583:4576] < btm_2[4591:4584]) ? 1 : 0;

assign detect_min[572][0] = (mid_1[4591:4584] < top_0[4583:4576]) ? 1 : 0;
assign detect_min[572][1] = (mid_1[4591:4584] < top_0[4591:4584]) ? 1 : 0;
assign detect_min[572][2] = (mid_1[4591:4584] < top_0[4599:4592]) ? 1 : 0;
assign detect_min[572][3] = (mid_1[4591:4584] < top_1[4583:4576]) ? 1 : 0;
assign detect_min[572][4] = (mid_1[4591:4584] < top_1[4591:4584]) ? 1 : 0;
assign detect_min[572][5] = (mid_1[4591:4584] < top_1[4599:4592]) ? 1 : 0;
assign detect_min[572][6] = (mid_1[4591:4584] < top_2[4583:4576]) ? 1 : 0;
assign detect_min[572][7] = (mid_1[4591:4584] < top_2[4591:4584]) ? 1 : 0;
assign detect_min[572][8] = (mid_1[4591:4584] < top_2[4599:4592]) ? 1 : 0;
assign detect_min[572][9] = (mid_1[4591:4584] < mid_0[4583:4576]) ? 1 : 0;
assign detect_min[572][10] = (mid_1[4591:4584] < mid_0[4591:4584]) ? 1 : 0;
assign detect_min[572][11] = (mid_1[4591:4584] < mid_0[4599:4592]) ? 1 : 0;
assign detect_min[572][12] = (mid_1[4591:4584] < mid_1[4583:4576]) ? 1 : 0;
assign detect_min[572][13] = (mid_1[4591:4584] < mid_1[4599:4592]) ? 1 : 0;
assign detect_min[572][14] = (mid_1[4591:4584] < mid_2[4583:4576]) ? 1 : 0;
assign detect_min[572][15] = (mid_1[4591:4584] < mid_2[4591:4584]) ? 1 : 0;
assign detect_min[572][16] = (mid_1[4591:4584] < mid_2[4599:4592]) ? 1 : 0;
assign detect_min[572][17] = (mid_1[4591:4584] < btm_0[4583:4576]) ? 1 : 0;
assign detect_min[572][18] = (mid_1[4591:4584] < btm_0[4591:4584]) ? 1 : 0;
assign detect_min[572][19] = (mid_1[4591:4584] < btm_0[4599:4592]) ? 1 : 0;
assign detect_min[572][20] = (mid_1[4591:4584] < btm_1[4583:4576]) ? 1 : 0;
assign detect_min[572][21] = (mid_1[4591:4584] < btm_1[4591:4584]) ? 1 : 0;
assign detect_min[572][22] = (mid_1[4591:4584] < btm_1[4599:4592]) ? 1 : 0;
assign detect_min[572][23] = (mid_1[4591:4584] < btm_2[4583:4576]) ? 1 : 0;
assign detect_min[572][24] = (mid_1[4591:4584] < btm_2[4591:4584]) ? 1 : 0;
assign detect_min[572][25] = (mid_1[4591:4584] < btm_2[4599:4592]) ? 1 : 0;

assign detect_min[573][0] = (mid_1[4599:4592] < top_0[4591:4584]) ? 1 : 0;
assign detect_min[573][1] = (mid_1[4599:4592] < top_0[4599:4592]) ? 1 : 0;
assign detect_min[573][2] = (mid_1[4599:4592] < top_0[4607:4600]) ? 1 : 0;
assign detect_min[573][3] = (mid_1[4599:4592] < top_1[4591:4584]) ? 1 : 0;
assign detect_min[573][4] = (mid_1[4599:4592] < top_1[4599:4592]) ? 1 : 0;
assign detect_min[573][5] = (mid_1[4599:4592] < top_1[4607:4600]) ? 1 : 0;
assign detect_min[573][6] = (mid_1[4599:4592] < top_2[4591:4584]) ? 1 : 0;
assign detect_min[573][7] = (mid_1[4599:4592] < top_2[4599:4592]) ? 1 : 0;
assign detect_min[573][8] = (mid_1[4599:4592] < top_2[4607:4600]) ? 1 : 0;
assign detect_min[573][9] = (mid_1[4599:4592] < mid_0[4591:4584]) ? 1 : 0;
assign detect_min[573][10] = (mid_1[4599:4592] < mid_0[4599:4592]) ? 1 : 0;
assign detect_min[573][11] = (mid_1[4599:4592] < mid_0[4607:4600]) ? 1 : 0;
assign detect_min[573][12] = (mid_1[4599:4592] < mid_1[4591:4584]) ? 1 : 0;
assign detect_min[573][13] = (mid_1[4599:4592] < mid_1[4607:4600]) ? 1 : 0;
assign detect_min[573][14] = (mid_1[4599:4592] < mid_2[4591:4584]) ? 1 : 0;
assign detect_min[573][15] = (mid_1[4599:4592] < mid_2[4599:4592]) ? 1 : 0;
assign detect_min[573][16] = (mid_1[4599:4592] < mid_2[4607:4600]) ? 1 : 0;
assign detect_min[573][17] = (mid_1[4599:4592] < btm_0[4591:4584]) ? 1 : 0;
assign detect_min[573][18] = (mid_1[4599:4592] < btm_0[4599:4592]) ? 1 : 0;
assign detect_min[573][19] = (mid_1[4599:4592] < btm_0[4607:4600]) ? 1 : 0;
assign detect_min[573][20] = (mid_1[4599:4592] < btm_1[4591:4584]) ? 1 : 0;
assign detect_min[573][21] = (mid_1[4599:4592] < btm_1[4599:4592]) ? 1 : 0;
assign detect_min[573][22] = (mid_1[4599:4592] < btm_1[4607:4600]) ? 1 : 0;
assign detect_min[573][23] = (mid_1[4599:4592] < btm_2[4591:4584]) ? 1 : 0;
assign detect_min[573][24] = (mid_1[4599:4592] < btm_2[4599:4592]) ? 1 : 0;
assign detect_min[573][25] = (mid_1[4599:4592] < btm_2[4607:4600]) ? 1 : 0;

assign detect_min[574][0] = (mid_1[4607:4600] < top_0[4599:4592]) ? 1 : 0;
assign detect_min[574][1] = (mid_1[4607:4600] < top_0[4607:4600]) ? 1 : 0;
assign detect_min[574][2] = (mid_1[4607:4600] < top_0[4615:4608]) ? 1 : 0;
assign detect_min[574][3] = (mid_1[4607:4600] < top_1[4599:4592]) ? 1 : 0;
assign detect_min[574][4] = (mid_1[4607:4600] < top_1[4607:4600]) ? 1 : 0;
assign detect_min[574][5] = (mid_1[4607:4600] < top_1[4615:4608]) ? 1 : 0;
assign detect_min[574][6] = (mid_1[4607:4600] < top_2[4599:4592]) ? 1 : 0;
assign detect_min[574][7] = (mid_1[4607:4600] < top_2[4607:4600]) ? 1 : 0;
assign detect_min[574][8] = (mid_1[4607:4600] < top_2[4615:4608]) ? 1 : 0;
assign detect_min[574][9] = (mid_1[4607:4600] < mid_0[4599:4592]) ? 1 : 0;
assign detect_min[574][10] = (mid_1[4607:4600] < mid_0[4607:4600]) ? 1 : 0;
assign detect_min[574][11] = (mid_1[4607:4600] < mid_0[4615:4608]) ? 1 : 0;
assign detect_min[574][12] = (mid_1[4607:4600] < mid_1[4599:4592]) ? 1 : 0;
assign detect_min[574][13] = (mid_1[4607:4600] < mid_1[4615:4608]) ? 1 : 0;
assign detect_min[574][14] = (mid_1[4607:4600] < mid_2[4599:4592]) ? 1 : 0;
assign detect_min[574][15] = (mid_1[4607:4600] < mid_2[4607:4600]) ? 1 : 0;
assign detect_min[574][16] = (mid_1[4607:4600] < mid_2[4615:4608]) ? 1 : 0;
assign detect_min[574][17] = (mid_1[4607:4600] < btm_0[4599:4592]) ? 1 : 0;
assign detect_min[574][18] = (mid_1[4607:4600] < btm_0[4607:4600]) ? 1 : 0;
assign detect_min[574][19] = (mid_1[4607:4600] < btm_0[4615:4608]) ? 1 : 0;
assign detect_min[574][20] = (mid_1[4607:4600] < btm_1[4599:4592]) ? 1 : 0;
assign detect_min[574][21] = (mid_1[4607:4600] < btm_1[4607:4600]) ? 1 : 0;
assign detect_min[574][22] = (mid_1[4607:4600] < btm_1[4615:4608]) ? 1 : 0;
assign detect_min[574][23] = (mid_1[4607:4600] < btm_2[4599:4592]) ? 1 : 0;
assign detect_min[574][24] = (mid_1[4607:4600] < btm_2[4607:4600]) ? 1 : 0;
assign detect_min[574][25] = (mid_1[4607:4600] < btm_2[4615:4608]) ? 1 : 0;

assign detect_min[575][0] = (mid_1[4615:4608] < top_0[4607:4600]) ? 1 : 0;
assign detect_min[575][1] = (mid_1[4615:4608] < top_0[4615:4608]) ? 1 : 0;
assign detect_min[575][2] = (mid_1[4615:4608] < top_0[4623:4616]) ? 1 : 0;
assign detect_min[575][3] = (mid_1[4615:4608] < top_1[4607:4600]) ? 1 : 0;
assign detect_min[575][4] = (mid_1[4615:4608] < top_1[4615:4608]) ? 1 : 0;
assign detect_min[575][5] = (mid_1[4615:4608] < top_1[4623:4616]) ? 1 : 0;
assign detect_min[575][6] = (mid_1[4615:4608] < top_2[4607:4600]) ? 1 : 0;
assign detect_min[575][7] = (mid_1[4615:4608] < top_2[4615:4608]) ? 1 : 0;
assign detect_min[575][8] = (mid_1[4615:4608] < top_2[4623:4616]) ? 1 : 0;
assign detect_min[575][9] = (mid_1[4615:4608] < mid_0[4607:4600]) ? 1 : 0;
assign detect_min[575][10] = (mid_1[4615:4608] < mid_0[4615:4608]) ? 1 : 0;
assign detect_min[575][11] = (mid_1[4615:4608] < mid_0[4623:4616]) ? 1 : 0;
assign detect_min[575][12] = (mid_1[4615:4608] < mid_1[4607:4600]) ? 1 : 0;
assign detect_min[575][13] = (mid_1[4615:4608] < mid_1[4623:4616]) ? 1 : 0;
assign detect_min[575][14] = (mid_1[4615:4608] < mid_2[4607:4600]) ? 1 : 0;
assign detect_min[575][15] = (mid_1[4615:4608] < mid_2[4615:4608]) ? 1 : 0;
assign detect_min[575][16] = (mid_1[4615:4608] < mid_2[4623:4616]) ? 1 : 0;
assign detect_min[575][17] = (mid_1[4615:4608] < btm_0[4607:4600]) ? 1 : 0;
assign detect_min[575][18] = (mid_1[4615:4608] < btm_0[4615:4608]) ? 1 : 0;
assign detect_min[575][19] = (mid_1[4615:4608] < btm_0[4623:4616]) ? 1 : 0;
assign detect_min[575][20] = (mid_1[4615:4608] < btm_1[4607:4600]) ? 1 : 0;
assign detect_min[575][21] = (mid_1[4615:4608] < btm_1[4615:4608]) ? 1 : 0;
assign detect_min[575][22] = (mid_1[4615:4608] < btm_1[4623:4616]) ? 1 : 0;
assign detect_min[575][23] = (mid_1[4615:4608] < btm_2[4607:4600]) ? 1 : 0;
assign detect_min[575][24] = (mid_1[4615:4608] < btm_2[4615:4608]) ? 1 : 0;
assign detect_min[575][25] = (mid_1[4615:4608] < btm_2[4623:4616]) ? 1 : 0;

assign detect_min[576][0] = (mid_1[4623:4616] < top_0[4615:4608]) ? 1 : 0;
assign detect_min[576][1] = (mid_1[4623:4616] < top_0[4623:4616]) ? 1 : 0;
assign detect_min[576][2] = (mid_1[4623:4616] < top_0[4631:4624]) ? 1 : 0;
assign detect_min[576][3] = (mid_1[4623:4616] < top_1[4615:4608]) ? 1 : 0;
assign detect_min[576][4] = (mid_1[4623:4616] < top_1[4623:4616]) ? 1 : 0;
assign detect_min[576][5] = (mid_1[4623:4616] < top_1[4631:4624]) ? 1 : 0;
assign detect_min[576][6] = (mid_1[4623:4616] < top_2[4615:4608]) ? 1 : 0;
assign detect_min[576][7] = (mid_1[4623:4616] < top_2[4623:4616]) ? 1 : 0;
assign detect_min[576][8] = (mid_1[4623:4616] < top_2[4631:4624]) ? 1 : 0;
assign detect_min[576][9] = (mid_1[4623:4616] < mid_0[4615:4608]) ? 1 : 0;
assign detect_min[576][10] = (mid_1[4623:4616] < mid_0[4623:4616]) ? 1 : 0;
assign detect_min[576][11] = (mid_1[4623:4616] < mid_0[4631:4624]) ? 1 : 0;
assign detect_min[576][12] = (mid_1[4623:4616] < mid_1[4615:4608]) ? 1 : 0;
assign detect_min[576][13] = (mid_1[4623:4616] < mid_1[4631:4624]) ? 1 : 0;
assign detect_min[576][14] = (mid_1[4623:4616] < mid_2[4615:4608]) ? 1 : 0;
assign detect_min[576][15] = (mid_1[4623:4616] < mid_2[4623:4616]) ? 1 : 0;
assign detect_min[576][16] = (mid_1[4623:4616] < mid_2[4631:4624]) ? 1 : 0;
assign detect_min[576][17] = (mid_1[4623:4616] < btm_0[4615:4608]) ? 1 : 0;
assign detect_min[576][18] = (mid_1[4623:4616] < btm_0[4623:4616]) ? 1 : 0;
assign detect_min[576][19] = (mid_1[4623:4616] < btm_0[4631:4624]) ? 1 : 0;
assign detect_min[576][20] = (mid_1[4623:4616] < btm_1[4615:4608]) ? 1 : 0;
assign detect_min[576][21] = (mid_1[4623:4616] < btm_1[4623:4616]) ? 1 : 0;
assign detect_min[576][22] = (mid_1[4623:4616] < btm_1[4631:4624]) ? 1 : 0;
assign detect_min[576][23] = (mid_1[4623:4616] < btm_2[4615:4608]) ? 1 : 0;
assign detect_min[576][24] = (mid_1[4623:4616] < btm_2[4623:4616]) ? 1 : 0;
assign detect_min[576][25] = (mid_1[4623:4616] < btm_2[4631:4624]) ? 1 : 0;

assign detect_min[577][0] = (mid_1[4631:4624] < top_0[4623:4616]) ? 1 : 0;
assign detect_min[577][1] = (mid_1[4631:4624] < top_0[4631:4624]) ? 1 : 0;
assign detect_min[577][2] = (mid_1[4631:4624] < top_0[4639:4632]) ? 1 : 0;
assign detect_min[577][3] = (mid_1[4631:4624] < top_1[4623:4616]) ? 1 : 0;
assign detect_min[577][4] = (mid_1[4631:4624] < top_1[4631:4624]) ? 1 : 0;
assign detect_min[577][5] = (mid_1[4631:4624] < top_1[4639:4632]) ? 1 : 0;
assign detect_min[577][6] = (mid_1[4631:4624] < top_2[4623:4616]) ? 1 : 0;
assign detect_min[577][7] = (mid_1[4631:4624] < top_2[4631:4624]) ? 1 : 0;
assign detect_min[577][8] = (mid_1[4631:4624] < top_2[4639:4632]) ? 1 : 0;
assign detect_min[577][9] = (mid_1[4631:4624] < mid_0[4623:4616]) ? 1 : 0;
assign detect_min[577][10] = (mid_1[4631:4624] < mid_0[4631:4624]) ? 1 : 0;
assign detect_min[577][11] = (mid_1[4631:4624] < mid_0[4639:4632]) ? 1 : 0;
assign detect_min[577][12] = (mid_1[4631:4624] < mid_1[4623:4616]) ? 1 : 0;
assign detect_min[577][13] = (mid_1[4631:4624] < mid_1[4639:4632]) ? 1 : 0;
assign detect_min[577][14] = (mid_1[4631:4624] < mid_2[4623:4616]) ? 1 : 0;
assign detect_min[577][15] = (mid_1[4631:4624] < mid_2[4631:4624]) ? 1 : 0;
assign detect_min[577][16] = (mid_1[4631:4624] < mid_2[4639:4632]) ? 1 : 0;
assign detect_min[577][17] = (mid_1[4631:4624] < btm_0[4623:4616]) ? 1 : 0;
assign detect_min[577][18] = (mid_1[4631:4624] < btm_0[4631:4624]) ? 1 : 0;
assign detect_min[577][19] = (mid_1[4631:4624] < btm_0[4639:4632]) ? 1 : 0;
assign detect_min[577][20] = (mid_1[4631:4624] < btm_1[4623:4616]) ? 1 : 0;
assign detect_min[577][21] = (mid_1[4631:4624] < btm_1[4631:4624]) ? 1 : 0;
assign detect_min[577][22] = (mid_1[4631:4624] < btm_1[4639:4632]) ? 1 : 0;
assign detect_min[577][23] = (mid_1[4631:4624] < btm_2[4623:4616]) ? 1 : 0;
assign detect_min[577][24] = (mid_1[4631:4624] < btm_2[4631:4624]) ? 1 : 0;
assign detect_min[577][25] = (mid_1[4631:4624] < btm_2[4639:4632]) ? 1 : 0;

assign detect_min[578][0] = (mid_1[4639:4632] < top_0[4631:4624]) ? 1 : 0;
assign detect_min[578][1] = (mid_1[4639:4632] < top_0[4639:4632]) ? 1 : 0;
assign detect_min[578][2] = (mid_1[4639:4632] < top_0[4647:4640]) ? 1 : 0;
assign detect_min[578][3] = (mid_1[4639:4632] < top_1[4631:4624]) ? 1 : 0;
assign detect_min[578][4] = (mid_1[4639:4632] < top_1[4639:4632]) ? 1 : 0;
assign detect_min[578][5] = (mid_1[4639:4632] < top_1[4647:4640]) ? 1 : 0;
assign detect_min[578][6] = (mid_1[4639:4632] < top_2[4631:4624]) ? 1 : 0;
assign detect_min[578][7] = (mid_1[4639:4632] < top_2[4639:4632]) ? 1 : 0;
assign detect_min[578][8] = (mid_1[4639:4632] < top_2[4647:4640]) ? 1 : 0;
assign detect_min[578][9] = (mid_1[4639:4632] < mid_0[4631:4624]) ? 1 : 0;
assign detect_min[578][10] = (mid_1[4639:4632] < mid_0[4639:4632]) ? 1 : 0;
assign detect_min[578][11] = (mid_1[4639:4632] < mid_0[4647:4640]) ? 1 : 0;
assign detect_min[578][12] = (mid_1[4639:4632] < mid_1[4631:4624]) ? 1 : 0;
assign detect_min[578][13] = (mid_1[4639:4632] < mid_1[4647:4640]) ? 1 : 0;
assign detect_min[578][14] = (mid_1[4639:4632] < mid_2[4631:4624]) ? 1 : 0;
assign detect_min[578][15] = (mid_1[4639:4632] < mid_2[4639:4632]) ? 1 : 0;
assign detect_min[578][16] = (mid_1[4639:4632] < mid_2[4647:4640]) ? 1 : 0;
assign detect_min[578][17] = (mid_1[4639:4632] < btm_0[4631:4624]) ? 1 : 0;
assign detect_min[578][18] = (mid_1[4639:4632] < btm_0[4639:4632]) ? 1 : 0;
assign detect_min[578][19] = (mid_1[4639:4632] < btm_0[4647:4640]) ? 1 : 0;
assign detect_min[578][20] = (mid_1[4639:4632] < btm_1[4631:4624]) ? 1 : 0;
assign detect_min[578][21] = (mid_1[4639:4632] < btm_1[4639:4632]) ? 1 : 0;
assign detect_min[578][22] = (mid_1[4639:4632] < btm_1[4647:4640]) ? 1 : 0;
assign detect_min[578][23] = (mid_1[4639:4632] < btm_2[4631:4624]) ? 1 : 0;
assign detect_min[578][24] = (mid_1[4639:4632] < btm_2[4639:4632]) ? 1 : 0;
assign detect_min[578][25] = (mid_1[4639:4632] < btm_2[4647:4640]) ? 1 : 0;

assign detect_min[579][0] = (mid_1[4647:4640] < top_0[4639:4632]) ? 1 : 0;
assign detect_min[579][1] = (mid_1[4647:4640] < top_0[4647:4640]) ? 1 : 0;
assign detect_min[579][2] = (mid_1[4647:4640] < top_0[4655:4648]) ? 1 : 0;
assign detect_min[579][3] = (mid_1[4647:4640] < top_1[4639:4632]) ? 1 : 0;
assign detect_min[579][4] = (mid_1[4647:4640] < top_1[4647:4640]) ? 1 : 0;
assign detect_min[579][5] = (mid_1[4647:4640] < top_1[4655:4648]) ? 1 : 0;
assign detect_min[579][6] = (mid_1[4647:4640] < top_2[4639:4632]) ? 1 : 0;
assign detect_min[579][7] = (mid_1[4647:4640] < top_2[4647:4640]) ? 1 : 0;
assign detect_min[579][8] = (mid_1[4647:4640] < top_2[4655:4648]) ? 1 : 0;
assign detect_min[579][9] = (mid_1[4647:4640] < mid_0[4639:4632]) ? 1 : 0;
assign detect_min[579][10] = (mid_1[4647:4640] < mid_0[4647:4640]) ? 1 : 0;
assign detect_min[579][11] = (mid_1[4647:4640] < mid_0[4655:4648]) ? 1 : 0;
assign detect_min[579][12] = (mid_1[4647:4640] < mid_1[4639:4632]) ? 1 : 0;
assign detect_min[579][13] = (mid_1[4647:4640] < mid_1[4655:4648]) ? 1 : 0;
assign detect_min[579][14] = (mid_1[4647:4640] < mid_2[4639:4632]) ? 1 : 0;
assign detect_min[579][15] = (mid_1[4647:4640] < mid_2[4647:4640]) ? 1 : 0;
assign detect_min[579][16] = (mid_1[4647:4640] < mid_2[4655:4648]) ? 1 : 0;
assign detect_min[579][17] = (mid_1[4647:4640] < btm_0[4639:4632]) ? 1 : 0;
assign detect_min[579][18] = (mid_1[4647:4640] < btm_0[4647:4640]) ? 1 : 0;
assign detect_min[579][19] = (mid_1[4647:4640] < btm_0[4655:4648]) ? 1 : 0;
assign detect_min[579][20] = (mid_1[4647:4640] < btm_1[4639:4632]) ? 1 : 0;
assign detect_min[579][21] = (mid_1[4647:4640] < btm_1[4647:4640]) ? 1 : 0;
assign detect_min[579][22] = (mid_1[4647:4640] < btm_1[4655:4648]) ? 1 : 0;
assign detect_min[579][23] = (mid_1[4647:4640] < btm_2[4639:4632]) ? 1 : 0;
assign detect_min[579][24] = (mid_1[4647:4640] < btm_2[4647:4640]) ? 1 : 0;
assign detect_min[579][25] = (mid_1[4647:4640] < btm_2[4655:4648]) ? 1 : 0;

assign detect_min[580][0] = (mid_1[4655:4648] < top_0[4647:4640]) ? 1 : 0;
assign detect_min[580][1] = (mid_1[4655:4648] < top_0[4655:4648]) ? 1 : 0;
assign detect_min[580][2] = (mid_1[4655:4648] < top_0[4663:4656]) ? 1 : 0;
assign detect_min[580][3] = (mid_1[4655:4648] < top_1[4647:4640]) ? 1 : 0;
assign detect_min[580][4] = (mid_1[4655:4648] < top_1[4655:4648]) ? 1 : 0;
assign detect_min[580][5] = (mid_1[4655:4648] < top_1[4663:4656]) ? 1 : 0;
assign detect_min[580][6] = (mid_1[4655:4648] < top_2[4647:4640]) ? 1 : 0;
assign detect_min[580][7] = (mid_1[4655:4648] < top_2[4655:4648]) ? 1 : 0;
assign detect_min[580][8] = (mid_1[4655:4648] < top_2[4663:4656]) ? 1 : 0;
assign detect_min[580][9] = (mid_1[4655:4648] < mid_0[4647:4640]) ? 1 : 0;
assign detect_min[580][10] = (mid_1[4655:4648] < mid_0[4655:4648]) ? 1 : 0;
assign detect_min[580][11] = (mid_1[4655:4648] < mid_0[4663:4656]) ? 1 : 0;
assign detect_min[580][12] = (mid_1[4655:4648] < mid_1[4647:4640]) ? 1 : 0;
assign detect_min[580][13] = (mid_1[4655:4648] < mid_1[4663:4656]) ? 1 : 0;
assign detect_min[580][14] = (mid_1[4655:4648] < mid_2[4647:4640]) ? 1 : 0;
assign detect_min[580][15] = (mid_1[4655:4648] < mid_2[4655:4648]) ? 1 : 0;
assign detect_min[580][16] = (mid_1[4655:4648] < mid_2[4663:4656]) ? 1 : 0;
assign detect_min[580][17] = (mid_1[4655:4648] < btm_0[4647:4640]) ? 1 : 0;
assign detect_min[580][18] = (mid_1[4655:4648] < btm_0[4655:4648]) ? 1 : 0;
assign detect_min[580][19] = (mid_1[4655:4648] < btm_0[4663:4656]) ? 1 : 0;
assign detect_min[580][20] = (mid_1[4655:4648] < btm_1[4647:4640]) ? 1 : 0;
assign detect_min[580][21] = (mid_1[4655:4648] < btm_1[4655:4648]) ? 1 : 0;
assign detect_min[580][22] = (mid_1[4655:4648] < btm_1[4663:4656]) ? 1 : 0;
assign detect_min[580][23] = (mid_1[4655:4648] < btm_2[4647:4640]) ? 1 : 0;
assign detect_min[580][24] = (mid_1[4655:4648] < btm_2[4655:4648]) ? 1 : 0;
assign detect_min[580][25] = (mid_1[4655:4648] < btm_2[4663:4656]) ? 1 : 0;

assign detect_min[581][0] = (mid_1[4663:4656] < top_0[4655:4648]) ? 1 : 0;
assign detect_min[581][1] = (mid_1[4663:4656] < top_0[4663:4656]) ? 1 : 0;
assign detect_min[581][2] = (mid_1[4663:4656] < top_0[4671:4664]) ? 1 : 0;
assign detect_min[581][3] = (mid_1[4663:4656] < top_1[4655:4648]) ? 1 : 0;
assign detect_min[581][4] = (mid_1[4663:4656] < top_1[4663:4656]) ? 1 : 0;
assign detect_min[581][5] = (mid_1[4663:4656] < top_1[4671:4664]) ? 1 : 0;
assign detect_min[581][6] = (mid_1[4663:4656] < top_2[4655:4648]) ? 1 : 0;
assign detect_min[581][7] = (mid_1[4663:4656] < top_2[4663:4656]) ? 1 : 0;
assign detect_min[581][8] = (mid_1[4663:4656] < top_2[4671:4664]) ? 1 : 0;
assign detect_min[581][9] = (mid_1[4663:4656] < mid_0[4655:4648]) ? 1 : 0;
assign detect_min[581][10] = (mid_1[4663:4656] < mid_0[4663:4656]) ? 1 : 0;
assign detect_min[581][11] = (mid_1[4663:4656] < mid_0[4671:4664]) ? 1 : 0;
assign detect_min[581][12] = (mid_1[4663:4656] < mid_1[4655:4648]) ? 1 : 0;
assign detect_min[581][13] = (mid_1[4663:4656] < mid_1[4671:4664]) ? 1 : 0;
assign detect_min[581][14] = (mid_1[4663:4656] < mid_2[4655:4648]) ? 1 : 0;
assign detect_min[581][15] = (mid_1[4663:4656] < mid_2[4663:4656]) ? 1 : 0;
assign detect_min[581][16] = (mid_1[4663:4656] < mid_2[4671:4664]) ? 1 : 0;
assign detect_min[581][17] = (mid_1[4663:4656] < btm_0[4655:4648]) ? 1 : 0;
assign detect_min[581][18] = (mid_1[4663:4656] < btm_0[4663:4656]) ? 1 : 0;
assign detect_min[581][19] = (mid_1[4663:4656] < btm_0[4671:4664]) ? 1 : 0;
assign detect_min[581][20] = (mid_1[4663:4656] < btm_1[4655:4648]) ? 1 : 0;
assign detect_min[581][21] = (mid_1[4663:4656] < btm_1[4663:4656]) ? 1 : 0;
assign detect_min[581][22] = (mid_1[4663:4656] < btm_1[4671:4664]) ? 1 : 0;
assign detect_min[581][23] = (mid_1[4663:4656] < btm_2[4655:4648]) ? 1 : 0;
assign detect_min[581][24] = (mid_1[4663:4656] < btm_2[4663:4656]) ? 1 : 0;
assign detect_min[581][25] = (mid_1[4663:4656] < btm_2[4671:4664]) ? 1 : 0;

assign detect_min[582][0] = (mid_1[4671:4664] < top_0[4663:4656]) ? 1 : 0;
assign detect_min[582][1] = (mid_1[4671:4664] < top_0[4671:4664]) ? 1 : 0;
assign detect_min[582][2] = (mid_1[4671:4664] < top_0[4679:4672]) ? 1 : 0;
assign detect_min[582][3] = (mid_1[4671:4664] < top_1[4663:4656]) ? 1 : 0;
assign detect_min[582][4] = (mid_1[4671:4664] < top_1[4671:4664]) ? 1 : 0;
assign detect_min[582][5] = (mid_1[4671:4664] < top_1[4679:4672]) ? 1 : 0;
assign detect_min[582][6] = (mid_1[4671:4664] < top_2[4663:4656]) ? 1 : 0;
assign detect_min[582][7] = (mid_1[4671:4664] < top_2[4671:4664]) ? 1 : 0;
assign detect_min[582][8] = (mid_1[4671:4664] < top_2[4679:4672]) ? 1 : 0;
assign detect_min[582][9] = (mid_1[4671:4664] < mid_0[4663:4656]) ? 1 : 0;
assign detect_min[582][10] = (mid_1[4671:4664] < mid_0[4671:4664]) ? 1 : 0;
assign detect_min[582][11] = (mid_1[4671:4664] < mid_0[4679:4672]) ? 1 : 0;
assign detect_min[582][12] = (mid_1[4671:4664] < mid_1[4663:4656]) ? 1 : 0;
assign detect_min[582][13] = (mid_1[4671:4664] < mid_1[4679:4672]) ? 1 : 0;
assign detect_min[582][14] = (mid_1[4671:4664] < mid_2[4663:4656]) ? 1 : 0;
assign detect_min[582][15] = (mid_1[4671:4664] < mid_2[4671:4664]) ? 1 : 0;
assign detect_min[582][16] = (mid_1[4671:4664] < mid_2[4679:4672]) ? 1 : 0;
assign detect_min[582][17] = (mid_1[4671:4664] < btm_0[4663:4656]) ? 1 : 0;
assign detect_min[582][18] = (mid_1[4671:4664] < btm_0[4671:4664]) ? 1 : 0;
assign detect_min[582][19] = (mid_1[4671:4664] < btm_0[4679:4672]) ? 1 : 0;
assign detect_min[582][20] = (mid_1[4671:4664] < btm_1[4663:4656]) ? 1 : 0;
assign detect_min[582][21] = (mid_1[4671:4664] < btm_1[4671:4664]) ? 1 : 0;
assign detect_min[582][22] = (mid_1[4671:4664] < btm_1[4679:4672]) ? 1 : 0;
assign detect_min[582][23] = (mid_1[4671:4664] < btm_2[4663:4656]) ? 1 : 0;
assign detect_min[582][24] = (mid_1[4671:4664] < btm_2[4671:4664]) ? 1 : 0;
assign detect_min[582][25] = (mid_1[4671:4664] < btm_2[4679:4672]) ? 1 : 0;

assign detect_min[583][0] = (mid_1[4679:4672] < top_0[4671:4664]) ? 1 : 0;
assign detect_min[583][1] = (mid_1[4679:4672] < top_0[4679:4672]) ? 1 : 0;
assign detect_min[583][2] = (mid_1[4679:4672] < top_0[4687:4680]) ? 1 : 0;
assign detect_min[583][3] = (mid_1[4679:4672] < top_1[4671:4664]) ? 1 : 0;
assign detect_min[583][4] = (mid_1[4679:4672] < top_1[4679:4672]) ? 1 : 0;
assign detect_min[583][5] = (mid_1[4679:4672] < top_1[4687:4680]) ? 1 : 0;
assign detect_min[583][6] = (mid_1[4679:4672] < top_2[4671:4664]) ? 1 : 0;
assign detect_min[583][7] = (mid_1[4679:4672] < top_2[4679:4672]) ? 1 : 0;
assign detect_min[583][8] = (mid_1[4679:4672] < top_2[4687:4680]) ? 1 : 0;
assign detect_min[583][9] = (mid_1[4679:4672] < mid_0[4671:4664]) ? 1 : 0;
assign detect_min[583][10] = (mid_1[4679:4672] < mid_0[4679:4672]) ? 1 : 0;
assign detect_min[583][11] = (mid_1[4679:4672] < mid_0[4687:4680]) ? 1 : 0;
assign detect_min[583][12] = (mid_1[4679:4672] < mid_1[4671:4664]) ? 1 : 0;
assign detect_min[583][13] = (mid_1[4679:4672] < mid_1[4687:4680]) ? 1 : 0;
assign detect_min[583][14] = (mid_1[4679:4672] < mid_2[4671:4664]) ? 1 : 0;
assign detect_min[583][15] = (mid_1[4679:4672] < mid_2[4679:4672]) ? 1 : 0;
assign detect_min[583][16] = (mid_1[4679:4672] < mid_2[4687:4680]) ? 1 : 0;
assign detect_min[583][17] = (mid_1[4679:4672] < btm_0[4671:4664]) ? 1 : 0;
assign detect_min[583][18] = (mid_1[4679:4672] < btm_0[4679:4672]) ? 1 : 0;
assign detect_min[583][19] = (mid_1[4679:4672] < btm_0[4687:4680]) ? 1 : 0;
assign detect_min[583][20] = (mid_1[4679:4672] < btm_1[4671:4664]) ? 1 : 0;
assign detect_min[583][21] = (mid_1[4679:4672] < btm_1[4679:4672]) ? 1 : 0;
assign detect_min[583][22] = (mid_1[4679:4672] < btm_1[4687:4680]) ? 1 : 0;
assign detect_min[583][23] = (mid_1[4679:4672] < btm_2[4671:4664]) ? 1 : 0;
assign detect_min[583][24] = (mid_1[4679:4672] < btm_2[4679:4672]) ? 1 : 0;
assign detect_min[583][25] = (mid_1[4679:4672] < btm_2[4687:4680]) ? 1 : 0;

assign detect_min[584][0] = (mid_1[4687:4680] < top_0[4679:4672]) ? 1 : 0;
assign detect_min[584][1] = (mid_1[4687:4680] < top_0[4687:4680]) ? 1 : 0;
assign detect_min[584][2] = (mid_1[4687:4680] < top_0[4695:4688]) ? 1 : 0;
assign detect_min[584][3] = (mid_1[4687:4680] < top_1[4679:4672]) ? 1 : 0;
assign detect_min[584][4] = (mid_1[4687:4680] < top_1[4687:4680]) ? 1 : 0;
assign detect_min[584][5] = (mid_1[4687:4680] < top_1[4695:4688]) ? 1 : 0;
assign detect_min[584][6] = (mid_1[4687:4680] < top_2[4679:4672]) ? 1 : 0;
assign detect_min[584][7] = (mid_1[4687:4680] < top_2[4687:4680]) ? 1 : 0;
assign detect_min[584][8] = (mid_1[4687:4680] < top_2[4695:4688]) ? 1 : 0;
assign detect_min[584][9] = (mid_1[4687:4680] < mid_0[4679:4672]) ? 1 : 0;
assign detect_min[584][10] = (mid_1[4687:4680] < mid_0[4687:4680]) ? 1 : 0;
assign detect_min[584][11] = (mid_1[4687:4680] < mid_0[4695:4688]) ? 1 : 0;
assign detect_min[584][12] = (mid_1[4687:4680] < mid_1[4679:4672]) ? 1 : 0;
assign detect_min[584][13] = (mid_1[4687:4680] < mid_1[4695:4688]) ? 1 : 0;
assign detect_min[584][14] = (mid_1[4687:4680] < mid_2[4679:4672]) ? 1 : 0;
assign detect_min[584][15] = (mid_1[4687:4680] < mid_2[4687:4680]) ? 1 : 0;
assign detect_min[584][16] = (mid_1[4687:4680] < mid_2[4695:4688]) ? 1 : 0;
assign detect_min[584][17] = (mid_1[4687:4680] < btm_0[4679:4672]) ? 1 : 0;
assign detect_min[584][18] = (mid_1[4687:4680] < btm_0[4687:4680]) ? 1 : 0;
assign detect_min[584][19] = (mid_1[4687:4680] < btm_0[4695:4688]) ? 1 : 0;
assign detect_min[584][20] = (mid_1[4687:4680] < btm_1[4679:4672]) ? 1 : 0;
assign detect_min[584][21] = (mid_1[4687:4680] < btm_1[4687:4680]) ? 1 : 0;
assign detect_min[584][22] = (mid_1[4687:4680] < btm_1[4695:4688]) ? 1 : 0;
assign detect_min[584][23] = (mid_1[4687:4680] < btm_2[4679:4672]) ? 1 : 0;
assign detect_min[584][24] = (mid_1[4687:4680] < btm_2[4687:4680]) ? 1 : 0;
assign detect_min[584][25] = (mid_1[4687:4680] < btm_2[4695:4688]) ? 1 : 0;

assign detect_min[585][0] = (mid_1[4695:4688] < top_0[4687:4680]) ? 1 : 0;
assign detect_min[585][1] = (mid_1[4695:4688] < top_0[4695:4688]) ? 1 : 0;
assign detect_min[585][2] = (mid_1[4695:4688] < top_0[4703:4696]) ? 1 : 0;
assign detect_min[585][3] = (mid_1[4695:4688] < top_1[4687:4680]) ? 1 : 0;
assign detect_min[585][4] = (mid_1[4695:4688] < top_1[4695:4688]) ? 1 : 0;
assign detect_min[585][5] = (mid_1[4695:4688] < top_1[4703:4696]) ? 1 : 0;
assign detect_min[585][6] = (mid_1[4695:4688] < top_2[4687:4680]) ? 1 : 0;
assign detect_min[585][7] = (mid_1[4695:4688] < top_2[4695:4688]) ? 1 : 0;
assign detect_min[585][8] = (mid_1[4695:4688] < top_2[4703:4696]) ? 1 : 0;
assign detect_min[585][9] = (mid_1[4695:4688] < mid_0[4687:4680]) ? 1 : 0;
assign detect_min[585][10] = (mid_1[4695:4688] < mid_0[4695:4688]) ? 1 : 0;
assign detect_min[585][11] = (mid_1[4695:4688] < mid_0[4703:4696]) ? 1 : 0;
assign detect_min[585][12] = (mid_1[4695:4688] < mid_1[4687:4680]) ? 1 : 0;
assign detect_min[585][13] = (mid_1[4695:4688] < mid_1[4703:4696]) ? 1 : 0;
assign detect_min[585][14] = (mid_1[4695:4688] < mid_2[4687:4680]) ? 1 : 0;
assign detect_min[585][15] = (mid_1[4695:4688] < mid_2[4695:4688]) ? 1 : 0;
assign detect_min[585][16] = (mid_1[4695:4688] < mid_2[4703:4696]) ? 1 : 0;
assign detect_min[585][17] = (mid_1[4695:4688] < btm_0[4687:4680]) ? 1 : 0;
assign detect_min[585][18] = (mid_1[4695:4688] < btm_0[4695:4688]) ? 1 : 0;
assign detect_min[585][19] = (mid_1[4695:4688] < btm_0[4703:4696]) ? 1 : 0;
assign detect_min[585][20] = (mid_1[4695:4688] < btm_1[4687:4680]) ? 1 : 0;
assign detect_min[585][21] = (mid_1[4695:4688] < btm_1[4695:4688]) ? 1 : 0;
assign detect_min[585][22] = (mid_1[4695:4688] < btm_1[4703:4696]) ? 1 : 0;
assign detect_min[585][23] = (mid_1[4695:4688] < btm_2[4687:4680]) ? 1 : 0;
assign detect_min[585][24] = (mid_1[4695:4688] < btm_2[4695:4688]) ? 1 : 0;
assign detect_min[585][25] = (mid_1[4695:4688] < btm_2[4703:4696]) ? 1 : 0;

assign detect_min[586][0] = (mid_1[4703:4696] < top_0[4695:4688]) ? 1 : 0;
assign detect_min[586][1] = (mid_1[4703:4696] < top_0[4703:4696]) ? 1 : 0;
assign detect_min[586][2] = (mid_1[4703:4696] < top_0[4711:4704]) ? 1 : 0;
assign detect_min[586][3] = (mid_1[4703:4696] < top_1[4695:4688]) ? 1 : 0;
assign detect_min[586][4] = (mid_1[4703:4696] < top_1[4703:4696]) ? 1 : 0;
assign detect_min[586][5] = (mid_1[4703:4696] < top_1[4711:4704]) ? 1 : 0;
assign detect_min[586][6] = (mid_1[4703:4696] < top_2[4695:4688]) ? 1 : 0;
assign detect_min[586][7] = (mid_1[4703:4696] < top_2[4703:4696]) ? 1 : 0;
assign detect_min[586][8] = (mid_1[4703:4696] < top_2[4711:4704]) ? 1 : 0;
assign detect_min[586][9] = (mid_1[4703:4696] < mid_0[4695:4688]) ? 1 : 0;
assign detect_min[586][10] = (mid_1[4703:4696] < mid_0[4703:4696]) ? 1 : 0;
assign detect_min[586][11] = (mid_1[4703:4696] < mid_0[4711:4704]) ? 1 : 0;
assign detect_min[586][12] = (mid_1[4703:4696] < mid_1[4695:4688]) ? 1 : 0;
assign detect_min[586][13] = (mid_1[4703:4696] < mid_1[4711:4704]) ? 1 : 0;
assign detect_min[586][14] = (mid_1[4703:4696] < mid_2[4695:4688]) ? 1 : 0;
assign detect_min[586][15] = (mid_1[4703:4696] < mid_2[4703:4696]) ? 1 : 0;
assign detect_min[586][16] = (mid_1[4703:4696] < mid_2[4711:4704]) ? 1 : 0;
assign detect_min[586][17] = (mid_1[4703:4696] < btm_0[4695:4688]) ? 1 : 0;
assign detect_min[586][18] = (mid_1[4703:4696] < btm_0[4703:4696]) ? 1 : 0;
assign detect_min[586][19] = (mid_1[4703:4696] < btm_0[4711:4704]) ? 1 : 0;
assign detect_min[586][20] = (mid_1[4703:4696] < btm_1[4695:4688]) ? 1 : 0;
assign detect_min[586][21] = (mid_1[4703:4696] < btm_1[4703:4696]) ? 1 : 0;
assign detect_min[586][22] = (mid_1[4703:4696] < btm_1[4711:4704]) ? 1 : 0;
assign detect_min[586][23] = (mid_1[4703:4696] < btm_2[4695:4688]) ? 1 : 0;
assign detect_min[586][24] = (mid_1[4703:4696] < btm_2[4703:4696]) ? 1 : 0;
assign detect_min[586][25] = (mid_1[4703:4696] < btm_2[4711:4704]) ? 1 : 0;

assign detect_min[587][0] = (mid_1[4711:4704] < top_0[4703:4696]) ? 1 : 0;
assign detect_min[587][1] = (mid_1[4711:4704] < top_0[4711:4704]) ? 1 : 0;
assign detect_min[587][2] = (mid_1[4711:4704] < top_0[4719:4712]) ? 1 : 0;
assign detect_min[587][3] = (mid_1[4711:4704] < top_1[4703:4696]) ? 1 : 0;
assign detect_min[587][4] = (mid_1[4711:4704] < top_1[4711:4704]) ? 1 : 0;
assign detect_min[587][5] = (mid_1[4711:4704] < top_1[4719:4712]) ? 1 : 0;
assign detect_min[587][6] = (mid_1[4711:4704] < top_2[4703:4696]) ? 1 : 0;
assign detect_min[587][7] = (mid_1[4711:4704] < top_2[4711:4704]) ? 1 : 0;
assign detect_min[587][8] = (mid_1[4711:4704] < top_2[4719:4712]) ? 1 : 0;
assign detect_min[587][9] = (mid_1[4711:4704] < mid_0[4703:4696]) ? 1 : 0;
assign detect_min[587][10] = (mid_1[4711:4704] < mid_0[4711:4704]) ? 1 : 0;
assign detect_min[587][11] = (mid_1[4711:4704] < mid_0[4719:4712]) ? 1 : 0;
assign detect_min[587][12] = (mid_1[4711:4704] < mid_1[4703:4696]) ? 1 : 0;
assign detect_min[587][13] = (mid_1[4711:4704] < mid_1[4719:4712]) ? 1 : 0;
assign detect_min[587][14] = (mid_1[4711:4704] < mid_2[4703:4696]) ? 1 : 0;
assign detect_min[587][15] = (mid_1[4711:4704] < mid_2[4711:4704]) ? 1 : 0;
assign detect_min[587][16] = (mid_1[4711:4704] < mid_2[4719:4712]) ? 1 : 0;
assign detect_min[587][17] = (mid_1[4711:4704] < btm_0[4703:4696]) ? 1 : 0;
assign detect_min[587][18] = (mid_1[4711:4704] < btm_0[4711:4704]) ? 1 : 0;
assign detect_min[587][19] = (mid_1[4711:4704] < btm_0[4719:4712]) ? 1 : 0;
assign detect_min[587][20] = (mid_1[4711:4704] < btm_1[4703:4696]) ? 1 : 0;
assign detect_min[587][21] = (mid_1[4711:4704] < btm_1[4711:4704]) ? 1 : 0;
assign detect_min[587][22] = (mid_1[4711:4704] < btm_1[4719:4712]) ? 1 : 0;
assign detect_min[587][23] = (mid_1[4711:4704] < btm_2[4703:4696]) ? 1 : 0;
assign detect_min[587][24] = (mid_1[4711:4704] < btm_2[4711:4704]) ? 1 : 0;
assign detect_min[587][25] = (mid_1[4711:4704] < btm_2[4719:4712]) ? 1 : 0;

assign detect_min[588][0] = (mid_1[4719:4712] < top_0[4711:4704]) ? 1 : 0;
assign detect_min[588][1] = (mid_1[4719:4712] < top_0[4719:4712]) ? 1 : 0;
assign detect_min[588][2] = (mid_1[4719:4712] < top_0[4727:4720]) ? 1 : 0;
assign detect_min[588][3] = (mid_1[4719:4712] < top_1[4711:4704]) ? 1 : 0;
assign detect_min[588][4] = (mid_1[4719:4712] < top_1[4719:4712]) ? 1 : 0;
assign detect_min[588][5] = (mid_1[4719:4712] < top_1[4727:4720]) ? 1 : 0;
assign detect_min[588][6] = (mid_1[4719:4712] < top_2[4711:4704]) ? 1 : 0;
assign detect_min[588][7] = (mid_1[4719:4712] < top_2[4719:4712]) ? 1 : 0;
assign detect_min[588][8] = (mid_1[4719:4712] < top_2[4727:4720]) ? 1 : 0;
assign detect_min[588][9] = (mid_1[4719:4712] < mid_0[4711:4704]) ? 1 : 0;
assign detect_min[588][10] = (mid_1[4719:4712] < mid_0[4719:4712]) ? 1 : 0;
assign detect_min[588][11] = (mid_1[4719:4712] < mid_0[4727:4720]) ? 1 : 0;
assign detect_min[588][12] = (mid_1[4719:4712] < mid_1[4711:4704]) ? 1 : 0;
assign detect_min[588][13] = (mid_1[4719:4712] < mid_1[4727:4720]) ? 1 : 0;
assign detect_min[588][14] = (mid_1[4719:4712] < mid_2[4711:4704]) ? 1 : 0;
assign detect_min[588][15] = (mid_1[4719:4712] < mid_2[4719:4712]) ? 1 : 0;
assign detect_min[588][16] = (mid_1[4719:4712] < mid_2[4727:4720]) ? 1 : 0;
assign detect_min[588][17] = (mid_1[4719:4712] < btm_0[4711:4704]) ? 1 : 0;
assign detect_min[588][18] = (mid_1[4719:4712] < btm_0[4719:4712]) ? 1 : 0;
assign detect_min[588][19] = (mid_1[4719:4712] < btm_0[4727:4720]) ? 1 : 0;
assign detect_min[588][20] = (mid_1[4719:4712] < btm_1[4711:4704]) ? 1 : 0;
assign detect_min[588][21] = (mid_1[4719:4712] < btm_1[4719:4712]) ? 1 : 0;
assign detect_min[588][22] = (mid_1[4719:4712] < btm_1[4727:4720]) ? 1 : 0;
assign detect_min[588][23] = (mid_1[4719:4712] < btm_2[4711:4704]) ? 1 : 0;
assign detect_min[588][24] = (mid_1[4719:4712] < btm_2[4719:4712]) ? 1 : 0;
assign detect_min[588][25] = (mid_1[4719:4712] < btm_2[4727:4720]) ? 1 : 0;

assign detect_min[589][0] = (mid_1[4727:4720] < top_0[4719:4712]) ? 1 : 0;
assign detect_min[589][1] = (mid_1[4727:4720] < top_0[4727:4720]) ? 1 : 0;
assign detect_min[589][2] = (mid_1[4727:4720] < top_0[4735:4728]) ? 1 : 0;
assign detect_min[589][3] = (mid_1[4727:4720] < top_1[4719:4712]) ? 1 : 0;
assign detect_min[589][4] = (mid_1[4727:4720] < top_1[4727:4720]) ? 1 : 0;
assign detect_min[589][5] = (mid_1[4727:4720] < top_1[4735:4728]) ? 1 : 0;
assign detect_min[589][6] = (mid_1[4727:4720] < top_2[4719:4712]) ? 1 : 0;
assign detect_min[589][7] = (mid_1[4727:4720] < top_2[4727:4720]) ? 1 : 0;
assign detect_min[589][8] = (mid_1[4727:4720] < top_2[4735:4728]) ? 1 : 0;
assign detect_min[589][9] = (mid_1[4727:4720] < mid_0[4719:4712]) ? 1 : 0;
assign detect_min[589][10] = (mid_1[4727:4720] < mid_0[4727:4720]) ? 1 : 0;
assign detect_min[589][11] = (mid_1[4727:4720] < mid_0[4735:4728]) ? 1 : 0;
assign detect_min[589][12] = (mid_1[4727:4720] < mid_1[4719:4712]) ? 1 : 0;
assign detect_min[589][13] = (mid_1[4727:4720] < mid_1[4735:4728]) ? 1 : 0;
assign detect_min[589][14] = (mid_1[4727:4720] < mid_2[4719:4712]) ? 1 : 0;
assign detect_min[589][15] = (mid_1[4727:4720] < mid_2[4727:4720]) ? 1 : 0;
assign detect_min[589][16] = (mid_1[4727:4720] < mid_2[4735:4728]) ? 1 : 0;
assign detect_min[589][17] = (mid_1[4727:4720] < btm_0[4719:4712]) ? 1 : 0;
assign detect_min[589][18] = (mid_1[4727:4720] < btm_0[4727:4720]) ? 1 : 0;
assign detect_min[589][19] = (mid_1[4727:4720] < btm_0[4735:4728]) ? 1 : 0;
assign detect_min[589][20] = (mid_1[4727:4720] < btm_1[4719:4712]) ? 1 : 0;
assign detect_min[589][21] = (mid_1[4727:4720] < btm_1[4727:4720]) ? 1 : 0;
assign detect_min[589][22] = (mid_1[4727:4720] < btm_1[4735:4728]) ? 1 : 0;
assign detect_min[589][23] = (mid_1[4727:4720] < btm_2[4719:4712]) ? 1 : 0;
assign detect_min[589][24] = (mid_1[4727:4720] < btm_2[4727:4720]) ? 1 : 0;
assign detect_min[589][25] = (mid_1[4727:4720] < btm_2[4735:4728]) ? 1 : 0;

assign detect_min[590][0] = (mid_1[4735:4728] < top_0[4727:4720]) ? 1 : 0;
assign detect_min[590][1] = (mid_1[4735:4728] < top_0[4735:4728]) ? 1 : 0;
assign detect_min[590][2] = (mid_1[4735:4728] < top_0[4743:4736]) ? 1 : 0;
assign detect_min[590][3] = (mid_1[4735:4728] < top_1[4727:4720]) ? 1 : 0;
assign detect_min[590][4] = (mid_1[4735:4728] < top_1[4735:4728]) ? 1 : 0;
assign detect_min[590][5] = (mid_1[4735:4728] < top_1[4743:4736]) ? 1 : 0;
assign detect_min[590][6] = (mid_1[4735:4728] < top_2[4727:4720]) ? 1 : 0;
assign detect_min[590][7] = (mid_1[4735:4728] < top_2[4735:4728]) ? 1 : 0;
assign detect_min[590][8] = (mid_1[4735:4728] < top_2[4743:4736]) ? 1 : 0;
assign detect_min[590][9] = (mid_1[4735:4728] < mid_0[4727:4720]) ? 1 : 0;
assign detect_min[590][10] = (mid_1[4735:4728] < mid_0[4735:4728]) ? 1 : 0;
assign detect_min[590][11] = (mid_1[4735:4728] < mid_0[4743:4736]) ? 1 : 0;
assign detect_min[590][12] = (mid_1[4735:4728] < mid_1[4727:4720]) ? 1 : 0;
assign detect_min[590][13] = (mid_1[4735:4728] < mid_1[4743:4736]) ? 1 : 0;
assign detect_min[590][14] = (mid_1[4735:4728] < mid_2[4727:4720]) ? 1 : 0;
assign detect_min[590][15] = (mid_1[4735:4728] < mid_2[4735:4728]) ? 1 : 0;
assign detect_min[590][16] = (mid_1[4735:4728] < mid_2[4743:4736]) ? 1 : 0;
assign detect_min[590][17] = (mid_1[4735:4728] < btm_0[4727:4720]) ? 1 : 0;
assign detect_min[590][18] = (mid_1[4735:4728] < btm_0[4735:4728]) ? 1 : 0;
assign detect_min[590][19] = (mid_1[4735:4728] < btm_0[4743:4736]) ? 1 : 0;
assign detect_min[590][20] = (mid_1[4735:4728] < btm_1[4727:4720]) ? 1 : 0;
assign detect_min[590][21] = (mid_1[4735:4728] < btm_1[4735:4728]) ? 1 : 0;
assign detect_min[590][22] = (mid_1[4735:4728] < btm_1[4743:4736]) ? 1 : 0;
assign detect_min[590][23] = (mid_1[4735:4728] < btm_2[4727:4720]) ? 1 : 0;
assign detect_min[590][24] = (mid_1[4735:4728] < btm_2[4735:4728]) ? 1 : 0;
assign detect_min[590][25] = (mid_1[4735:4728] < btm_2[4743:4736]) ? 1 : 0;

assign detect_min[591][0] = (mid_1[4743:4736] < top_0[4735:4728]) ? 1 : 0;
assign detect_min[591][1] = (mid_1[4743:4736] < top_0[4743:4736]) ? 1 : 0;
assign detect_min[591][2] = (mid_1[4743:4736] < top_0[4751:4744]) ? 1 : 0;
assign detect_min[591][3] = (mid_1[4743:4736] < top_1[4735:4728]) ? 1 : 0;
assign detect_min[591][4] = (mid_1[4743:4736] < top_1[4743:4736]) ? 1 : 0;
assign detect_min[591][5] = (mid_1[4743:4736] < top_1[4751:4744]) ? 1 : 0;
assign detect_min[591][6] = (mid_1[4743:4736] < top_2[4735:4728]) ? 1 : 0;
assign detect_min[591][7] = (mid_1[4743:4736] < top_2[4743:4736]) ? 1 : 0;
assign detect_min[591][8] = (mid_1[4743:4736] < top_2[4751:4744]) ? 1 : 0;
assign detect_min[591][9] = (mid_1[4743:4736] < mid_0[4735:4728]) ? 1 : 0;
assign detect_min[591][10] = (mid_1[4743:4736] < mid_0[4743:4736]) ? 1 : 0;
assign detect_min[591][11] = (mid_1[4743:4736] < mid_0[4751:4744]) ? 1 : 0;
assign detect_min[591][12] = (mid_1[4743:4736] < mid_1[4735:4728]) ? 1 : 0;
assign detect_min[591][13] = (mid_1[4743:4736] < mid_1[4751:4744]) ? 1 : 0;
assign detect_min[591][14] = (mid_1[4743:4736] < mid_2[4735:4728]) ? 1 : 0;
assign detect_min[591][15] = (mid_1[4743:4736] < mid_2[4743:4736]) ? 1 : 0;
assign detect_min[591][16] = (mid_1[4743:4736] < mid_2[4751:4744]) ? 1 : 0;
assign detect_min[591][17] = (mid_1[4743:4736] < btm_0[4735:4728]) ? 1 : 0;
assign detect_min[591][18] = (mid_1[4743:4736] < btm_0[4743:4736]) ? 1 : 0;
assign detect_min[591][19] = (mid_1[4743:4736] < btm_0[4751:4744]) ? 1 : 0;
assign detect_min[591][20] = (mid_1[4743:4736] < btm_1[4735:4728]) ? 1 : 0;
assign detect_min[591][21] = (mid_1[4743:4736] < btm_1[4743:4736]) ? 1 : 0;
assign detect_min[591][22] = (mid_1[4743:4736] < btm_1[4751:4744]) ? 1 : 0;
assign detect_min[591][23] = (mid_1[4743:4736] < btm_2[4735:4728]) ? 1 : 0;
assign detect_min[591][24] = (mid_1[4743:4736] < btm_2[4743:4736]) ? 1 : 0;
assign detect_min[591][25] = (mid_1[4743:4736] < btm_2[4751:4744]) ? 1 : 0;

assign detect_min[592][0] = (mid_1[4751:4744] < top_0[4743:4736]) ? 1 : 0;
assign detect_min[592][1] = (mid_1[4751:4744] < top_0[4751:4744]) ? 1 : 0;
assign detect_min[592][2] = (mid_1[4751:4744] < top_0[4759:4752]) ? 1 : 0;
assign detect_min[592][3] = (mid_1[4751:4744] < top_1[4743:4736]) ? 1 : 0;
assign detect_min[592][4] = (mid_1[4751:4744] < top_1[4751:4744]) ? 1 : 0;
assign detect_min[592][5] = (mid_1[4751:4744] < top_1[4759:4752]) ? 1 : 0;
assign detect_min[592][6] = (mid_1[4751:4744] < top_2[4743:4736]) ? 1 : 0;
assign detect_min[592][7] = (mid_1[4751:4744] < top_2[4751:4744]) ? 1 : 0;
assign detect_min[592][8] = (mid_1[4751:4744] < top_2[4759:4752]) ? 1 : 0;
assign detect_min[592][9] = (mid_1[4751:4744] < mid_0[4743:4736]) ? 1 : 0;
assign detect_min[592][10] = (mid_1[4751:4744] < mid_0[4751:4744]) ? 1 : 0;
assign detect_min[592][11] = (mid_1[4751:4744] < mid_0[4759:4752]) ? 1 : 0;
assign detect_min[592][12] = (mid_1[4751:4744] < mid_1[4743:4736]) ? 1 : 0;
assign detect_min[592][13] = (mid_1[4751:4744] < mid_1[4759:4752]) ? 1 : 0;
assign detect_min[592][14] = (mid_1[4751:4744] < mid_2[4743:4736]) ? 1 : 0;
assign detect_min[592][15] = (mid_1[4751:4744] < mid_2[4751:4744]) ? 1 : 0;
assign detect_min[592][16] = (mid_1[4751:4744] < mid_2[4759:4752]) ? 1 : 0;
assign detect_min[592][17] = (mid_1[4751:4744] < btm_0[4743:4736]) ? 1 : 0;
assign detect_min[592][18] = (mid_1[4751:4744] < btm_0[4751:4744]) ? 1 : 0;
assign detect_min[592][19] = (mid_1[4751:4744] < btm_0[4759:4752]) ? 1 : 0;
assign detect_min[592][20] = (mid_1[4751:4744] < btm_1[4743:4736]) ? 1 : 0;
assign detect_min[592][21] = (mid_1[4751:4744] < btm_1[4751:4744]) ? 1 : 0;
assign detect_min[592][22] = (mid_1[4751:4744] < btm_1[4759:4752]) ? 1 : 0;
assign detect_min[592][23] = (mid_1[4751:4744] < btm_2[4743:4736]) ? 1 : 0;
assign detect_min[592][24] = (mid_1[4751:4744] < btm_2[4751:4744]) ? 1 : 0;
assign detect_min[592][25] = (mid_1[4751:4744] < btm_2[4759:4752]) ? 1 : 0;

assign detect_min[593][0] = (mid_1[4759:4752] < top_0[4751:4744]) ? 1 : 0;
assign detect_min[593][1] = (mid_1[4759:4752] < top_0[4759:4752]) ? 1 : 0;
assign detect_min[593][2] = (mid_1[4759:4752] < top_0[4767:4760]) ? 1 : 0;
assign detect_min[593][3] = (mid_1[4759:4752] < top_1[4751:4744]) ? 1 : 0;
assign detect_min[593][4] = (mid_1[4759:4752] < top_1[4759:4752]) ? 1 : 0;
assign detect_min[593][5] = (mid_1[4759:4752] < top_1[4767:4760]) ? 1 : 0;
assign detect_min[593][6] = (mid_1[4759:4752] < top_2[4751:4744]) ? 1 : 0;
assign detect_min[593][7] = (mid_1[4759:4752] < top_2[4759:4752]) ? 1 : 0;
assign detect_min[593][8] = (mid_1[4759:4752] < top_2[4767:4760]) ? 1 : 0;
assign detect_min[593][9] = (mid_1[4759:4752] < mid_0[4751:4744]) ? 1 : 0;
assign detect_min[593][10] = (mid_1[4759:4752] < mid_0[4759:4752]) ? 1 : 0;
assign detect_min[593][11] = (mid_1[4759:4752] < mid_0[4767:4760]) ? 1 : 0;
assign detect_min[593][12] = (mid_1[4759:4752] < mid_1[4751:4744]) ? 1 : 0;
assign detect_min[593][13] = (mid_1[4759:4752] < mid_1[4767:4760]) ? 1 : 0;
assign detect_min[593][14] = (mid_1[4759:4752] < mid_2[4751:4744]) ? 1 : 0;
assign detect_min[593][15] = (mid_1[4759:4752] < mid_2[4759:4752]) ? 1 : 0;
assign detect_min[593][16] = (mid_1[4759:4752] < mid_2[4767:4760]) ? 1 : 0;
assign detect_min[593][17] = (mid_1[4759:4752] < btm_0[4751:4744]) ? 1 : 0;
assign detect_min[593][18] = (mid_1[4759:4752] < btm_0[4759:4752]) ? 1 : 0;
assign detect_min[593][19] = (mid_1[4759:4752] < btm_0[4767:4760]) ? 1 : 0;
assign detect_min[593][20] = (mid_1[4759:4752] < btm_1[4751:4744]) ? 1 : 0;
assign detect_min[593][21] = (mid_1[4759:4752] < btm_1[4759:4752]) ? 1 : 0;
assign detect_min[593][22] = (mid_1[4759:4752] < btm_1[4767:4760]) ? 1 : 0;
assign detect_min[593][23] = (mid_1[4759:4752] < btm_2[4751:4744]) ? 1 : 0;
assign detect_min[593][24] = (mid_1[4759:4752] < btm_2[4759:4752]) ? 1 : 0;
assign detect_min[593][25] = (mid_1[4759:4752] < btm_2[4767:4760]) ? 1 : 0;

assign detect_min[594][0] = (mid_1[4767:4760] < top_0[4759:4752]) ? 1 : 0;
assign detect_min[594][1] = (mid_1[4767:4760] < top_0[4767:4760]) ? 1 : 0;
assign detect_min[594][2] = (mid_1[4767:4760] < top_0[4775:4768]) ? 1 : 0;
assign detect_min[594][3] = (mid_1[4767:4760] < top_1[4759:4752]) ? 1 : 0;
assign detect_min[594][4] = (mid_1[4767:4760] < top_1[4767:4760]) ? 1 : 0;
assign detect_min[594][5] = (mid_1[4767:4760] < top_1[4775:4768]) ? 1 : 0;
assign detect_min[594][6] = (mid_1[4767:4760] < top_2[4759:4752]) ? 1 : 0;
assign detect_min[594][7] = (mid_1[4767:4760] < top_2[4767:4760]) ? 1 : 0;
assign detect_min[594][8] = (mid_1[4767:4760] < top_2[4775:4768]) ? 1 : 0;
assign detect_min[594][9] = (mid_1[4767:4760] < mid_0[4759:4752]) ? 1 : 0;
assign detect_min[594][10] = (mid_1[4767:4760] < mid_0[4767:4760]) ? 1 : 0;
assign detect_min[594][11] = (mid_1[4767:4760] < mid_0[4775:4768]) ? 1 : 0;
assign detect_min[594][12] = (mid_1[4767:4760] < mid_1[4759:4752]) ? 1 : 0;
assign detect_min[594][13] = (mid_1[4767:4760] < mid_1[4775:4768]) ? 1 : 0;
assign detect_min[594][14] = (mid_1[4767:4760] < mid_2[4759:4752]) ? 1 : 0;
assign detect_min[594][15] = (mid_1[4767:4760] < mid_2[4767:4760]) ? 1 : 0;
assign detect_min[594][16] = (mid_1[4767:4760] < mid_2[4775:4768]) ? 1 : 0;
assign detect_min[594][17] = (mid_1[4767:4760] < btm_0[4759:4752]) ? 1 : 0;
assign detect_min[594][18] = (mid_1[4767:4760] < btm_0[4767:4760]) ? 1 : 0;
assign detect_min[594][19] = (mid_1[4767:4760] < btm_0[4775:4768]) ? 1 : 0;
assign detect_min[594][20] = (mid_1[4767:4760] < btm_1[4759:4752]) ? 1 : 0;
assign detect_min[594][21] = (mid_1[4767:4760] < btm_1[4767:4760]) ? 1 : 0;
assign detect_min[594][22] = (mid_1[4767:4760] < btm_1[4775:4768]) ? 1 : 0;
assign detect_min[594][23] = (mid_1[4767:4760] < btm_2[4759:4752]) ? 1 : 0;
assign detect_min[594][24] = (mid_1[4767:4760] < btm_2[4767:4760]) ? 1 : 0;
assign detect_min[594][25] = (mid_1[4767:4760] < btm_2[4775:4768]) ? 1 : 0;

assign detect_min[595][0] = (mid_1[4775:4768] < top_0[4767:4760]) ? 1 : 0;
assign detect_min[595][1] = (mid_1[4775:4768] < top_0[4775:4768]) ? 1 : 0;
assign detect_min[595][2] = (mid_1[4775:4768] < top_0[4783:4776]) ? 1 : 0;
assign detect_min[595][3] = (mid_1[4775:4768] < top_1[4767:4760]) ? 1 : 0;
assign detect_min[595][4] = (mid_1[4775:4768] < top_1[4775:4768]) ? 1 : 0;
assign detect_min[595][5] = (mid_1[4775:4768] < top_1[4783:4776]) ? 1 : 0;
assign detect_min[595][6] = (mid_1[4775:4768] < top_2[4767:4760]) ? 1 : 0;
assign detect_min[595][7] = (mid_1[4775:4768] < top_2[4775:4768]) ? 1 : 0;
assign detect_min[595][8] = (mid_1[4775:4768] < top_2[4783:4776]) ? 1 : 0;
assign detect_min[595][9] = (mid_1[4775:4768] < mid_0[4767:4760]) ? 1 : 0;
assign detect_min[595][10] = (mid_1[4775:4768] < mid_0[4775:4768]) ? 1 : 0;
assign detect_min[595][11] = (mid_1[4775:4768] < mid_0[4783:4776]) ? 1 : 0;
assign detect_min[595][12] = (mid_1[4775:4768] < mid_1[4767:4760]) ? 1 : 0;
assign detect_min[595][13] = (mid_1[4775:4768] < mid_1[4783:4776]) ? 1 : 0;
assign detect_min[595][14] = (mid_1[4775:4768] < mid_2[4767:4760]) ? 1 : 0;
assign detect_min[595][15] = (mid_1[4775:4768] < mid_2[4775:4768]) ? 1 : 0;
assign detect_min[595][16] = (mid_1[4775:4768] < mid_2[4783:4776]) ? 1 : 0;
assign detect_min[595][17] = (mid_1[4775:4768] < btm_0[4767:4760]) ? 1 : 0;
assign detect_min[595][18] = (mid_1[4775:4768] < btm_0[4775:4768]) ? 1 : 0;
assign detect_min[595][19] = (mid_1[4775:4768] < btm_0[4783:4776]) ? 1 : 0;
assign detect_min[595][20] = (mid_1[4775:4768] < btm_1[4767:4760]) ? 1 : 0;
assign detect_min[595][21] = (mid_1[4775:4768] < btm_1[4775:4768]) ? 1 : 0;
assign detect_min[595][22] = (mid_1[4775:4768] < btm_1[4783:4776]) ? 1 : 0;
assign detect_min[595][23] = (mid_1[4775:4768] < btm_2[4767:4760]) ? 1 : 0;
assign detect_min[595][24] = (mid_1[4775:4768] < btm_2[4775:4768]) ? 1 : 0;
assign detect_min[595][25] = (mid_1[4775:4768] < btm_2[4783:4776]) ? 1 : 0;

assign detect_min[596][0] = (mid_1[4783:4776] < top_0[4775:4768]) ? 1 : 0;
assign detect_min[596][1] = (mid_1[4783:4776] < top_0[4783:4776]) ? 1 : 0;
assign detect_min[596][2] = (mid_1[4783:4776] < top_0[4791:4784]) ? 1 : 0;
assign detect_min[596][3] = (mid_1[4783:4776] < top_1[4775:4768]) ? 1 : 0;
assign detect_min[596][4] = (mid_1[4783:4776] < top_1[4783:4776]) ? 1 : 0;
assign detect_min[596][5] = (mid_1[4783:4776] < top_1[4791:4784]) ? 1 : 0;
assign detect_min[596][6] = (mid_1[4783:4776] < top_2[4775:4768]) ? 1 : 0;
assign detect_min[596][7] = (mid_1[4783:4776] < top_2[4783:4776]) ? 1 : 0;
assign detect_min[596][8] = (mid_1[4783:4776] < top_2[4791:4784]) ? 1 : 0;
assign detect_min[596][9] = (mid_1[4783:4776] < mid_0[4775:4768]) ? 1 : 0;
assign detect_min[596][10] = (mid_1[4783:4776] < mid_0[4783:4776]) ? 1 : 0;
assign detect_min[596][11] = (mid_1[4783:4776] < mid_0[4791:4784]) ? 1 : 0;
assign detect_min[596][12] = (mid_1[4783:4776] < mid_1[4775:4768]) ? 1 : 0;
assign detect_min[596][13] = (mid_1[4783:4776] < mid_1[4791:4784]) ? 1 : 0;
assign detect_min[596][14] = (mid_1[4783:4776] < mid_2[4775:4768]) ? 1 : 0;
assign detect_min[596][15] = (mid_1[4783:4776] < mid_2[4783:4776]) ? 1 : 0;
assign detect_min[596][16] = (mid_1[4783:4776] < mid_2[4791:4784]) ? 1 : 0;
assign detect_min[596][17] = (mid_1[4783:4776] < btm_0[4775:4768]) ? 1 : 0;
assign detect_min[596][18] = (mid_1[4783:4776] < btm_0[4783:4776]) ? 1 : 0;
assign detect_min[596][19] = (mid_1[4783:4776] < btm_0[4791:4784]) ? 1 : 0;
assign detect_min[596][20] = (mid_1[4783:4776] < btm_1[4775:4768]) ? 1 : 0;
assign detect_min[596][21] = (mid_1[4783:4776] < btm_1[4783:4776]) ? 1 : 0;
assign detect_min[596][22] = (mid_1[4783:4776] < btm_1[4791:4784]) ? 1 : 0;
assign detect_min[596][23] = (mid_1[4783:4776] < btm_2[4775:4768]) ? 1 : 0;
assign detect_min[596][24] = (mid_1[4783:4776] < btm_2[4783:4776]) ? 1 : 0;
assign detect_min[596][25] = (mid_1[4783:4776] < btm_2[4791:4784]) ? 1 : 0;

assign detect_min[597][0] = (mid_1[4791:4784] < top_0[4783:4776]) ? 1 : 0;
assign detect_min[597][1] = (mid_1[4791:4784] < top_0[4791:4784]) ? 1 : 0;
assign detect_min[597][2] = (mid_1[4791:4784] < top_0[4799:4792]) ? 1 : 0;
assign detect_min[597][3] = (mid_1[4791:4784] < top_1[4783:4776]) ? 1 : 0;
assign detect_min[597][4] = (mid_1[4791:4784] < top_1[4791:4784]) ? 1 : 0;
assign detect_min[597][5] = (mid_1[4791:4784] < top_1[4799:4792]) ? 1 : 0;
assign detect_min[597][6] = (mid_1[4791:4784] < top_2[4783:4776]) ? 1 : 0;
assign detect_min[597][7] = (mid_1[4791:4784] < top_2[4791:4784]) ? 1 : 0;
assign detect_min[597][8] = (mid_1[4791:4784] < top_2[4799:4792]) ? 1 : 0;
assign detect_min[597][9] = (mid_1[4791:4784] < mid_0[4783:4776]) ? 1 : 0;
assign detect_min[597][10] = (mid_1[4791:4784] < mid_0[4791:4784]) ? 1 : 0;
assign detect_min[597][11] = (mid_1[4791:4784] < mid_0[4799:4792]) ? 1 : 0;
assign detect_min[597][12] = (mid_1[4791:4784] < mid_1[4783:4776]) ? 1 : 0;
assign detect_min[597][13] = (mid_1[4791:4784] < mid_1[4799:4792]) ? 1 : 0;
assign detect_min[597][14] = (mid_1[4791:4784] < mid_2[4783:4776]) ? 1 : 0;
assign detect_min[597][15] = (mid_1[4791:4784] < mid_2[4791:4784]) ? 1 : 0;
assign detect_min[597][16] = (mid_1[4791:4784] < mid_2[4799:4792]) ? 1 : 0;
assign detect_min[597][17] = (mid_1[4791:4784] < btm_0[4783:4776]) ? 1 : 0;
assign detect_min[597][18] = (mid_1[4791:4784] < btm_0[4791:4784]) ? 1 : 0;
assign detect_min[597][19] = (mid_1[4791:4784] < btm_0[4799:4792]) ? 1 : 0;
assign detect_min[597][20] = (mid_1[4791:4784] < btm_1[4783:4776]) ? 1 : 0;
assign detect_min[597][21] = (mid_1[4791:4784] < btm_1[4791:4784]) ? 1 : 0;
assign detect_min[597][22] = (mid_1[4791:4784] < btm_1[4799:4792]) ? 1 : 0;
assign detect_min[597][23] = (mid_1[4791:4784] < btm_2[4783:4776]) ? 1 : 0;
assign detect_min[597][24] = (mid_1[4791:4784] < btm_2[4791:4784]) ? 1 : 0;
assign detect_min[597][25] = (mid_1[4791:4784] < btm_2[4799:4792]) ? 1 : 0;

assign detect_min[598][0] = (mid_1[4799:4792] < top_0[4791:4784]) ? 1 : 0;
assign detect_min[598][1] = (mid_1[4799:4792] < top_0[4799:4792]) ? 1 : 0;
assign detect_min[598][2] = (mid_1[4799:4792] < top_0[4807:4800]) ? 1 : 0;
assign detect_min[598][3] = (mid_1[4799:4792] < top_1[4791:4784]) ? 1 : 0;
assign detect_min[598][4] = (mid_1[4799:4792] < top_1[4799:4792]) ? 1 : 0;
assign detect_min[598][5] = (mid_1[4799:4792] < top_1[4807:4800]) ? 1 : 0;
assign detect_min[598][6] = (mid_1[4799:4792] < top_2[4791:4784]) ? 1 : 0;
assign detect_min[598][7] = (mid_1[4799:4792] < top_2[4799:4792]) ? 1 : 0;
assign detect_min[598][8] = (mid_1[4799:4792] < top_2[4807:4800]) ? 1 : 0;
assign detect_min[598][9] = (mid_1[4799:4792] < mid_0[4791:4784]) ? 1 : 0;
assign detect_min[598][10] = (mid_1[4799:4792] < mid_0[4799:4792]) ? 1 : 0;
assign detect_min[598][11] = (mid_1[4799:4792] < mid_0[4807:4800]) ? 1 : 0;
assign detect_min[598][12] = (mid_1[4799:4792] < mid_1[4791:4784]) ? 1 : 0;
assign detect_min[598][13] = (mid_1[4799:4792] < mid_1[4807:4800]) ? 1 : 0;
assign detect_min[598][14] = (mid_1[4799:4792] < mid_2[4791:4784]) ? 1 : 0;
assign detect_min[598][15] = (mid_1[4799:4792] < mid_2[4799:4792]) ? 1 : 0;
assign detect_min[598][16] = (mid_1[4799:4792] < mid_2[4807:4800]) ? 1 : 0;
assign detect_min[598][17] = (mid_1[4799:4792] < btm_0[4791:4784]) ? 1 : 0;
assign detect_min[598][18] = (mid_1[4799:4792] < btm_0[4799:4792]) ? 1 : 0;
assign detect_min[598][19] = (mid_1[4799:4792] < btm_0[4807:4800]) ? 1 : 0;
assign detect_min[598][20] = (mid_1[4799:4792] < btm_1[4791:4784]) ? 1 : 0;
assign detect_min[598][21] = (mid_1[4799:4792] < btm_1[4799:4792]) ? 1 : 0;
assign detect_min[598][22] = (mid_1[4799:4792] < btm_1[4807:4800]) ? 1 : 0;
assign detect_min[598][23] = (mid_1[4799:4792] < btm_2[4791:4784]) ? 1 : 0;
assign detect_min[598][24] = (mid_1[4799:4792] < btm_2[4799:4792]) ? 1 : 0;
assign detect_min[598][25] = (mid_1[4799:4792] < btm_2[4807:4800]) ? 1 : 0;

assign detect_min[599][0] = (mid_1[4807:4800] < top_0[4799:4792]) ? 1 : 0;
assign detect_min[599][1] = (mid_1[4807:4800] < top_0[4807:4800]) ? 1 : 0;
assign detect_min[599][2] = (mid_1[4807:4800] < top_0[4815:4808]) ? 1 : 0;
assign detect_min[599][3] = (mid_1[4807:4800] < top_1[4799:4792]) ? 1 : 0;
assign detect_min[599][4] = (mid_1[4807:4800] < top_1[4807:4800]) ? 1 : 0;
assign detect_min[599][5] = (mid_1[4807:4800] < top_1[4815:4808]) ? 1 : 0;
assign detect_min[599][6] = (mid_1[4807:4800] < top_2[4799:4792]) ? 1 : 0;
assign detect_min[599][7] = (mid_1[4807:4800] < top_2[4807:4800]) ? 1 : 0;
assign detect_min[599][8] = (mid_1[4807:4800] < top_2[4815:4808]) ? 1 : 0;
assign detect_min[599][9] = (mid_1[4807:4800] < mid_0[4799:4792]) ? 1 : 0;
assign detect_min[599][10] = (mid_1[4807:4800] < mid_0[4807:4800]) ? 1 : 0;
assign detect_min[599][11] = (mid_1[4807:4800] < mid_0[4815:4808]) ? 1 : 0;
assign detect_min[599][12] = (mid_1[4807:4800] < mid_1[4799:4792]) ? 1 : 0;
assign detect_min[599][13] = (mid_1[4807:4800] < mid_1[4815:4808]) ? 1 : 0;
assign detect_min[599][14] = (mid_1[4807:4800] < mid_2[4799:4792]) ? 1 : 0;
assign detect_min[599][15] = (mid_1[4807:4800] < mid_2[4807:4800]) ? 1 : 0;
assign detect_min[599][16] = (mid_1[4807:4800] < mid_2[4815:4808]) ? 1 : 0;
assign detect_min[599][17] = (mid_1[4807:4800] < btm_0[4799:4792]) ? 1 : 0;
assign detect_min[599][18] = (mid_1[4807:4800] < btm_0[4807:4800]) ? 1 : 0;
assign detect_min[599][19] = (mid_1[4807:4800] < btm_0[4815:4808]) ? 1 : 0;
assign detect_min[599][20] = (mid_1[4807:4800] < btm_1[4799:4792]) ? 1 : 0;
assign detect_min[599][21] = (mid_1[4807:4800] < btm_1[4807:4800]) ? 1 : 0;
assign detect_min[599][22] = (mid_1[4807:4800] < btm_1[4815:4808]) ? 1 : 0;
assign detect_min[599][23] = (mid_1[4807:4800] < btm_2[4799:4792]) ? 1 : 0;
assign detect_min[599][24] = (mid_1[4807:4800] < btm_2[4807:4800]) ? 1 : 0;
assign detect_min[599][25] = (mid_1[4807:4800] < btm_2[4815:4808]) ? 1 : 0;

assign detect_min[600][0] = (mid_1[4815:4808] < top_0[4807:4800]) ? 1 : 0;
assign detect_min[600][1] = (mid_1[4815:4808] < top_0[4815:4808]) ? 1 : 0;
assign detect_min[600][2] = (mid_1[4815:4808] < top_0[4823:4816]) ? 1 : 0;
assign detect_min[600][3] = (mid_1[4815:4808] < top_1[4807:4800]) ? 1 : 0;
assign detect_min[600][4] = (mid_1[4815:4808] < top_1[4815:4808]) ? 1 : 0;
assign detect_min[600][5] = (mid_1[4815:4808] < top_1[4823:4816]) ? 1 : 0;
assign detect_min[600][6] = (mid_1[4815:4808] < top_2[4807:4800]) ? 1 : 0;
assign detect_min[600][7] = (mid_1[4815:4808] < top_2[4815:4808]) ? 1 : 0;
assign detect_min[600][8] = (mid_1[4815:4808] < top_2[4823:4816]) ? 1 : 0;
assign detect_min[600][9] = (mid_1[4815:4808] < mid_0[4807:4800]) ? 1 : 0;
assign detect_min[600][10] = (mid_1[4815:4808] < mid_0[4815:4808]) ? 1 : 0;
assign detect_min[600][11] = (mid_1[4815:4808] < mid_0[4823:4816]) ? 1 : 0;
assign detect_min[600][12] = (mid_1[4815:4808] < mid_1[4807:4800]) ? 1 : 0;
assign detect_min[600][13] = (mid_1[4815:4808] < mid_1[4823:4816]) ? 1 : 0;
assign detect_min[600][14] = (mid_1[4815:4808] < mid_2[4807:4800]) ? 1 : 0;
assign detect_min[600][15] = (mid_1[4815:4808] < mid_2[4815:4808]) ? 1 : 0;
assign detect_min[600][16] = (mid_1[4815:4808] < mid_2[4823:4816]) ? 1 : 0;
assign detect_min[600][17] = (mid_1[4815:4808] < btm_0[4807:4800]) ? 1 : 0;
assign detect_min[600][18] = (mid_1[4815:4808] < btm_0[4815:4808]) ? 1 : 0;
assign detect_min[600][19] = (mid_1[4815:4808] < btm_0[4823:4816]) ? 1 : 0;
assign detect_min[600][20] = (mid_1[4815:4808] < btm_1[4807:4800]) ? 1 : 0;
assign detect_min[600][21] = (mid_1[4815:4808] < btm_1[4815:4808]) ? 1 : 0;
assign detect_min[600][22] = (mid_1[4815:4808] < btm_1[4823:4816]) ? 1 : 0;
assign detect_min[600][23] = (mid_1[4815:4808] < btm_2[4807:4800]) ? 1 : 0;
assign detect_min[600][24] = (mid_1[4815:4808] < btm_2[4815:4808]) ? 1 : 0;
assign detect_min[600][25] = (mid_1[4815:4808] < btm_2[4823:4816]) ? 1 : 0;

assign detect_min[601][0] = (mid_1[4823:4816] < top_0[4815:4808]) ? 1 : 0;
assign detect_min[601][1] = (mid_1[4823:4816] < top_0[4823:4816]) ? 1 : 0;
assign detect_min[601][2] = (mid_1[4823:4816] < top_0[4831:4824]) ? 1 : 0;
assign detect_min[601][3] = (mid_1[4823:4816] < top_1[4815:4808]) ? 1 : 0;
assign detect_min[601][4] = (mid_1[4823:4816] < top_1[4823:4816]) ? 1 : 0;
assign detect_min[601][5] = (mid_1[4823:4816] < top_1[4831:4824]) ? 1 : 0;
assign detect_min[601][6] = (mid_1[4823:4816] < top_2[4815:4808]) ? 1 : 0;
assign detect_min[601][7] = (mid_1[4823:4816] < top_2[4823:4816]) ? 1 : 0;
assign detect_min[601][8] = (mid_1[4823:4816] < top_2[4831:4824]) ? 1 : 0;
assign detect_min[601][9] = (mid_1[4823:4816] < mid_0[4815:4808]) ? 1 : 0;
assign detect_min[601][10] = (mid_1[4823:4816] < mid_0[4823:4816]) ? 1 : 0;
assign detect_min[601][11] = (mid_1[4823:4816] < mid_0[4831:4824]) ? 1 : 0;
assign detect_min[601][12] = (mid_1[4823:4816] < mid_1[4815:4808]) ? 1 : 0;
assign detect_min[601][13] = (mid_1[4823:4816] < mid_1[4831:4824]) ? 1 : 0;
assign detect_min[601][14] = (mid_1[4823:4816] < mid_2[4815:4808]) ? 1 : 0;
assign detect_min[601][15] = (mid_1[4823:4816] < mid_2[4823:4816]) ? 1 : 0;
assign detect_min[601][16] = (mid_1[4823:4816] < mid_2[4831:4824]) ? 1 : 0;
assign detect_min[601][17] = (mid_1[4823:4816] < btm_0[4815:4808]) ? 1 : 0;
assign detect_min[601][18] = (mid_1[4823:4816] < btm_0[4823:4816]) ? 1 : 0;
assign detect_min[601][19] = (mid_1[4823:4816] < btm_0[4831:4824]) ? 1 : 0;
assign detect_min[601][20] = (mid_1[4823:4816] < btm_1[4815:4808]) ? 1 : 0;
assign detect_min[601][21] = (mid_1[4823:4816] < btm_1[4823:4816]) ? 1 : 0;
assign detect_min[601][22] = (mid_1[4823:4816] < btm_1[4831:4824]) ? 1 : 0;
assign detect_min[601][23] = (mid_1[4823:4816] < btm_2[4815:4808]) ? 1 : 0;
assign detect_min[601][24] = (mid_1[4823:4816] < btm_2[4823:4816]) ? 1 : 0;
assign detect_min[601][25] = (mid_1[4823:4816] < btm_2[4831:4824]) ? 1 : 0;

assign detect_min[602][0] = (mid_1[4831:4824] < top_0[4823:4816]) ? 1 : 0;
assign detect_min[602][1] = (mid_1[4831:4824] < top_0[4831:4824]) ? 1 : 0;
assign detect_min[602][2] = (mid_1[4831:4824] < top_0[4839:4832]) ? 1 : 0;
assign detect_min[602][3] = (mid_1[4831:4824] < top_1[4823:4816]) ? 1 : 0;
assign detect_min[602][4] = (mid_1[4831:4824] < top_1[4831:4824]) ? 1 : 0;
assign detect_min[602][5] = (mid_1[4831:4824] < top_1[4839:4832]) ? 1 : 0;
assign detect_min[602][6] = (mid_1[4831:4824] < top_2[4823:4816]) ? 1 : 0;
assign detect_min[602][7] = (mid_1[4831:4824] < top_2[4831:4824]) ? 1 : 0;
assign detect_min[602][8] = (mid_1[4831:4824] < top_2[4839:4832]) ? 1 : 0;
assign detect_min[602][9] = (mid_1[4831:4824] < mid_0[4823:4816]) ? 1 : 0;
assign detect_min[602][10] = (mid_1[4831:4824] < mid_0[4831:4824]) ? 1 : 0;
assign detect_min[602][11] = (mid_1[4831:4824] < mid_0[4839:4832]) ? 1 : 0;
assign detect_min[602][12] = (mid_1[4831:4824] < mid_1[4823:4816]) ? 1 : 0;
assign detect_min[602][13] = (mid_1[4831:4824] < mid_1[4839:4832]) ? 1 : 0;
assign detect_min[602][14] = (mid_1[4831:4824] < mid_2[4823:4816]) ? 1 : 0;
assign detect_min[602][15] = (mid_1[4831:4824] < mid_2[4831:4824]) ? 1 : 0;
assign detect_min[602][16] = (mid_1[4831:4824] < mid_2[4839:4832]) ? 1 : 0;
assign detect_min[602][17] = (mid_1[4831:4824] < btm_0[4823:4816]) ? 1 : 0;
assign detect_min[602][18] = (mid_1[4831:4824] < btm_0[4831:4824]) ? 1 : 0;
assign detect_min[602][19] = (mid_1[4831:4824] < btm_0[4839:4832]) ? 1 : 0;
assign detect_min[602][20] = (mid_1[4831:4824] < btm_1[4823:4816]) ? 1 : 0;
assign detect_min[602][21] = (mid_1[4831:4824] < btm_1[4831:4824]) ? 1 : 0;
assign detect_min[602][22] = (mid_1[4831:4824] < btm_1[4839:4832]) ? 1 : 0;
assign detect_min[602][23] = (mid_1[4831:4824] < btm_2[4823:4816]) ? 1 : 0;
assign detect_min[602][24] = (mid_1[4831:4824] < btm_2[4831:4824]) ? 1 : 0;
assign detect_min[602][25] = (mid_1[4831:4824] < btm_2[4839:4832]) ? 1 : 0;

assign detect_min[603][0] = (mid_1[4839:4832] < top_0[4831:4824]) ? 1 : 0;
assign detect_min[603][1] = (mid_1[4839:4832] < top_0[4839:4832]) ? 1 : 0;
assign detect_min[603][2] = (mid_1[4839:4832] < top_0[4847:4840]) ? 1 : 0;
assign detect_min[603][3] = (mid_1[4839:4832] < top_1[4831:4824]) ? 1 : 0;
assign detect_min[603][4] = (mid_1[4839:4832] < top_1[4839:4832]) ? 1 : 0;
assign detect_min[603][5] = (mid_1[4839:4832] < top_1[4847:4840]) ? 1 : 0;
assign detect_min[603][6] = (mid_1[4839:4832] < top_2[4831:4824]) ? 1 : 0;
assign detect_min[603][7] = (mid_1[4839:4832] < top_2[4839:4832]) ? 1 : 0;
assign detect_min[603][8] = (mid_1[4839:4832] < top_2[4847:4840]) ? 1 : 0;
assign detect_min[603][9] = (mid_1[4839:4832] < mid_0[4831:4824]) ? 1 : 0;
assign detect_min[603][10] = (mid_1[4839:4832] < mid_0[4839:4832]) ? 1 : 0;
assign detect_min[603][11] = (mid_1[4839:4832] < mid_0[4847:4840]) ? 1 : 0;
assign detect_min[603][12] = (mid_1[4839:4832] < mid_1[4831:4824]) ? 1 : 0;
assign detect_min[603][13] = (mid_1[4839:4832] < mid_1[4847:4840]) ? 1 : 0;
assign detect_min[603][14] = (mid_1[4839:4832] < mid_2[4831:4824]) ? 1 : 0;
assign detect_min[603][15] = (mid_1[4839:4832] < mid_2[4839:4832]) ? 1 : 0;
assign detect_min[603][16] = (mid_1[4839:4832] < mid_2[4847:4840]) ? 1 : 0;
assign detect_min[603][17] = (mid_1[4839:4832] < btm_0[4831:4824]) ? 1 : 0;
assign detect_min[603][18] = (mid_1[4839:4832] < btm_0[4839:4832]) ? 1 : 0;
assign detect_min[603][19] = (mid_1[4839:4832] < btm_0[4847:4840]) ? 1 : 0;
assign detect_min[603][20] = (mid_1[4839:4832] < btm_1[4831:4824]) ? 1 : 0;
assign detect_min[603][21] = (mid_1[4839:4832] < btm_1[4839:4832]) ? 1 : 0;
assign detect_min[603][22] = (mid_1[4839:4832] < btm_1[4847:4840]) ? 1 : 0;
assign detect_min[603][23] = (mid_1[4839:4832] < btm_2[4831:4824]) ? 1 : 0;
assign detect_min[603][24] = (mid_1[4839:4832] < btm_2[4839:4832]) ? 1 : 0;
assign detect_min[603][25] = (mid_1[4839:4832] < btm_2[4847:4840]) ? 1 : 0;

assign detect_min[604][0] = (mid_1[4847:4840] < top_0[4839:4832]) ? 1 : 0;
assign detect_min[604][1] = (mid_1[4847:4840] < top_0[4847:4840]) ? 1 : 0;
assign detect_min[604][2] = (mid_1[4847:4840] < top_0[4855:4848]) ? 1 : 0;
assign detect_min[604][3] = (mid_1[4847:4840] < top_1[4839:4832]) ? 1 : 0;
assign detect_min[604][4] = (mid_1[4847:4840] < top_1[4847:4840]) ? 1 : 0;
assign detect_min[604][5] = (mid_1[4847:4840] < top_1[4855:4848]) ? 1 : 0;
assign detect_min[604][6] = (mid_1[4847:4840] < top_2[4839:4832]) ? 1 : 0;
assign detect_min[604][7] = (mid_1[4847:4840] < top_2[4847:4840]) ? 1 : 0;
assign detect_min[604][8] = (mid_1[4847:4840] < top_2[4855:4848]) ? 1 : 0;
assign detect_min[604][9] = (mid_1[4847:4840] < mid_0[4839:4832]) ? 1 : 0;
assign detect_min[604][10] = (mid_1[4847:4840] < mid_0[4847:4840]) ? 1 : 0;
assign detect_min[604][11] = (mid_1[4847:4840] < mid_0[4855:4848]) ? 1 : 0;
assign detect_min[604][12] = (mid_1[4847:4840] < mid_1[4839:4832]) ? 1 : 0;
assign detect_min[604][13] = (mid_1[4847:4840] < mid_1[4855:4848]) ? 1 : 0;
assign detect_min[604][14] = (mid_1[4847:4840] < mid_2[4839:4832]) ? 1 : 0;
assign detect_min[604][15] = (mid_1[4847:4840] < mid_2[4847:4840]) ? 1 : 0;
assign detect_min[604][16] = (mid_1[4847:4840] < mid_2[4855:4848]) ? 1 : 0;
assign detect_min[604][17] = (mid_1[4847:4840] < btm_0[4839:4832]) ? 1 : 0;
assign detect_min[604][18] = (mid_1[4847:4840] < btm_0[4847:4840]) ? 1 : 0;
assign detect_min[604][19] = (mid_1[4847:4840] < btm_0[4855:4848]) ? 1 : 0;
assign detect_min[604][20] = (mid_1[4847:4840] < btm_1[4839:4832]) ? 1 : 0;
assign detect_min[604][21] = (mid_1[4847:4840] < btm_1[4847:4840]) ? 1 : 0;
assign detect_min[604][22] = (mid_1[4847:4840] < btm_1[4855:4848]) ? 1 : 0;
assign detect_min[604][23] = (mid_1[4847:4840] < btm_2[4839:4832]) ? 1 : 0;
assign detect_min[604][24] = (mid_1[4847:4840] < btm_2[4847:4840]) ? 1 : 0;
assign detect_min[604][25] = (mid_1[4847:4840] < btm_2[4855:4848]) ? 1 : 0;

assign detect_min[605][0] = (mid_1[4855:4848] < top_0[4847:4840]) ? 1 : 0;
assign detect_min[605][1] = (mid_1[4855:4848] < top_0[4855:4848]) ? 1 : 0;
assign detect_min[605][2] = (mid_1[4855:4848] < top_0[4863:4856]) ? 1 : 0;
assign detect_min[605][3] = (mid_1[4855:4848] < top_1[4847:4840]) ? 1 : 0;
assign detect_min[605][4] = (mid_1[4855:4848] < top_1[4855:4848]) ? 1 : 0;
assign detect_min[605][5] = (mid_1[4855:4848] < top_1[4863:4856]) ? 1 : 0;
assign detect_min[605][6] = (mid_1[4855:4848] < top_2[4847:4840]) ? 1 : 0;
assign detect_min[605][7] = (mid_1[4855:4848] < top_2[4855:4848]) ? 1 : 0;
assign detect_min[605][8] = (mid_1[4855:4848] < top_2[4863:4856]) ? 1 : 0;
assign detect_min[605][9] = (mid_1[4855:4848] < mid_0[4847:4840]) ? 1 : 0;
assign detect_min[605][10] = (mid_1[4855:4848] < mid_0[4855:4848]) ? 1 : 0;
assign detect_min[605][11] = (mid_1[4855:4848] < mid_0[4863:4856]) ? 1 : 0;
assign detect_min[605][12] = (mid_1[4855:4848] < mid_1[4847:4840]) ? 1 : 0;
assign detect_min[605][13] = (mid_1[4855:4848] < mid_1[4863:4856]) ? 1 : 0;
assign detect_min[605][14] = (mid_1[4855:4848] < mid_2[4847:4840]) ? 1 : 0;
assign detect_min[605][15] = (mid_1[4855:4848] < mid_2[4855:4848]) ? 1 : 0;
assign detect_min[605][16] = (mid_1[4855:4848] < mid_2[4863:4856]) ? 1 : 0;
assign detect_min[605][17] = (mid_1[4855:4848] < btm_0[4847:4840]) ? 1 : 0;
assign detect_min[605][18] = (mid_1[4855:4848] < btm_0[4855:4848]) ? 1 : 0;
assign detect_min[605][19] = (mid_1[4855:4848] < btm_0[4863:4856]) ? 1 : 0;
assign detect_min[605][20] = (mid_1[4855:4848] < btm_1[4847:4840]) ? 1 : 0;
assign detect_min[605][21] = (mid_1[4855:4848] < btm_1[4855:4848]) ? 1 : 0;
assign detect_min[605][22] = (mid_1[4855:4848] < btm_1[4863:4856]) ? 1 : 0;
assign detect_min[605][23] = (mid_1[4855:4848] < btm_2[4847:4840]) ? 1 : 0;
assign detect_min[605][24] = (mid_1[4855:4848] < btm_2[4855:4848]) ? 1 : 0;
assign detect_min[605][25] = (mid_1[4855:4848] < btm_2[4863:4856]) ? 1 : 0;

assign detect_min[606][0] = (mid_1[4863:4856] < top_0[4855:4848]) ? 1 : 0;
assign detect_min[606][1] = (mid_1[4863:4856] < top_0[4863:4856]) ? 1 : 0;
assign detect_min[606][2] = (mid_1[4863:4856] < top_0[4871:4864]) ? 1 : 0;
assign detect_min[606][3] = (mid_1[4863:4856] < top_1[4855:4848]) ? 1 : 0;
assign detect_min[606][4] = (mid_1[4863:4856] < top_1[4863:4856]) ? 1 : 0;
assign detect_min[606][5] = (mid_1[4863:4856] < top_1[4871:4864]) ? 1 : 0;
assign detect_min[606][6] = (mid_1[4863:4856] < top_2[4855:4848]) ? 1 : 0;
assign detect_min[606][7] = (mid_1[4863:4856] < top_2[4863:4856]) ? 1 : 0;
assign detect_min[606][8] = (mid_1[4863:4856] < top_2[4871:4864]) ? 1 : 0;
assign detect_min[606][9] = (mid_1[4863:4856] < mid_0[4855:4848]) ? 1 : 0;
assign detect_min[606][10] = (mid_1[4863:4856] < mid_0[4863:4856]) ? 1 : 0;
assign detect_min[606][11] = (mid_1[4863:4856] < mid_0[4871:4864]) ? 1 : 0;
assign detect_min[606][12] = (mid_1[4863:4856] < mid_1[4855:4848]) ? 1 : 0;
assign detect_min[606][13] = (mid_1[4863:4856] < mid_1[4871:4864]) ? 1 : 0;
assign detect_min[606][14] = (mid_1[4863:4856] < mid_2[4855:4848]) ? 1 : 0;
assign detect_min[606][15] = (mid_1[4863:4856] < mid_2[4863:4856]) ? 1 : 0;
assign detect_min[606][16] = (mid_1[4863:4856] < mid_2[4871:4864]) ? 1 : 0;
assign detect_min[606][17] = (mid_1[4863:4856] < btm_0[4855:4848]) ? 1 : 0;
assign detect_min[606][18] = (mid_1[4863:4856] < btm_0[4863:4856]) ? 1 : 0;
assign detect_min[606][19] = (mid_1[4863:4856] < btm_0[4871:4864]) ? 1 : 0;
assign detect_min[606][20] = (mid_1[4863:4856] < btm_1[4855:4848]) ? 1 : 0;
assign detect_min[606][21] = (mid_1[4863:4856] < btm_1[4863:4856]) ? 1 : 0;
assign detect_min[606][22] = (mid_1[4863:4856] < btm_1[4871:4864]) ? 1 : 0;
assign detect_min[606][23] = (mid_1[4863:4856] < btm_2[4855:4848]) ? 1 : 0;
assign detect_min[606][24] = (mid_1[4863:4856] < btm_2[4863:4856]) ? 1 : 0;
assign detect_min[606][25] = (mid_1[4863:4856] < btm_2[4871:4864]) ? 1 : 0;

assign detect_min[607][0] = (mid_1[4871:4864] < top_0[4863:4856]) ? 1 : 0;
assign detect_min[607][1] = (mid_1[4871:4864] < top_0[4871:4864]) ? 1 : 0;
assign detect_min[607][2] = (mid_1[4871:4864] < top_0[4879:4872]) ? 1 : 0;
assign detect_min[607][3] = (mid_1[4871:4864] < top_1[4863:4856]) ? 1 : 0;
assign detect_min[607][4] = (mid_1[4871:4864] < top_1[4871:4864]) ? 1 : 0;
assign detect_min[607][5] = (mid_1[4871:4864] < top_1[4879:4872]) ? 1 : 0;
assign detect_min[607][6] = (mid_1[4871:4864] < top_2[4863:4856]) ? 1 : 0;
assign detect_min[607][7] = (mid_1[4871:4864] < top_2[4871:4864]) ? 1 : 0;
assign detect_min[607][8] = (mid_1[4871:4864] < top_2[4879:4872]) ? 1 : 0;
assign detect_min[607][9] = (mid_1[4871:4864] < mid_0[4863:4856]) ? 1 : 0;
assign detect_min[607][10] = (mid_1[4871:4864] < mid_0[4871:4864]) ? 1 : 0;
assign detect_min[607][11] = (mid_1[4871:4864] < mid_0[4879:4872]) ? 1 : 0;
assign detect_min[607][12] = (mid_1[4871:4864] < mid_1[4863:4856]) ? 1 : 0;
assign detect_min[607][13] = (mid_1[4871:4864] < mid_1[4879:4872]) ? 1 : 0;
assign detect_min[607][14] = (mid_1[4871:4864] < mid_2[4863:4856]) ? 1 : 0;
assign detect_min[607][15] = (mid_1[4871:4864] < mid_2[4871:4864]) ? 1 : 0;
assign detect_min[607][16] = (mid_1[4871:4864] < mid_2[4879:4872]) ? 1 : 0;
assign detect_min[607][17] = (mid_1[4871:4864] < btm_0[4863:4856]) ? 1 : 0;
assign detect_min[607][18] = (mid_1[4871:4864] < btm_0[4871:4864]) ? 1 : 0;
assign detect_min[607][19] = (mid_1[4871:4864] < btm_0[4879:4872]) ? 1 : 0;
assign detect_min[607][20] = (mid_1[4871:4864] < btm_1[4863:4856]) ? 1 : 0;
assign detect_min[607][21] = (mid_1[4871:4864] < btm_1[4871:4864]) ? 1 : 0;
assign detect_min[607][22] = (mid_1[4871:4864] < btm_1[4879:4872]) ? 1 : 0;
assign detect_min[607][23] = (mid_1[4871:4864] < btm_2[4863:4856]) ? 1 : 0;
assign detect_min[607][24] = (mid_1[4871:4864] < btm_2[4871:4864]) ? 1 : 0;
assign detect_min[607][25] = (mid_1[4871:4864] < btm_2[4879:4872]) ? 1 : 0;

assign detect_min[608][0] = (mid_1[4879:4872] < top_0[4871:4864]) ? 1 : 0;
assign detect_min[608][1] = (mid_1[4879:4872] < top_0[4879:4872]) ? 1 : 0;
assign detect_min[608][2] = (mid_1[4879:4872] < top_0[4887:4880]) ? 1 : 0;
assign detect_min[608][3] = (mid_1[4879:4872] < top_1[4871:4864]) ? 1 : 0;
assign detect_min[608][4] = (mid_1[4879:4872] < top_1[4879:4872]) ? 1 : 0;
assign detect_min[608][5] = (mid_1[4879:4872] < top_1[4887:4880]) ? 1 : 0;
assign detect_min[608][6] = (mid_1[4879:4872] < top_2[4871:4864]) ? 1 : 0;
assign detect_min[608][7] = (mid_1[4879:4872] < top_2[4879:4872]) ? 1 : 0;
assign detect_min[608][8] = (mid_1[4879:4872] < top_2[4887:4880]) ? 1 : 0;
assign detect_min[608][9] = (mid_1[4879:4872] < mid_0[4871:4864]) ? 1 : 0;
assign detect_min[608][10] = (mid_1[4879:4872] < mid_0[4879:4872]) ? 1 : 0;
assign detect_min[608][11] = (mid_1[4879:4872] < mid_0[4887:4880]) ? 1 : 0;
assign detect_min[608][12] = (mid_1[4879:4872] < mid_1[4871:4864]) ? 1 : 0;
assign detect_min[608][13] = (mid_1[4879:4872] < mid_1[4887:4880]) ? 1 : 0;
assign detect_min[608][14] = (mid_1[4879:4872] < mid_2[4871:4864]) ? 1 : 0;
assign detect_min[608][15] = (mid_1[4879:4872] < mid_2[4879:4872]) ? 1 : 0;
assign detect_min[608][16] = (mid_1[4879:4872] < mid_2[4887:4880]) ? 1 : 0;
assign detect_min[608][17] = (mid_1[4879:4872] < btm_0[4871:4864]) ? 1 : 0;
assign detect_min[608][18] = (mid_1[4879:4872] < btm_0[4879:4872]) ? 1 : 0;
assign detect_min[608][19] = (mid_1[4879:4872] < btm_0[4887:4880]) ? 1 : 0;
assign detect_min[608][20] = (mid_1[4879:4872] < btm_1[4871:4864]) ? 1 : 0;
assign detect_min[608][21] = (mid_1[4879:4872] < btm_1[4879:4872]) ? 1 : 0;
assign detect_min[608][22] = (mid_1[4879:4872] < btm_1[4887:4880]) ? 1 : 0;
assign detect_min[608][23] = (mid_1[4879:4872] < btm_2[4871:4864]) ? 1 : 0;
assign detect_min[608][24] = (mid_1[4879:4872] < btm_2[4879:4872]) ? 1 : 0;
assign detect_min[608][25] = (mid_1[4879:4872] < btm_2[4887:4880]) ? 1 : 0;

assign detect_min[609][0] = (mid_1[4887:4880] < top_0[4879:4872]) ? 1 : 0;
assign detect_min[609][1] = (mid_1[4887:4880] < top_0[4887:4880]) ? 1 : 0;
assign detect_min[609][2] = (mid_1[4887:4880] < top_0[4895:4888]) ? 1 : 0;
assign detect_min[609][3] = (mid_1[4887:4880] < top_1[4879:4872]) ? 1 : 0;
assign detect_min[609][4] = (mid_1[4887:4880] < top_1[4887:4880]) ? 1 : 0;
assign detect_min[609][5] = (mid_1[4887:4880] < top_1[4895:4888]) ? 1 : 0;
assign detect_min[609][6] = (mid_1[4887:4880] < top_2[4879:4872]) ? 1 : 0;
assign detect_min[609][7] = (mid_1[4887:4880] < top_2[4887:4880]) ? 1 : 0;
assign detect_min[609][8] = (mid_1[4887:4880] < top_2[4895:4888]) ? 1 : 0;
assign detect_min[609][9] = (mid_1[4887:4880] < mid_0[4879:4872]) ? 1 : 0;
assign detect_min[609][10] = (mid_1[4887:4880] < mid_0[4887:4880]) ? 1 : 0;
assign detect_min[609][11] = (mid_1[4887:4880] < mid_0[4895:4888]) ? 1 : 0;
assign detect_min[609][12] = (mid_1[4887:4880] < mid_1[4879:4872]) ? 1 : 0;
assign detect_min[609][13] = (mid_1[4887:4880] < mid_1[4895:4888]) ? 1 : 0;
assign detect_min[609][14] = (mid_1[4887:4880] < mid_2[4879:4872]) ? 1 : 0;
assign detect_min[609][15] = (mid_1[4887:4880] < mid_2[4887:4880]) ? 1 : 0;
assign detect_min[609][16] = (mid_1[4887:4880] < mid_2[4895:4888]) ? 1 : 0;
assign detect_min[609][17] = (mid_1[4887:4880] < btm_0[4879:4872]) ? 1 : 0;
assign detect_min[609][18] = (mid_1[4887:4880] < btm_0[4887:4880]) ? 1 : 0;
assign detect_min[609][19] = (mid_1[4887:4880] < btm_0[4895:4888]) ? 1 : 0;
assign detect_min[609][20] = (mid_1[4887:4880] < btm_1[4879:4872]) ? 1 : 0;
assign detect_min[609][21] = (mid_1[4887:4880] < btm_1[4887:4880]) ? 1 : 0;
assign detect_min[609][22] = (mid_1[4887:4880] < btm_1[4895:4888]) ? 1 : 0;
assign detect_min[609][23] = (mid_1[4887:4880] < btm_2[4879:4872]) ? 1 : 0;
assign detect_min[609][24] = (mid_1[4887:4880] < btm_2[4887:4880]) ? 1 : 0;
assign detect_min[609][25] = (mid_1[4887:4880] < btm_2[4895:4888]) ? 1 : 0;

assign detect_min[610][0] = (mid_1[4895:4888] < top_0[4887:4880]) ? 1 : 0;
assign detect_min[610][1] = (mid_1[4895:4888] < top_0[4895:4888]) ? 1 : 0;
assign detect_min[610][2] = (mid_1[4895:4888] < top_0[4903:4896]) ? 1 : 0;
assign detect_min[610][3] = (mid_1[4895:4888] < top_1[4887:4880]) ? 1 : 0;
assign detect_min[610][4] = (mid_1[4895:4888] < top_1[4895:4888]) ? 1 : 0;
assign detect_min[610][5] = (mid_1[4895:4888] < top_1[4903:4896]) ? 1 : 0;
assign detect_min[610][6] = (mid_1[4895:4888] < top_2[4887:4880]) ? 1 : 0;
assign detect_min[610][7] = (mid_1[4895:4888] < top_2[4895:4888]) ? 1 : 0;
assign detect_min[610][8] = (mid_1[4895:4888] < top_2[4903:4896]) ? 1 : 0;
assign detect_min[610][9] = (mid_1[4895:4888] < mid_0[4887:4880]) ? 1 : 0;
assign detect_min[610][10] = (mid_1[4895:4888] < mid_0[4895:4888]) ? 1 : 0;
assign detect_min[610][11] = (mid_1[4895:4888] < mid_0[4903:4896]) ? 1 : 0;
assign detect_min[610][12] = (mid_1[4895:4888] < mid_1[4887:4880]) ? 1 : 0;
assign detect_min[610][13] = (mid_1[4895:4888] < mid_1[4903:4896]) ? 1 : 0;
assign detect_min[610][14] = (mid_1[4895:4888] < mid_2[4887:4880]) ? 1 : 0;
assign detect_min[610][15] = (mid_1[4895:4888] < mid_2[4895:4888]) ? 1 : 0;
assign detect_min[610][16] = (mid_1[4895:4888] < mid_2[4903:4896]) ? 1 : 0;
assign detect_min[610][17] = (mid_1[4895:4888] < btm_0[4887:4880]) ? 1 : 0;
assign detect_min[610][18] = (mid_1[4895:4888] < btm_0[4895:4888]) ? 1 : 0;
assign detect_min[610][19] = (mid_1[4895:4888] < btm_0[4903:4896]) ? 1 : 0;
assign detect_min[610][20] = (mid_1[4895:4888] < btm_1[4887:4880]) ? 1 : 0;
assign detect_min[610][21] = (mid_1[4895:4888] < btm_1[4895:4888]) ? 1 : 0;
assign detect_min[610][22] = (mid_1[4895:4888] < btm_1[4903:4896]) ? 1 : 0;
assign detect_min[610][23] = (mid_1[4895:4888] < btm_2[4887:4880]) ? 1 : 0;
assign detect_min[610][24] = (mid_1[4895:4888] < btm_2[4895:4888]) ? 1 : 0;
assign detect_min[610][25] = (mid_1[4895:4888] < btm_2[4903:4896]) ? 1 : 0;

assign detect_min[611][0] = (mid_1[4903:4896] < top_0[4895:4888]) ? 1 : 0;
assign detect_min[611][1] = (mid_1[4903:4896] < top_0[4903:4896]) ? 1 : 0;
assign detect_min[611][2] = (mid_1[4903:4896] < top_0[4911:4904]) ? 1 : 0;
assign detect_min[611][3] = (mid_1[4903:4896] < top_1[4895:4888]) ? 1 : 0;
assign detect_min[611][4] = (mid_1[4903:4896] < top_1[4903:4896]) ? 1 : 0;
assign detect_min[611][5] = (mid_1[4903:4896] < top_1[4911:4904]) ? 1 : 0;
assign detect_min[611][6] = (mid_1[4903:4896] < top_2[4895:4888]) ? 1 : 0;
assign detect_min[611][7] = (mid_1[4903:4896] < top_2[4903:4896]) ? 1 : 0;
assign detect_min[611][8] = (mid_1[4903:4896] < top_2[4911:4904]) ? 1 : 0;
assign detect_min[611][9] = (mid_1[4903:4896] < mid_0[4895:4888]) ? 1 : 0;
assign detect_min[611][10] = (mid_1[4903:4896] < mid_0[4903:4896]) ? 1 : 0;
assign detect_min[611][11] = (mid_1[4903:4896] < mid_0[4911:4904]) ? 1 : 0;
assign detect_min[611][12] = (mid_1[4903:4896] < mid_1[4895:4888]) ? 1 : 0;
assign detect_min[611][13] = (mid_1[4903:4896] < mid_1[4911:4904]) ? 1 : 0;
assign detect_min[611][14] = (mid_1[4903:4896] < mid_2[4895:4888]) ? 1 : 0;
assign detect_min[611][15] = (mid_1[4903:4896] < mid_2[4903:4896]) ? 1 : 0;
assign detect_min[611][16] = (mid_1[4903:4896] < mid_2[4911:4904]) ? 1 : 0;
assign detect_min[611][17] = (mid_1[4903:4896] < btm_0[4895:4888]) ? 1 : 0;
assign detect_min[611][18] = (mid_1[4903:4896] < btm_0[4903:4896]) ? 1 : 0;
assign detect_min[611][19] = (mid_1[4903:4896] < btm_0[4911:4904]) ? 1 : 0;
assign detect_min[611][20] = (mid_1[4903:4896] < btm_1[4895:4888]) ? 1 : 0;
assign detect_min[611][21] = (mid_1[4903:4896] < btm_1[4903:4896]) ? 1 : 0;
assign detect_min[611][22] = (mid_1[4903:4896] < btm_1[4911:4904]) ? 1 : 0;
assign detect_min[611][23] = (mid_1[4903:4896] < btm_2[4895:4888]) ? 1 : 0;
assign detect_min[611][24] = (mid_1[4903:4896] < btm_2[4903:4896]) ? 1 : 0;
assign detect_min[611][25] = (mid_1[4903:4896] < btm_2[4911:4904]) ? 1 : 0;

assign detect_min[612][0] = (mid_1[4911:4904] < top_0[4903:4896]) ? 1 : 0;
assign detect_min[612][1] = (mid_1[4911:4904] < top_0[4911:4904]) ? 1 : 0;
assign detect_min[612][2] = (mid_1[4911:4904] < top_0[4919:4912]) ? 1 : 0;
assign detect_min[612][3] = (mid_1[4911:4904] < top_1[4903:4896]) ? 1 : 0;
assign detect_min[612][4] = (mid_1[4911:4904] < top_1[4911:4904]) ? 1 : 0;
assign detect_min[612][5] = (mid_1[4911:4904] < top_1[4919:4912]) ? 1 : 0;
assign detect_min[612][6] = (mid_1[4911:4904] < top_2[4903:4896]) ? 1 : 0;
assign detect_min[612][7] = (mid_1[4911:4904] < top_2[4911:4904]) ? 1 : 0;
assign detect_min[612][8] = (mid_1[4911:4904] < top_2[4919:4912]) ? 1 : 0;
assign detect_min[612][9] = (mid_1[4911:4904] < mid_0[4903:4896]) ? 1 : 0;
assign detect_min[612][10] = (mid_1[4911:4904] < mid_0[4911:4904]) ? 1 : 0;
assign detect_min[612][11] = (mid_1[4911:4904] < mid_0[4919:4912]) ? 1 : 0;
assign detect_min[612][12] = (mid_1[4911:4904] < mid_1[4903:4896]) ? 1 : 0;
assign detect_min[612][13] = (mid_1[4911:4904] < mid_1[4919:4912]) ? 1 : 0;
assign detect_min[612][14] = (mid_1[4911:4904] < mid_2[4903:4896]) ? 1 : 0;
assign detect_min[612][15] = (mid_1[4911:4904] < mid_2[4911:4904]) ? 1 : 0;
assign detect_min[612][16] = (mid_1[4911:4904] < mid_2[4919:4912]) ? 1 : 0;
assign detect_min[612][17] = (mid_1[4911:4904] < btm_0[4903:4896]) ? 1 : 0;
assign detect_min[612][18] = (mid_1[4911:4904] < btm_0[4911:4904]) ? 1 : 0;
assign detect_min[612][19] = (mid_1[4911:4904] < btm_0[4919:4912]) ? 1 : 0;
assign detect_min[612][20] = (mid_1[4911:4904] < btm_1[4903:4896]) ? 1 : 0;
assign detect_min[612][21] = (mid_1[4911:4904] < btm_1[4911:4904]) ? 1 : 0;
assign detect_min[612][22] = (mid_1[4911:4904] < btm_1[4919:4912]) ? 1 : 0;
assign detect_min[612][23] = (mid_1[4911:4904] < btm_2[4903:4896]) ? 1 : 0;
assign detect_min[612][24] = (mid_1[4911:4904] < btm_2[4911:4904]) ? 1 : 0;
assign detect_min[612][25] = (mid_1[4911:4904] < btm_2[4919:4912]) ? 1 : 0;

assign detect_min[613][0] = (mid_1[4919:4912] < top_0[4911:4904]) ? 1 : 0;
assign detect_min[613][1] = (mid_1[4919:4912] < top_0[4919:4912]) ? 1 : 0;
assign detect_min[613][2] = (mid_1[4919:4912] < top_0[4927:4920]) ? 1 : 0;
assign detect_min[613][3] = (mid_1[4919:4912] < top_1[4911:4904]) ? 1 : 0;
assign detect_min[613][4] = (mid_1[4919:4912] < top_1[4919:4912]) ? 1 : 0;
assign detect_min[613][5] = (mid_1[4919:4912] < top_1[4927:4920]) ? 1 : 0;
assign detect_min[613][6] = (mid_1[4919:4912] < top_2[4911:4904]) ? 1 : 0;
assign detect_min[613][7] = (mid_1[4919:4912] < top_2[4919:4912]) ? 1 : 0;
assign detect_min[613][8] = (mid_1[4919:4912] < top_2[4927:4920]) ? 1 : 0;
assign detect_min[613][9] = (mid_1[4919:4912] < mid_0[4911:4904]) ? 1 : 0;
assign detect_min[613][10] = (mid_1[4919:4912] < mid_0[4919:4912]) ? 1 : 0;
assign detect_min[613][11] = (mid_1[4919:4912] < mid_0[4927:4920]) ? 1 : 0;
assign detect_min[613][12] = (mid_1[4919:4912] < mid_1[4911:4904]) ? 1 : 0;
assign detect_min[613][13] = (mid_1[4919:4912] < mid_1[4927:4920]) ? 1 : 0;
assign detect_min[613][14] = (mid_1[4919:4912] < mid_2[4911:4904]) ? 1 : 0;
assign detect_min[613][15] = (mid_1[4919:4912] < mid_2[4919:4912]) ? 1 : 0;
assign detect_min[613][16] = (mid_1[4919:4912] < mid_2[4927:4920]) ? 1 : 0;
assign detect_min[613][17] = (mid_1[4919:4912] < btm_0[4911:4904]) ? 1 : 0;
assign detect_min[613][18] = (mid_1[4919:4912] < btm_0[4919:4912]) ? 1 : 0;
assign detect_min[613][19] = (mid_1[4919:4912] < btm_0[4927:4920]) ? 1 : 0;
assign detect_min[613][20] = (mid_1[4919:4912] < btm_1[4911:4904]) ? 1 : 0;
assign detect_min[613][21] = (mid_1[4919:4912] < btm_1[4919:4912]) ? 1 : 0;
assign detect_min[613][22] = (mid_1[4919:4912] < btm_1[4927:4920]) ? 1 : 0;
assign detect_min[613][23] = (mid_1[4919:4912] < btm_2[4911:4904]) ? 1 : 0;
assign detect_min[613][24] = (mid_1[4919:4912] < btm_2[4919:4912]) ? 1 : 0;
assign detect_min[613][25] = (mid_1[4919:4912] < btm_2[4927:4920]) ? 1 : 0;

assign detect_min[614][0] = (mid_1[4927:4920] < top_0[4919:4912]) ? 1 : 0;
assign detect_min[614][1] = (mid_1[4927:4920] < top_0[4927:4920]) ? 1 : 0;
assign detect_min[614][2] = (mid_1[4927:4920] < top_0[4935:4928]) ? 1 : 0;
assign detect_min[614][3] = (mid_1[4927:4920] < top_1[4919:4912]) ? 1 : 0;
assign detect_min[614][4] = (mid_1[4927:4920] < top_1[4927:4920]) ? 1 : 0;
assign detect_min[614][5] = (mid_1[4927:4920] < top_1[4935:4928]) ? 1 : 0;
assign detect_min[614][6] = (mid_1[4927:4920] < top_2[4919:4912]) ? 1 : 0;
assign detect_min[614][7] = (mid_1[4927:4920] < top_2[4927:4920]) ? 1 : 0;
assign detect_min[614][8] = (mid_1[4927:4920] < top_2[4935:4928]) ? 1 : 0;
assign detect_min[614][9] = (mid_1[4927:4920] < mid_0[4919:4912]) ? 1 : 0;
assign detect_min[614][10] = (mid_1[4927:4920] < mid_0[4927:4920]) ? 1 : 0;
assign detect_min[614][11] = (mid_1[4927:4920] < mid_0[4935:4928]) ? 1 : 0;
assign detect_min[614][12] = (mid_1[4927:4920] < mid_1[4919:4912]) ? 1 : 0;
assign detect_min[614][13] = (mid_1[4927:4920] < mid_1[4935:4928]) ? 1 : 0;
assign detect_min[614][14] = (mid_1[4927:4920] < mid_2[4919:4912]) ? 1 : 0;
assign detect_min[614][15] = (mid_1[4927:4920] < mid_2[4927:4920]) ? 1 : 0;
assign detect_min[614][16] = (mid_1[4927:4920] < mid_2[4935:4928]) ? 1 : 0;
assign detect_min[614][17] = (mid_1[4927:4920] < btm_0[4919:4912]) ? 1 : 0;
assign detect_min[614][18] = (mid_1[4927:4920] < btm_0[4927:4920]) ? 1 : 0;
assign detect_min[614][19] = (mid_1[4927:4920] < btm_0[4935:4928]) ? 1 : 0;
assign detect_min[614][20] = (mid_1[4927:4920] < btm_1[4919:4912]) ? 1 : 0;
assign detect_min[614][21] = (mid_1[4927:4920] < btm_1[4927:4920]) ? 1 : 0;
assign detect_min[614][22] = (mid_1[4927:4920] < btm_1[4935:4928]) ? 1 : 0;
assign detect_min[614][23] = (mid_1[4927:4920] < btm_2[4919:4912]) ? 1 : 0;
assign detect_min[614][24] = (mid_1[4927:4920] < btm_2[4927:4920]) ? 1 : 0;
assign detect_min[614][25] = (mid_1[4927:4920] < btm_2[4935:4928]) ? 1 : 0;

assign detect_min[615][0] = (mid_1[4935:4928] < top_0[4927:4920]) ? 1 : 0;
assign detect_min[615][1] = (mid_1[4935:4928] < top_0[4935:4928]) ? 1 : 0;
assign detect_min[615][2] = (mid_1[4935:4928] < top_0[4943:4936]) ? 1 : 0;
assign detect_min[615][3] = (mid_1[4935:4928] < top_1[4927:4920]) ? 1 : 0;
assign detect_min[615][4] = (mid_1[4935:4928] < top_1[4935:4928]) ? 1 : 0;
assign detect_min[615][5] = (mid_1[4935:4928] < top_1[4943:4936]) ? 1 : 0;
assign detect_min[615][6] = (mid_1[4935:4928] < top_2[4927:4920]) ? 1 : 0;
assign detect_min[615][7] = (mid_1[4935:4928] < top_2[4935:4928]) ? 1 : 0;
assign detect_min[615][8] = (mid_1[4935:4928] < top_2[4943:4936]) ? 1 : 0;
assign detect_min[615][9] = (mid_1[4935:4928] < mid_0[4927:4920]) ? 1 : 0;
assign detect_min[615][10] = (mid_1[4935:4928] < mid_0[4935:4928]) ? 1 : 0;
assign detect_min[615][11] = (mid_1[4935:4928] < mid_0[4943:4936]) ? 1 : 0;
assign detect_min[615][12] = (mid_1[4935:4928] < mid_1[4927:4920]) ? 1 : 0;
assign detect_min[615][13] = (mid_1[4935:4928] < mid_1[4943:4936]) ? 1 : 0;
assign detect_min[615][14] = (mid_1[4935:4928] < mid_2[4927:4920]) ? 1 : 0;
assign detect_min[615][15] = (mid_1[4935:4928] < mid_2[4935:4928]) ? 1 : 0;
assign detect_min[615][16] = (mid_1[4935:4928] < mid_2[4943:4936]) ? 1 : 0;
assign detect_min[615][17] = (mid_1[4935:4928] < btm_0[4927:4920]) ? 1 : 0;
assign detect_min[615][18] = (mid_1[4935:4928] < btm_0[4935:4928]) ? 1 : 0;
assign detect_min[615][19] = (mid_1[4935:4928] < btm_0[4943:4936]) ? 1 : 0;
assign detect_min[615][20] = (mid_1[4935:4928] < btm_1[4927:4920]) ? 1 : 0;
assign detect_min[615][21] = (mid_1[4935:4928] < btm_1[4935:4928]) ? 1 : 0;
assign detect_min[615][22] = (mid_1[4935:4928] < btm_1[4943:4936]) ? 1 : 0;
assign detect_min[615][23] = (mid_1[4935:4928] < btm_2[4927:4920]) ? 1 : 0;
assign detect_min[615][24] = (mid_1[4935:4928] < btm_2[4935:4928]) ? 1 : 0;
assign detect_min[615][25] = (mid_1[4935:4928] < btm_2[4943:4936]) ? 1 : 0;

assign detect_min[616][0] = (mid_1[4943:4936] < top_0[4935:4928]) ? 1 : 0;
assign detect_min[616][1] = (mid_1[4943:4936] < top_0[4943:4936]) ? 1 : 0;
assign detect_min[616][2] = (mid_1[4943:4936] < top_0[4951:4944]) ? 1 : 0;
assign detect_min[616][3] = (mid_1[4943:4936] < top_1[4935:4928]) ? 1 : 0;
assign detect_min[616][4] = (mid_1[4943:4936] < top_1[4943:4936]) ? 1 : 0;
assign detect_min[616][5] = (mid_1[4943:4936] < top_1[4951:4944]) ? 1 : 0;
assign detect_min[616][6] = (mid_1[4943:4936] < top_2[4935:4928]) ? 1 : 0;
assign detect_min[616][7] = (mid_1[4943:4936] < top_2[4943:4936]) ? 1 : 0;
assign detect_min[616][8] = (mid_1[4943:4936] < top_2[4951:4944]) ? 1 : 0;
assign detect_min[616][9] = (mid_1[4943:4936] < mid_0[4935:4928]) ? 1 : 0;
assign detect_min[616][10] = (mid_1[4943:4936] < mid_0[4943:4936]) ? 1 : 0;
assign detect_min[616][11] = (mid_1[4943:4936] < mid_0[4951:4944]) ? 1 : 0;
assign detect_min[616][12] = (mid_1[4943:4936] < mid_1[4935:4928]) ? 1 : 0;
assign detect_min[616][13] = (mid_1[4943:4936] < mid_1[4951:4944]) ? 1 : 0;
assign detect_min[616][14] = (mid_1[4943:4936] < mid_2[4935:4928]) ? 1 : 0;
assign detect_min[616][15] = (mid_1[4943:4936] < mid_2[4943:4936]) ? 1 : 0;
assign detect_min[616][16] = (mid_1[4943:4936] < mid_2[4951:4944]) ? 1 : 0;
assign detect_min[616][17] = (mid_1[4943:4936] < btm_0[4935:4928]) ? 1 : 0;
assign detect_min[616][18] = (mid_1[4943:4936] < btm_0[4943:4936]) ? 1 : 0;
assign detect_min[616][19] = (mid_1[4943:4936] < btm_0[4951:4944]) ? 1 : 0;
assign detect_min[616][20] = (mid_1[4943:4936] < btm_1[4935:4928]) ? 1 : 0;
assign detect_min[616][21] = (mid_1[4943:4936] < btm_1[4943:4936]) ? 1 : 0;
assign detect_min[616][22] = (mid_1[4943:4936] < btm_1[4951:4944]) ? 1 : 0;
assign detect_min[616][23] = (mid_1[4943:4936] < btm_2[4935:4928]) ? 1 : 0;
assign detect_min[616][24] = (mid_1[4943:4936] < btm_2[4943:4936]) ? 1 : 0;
assign detect_min[616][25] = (mid_1[4943:4936] < btm_2[4951:4944]) ? 1 : 0;

assign detect_min[617][0] = (mid_1[4951:4944] < top_0[4943:4936]) ? 1 : 0;
assign detect_min[617][1] = (mid_1[4951:4944] < top_0[4951:4944]) ? 1 : 0;
assign detect_min[617][2] = (mid_1[4951:4944] < top_0[4959:4952]) ? 1 : 0;
assign detect_min[617][3] = (mid_1[4951:4944] < top_1[4943:4936]) ? 1 : 0;
assign detect_min[617][4] = (mid_1[4951:4944] < top_1[4951:4944]) ? 1 : 0;
assign detect_min[617][5] = (mid_1[4951:4944] < top_1[4959:4952]) ? 1 : 0;
assign detect_min[617][6] = (mid_1[4951:4944] < top_2[4943:4936]) ? 1 : 0;
assign detect_min[617][7] = (mid_1[4951:4944] < top_2[4951:4944]) ? 1 : 0;
assign detect_min[617][8] = (mid_1[4951:4944] < top_2[4959:4952]) ? 1 : 0;
assign detect_min[617][9] = (mid_1[4951:4944] < mid_0[4943:4936]) ? 1 : 0;
assign detect_min[617][10] = (mid_1[4951:4944] < mid_0[4951:4944]) ? 1 : 0;
assign detect_min[617][11] = (mid_1[4951:4944] < mid_0[4959:4952]) ? 1 : 0;
assign detect_min[617][12] = (mid_1[4951:4944] < mid_1[4943:4936]) ? 1 : 0;
assign detect_min[617][13] = (mid_1[4951:4944] < mid_1[4959:4952]) ? 1 : 0;
assign detect_min[617][14] = (mid_1[4951:4944] < mid_2[4943:4936]) ? 1 : 0;
assign detect_min[617][15] = (mid_1[4951:4944] < mid_2[4951:4944]) ? 1 : 0;
assign detect_min[617][16] = (mid_1[4951:4944] < mid_2[4959:4952]) ? 1 : 0;
assign detect_min[617][17] = (mid_1[4951:4944] < btm_0[4943:4936]) ? 1 : 0;
assign detect_min[617][18] = (mid_1[4951:4944] < btm_0[4951:4944]) ? 1 : 0;
assign detect_min[617][19] = (mid_1[4951:4944] < btm_0[4959:4952]) ? 1 : 0;
assign detect_min[617][20] = (mid_1[4951:4944] < btm_1[4943:4936]) ? 1 : 0;
assign detect_min[617][21] = (mid_1[4951:4944] < btm_1[4951:4944]) ? 1 : 0;
assign detect_min[617][22] = (mid_1[4951:4944] < btm_1[4959:4952]) ? 1 : 0;
assign detect_min[617][23] = (mid_1[4951:4944] < btm_2[4943:4936]) ? 1 : 0;
assign detect_min[617][24] = (mid_1[4951:4944] < btm_2[4951:4944]) ? 1 : 0;
assign detect_min[617][25] = (mid_1[4951:4944] < btm_2[4959:4952]) ? 1 : 0;

assign detect_min[618][0] = (mid_1[4959:4952] < top_0[4951:4944]) ? 1 : 0;
assign detect_min[618][1] = (mid_1[4959:4952] < top_0[4959:4952]) ? 1 : 0;
assign detect_min[618][2] = (mid_1[4959:4952] < top_0[4967:4960]) ? 1 : 0;
assign detect_min[618][3] = (mid_1[4959:4952] < top_1[4951:4944]) ? 1 : 0;
assign detect_min[618][4] = (mid_1[4959:4952] < top_1[4959:4952]) ? 1 : 0;
assign detect_min[618][5] = (mid_1[4959:4952] < top_1[4967:4960]) ? 1 : 0;
assign detect_min[618][6] = (mid_1[4959:4952] < top_2[4951:4944]) ? 1 : 0;
assign detect_min[618][7] = (mid_1[4959:4952] < top_2[4959:4952]) ? 1 : 0;
assign detect_min[618][8] = (mid_1[4959:4952] < top_2[4967:4960]) ? 1 : 0;
assign detect_min[618][9] = (mid_1[4959:4952] < mid_0[4951:4944]) ? 1 : 0;
assign detect_min[618][10] = (mid_1[4959:4952] < mid_0[4959:4952]) ? 1 : 0;
assign detect_min[618][11] = (mid_1[4959:4952] < mid_0[4967:4960]) ? 1 : 0;
assign detect_min[618][12] = (mid_1[4959:4952] < mid_1[4951:4944]) ? 1 : 0;
assign detect_min[618][13] = (mid_1[4959:4952] < mid_1[4967:4960]) ? 1 : 0;
assign detect_min[618][14] = (mid_1[4959:4952] < mid_2[4951:4944]) ? 1 : 0;
assign detect_min[618][15] = (mid_1[4959:4952] < mid_2[4959:4952]) ? 1 : 0;
assign detect_min[618][16] = (mid_1[4959:4952] < mid_2[4967:4960]) ? 1 : 0;
assign detect_min[618][17] = (mid_1[4959:4952] < btm_0[4951:4944]) ? 1 : 0;
assign detect_min[618][18] = (mid_1[4959:4952] < btm_0[4959:4952]) ? 1 : 0;
assign detect_min[618][19] = (mid_1[4959:4952] < btm_0[4967:4960]) ? 1 : 0;
assign detect_min[618][20] = (mid_1[4959:4952] < btm_1[4951:4944]) ? 1 : 0;
assign detect_min[618][21] = (mid_1[4959:4952] < btm_1[4959:4952]) ? 1 : 0;
assign detect_min[618][22] = (mid_1[4959:4952] < btm_1[4967:4960]) ? 1 : 0;
assign detect_min[618][23] = (mid_1[4959:4952] < btm_2[4951:4944]) ? 1 : 0;
assign detect_min[618][24] = (mid_1[4959:4952] < btm_2[4959:4952]) ? 1 : 0;
assign detect_min[618][25] = (mid_1[4959:4952] < btm_2[4967:4960]) ? 1 : 0;

assign detect_min[619][0] = (mid_1[4967:4960] < top_0[4959:4952]) ? 1 : 0;
assign detect_min[619][1] = (mid_1[4967:4960] < top_0[4967:4960]) ? 1 : 0;
assign detect_min[619][2] = (mid_1[4967:4960] < top_0[4975:4968]) ? 1 : 0;
assign detect_min[619][3] = (mid_1[4967:4960] < top_1[4959:4952]) ? 1 : 0;
assign detect_min[619][4] = (mid_1[4967:4960] < top_1[4967:4960]) ? 1 : 0;
assign detect_min[619][5] = (mid_1[4967:4960] < top_1[4975:4968]) ? 1 : 0;
assign detect_min[619][6] = (mid_1[4967:4960] < top_2[4959:4952]) ? 1 : 0;
assign detect_min[619][7] = (mid_1[4967:4960] < top_2[4967:4960]) ? 1 : 0;
assign detect_min[619][8] = (mid_1[4967:4960] < top_2[4975:4968]) ? 1 : 0;
assign detect_min[619][9] = (mid_1[4967:4960] < mid_0[4959:4952]) ? 1 : 0;
assign detect_min[619][10] = (mid_1[4967:4960] < mid_0[4967:4960]) ? 1 : 0;
assign detect_min[619][11] = (mid_1[4967:4960] < mid_0[4975:4968]) ? 1 : 0;
assign detect_min[619][12] = (mid_1[4967:4960] < mid_1[4959:4952]) ? 1 : 0;
assign detect_min[619][13] = (mid_1[4967:4960] < mid_1[4975:4968]) ? 1 : 0;
assign detect_min[619][14] = (mid_1[4967:4960] < mid_2[4959:4952]) ? 1 : 0;
assign detect_min[619][15] = (mid_1[4967:4960] < mid_2[4967:4960]) ? 1 : 0;
assign detect_min[619][16] = (mid_1[4967:4960] < mid_2[4975:4968]) ? 1 : 0;
assign detect_min[619][17] = (mid_1[4967:4960] < btm_0[4959:4952]) ? 1 : 0;
assign detect_min[619][18] = (mid_1[4967:4960] < btm_0[4967:4960]) ? 1 : 0;
assign detect_min[619][19] = (mid_1[4967:4960] < btm_0[4975:4968]) ? 1 : 0;
assign detect_min[619][20] = (mid_1[4967:4960] < btm_1[4959:4952]) ? 1 : 0;
assign detect_min[619][21] = (mid_1[4967:4960] < btm_1[4967:4960]) ? 1 : 0;
assign detect_min[619][22] = (mid_1[4967:4960] < btm_1[4975:4968]) ? 1 : 0;
assign detect_min[619][23] = (mid_1[4967:4960] < btm_2[4959:4952]) ? 1 : 0;
assign detect_min[619][24] = (mid_1[4967:4960] < btm_2[4967:4960]) ? 1 : 0;
assign detect_min[619][25] = (mid_1[4967:4960] < btm_2[4975:4968]) ? 1 : 0;

assign detect_min[620][0] = (mid_1[4975:4968] < top_0[4967:4960]) ? 1 : 0;
assign detect_min[620][1] = (mid_1[4975:4968] < top_0[4975:4968]) ? 1 : 0;
assign detect_min[620][2] = (mid_1[4975:4968] < top_0[4983:4976]) ? 1 : 0;
assign detect_min[620][3] = (mid_1[4975:4968] < top_1[4967:4960]) ? 1 : 0;
assign detect_min[620][4] = (mid_1[4975:4968] < top_1[4975:4968]) ? 1 : 0;
assign detect_min[620][5] = (mid_1[4975:4968] < top_1[4983:4976]) ? 1 : 0;
assign detect_min[620][6] = (mid_1[4975:4968] < top_2[4967:4960]) ? 1 : 0;
assign detect_min[620][7] = (mid_1[4975:4968] < top_2[4975:4968]) ? 1 : 0;
assign detect_min[620][8] = (mid_1[4975:4968] < top_2[4983:4976]) ? 1 : 0;
assign detect_min[620][9] = (mid_1[4975:4968] < mid_0[4967:4960]) ? 1 : 0;
assign detect_min[620][10] = (mid_1[4975:4968] < mid_0[4975:4968]) ? 1 : 0;
assign detect_min[620][11] = (mid_1[4975:4968] < mid_0[4983:4976]) ? 1 : 0;
assign detect_min[620][12] = (mid_1[4975:4968] < mid_1[4967:4960]) ? 1 : 0;
assign detect_min[620][13] = (mid_1[4975:4968] < mid_1[4983:4976]) ? 1 : 0;
assign detect_min[620][14] = (mid_1[4975:4968] < mid_2[4967:4960]) ? 1 : 0;
assign detect_min[620][15] = (mid_1[4975:4968] < mid_2[4975:4968]) ? 1 : 0;
assign detect_min[620][16] = (mid_1[4975:4968] < mid_2[4983:4976]) ? 1 : 0;
assign detect_min[620][17] = (mid_1[4975:4968] < btm_0[4967:4960]) ? 1 : 0;
assign detect_min[620][18] = (mid_1[4975:4968] < btm_0[4975:4968]) ? 1 : 0;
assign detect_min[620][19] = (mid_1[4975:4968] < btm_0[4983:4976]) ? 1 : 0;
assign detect_min[620][20] = (mid_1[4975:4968] < btm_1[4967:4960]) ? 1 : 0;
assign detect_min[620][21] = (mid_1[4975:4968] < btm_1[4975:4968]) ? 1 : 0;
assign detect_min[620][22] = (mid_1[4975:4968] < btm_1[4983:4976]) ? 1 : 0;
assign detect_min[620][23] = (mid_1[4975:4968] < btm_2[4967:4960]) ? 1 : 0;
assign detect_min[620][24] = (mid_1[4975:4968] < btm_2[4975:4968]) ? 1 : 0;
assign detect_min[620][25] = (mid_1[4975:4968] < btm_2[4983:4976]) ? 1 : 0;

assign detect_min[621][0] = (mid_1[4983:4976] < top_0[4975:4968]) ? 1 : 0;
assign detect_min[621][1] = (mid_1[4983:4976] < top_0[4983:4976]) ? 1 : 0;
assign detect_min[621][2] = (mid_1[4983:4976] < top_0[4991:4984]) ? 1 : 0;
assign detect_min[621][3] = (mid_1[4983:4976] < top_1[4975:4968]) ? 1 : 0;
assign detect_min[621][4] = (mid_1[4983:4976] < top_1[4983:4976]) ? 1 : 0;
assign detect_min[621][5] = (mid_1[4983:4976] < top_1[4991:4984]) ? 1 : 0;
assign detect_min[621][6] = (mid_1[4983:4976] < top_2[4975:4968]) ? 1 : 0;
assign detect_min[621][7] = (mid_1[4983:4976] < top_2[4983:4976]) ? 1 : 0;
assign detect_min[621][8] = (mid_1[4983:4976] < top_2[4991:4984]) ? 1 : 0;
assign detect_min[621][9] = (mid_1[4983:4976] < mid_0[4975:4968]) ? 1 : 0;
assign detect_min[621][10] = (mid_1[4983:4976] < mid_0[4983:4976]) ? 1 : 0;
assign detect_min[621][11] = (mid_1[4983:4976] < mid_0[4991:4984]) ? 1 : 0;
assign detect_min[621][12] = (mid_1[4983:4976] < mid_1[4975:4968]) ? 1 : 0;
assign detect_min[621][13] = (mid_1[4983:4976] < mid_1[4991:4984]) ? 1 : 0;
assign detect_min[621][14] = (mid_1[4983:4976] < mid_2[4975:4968]) ? 1 : 0;
assign detect_min[621][15] = (mid_1[4983:4976] < mid_2[4983:4976]) ? 1 : 0;
assign detect_min[621][16] = (mid_1[4983:4976] < mid_2[4991:4984]) ? 1 : 0;
assign detect_min[621][17] = (mid_1[4983:4976] < btm_0[4975:4968]) ? 1 : 0;
assign detect_min[621][18] = (mid_1[4983:4976] < btm_0[4983:4976]) ? 1 : 0;
assign detect_min[621][19] = (mid_1[4983:4976] < btm_0[4991:4984]) ? 1 : 0;
assign detect_min[621][20] = (mid_1[4983:4976] < btm_1[4975:4968]) ? 1 : 0;
assign detect_min[621][21] = (mid_1[4983:4976] < btm_1[4983:4976]) ? 1 : 0;
assign detect_min[621][22] = (mid_1[4983:4976] < btm_1[4991:4984]) ? 1 : 0;
assign detect_min[621][23] = (mid_1[4983:4976] < btm_2[4975:4968]) ? 1 : 0;
assign detect_min[621][24] = (mid_1[4983:4976] < btm_2[4983:4976]) ? 1 : 0;
assign detect_min[621][25] = (mid_1[4983:4976] < btm_2[4991:4984]) ? 1 : 0;

assign detect_min[622][0] = (mid_1[4991:4984] < top_0[4983:4976]) ? 1 : 0;
assign detect_min[622][1] = (mid_1[4991:4984] < top_0[4991:4984]) ? 1 : 0;
assign detect_min[622][2] = (mid_1[4991:4984] < top_0[4999:4992]) ? 1 : 0;
assign detect_min[622][3] = (mid_1[4991:4984] < top_1[4983:4976]) ? 1 : 0;
assign detect_min[622][4] = (mid_1[4991:4984] < top_1[4991:4984]) ? 1 : 0;
assign detect_min[622][5] = (mid_1[4991:4984] < top_1[4999:4992]) ? 1 : 0;
assign detect_min[622][6] = (mid_1[4991:4984] < top_2[4983:4976]) ? 1 : 0;
assign detect_min[622][7] = (mid_1[4991:4984] < top_2[4991:4984]) ? 1 : 0;
assign detect_min[622][8] = (mid_1[4991:4984] < top_2[4999:4992]) ? 1 : 0;
assign detect_min[622][9] = (mid_1[4991:4984] < mid_0[4983:4976]) ? 1 : 0;
assign detect_min[622][10] = (mid_1[4991:4984] < mid_0[4991:4984]) ? 1 : 0;
assign detect_min[622][11] = (mid_1[4991:4984] < mid_0[4999:4992]) ? 1 : 0;
assign detect_min[622][12] = (mid_1[4991:4984] < mid_1[4983:4976]) ? 1 : 0;
assign detect_min[622][13] = (mid_1[4991:4984] < mid_1[4999:4992]) ? 1 : 0;
assign detect_min[622][14] = (mid_1[4991:4984] < mid_2[4983:4976]) ? 1 : 0;
assign detect_min[622][15] = (mid_1[4991:4984] < mid_2[4991:4984]) ? 1 : 0;
assign detect_min[622][16] = (mid_1[4991:4984] < mid_2[4999:4992]) ? 1 : 0;
assign detect_min[622][17] = (mid_1[4991:4984] < btm_0[4983:4976]) ? 1 : 0;
assign detect_min[622][18] = (mid_1[4991:4984] < btm_0[4991:4984]) ? 1 : 0;
assign detect_min[622][19] = (mid_1[4991:4984] < btm_0[4999:4992]) ? 1 : 0;
assign detect_min[622][20] = (mid_1[4991:4984] < btm_1[4983:4976]) ? 1 : 0;
assign detect_min[622][21] = (mid_1[4991:4984] < btm_1[4991:4984]) ? 1 : 0;
assign detect_min[622][22] = (mid_1[4991:4984] < btm_1[4999:4992]) ? 1 : 0;
assign detect_min[622][23] = (mid_1[4991:4984] < btm_2[4983:4976]) ? 1 : 0;
assign detect_min[622][24] = (mid_1[4991:4984] < btm_2[4991:4984]) ? 1 : 0;
assign detect_min[622][25] = (mid_1[4991:4984] < btm_2[4999:4992]) ? 1 : 0;

assign detect_min[623][0] = (mid_1[4999:4992] < top_0[4991:4984]) ? 1 : 0;
assign detect_min[623][1] = (mid_1[4999:4992] < top_0[4999:4992]) ? 1 : 0;
assign detect_min[623][2] = (mid_1[4999:4992] < top_0[5007:5000]) ? 1 : 0;
assign detect_min[623][3] = (mid_1[4999:4992] < top_1[4991:4984]) ? 1 : 0;
assign detect_min[623][4] = (mid_1[4999:4992] < top_1[4999:4992]) ? 1 : 0;
assign detect_min[623][5] = (mid_1[4999:4992] < top_1[5007:5000]) ? 1 : 0;
assign detect_min[623][6] = (mid_1[4999:4992] < top_2[4991:4984]) ? 1 : 0;
assign detect_min[623][7] = (mid_1[4999:4992] < top_2[4999:4992]) ? 1 : 0;
assign detect_min[623][8] = (mid_1[4999:4992] < top_2[5007:5000]) ? 1 : 0;
assign detect_min[623][9] = (mid_1[4999:4992] < mid_0[4991:4984]) ? 1 : 0;
assign detect_min[623][10] = (mid_1[4999:4992] < mid_0[4999:4992]) ? 1 : 0;
assign detect_min[623][11] = (mid_1[4999:4992] < mid_0[5007:5000]) ? 1 : 0;
assign detect_min[623][12] = (mid_1[4999:4992] < mid_1[4991:4984]) ? 1 : 0;
assign detect_min[623][13] = (mid_1[4999:4992] < mid_1[5007:5000]) ? 1 : 0;
assign detect_min[623][14] = (mid_1[4999:4992] < mid_2[4991:4984]) ? 1 : 0;
assign detect_min[623][15] = (mid_1[4999:4992] < mid_2[4999:4992]) ? 1 : 0;
assign detect_min[623][16] = (mid_1[4999:4992] < mid_2[5007:5000]) ? 1 : 0;
assign detect_min[623][17] = (mid_1[4999:4992] < btm_0[4991:4984]) ? 1 : 0;
assign detect_min[623][18] = (mid_1[4999:4992] < btm_0[4999:4992]) ? 1 : 0;
assign detect_min[623][19] = (mid_1[4999:4992] < btm_0[5007:5000]) ? 1 : 0;
assign detect_min[623][20] = (mid_1[4999:4992] < btm_1[4991:4984]) ? 1 : 0;
assign detect_min[623][21] = (mid_1[4999:4992] < btm_1[4999:4992]) ? 1 : 0;
assign detect_min[623][22] = (mid_1[4999:4992] < btm_1[5007:5000]) ? 1 : 0;
assign detect_min[623][23] = (mid_1[4999:4992] < btm_2[4991:4984]) ? 1 : 0;
assign detect_min[623][24] = (mid_1[4999:4992] < btm_2[4999:4992]) ? 1 : 0;
assign detect_min[623][25] = (mid_1[4999:4992] < btm_2[5007:5000]) ? 1 : 0;

assign detect_min[624][0] = (mid_1[5007:5000] < top_0[4999:4992]) ? 1 : 0;
assign detect_min[624][1] = (mid_1[5007:5000] < top_0[5007:5000]) ? 1 : 0;
assign detect_min[624][2] = (mid_1[5007:5000] < top_0[5015:5008]) ? 1 : 0;
assign detect_min[624][3] = (mid_1[5007:5000] < top_1[4999:4992]) ? 1 : 0;
assign detect_min[624][4] = (mid_1[5007:5000] < top_1[5007:5000]) ? 1 : 0;
assign detect_min[624][5] = (mid_1[5007:5000] < top_1[5015:5008]) ? 1 : 0;
assign detect_min[624][6] = (mid_1[5007:5000] < top_2[4999:4992]) ? 1 : 0;
assign detect_min[624][7] = (mid_1[5007:5000] < top_2[5007:5000]) ? 1 : 0;
assign detect_min[624][8] = (mid_1[5007:5000] < top_2[5015:5008]) ? 1 : 0;
assign detect_min[624][9] = (mid_1[5007:5000] < mid_0[4999:4992]) ? 1 : 0;
assign detect_min[624][10] = (mid_1[5007:5000] < mid_0[5007:5000]) ? 1 : 0;
assign detect_min[624][11] = (mid_1[5007:5000] < mid_0[5015:5008]) ? 1 : 0;
assign detect_min[624][12] = (mid_1[5007:5000] < mid_1[4999:4992]) ? 1 : 0;
assign detect_min[624][13] = (mid_1[5007:5000] < mid_1[5015:5008]) ? 1 : 0;
assign detect_min[624][14] = (mid_1[5007:5000] < mid_2[4999:4992]) ? 1 : 0;
assign detect_min[624][15] = (mid_1[5007:5000] < mid_2[5007:5000]) ? 1 : 0;
assign detect_min[624][16] = (mid_1[5007:5000] < mid_2[5015:5008]) ? 1 : 0;
assign detect_min[624][17] = (mid_1[5007:5000] < btm_0[4999:4992]) ? 1 : 0;
assign detect_min[624][18] = (mid_1[5007:5000] < btm_0[5007:5000]) ? 1 : 0;
assign detect_min[624][19] = (mid_1[5007:5000] < btm_0[5015:5008]) ? 1 : 0;
assign detect_min[624][20] = (mid_1[5007:5000] < btm_1[4999:4992]) ? 1 : 0;
assign detect_min[624][21] = (mid_1[5007:5000] < btm_1[5007:5000]) ? 1 : 0;
assign detect_min[624][22] = (mid_1[5007:5000] < btm_1[5015:5008]) ? 1 : 0;
assign detect_min[624][23] = (mid_1[5007:5000] < btm_2[4999:4992]) ? 1 : 0;
assign detect_min[624][24] = (mid_1[5007:5000] < btm_2[5007:5000]) ? 1 : 0;
assign detect_min[624][25] = (mid_1[5007:5000] < btm_2[5015:5008]) ? 1 : 0;

assign detect_min[625][0] = (mid_1[5015:5008] < top_0[5007:5000]) ? 1 : 0;
assign detect_min[625][1] = (mid_1[5015:5008] < top_0[5015:5008]) ? 1 : 0;
assign detect_min[625][2] = (mid_1[5015:5008] < top_0[5023:5016]) ? 1 : 0;
assign detect_min[625][3] = (mid_1[5015:5008] < top_1[5007:5000]) ? 1 : 0;
assign detect_min[625][4] = (mid_1[5015:5008] < top_1[5015:5008]) ? 1 : 0;
assign detect_min[625][5] = (mid_1[5015:5008] < top_1[5023:5016]) ? 1 : 0;
assign detect_min[625][6] = (mid_1[5015:5008] < top_2[5007:5000]) ? 1 : 0;
assign detect_min[625][7] = (mid_1[5015:5008] < top_2[5015:5008]) ? 1 : 0;
assign detect_min[625][8] = (mid_1[5015:5008] < top_2[5023:5016]) ? 1 : 0;
assign detect_min[625][9] = (mid_1[5015:5008] < mid_0[5007:5000]) ? 1 : 0;
assign detect_min[625][10] = (mid_1[5015:5008] < mid_0[5015:5008]) ? 1 : 0;
assign detect_min[625][11] = (mid_1[5015:5008] < mid_0[5023:5016]) ? 1 : 0;
assign detect_min[625][12] = (mid_1[5015:5008] < mid_1[5007:5000]) ? 1 : 0;
assign detect_min[625][13] = (mid_1[5015:5008] < mid_1[5023:5016]) ? 1 : 0;
assign detect_min[625][14] = (mid_1[5015:5008] < mid_2[5007:5000]) ? 1 : 0;
assign detect_min[625][15] = (mid_1[5015:5008] < mid_2[5015:5008]) ? 1 : 0;
assign detect_min[625][16] = (mid_1[5015:5008] < mid_2[5023:5016]) ? 1 : 0;
assign detect_min[625][17] = (mid_1[5015:5008] < btm_0[5007:5000]) ? 1 : 0;
assign detect_min[625][18] = (mid_1[5015:5008] < btm_0[5015:5008]) ? 1 : 0;
assign detect_min[625][19] = (mid_1[5015:5008] < btm_0[5023:5016]) ? 1 : 0;
assign detect_min[625][20] = (mid_1[5015:5008] < btm_1[5007:5000]) ? 1 : 0;
assign detect_min[625][21] = (mid_1[5015:5008] < btm_1[5015:5008]) ? 1 : 0;
assign detect_min[625][22] = (mid_1[5015:5008] < btm_1[5023:5016]) ? 1 : 0;
assign detect_min[625][23] = (mid_1[5015:5008] < btm_2[5007:5000]) ? 1 : 0;
assign detect_min[625][24] = (mid_1[5015:5008] < btm_2[5015:5008]) ? 1 : 0;
assign detect_min[625][25] = (mid_1[5015:5008] < btm_2[5023:5016]) ? 1 : 0;

assign detect_min[626][0] = (mid_1[5023:5016] < top_0[5015:5008]) ? 1 : 0;
assign detect_min[626][1] = (mid_1[5023:5016] < top_0[5023:5016]) ? 1 : 0;
assign detect_min[626][2] = (mid_1[5023:5016] < top_0[5031:5024]) ? 1 : 0;
assign detect_min[626][3] = (mid_1[5023:5016] < top_1[5015:5008]) ? 1 : 0;
assign detect_min[626][4] = (mid_1[5023:5016] < top_1[5023:5016]) ? 1 : 0;
assign detect_min[626][5] = (mid_1[5023:5016] < top_1[5031:5024]) ? 1 : 0;
assign detect_min[626][6] = (mid_1[5023:5016] < top_2[5015:5008]) ? 1 : 0;
assign detect_min[626][7] = (mid_1[5023:5016] < top_2[5023:5016]) ? 1 : 0;
assign detect_min[626][8] = (mid_1[5023:5016] < top_2[5031:5024]) ? 1 : 0;
assign detect_min[626][9] = (mid_1[5023:5016] < mid_0[5015:5008]) ? 1 : 0;
assign detect_min[626][10] = (mid_1[5023:5016] < mid_0[5023:5016]) ? 1 : 0;
assign detect_min[626][11] = (mid_1[5023:5016] < mid_0[5031:5024]) ? 1 : 0;
assign detect_min[626][12] = (mid_1[5023:5016] < mid_1[5015:5008]) ? 1 : 0;
assign detect_min[626][13] = (mid_1[5023:5016] < mid_1[5031:5024]) ? 1 : 0;
assign detect_min[626][14] = (mid_1[5023:5016] < mid_2[5015:5008]) ? 1 : 0;
assign detect_min[626][15] = (mid_1[5023:5016] < mid_2[5023:5016]) ? 1 : 0;
assign detect_min[626][16] = (mid_1[5023:5016] < mid_2[5031:5024]) ? 1 : 0;
assign detect_min[626][17] = (mid_1[5023:5016] < btm_0[5015:5008]) ? 1 : 0;
assign detect_min[626][18] = (mid_1[5023:5016] < btm_0[5023:5016]) ? 1 : 0;
assign detect_min[626][19] = (mid_1[5023:5016] < btm_0[5031:5024]) ? 1 : 0;
assign detect_min[626][20] = (mid_1[5023:5016] < btm_1[5015:5008]) ? 1 : 0;
assign detect_min[626][21] = (mid_1[5023:5016] < btm_1[5023:5016]) ? 1 : 0;
assign detect_min[626][22] = (mid_1[5023:5016] < btm_1[5031:5024]) ? 1 : 0;
assign detect_min[626][23] = (mid_1[5023:5016] < btm_2[5015:5008]) ? 1 : 0;
assign detect_min[626][24] = (mid_1[5023:5016] < btm_2[5023:5016]) ? 1 : 0;
assign detect_min[626][25] = (mid_1[5023:5016] < btm_2[5031:5024]) ? 1 : 0;

assign detect_min[627][0] = (mid_1[5031:5024] < top_0[5023:5016]) ? 1 : 0;
assign detect_min[627][1] = (mid_1[5031:5024] < top_0[5031:5024]) ? 1 : 0;
assign detect_min[627][2] = (mid_1[5031:5024] < top_0[5039:5032]) ? 1 : 0;
assign detect_min[627][3] = (mid_1[5031:5024] < top_1[5023:5016]) ? 1 : 0;
assign detect_min[627][4] = (mid_1[5031:5024] < top_1[5031:5024]) ? 1 : 0;
assign detect_min[627][5] = (mid_1[5031:5024] < top_1[5039:5032]) ? 1 : 0;
assign detect_min[627][6] = (mid_1[5031:5024] < top_2[5023:5016]) ? 1 : 0;
assign detect_min[627][7] = (mid_1[5031:5024] < top_2[5031:5024]) ? 1 : 0;
assign detect_min[627][8] = (mid_1[5031:5024] < top_2[5039:5032]) ? 1 : 0;
assign detect_min[627][9] = (mid_1[5031:5024] < mid_0[5023:5016]) ? 1 : 0;
assign detect_min[627][10] = (mid_1[5031:5024] < mid_0[5031:5024]) ? 1 : 0;
assign detect_min[627][11] = (mid_1[5031:5024] < mid_0[5039:5032]) ? 1 : 0;
assign detect_min[627][12] = (mid_1[5031:5024] < mid_1[5023:5016]) ? 1 : 0;
assign detect_min[627][13] = (mid_1[5031:5024] < mid_1[5039:5032]) ? 1 : 0;
assign detect_min[627][14] = (mid_1[5031:5024] < mid_2[5023:5016]) ? 1 : 0;
assign detect_min[627][15] = (mid_1[5031:5024] < mid_2[5031:5024]) ? 1 : 0;
assign detect_min[627][16] = (mid_1[5031:5024] < mid_2[5039:5032]) ? 1 : 0;
assign detect_min[627][17] = (mid_1[5031:5024] < btm_0[5023:5016]) ? 1 : 0;
assign detect_min[627][18] = (mid_1[5031:5024] < btm_0[5031:5024]) ? 1 : 0;
assign detect_min[627][19] = (mid_1[5031:5024] < btm_0[5039:5032]) ? 1 : 0;
assign detect_min[627][20] = (mid_1[5031:5024] < btm_1[5023:5016]) ? 1 : 0;
assign detect_min[627][21] = (mid_1[5031:5024] < btm_1[5031:5024]) ? 1 : 0;
assign detect_min[627][22] = (mid_1[5031:5024] < btm_1[5039:5032]) ? 1 : 0;
assign detect_min[627][23] = (mid_1[5031:5024] < btm_2[5023:5016]) ? 1 : 0;
assign detect_min[627][24] = (mid_1[5031:5024] < btm_2[5031:5024]) ? 1 : 0;
assign detect_min[627][25] = (mid_1[5031:5024] < btm_2[5039:5032]) ? 1 : 0;

assign detect_min[628][0] = (mid_1[5039:5032] < top_0[5031:5024]) ? 1 : 0;
assign detect_min[628][1] = (mid_1[5039:5032] < top_0[5039:5032]) ? 1 : 0;
assign detect_min[628][2] = (mid_1[5039:5032] < top_0[5047:5040]) ? 1 : 0;
assign detect_min[628][3] = (mid_1[5039:5032] < top_1[5031:5024]) ? 1 : 0;
assign detect_min[628][4] = (mid_1[5039:5032] < top_1[5039:5032]) ? 1 : 0;
assign detect_min[628][5] = (mid_1[5039:5032] < top_1[5047:5040]) ? 1 : 0;
assign detect_min[628][6] = (mid_1[5039:5032] < top_2[5031:5024]) ? 1 : 0;
assign detect_min[628][7] = (mid_1[5039:5032] < top_2[5039:5032]) ? 1 : 0;
assign detect_min[628][8] = (mid_1[5039:5032] < top_2[5047:5040]) ? 1 : 0;
assign detect_min[628][9] = (mid_1[5039:5032] < mid_0[5031:5024]) ? 1 : 0;
assign detect_min[628][10] = (mid_1[5039:5032] < mid_0[5039:5032]) ? 1 : 0;
assign detect_min[628][11] = (mid_1[5039:5032] < mid_0[5047:5040]) ? 1 : 0;
assign detect_min[628][12] = (mid_1[5039:5032] < mid_1[5031:5024]) ? 1 : 0;
assign detect_min[628][13] = (mid_1[5039:5032] < mid_1[5047:5040]) ? 1 : 0;
assign detect_min[628][14] = (mid_1[5039:5032] < mid_2[5031:5024]) ? 1 : 0;
assign detect_min[628][15] = (mid_1[5039:5032] < mid_2[5039:5032]) ? 1 : 0;
assign detect_min[628][16] = (mid_1[5039:5032] < mid_2[5047:5040]) ? 1 : 0;
assign detect_min[628][17] = (mid_1[5039:5032] < btm_0[5031:5024]) ? 1 : 0;
assign detect_min[628][18] = (mid_1[5039:5032] < btm_0[5039:5032]) ? 1 : 0;
assign detect_min[628][19] = (mid_1[5039:5032] < btm_0[5047:5040]) ? 1 : 0;
assign detect_min[628][20] = (mid_1[5039:5032] < btm_1[5031:5024]) ? 1 : 0;
assign detect_min[628][21] = (mid_1[5039:5032] < btm_1[5039:5032]) ? 1 : 0;
assign detect_min[628][22] = (mid_1[5039:5032] < btm_1[5047:5040]) ? 1 : 0;
assign detect_min[628][23] = (mid_1[5039:5032] < btm_2[5031:5024]) ? 1 : 0;
assign detect_min[628][24] = (mid_1[5039:5032] < btm_2[5039:5032]) ? 1 : 0;
assign detect_min[628][25] = (mid_1[5039:5032] < btm_2[5047:5040]) ? 1 : 0;

assign detect_min[629][0] = (mid_1[5047:5040] < top_0[5039:5032]) ? 1 : 0;
assign detect_min[629][1] = (mid_1[5047:5040] < top_0[5047:5040]) ? 1 : 0;
assign detect_min[629][2] = (mid_1[5047:5040] < top_0[5055:5048]) ? 1 : 0;
assign detect_min[629][3] = (mid_1[5047:5040] < top_1[5039:5032]) ? 1 : 0;
assign detect_min[629][4] = (mid_1[5047:5040] < top_1[5047:5040]) ? 1 : 0;
assign detect_min[629][5] = (mid_1[5047:5040] < top_1[5055:5048]) ? 1 : 0;
assign detect_min[629][6] = (mid_1[5047:5040] < top_2[5039:5032]) ? 1 : 0;
assign detect_min[629][7] = (mid_1[5047:5040] < top_2[5047:5040]) ? 1 : 0;
assign detect_min[629][8] = (mid_1[5047:5040] < top_2[5055:5048]) ? 1 : 0;
assign detect_min[629][9] = (mid_1[5047:5040] < mid_0[5039:5032]) ? 1 : 0;
assign detect_min[629][10] = (mid_1[5047:5040] < mid_0[5047:5040]) ? 1 : 0;
assign detect_min[629][11] = (mid_1[5047:5040] < mid_0[5055:5048]) ? 1 : 0;
assign detect_min[629][12] = (mid_1[5047:5040] < mid_1[5039:5032]) ? 1 : 0;
assign detect_min[629][13] = (mid_1[5047:5040] < mid_1[5055:5048]) ? 1 : 0;
assign detect_min[629][14] = (mid_1[5047:5040] < mid_2[5039:5032]) ? 1 : 0;
assign detect_min[629][15] = (mid_1[5047:5040] < mid_2[5047:5040]) ? 1 : 0;
assign detect_min[629][16] = (mid_1[5047:5040] < mid_2[5055:5048]) ? 1 : 0;
assign detect_min[629][17] = (mid_1[5047:5040] < btm_0[5039:5032]) ? 1 : 0;
assign detect_min[629][18] = (mid_1[5047:5040] < btm_0[5047:5040]) ? 1 : 0;
assign detect_min[629][19] = (mid_1[5047:5040] < btm_0[5055:5048]) ? 1 : 0;
assign detect_min[629][20] = (mid_1[5047:5040] < btm_1[5039:5032]) ? 1 : 0;
assign detect_min[629][21] = (mid_1[5047:5040] < btm_1[5047:5040]) ? 1 : 0;
assign detect_min[629][22] = (mid_1[5047:5040] < btm_1[5055:5048]) ? 1 : 0;
assign detect_min[629][23] = (mid_1[5047:5040] < btm_2[5039:5032]) ? 1 : 0;
assign detect_min[629][24] = (mid_1[5047:5040] < btm_2[5047:5040]) ? 1 : 0;
assign detect_min[629][25] = (mid_1[5047:5040] < btm_2[5055:5048]) ? 1 : 0;

assign detect_min[630][0] = (mid_1[5055:5048] < top_0[5047:5040]) ? 1 : 0;
assign detect_min[630][1] = (mid_1[5055:5048] < top_0[5055:5048]) ? 1 : 0;
assign detect_min[630][2] = (mid_1[5055:5048] < top_0[5063:5056]) ? 1 : 0;
assign detect_min[630][3] = (mid_1[5055:5048] < top_1[5047:5040]) ? 1 : 0;
assign detect_min[630][4] = (mid_1[5055:5048] < top_1[5055:5048]) ? 1 : 0;
assign detect_min[630][5] = (mid_1[5055:5048] < top_1[5063:5056]) ? 1 : 0;
assign detect_min[630][6] = (mid_1[5055:5048] < top_2[5047:5040]) ? 1 : 0;
assign detect_min[630][7] = (mid_1[5055:5048] < top_2[5055:5048]) ? 1 : 0;
assign detect_min[630][8] = (mid_1[5055:5048] < top_2[5063:5056]) ? 1 : 0;
assign detect_min[630][9] = (mid_1[5055:5048] < mid_0[5047:5040]) ? 1 : 0;
assign detect_min[630][10] = (mid_1[5055:5048] < mid_0[5055:5048]) ? 1 : 0;
assign detect_min[630][11] = (mid_1[5055:5048] < mid_0[5063:5056]) ? 1 : 0;
assign detect_min[630][12] = (mid_1[5055:5048] < mid_1[5047:5040]) ? 1 : 0;
assign detect_min[630][13] = (mid_1[5055:5048] < mid_1[5063:5056]) ? 1 : 0;
assign detect_min[630][14] = (mid_1[5055:5048] < mid_2[5047:5040]) ? 1 : 0;
assign detect_min[630][15] = (mid_1[5055:5048] < mid_2[5055:5048]) ? 1 : 0;
assign detect_min[630][16] = (mid_1[5055:5048] < mid_2[5063:5056]) ? 1 : 0;
assign detect_min[630][17] = (mid_1[5055:5048] < btm_0[5047:5040]) ? 1 : 0;
assign detect_min[630][18] = (mid_1[5055:5048] < btm_0[5055:5048]) ? 1 : 0;
assign detect_min[630][19] = (mid_1[5055:5048] < btm_0[5063:5056]) ? 1 : 0;
assign detect_min[630][20] = (mid_1[5055:5048] < btm_1[5047:5040]) ? 1 : 0;
assign detect_min[630][21] = (mid_1[5055:5048] < btm_1[5055:5048]) ? 1 : 0;
assign detect_min[630][22] = (mid_1[5055:5048] < btm_1[5063:5056]) ? 1 : 0;
assign detect_min[630][23] = (mid_1[5055:5048] < btm_2[5047:5040]) ? 1 : 0;
assign detect_min[630][24] = (mid_1[5055:5048] < btm_2[5055:5048]) ? 1 : 0;
assign detect_min[630][25] = (mid_1[5055:5048] < btm_2[5063:5056]) ? 1 : 0;

assign detect_min[631][0] = (mid_1[5063:5056] < top_0[5055:5048]) ? 1 : 0;
assign detect_min[631][1] = (mid_1[5063:5056] < top_0[5063:5056]) ? 1 : 0;
assign detect_min[631][2] = (mid_1[5063:5056] < top_0[5071:5064]) ? 1 : 0;
assign detect_min[631][3] = (mid_1[5063:5056] < top_1[5055:5048]) ? 1 : 0;
assign detect_min[631][4] = (mid_1[5063:5056] < top_1[5063:5056]) ? 1 : 0;
assign detect_min[631][5] = (mid_1[5063:5056] < top_1[5071:5064]) ? 1 : 0;
assign detect_min[631][6] = (mid_1[5063:5056] < top_2[5055:5048]) ? 1 : 0;
assign detect_min[631][7] = (mid_1[5063:5056] < top_2[5063:5056]) ? 1 : 0;
assign detect_min[631][8] = (mid_1[5063:5056] < top_2[5071:5064]) ? 1 : 0;
assign detect_min[631][9] = (mid_1[5063:5056] < mid_0[5055:5048]) ? 1 : 0;
assign detect_min[631][10] = (mid_1[5063:5056] < mid_0[5063:5056]) ? 1 : 0;
assign detect_min[631][11] = (mid_1[5063:5056] < mid_0[5071:5064]) ? 1 : 0;
assign detect_min[631][12] = (mid_1[5063:5056] < mid_1[5055:5048]) ? 1 : 0;
assign detect_min[631][13] = (mid_1[5063:5056] < mid_1[5071:5064]) ? 1 : 0;
assign detect_min[631][14] = (mid_1[5063:5056] < mid_2[5055:5048]) ? 1 : 0;
assign detect_min[631][15] = (mid_1[5063:5056] < mid_2[5063:5056]) ? 1 : 0;
assign detect_min[631][16] = (mid_1[5063:5056] < mid_2[5071:5064]) ? 1 : 0;
assign detect_min[631][17] = (mid_1[5063:5056] < btm_0[5055:5048]) ? 1 : 0;
assign detect_min[631][18] = (mid_1[5063:5056] < btm_0[5063:5056]) ? 1 : 0;
assign detect_min[631][19] = (mid_1[5063:5056] < btm_0[5071:5064]) ? 1 : 0;
assign detect_min[631][20] = (mid_1[5063:5056] < btm_1[5055:5048]) ? 1 : 0;
assign detect_min[631][21] = (mid_1[5063:5056] < btm_1[5063:5056]) ? 1 : 0;
assign detect_min[631][22] = (mid_1[5063:5056] < btm_1[5071:5064]) ? 1 : 0;
assign detect_min[631][23] = (mid_1[5063:5056] < btm_2[5055:5048]) ? 1 : 0;
assign detect_min[631][24] = (mid_1[5063:5056] < btm_2[5063:5056]) ? 1 : 0;
assign detect_min[631][25] = (mid_1[5063:5056] < btm_2[5071:5064]) ? 1 : 0;

assign detect_min[632][0] = (mid_1[5071:5064] < top_0[5063:5056]) ? 1 : 0;
assign detect_min[632][1] = (mid_1[5071:5064] < top_0[5071:5064]) ? 1 : 0;
assign detect_min[632][2] = (mid_1[5071:5064] < top_0[5079:5072]) ? 1 : 0;
assign detect_min[632][3] = (mid_1[5071:5064] < top_1[5063:5056]) ? 1 : 0;
assign detect_min[632][4] = (mid_1[5071:5064] < top_1[5071:5064]) ? 1 : 0;
assign detect_min[632][5] = (mid_1[5071:5064] < top_1[5079:5072]) ? 1 : 0;
assign detect_min[632][6] = (mid_1[5071:5064] < top_2[5063:5056]) ? 1 : 0;
assign detect_min[632][7] = (mid_1[5071:5064] < top_2[5071:5064]) ? 1 : 0;
assign detect_min[632][8] = (mid_1[5071:5064] < top_2[5079:5072]) ? 1 : 0;
assign detect_min[632][9] = (mid_1[5071:5064] < mid_0[5063:5056]) ? 1 : 0;
assign detect_min[632][10] = (mid_1[5071:5064] < mid_0[5071:5064]) ? 1 : 0;
assign detect_min[632][11] = (mid_1[5071:5064] < mid_0[5079:5072]) ? 1 : 0;
assign detect_min[632][12] = (mid_1[5071:5064] < mid_1[5063:5056]) ? 1 : 0;
assign detect_min[632][13] = (mid_1[5071:5064] < mid_1[5079:5072]) ? 1 : 0;
assign detect_min[632][14] = (mid_1[5071:5064] < mid_2[5063:5056]) ? 1 : 0;
assign detect_min[632][15] = (mid_1[5071:5064] < mid_2[5071:5064]) ? 1 : 0;
assign detect_min[632][16] = (mid_1[5071:5064] < mid_2[5079:5072]) ? 1 : 0;
assign detect_min[632][17] = (mid_1[5071:5064] < btm_0[5063:5056]) ? 1 : 0;
assign detect_min[632][18] = (mid_1[5071:5064] < btm_0[5071:5064]) ? 1 : 0;
assign detect_min[632][19] = (mid_1[5071:5064] < btm_0[5079:5072]) ? 1 : 0;
assign detect_min[632][20] = (mid_1[5071:5064] < btm_1[5063:5056]) ? 1 : 0;
assign detect_min[632][21] = (mid_1[5071:5064] < btm_1[5071:5064]) ? 1 : 0;
assign detect_min[632][22] = (mid_1[5071:5064] < btm_1[5079:5072]) ? 1 : 0;
assign detect_min[632][23] = (mid_1[5071:5064] < btm_2[5063:5056]) ? 1 : 0;
assign detect_min[632][24] = (mid_1[5071:5064] < btm_2[5071:5064]) ? 1 : 0;
assign detect_min[632][25] = (mid_1[5071:5064] < btm_2[5079:5072]) ? 1 : 0;

assign detect_min[633][0] = (mid_1[5079:5072] < top_0[5071:5064]) ? 1 : 0;
assign detect_min[633][1] = (mid_1[5079:5072] < top_0[5079:5072]) ? 1 : 0;
assign detect_min[633][2] = (mid_1[5079:5072] < top_0[5087:5080]) ? 1 : 0;
assign detect_min[633][3] = (mid_1[5079:5072] < top_1[5071:5064]) ? 1 : 0;
assign detect_min[633][4] = (mid_1[5079:5072] < top_1[5079:5072]) ? 1 : 0;
assign detect_min[633][5] = (mid_1[5079:5072] < top_1[5087:5080]) ? 1 : 0;
assign detect_min[633][6] = (mid_1[5079:5072] < top_2[5071:5064]) ? 1 : 0;
assign detect_min[633][7] = (mid_1[5079:5072] < top_2[5079:5072]) ? 1 : 0;
assign detect_min[633][8] = (mid_1[5079:5072] < top_2[5087:5080]) ? 1 : 0;
assign detect_min[633][9] = (mid_1[5079:5072] < mid_0[5071:5064]) ? 1 : 0;
assign detect_min[633][10] = (mid_1[5079:5072] < mid_0[5079:5072]) ? 1 : 0;
assign detect_min[633][11] = (mid_1[5079:5072] < mid_0[5087:5080]) ? 1 : 0;
assign detect_min[633][12] = (mid_1[5079:5072] < mid_1[5071:5064]) ? 1 : 0;
assign detect_min[633][13] = (mid_1[5079:5072] < mid_1[5087:5080]) ? 1 : 0;
assign detect_min[633][14] = (mid_1[5079:5072] < mid_2[5071:5064]) ? 1 : 0;
assign detect_min[633][15] = (mid_1[5079:5072] < mid_2[5079:5072]) ? 1 : 0;
assign detect_min[633][16] = (mid_1[5079:5072] < mid_2[5087:5080]) ? 1 : 0;
assign detect_min[633][17] = (mid_1[5079:5072] < btm_0[5071:5064]) ? 1 : 0;
assign detect_min[633][18] = (mid_1[5079:5072] < btm_0[5079:5072]) ? 1 : 0;
assign detect_min[633][19] = (mid_1[5079:5072] < btm_0[5087:5080]) ? 1 : 0;
assign detect_min[633][20] = (mid_1[5079:5072] < btm_1[5071:5064]) ? 1 : 0;
assign detect_min[633][21] = (mid_1[5079:5072] < btm_1[5079:5072]) ? 1 : 0;
assign detect_min[633][22] = (mid_1[5079:5072] < btm_1[5087:5080]) ? 1 : 0;
assign detect_min[633][23] = (mid_1[5079:5072] < btm_2[5071:5064]) ? 1 : 0;
assign detect_min[633][24] = (mid_1[5079:5072] < btm_2[5079:5072]) ? 1 : 0;
assign detect_min[633][25] = (mid_1[5079:5072] < btm_2[5087:5080]) ? 1 : 0;

assign detect_min[634][0] = (mid_1[5087:5080] < top_0[5079:5072]) ? 1 : 0;
assign detect_min[634][1] = (mid_1[5087:5080] < top_0[5087:5080]) ? 1 : 0;
assign detect_min[634][2] = (mid_1[5087:5080] < top_0[5095:5088]) ? 1 : 0;
assign detect_min[634][3] = (mid_1[5087:5080] < top_1[5079:5072]) ? 1 : 0;
assign detect_min[634][4] = (mid_1[5087:5080] < top_1[5087:5080]) ? 1 : 0;
assign detect_min[634][5] = (mid_1[5087:5080] < top_1[5095:5088]) ? 1 : 0;
assign detect_min[634][6] = (mid_1[5087:5080] < top_2[5079:5072]) ? 1 : 0;
assign detect_min[634][7] = (mid_1[5087:5080] < top_2[5087:5080]) ? 1 : 0;
assign detect_min[634][8] = (mid_1[5087:5080] < top_2[5095:5088]) ? 1 : 0;
assign detect_min[634][9] = (mid_1[5087:5080] < mid_0[5079:5072]) ? 1 : 0;
assign detect_min[634][10] = (mid_1[5087:5080] < mid_0[5087:5080]) ? 1 : 0;
assign detect_min[634][11] = (mid_1[5087:5080] < mid_0[5095:5088]) ? 1 : 0;
assign detect_min[634][12] = (mid_1[5087:5080] < mid_1[5079:5072]) ? 1 : 0;
assign detect_min[634][13] = (mid_1[5087:5080] < mid_1[5095:5088]) ? 1 : 0;
assign detect_min[634][14] = (mid_1[5087:5080] < mid_2[5079:5072]) ? 1 : 0;
assign detect_min[634][15] = (mid_1[5087:5080] < mid_2[5087:5080]) ? 1 : 0;
assign detect_min[634][16] = (mid_1[5087:5080] < mid_2[5095:5088]) ? 1 : 0;
assign detect_min[634][17] = (mid_1[5087:5080] < btm_0[5079:5072]) ? 1 : 0;
assign detect_min[634][18] = (mid_1[5087:5080] < btm_0[5087:5080]) ? 1 : 0;
assign detect_min[634][19] = (mid_1[5087:5080] < btm_0[5095:5088]) ? 1 : 0;
assign detect_min[634][20] = (mid_1[5087:5080] < btm_1[5079:5072]) ? 1 : 0;
assign detect_min[634][21] = (mid_1[5087:5080] < btm_1[5087:5080]) ? 1 : 0;
assign detect_min[634][22] = (mid_1[5087:5080] < btm_1[5095:5088]) ? 1 : 0;
assign detect_min[634][23] = (mid_1[5087:5080] < btm_2[5079:5072]) ? 1 : 0;
assign detect_min[634][24] = (mid_1[5087:5080] < btm_2[5087:5080]) ? 1 : 0;
assign detect_min[634][25] = (mid_1[5087:5080] < btm_2[5095:5088]) ? 1 : 0;

assign detect_min[635][0] = (mid_1[5095:5088] < top_0[5087:5080]) ? 1 : 0;
assign detect_min[635][1] = (mid_1[5095:5088] < top_0[5095:5088]) ? 1 : 0;
assign detect_min[635][2] = (mid_1[5095:5088] < top_0[5103:5096]) ? 1 : 0;
assign detect_min[635][3] = (mid_1[5095:5088] < top_1[5087:5080]) ? 1 : 0;
assign detect_min[635][4] = (mid_1[5095:5088] < top_1[5095:5088]) ? 1 : 0;
assign detect_min[635][5] = (mid_1[5095:5088] < top_1[5103:5096]) ? 1 : 0;
assign detect_min[635][6] = (mid_1[5095:5088] < top_2[5087:5080]) ? 1 : 0;
assign detect_min[635][7] = (mid_1[5095:5088] < top_2[5095:5088]) ? 1 : 0;
assign detect_min[635][8] = (mid_1[5095:5088] < top_2[5103:5096]) ? 1 : 0;
assign detect_min[635][9] = (mid_1[5095:5088] < mid_0[5087:5080]) ? 1 : 0;
assign detect_min[635][10] = (mid_1[5095:5088] < mid_0[5095:5088]) ? 1 : 0;
assign detect_min[635][11] = (mid_1[5095:5088] < mid_0[5103:5096]) ? 1 : 0;
assign detect_min[635][12] = (mid_1[5095:5088] < mid_1[5087:5080]) ? 1 : 0;
assign detect_min[635][13] = (mid_1[5095:5088] < mid_1[5103:5096]) ? 1 : 0;
assign detect_min[635][14] = (mid_1[5095:5088] < mid_2[5087:5080]) ? 1 : 0;
assign detect_min[635][15] = (mid_1[5095:5088] < mid_2[5095:5088]) ? 1 : 0;
assign detect_min[635][16] = (mid_1[5095:5088] < mid_2[5103:5096]) ? 1 : 0;
assign detect_min[635][17] = (mid_1[5095:5088] < btm_0[5087:5080]) ? 1 : 0;
assign detect_min[635][18] = (mid_1[5095:5088] < btm_0[5095:5088]) ? 1 : 0;
assign detect_min[635][19] = (mid_1[5095:5088] < btm_0[5103:5096]) ? 1 : 0;
assign detect_min[635][20] = (mid_1[5095:5088] < btm_1[5087:5080]) ? 1 : 0;
assign detect_min[635][21] = (mid_1[5095:5088] < btm_1[5095:5088]) ? 1 : 0;
assign detect_min[635][22] = (mid_1[5095:5088] < btm_1[5103:5096]) ? 1 : 0;
assign detect_min[635][23] = (mid_1[5095:5088] < btm_2[5087:5080]) ? 1 : 0;
assign detect_min[635][24] = (mid_1[5095:5088] < btm_2[5095:5088]) ? 1 : 0;
assign detect_min[635][25] = (mid_1[5095:5088] < btm_2[5103:5096]) ? 1 : 0;

assign detect_min[636][0] = (mid_1[5103:5096] < top_0[5095:5088]) ? 1 : 0;
assign detect_min[636][1] = (mid_1[5103:5096] < top_0[5103:5096]) ? 1 : 0;
assign detect_min[636][2] = (mid_1[5103:5096] < top_0[5111:5104]) ? 1 : 0;
assign detect_min[636][3] = (mid_1[5103:5096] < top_1[5095:5088]) ? 1 : 0;
assign detect_min[636][4] = (mid_1[5103:5096] < top_1[5103:5096]) ? 1 : 0;
assign detect_min[636][5] = (mid_1[5103:5096] < top_1[5111:5104]) ? 1 : 0;
assign detect_min[636][6] = (mid_1[5103:5096] < top_2[5095:5088]) ? 1 : 0;
assign detect_min[636][7] = (mid_1[5103:5096] < top_2[5103:5096]) ? 1 : 0;
assign detect_min[636][8] = (mid_1[5103:5096] < top_2[5111:5104]) ? 1 : 0;
assign detect_min[636][9] = (mid_1[5103:5096] < mid_0[5095:5088]) ? 1 : 0;
assign detect_min[636][10] = (mid_1[5103:5096] < mid_0[5103:5096]) ? 1 : 0;
assign detect_min[636][11] = (mid_1[5103:5096] < mid_0[5111:5104]) ? 1 : 0;
assign detect_min[636][12] = (mid_1[5103:5096] < mid_1[5095:5088]) ? 1 : 0;
assign detect_min[636][13] = (mid_1[5103:5096] < mid_1[5111:5104]) ? 1 : 0;
assign detect_min[636][14] = (mid_1[5103:5096] < mid_2[5095:5088]) ? 1 : 0;
assign detect_min[636][15] = (mid_1[5103:5096] < mid_2[5103:5096]) ? 1 : 0;
assign detect_min[636][16] = (mid_1[5103:5096] < mid_2[5111:5104]) ? 1 : 0;
assign detect_min[636][17] = (mid_1[5103:5096] < btm_0[5095:5088]) ? 1 : 0;
assign detect_min[636][18] = (mid_1[5103:5096] < btm_0[5103:5096]) ? 1 : 0;
assign detect_min[636][19] = (mid_1[5103:5096] < btm_0[5111:5104]) ? 1 : 0;
assign detect_min[636][20] = (mid_1[5103:5096] < btm_1[5095:5088]) ? 1 : 0;
assign detect_min[636][21] = (mid_1[5103:5096] < btm_1[5103:5096]) ? 1 : 0;
assign detect_min[636][22] = (mid_1[5103:5096] < btm_1[5111:5104]) ? 1 : 0;
assign detect_min[636][23] = (mid_1[5103:5096] < btm_2[5095:5088]) ? 1 : 0;
assign detect_min[636][24] = (mid_1[5103:5096] < btm_2[5103:5096]) ? 1 : 0;
assign detect_min[636][25] = (mid_1[5103:5096] < btm_2[5111:5104]) ? 1 : 0;

assign detect_min[637][0] = (mid_1[5111:5104] < top_0[5103:5096]) ? 1 : 0;
assign detect_min[637][1] = (mid_1[5111:5104] < top_0[5111:5104]) ? 1 : 0;
assign detect_min[637][2] = (mid_1[5111:5104] < top_0[5119:5112]) ? 1 : 0;
assign detect_min[637][3] = (mid_1[5111:5104] < top_1[5103:5096]) ? 1 : 0;
assign detect_min[637][4] = (mid_1[5111:5104] < top_1[5111:5104]) ? 1 : 0;
assign detect_min[637][5] = (mid_1[5111:5104] < top_1[5119:5112]) ? 1 : 0;
assign detect_min[637][6] = (mid_1[5111:5104] < top_2[5103:5096]) ? 1 : 0;
assign detect_min[637][7] = (mid_1[5111:5104] < top_2[5111:5104]) ? 1 : 0;
assign detect_min[637][8] = (mid_1[5111:5104] < top_2[5119:5112]) ? 1 : 0;
assign detect_min[637][9] = (mid_1[5111:5104] < mid_0[5103:5096]) ? 1 : 0;
assign detect_min[637][10] = (mid_1[5111:5104] < mid_0[5111:5104]) ? 1 : 0;
assign detect_min[637][11] = (mid_1[5111:5104] < mid_0[5119:5112]) ? 1 : 0;
assign detect_min[637][12] = (mid_1[5111:5104] < mid_1[5103:5096]) ? 1 : 0;
assign detect_min[637][13] = (mid_1[5111:5104] < mid_1[5119:5112]) ? 1 : 0;
assign detect_min[637][14] = (mid_1[5111:5104] < mid_2[5103:5096]) ? 1 : 0;
assign detect_min[637][15] = (mid_1[5111:5104] < mid_2[5111:5104]) ? 1 : 0;
assign detect_min[637][16] = (mid_1[5111:5104] < mid_2[5119:5112]) ? 1 : 0;
assign detect_min[637][17] = (mid_1[5111:5104] < btm_0[5103:5096]) ? 1 : 0;
assign detect_min[637][18] = (mid_1[5111:5104] < btm_0[5111:5104]) ? 1 : 0;
assign detect_min[637][19] = (mid_1[5111:5104] < btm_0[5119:5112]) ? 1 : 0;
assign detect_min[637][20] = (mid_1[5111:5104] < btm_1[5103:5096]) ? 1 : 0;
assign detect_min[637][21] = (mid_1[5111:5104] < btm_1[5111:5104]) ? 1 : 0;
assign detect_min[637][22] = (mid_1[5111:5104] < btm_1[5119:5112]) ? 1 : 0;
assign detect_min[637][23] = (mid_1[5111:5104] < btm_2[5103:5096]) ? 1 : 0;
assign detect_min[637][24] = (mid_1[5111:5104] < btm_2[5111:5104]) ? 1 : 0;
assign detect_min[637][25] = (mid_1[5111:5104] < btm_2[5119:5112]) ? 1 : 0;

wire [637:0] is_min;
assign is_min[0] = (&detect_min[0]) ? 1:0;
assign is_min[1] = (&detect_min[1]) ? 1:0;
assign is_min[2] = (&detect_min[2]) ? 1:0;
assign is_min[3] = (&detect_min[3]) ? 1:0;
assign is_min[4] = (&detect_min[4]) ? 1:0;
assign is_min[5] = (&detect_min[5]) ? 1:0;
assign is_min[6] = (&detect_min[6]) ? 1:0;
assign is_min[7] = (&detect_min[7]) ? 1:0;
assign is_min[8] = (&detect_min[8]) ? 1:0;
assign is_min[9] = (&detect_min[9]) ? 1:0;
assign is_min[10] = (&detect_min[10]) ? 1:0;
assign is_min[11] = (&detect_min[11]) ? 1:0;
assign is_min[12] = (&detect_min[12]) ? 1:0;
assign is_min[13] = (&detect_min[13]) ? 1:0;
assign is_min[14] = (&detect_min[14]) ? 1:0;
assign is_min[15] = (&detect_min[15]) ? 1:0;
assign is_min[16] = (&detect_min[16]) ? 1:0;
assign is_min[17] = (&detect_min[17]) ? 1:0;
assign is_min[18] = (&detect_min[18]) ? 1:0;
assign is_min[19] = (&detect_min[19]) ? 1:0;
assign is_min[20] = (&detect_min[20]) ? 1:0;
assign is_min[21] = (&detect_min[21]) ? 1:0;
assign is_min[22] = (&detect_min[22]) ? 1:0;
assign is_min[23] = (&detect_min[23]) ? 1:0;
assign is_min[24] = (&detect_min[24]) ? 1:0;
assign is_min[25] = (&detect_min[25]) ? 1:0;
assign is_min[26] = (&detect_min[26]) ? 1:0;
assign is_min[27] = (&detect_min[27]) ? 1:0;
assign is_min[28] = (&detect_min[28]) ? 1:0;
assign is_min[29] = (&detect_min[29]) ? 1:0;
assign is_min[30] = (&detect_min[30]) ? 1:0;
assign is_min[31] = (&detect_min[31]) ? 1:0;
assign is_min[32] = (&detect_min[32]) ? 1:0;
assign is_min[33] = (&detect_min[33]) ? 1:0;
assign is_min[34] = (&detect_min[34]) ? 1:0;
assign is_min[35] = (&detect_min[35]) ? 1:0;
assign is_min[36] = (&detect_min[36]) ? 1:0;
assign is_min[37] = (&detect_min[37]) ? 1:0;
assign is_min[38] = (&detect_min[38]) ? 1:0;
assign is_min[39] = (&detect_min[39]) ? 1:0;
assign is_min[40] = (&detect_min[40]) ? 1:0;
assign is_min[41] = (&detect_min[41]) ? 1:0;
assign is_min[42] = (&detect_min[42]) ? 1:0;
assign is_min[43] = (&detect_min[43]) ? 1:0;
assign is_min[44] = (&detect_min[44]) ? 1:0;
assign is_min[45] = (&detect_min[45]) ? 1:0;
assign is_min[46] = (&detect_min[46]) ? 1:0;
assign is_min[47] = (&detect_min[47]) ? 1:0;
assign is_min[48] = (&detect_min[48]) ? 1:0;
assign is_min[49] = (&detect_min[49]) ? 1:0;
assign is_min[50] = (&detect_min[50]) ? 1:0;
assign is_min[51] = (&detect_min[51]) ? 1:0;
assign is_min[52] = (&detect_min[52]) ? 1:0;
assign is_min[53] = (&detect_min[53]) ? 1:0;
assign is_min[54] = (&detect_min[54]) ? 1:0;
assign is_min[55] = (&detect_min[55]) ? 1:0;
assign is_min[56] = (&detect_min[56]) ? 1:0;
assign is_min[57] = (&detect_min[57]) ? 1:0;
assign is_min[58] = (&detect_min[58]) ? 1:0;
assign is_min[59] = (&detect_min[59]) ? 1:0;
assign is_min[60] = (&detect_min[60]) ? 1:0;
assign is_min[61] = (&detect_min[61]) ? 1:0;
assign is_min[62] = (&detect_min[62]) ? 1:0;
assign is_min[63] = (&detect_min[63]) ? 1:0;
assign is_min[64] = (&detect_min[64]) ? 1:0;
assign is_min[65] = (&detect_min[65]) ? 1:0;
assign is_min[66] = (&detect_min[66]) ? 1:0;
assign is_min[67] = (&detect_min[67]) ? 1:0;
assign is_min[68] = (&detect_min[68]) ? 1:0;
assign is_min[69] = (&detect_min[69]) ? 1:0;
assign is_min[70] = (&detect_min[70]) ? 1:0;
assign is_min[71] = (&detect_min[71]) ? 1:0;
assign is_min[72] = (&detect_min[72]) ? 1:0;
assign is_min[73] = (&detect_min[73]) ? 1:0;
assign is_min[74] = (&detect_min[74]) ? 1:0;
assign is_min[75] = (&detect_min[75]) ? 1:0;
assign is_min[76] = (&detect_min[76]) ? 1:0;
assign is_min[77] = (&detect_min[77]) ? 1:0;
assign is_min[78] = (&detect_min[78]) ? 1:0;
assign is_min[79] = (&detect_min[79]) ? 1:0;
assign is_min[80] = (&detect_min[80]) ? 1:0;
assign is_min[81] = (&detect_min[81]) ? 1:0;
assign is_min[82] = (&detect_min[82]) ? 1:0;
assign is_min[83] = (&detect_min[83]) ? 1:0;
assign is_min[84] = (&detect_min[84]) ? 1:0;
assign is_min[85] = (&detect_min[85]) ? 1:0;
assign is_min[86] = (&detect_min[86]) ? 1:0;
assign is_min[87] = (&detect_min[87]) ? 1:0;
assign is_min[88] = (&detect_min[88]) ? 1:0;
assign is_min[89] = (&detect_min[89]) ? 1:0;
assign is_min[90] = (&detect_min[90]) ? 1:0;
assign is_min[91] = (&detect_min[91]) ? 1:0;
assign is_min[92] = (&detect_min[92]) ? 1:0;
assign is_min[93] = (&detect_min[93]) ? 1:0;
assign is_min[94] = (&detect_min[94]) ? 1:0;
assign is_min[95] = (&detect_min[95]) ? 1:0;
assign is_min[96] = (&detect_min[96]) ? 1:0;
assign is_min[97] = (&detect_min[97]) ? 1:0;
assign is_min[98] = (&detect_min[98]) ? 1:0;
assign is_min[99] = (&detect_min[99]) ? 1:0;
assign is_min[100] = (&detect_min[100]) ? 1:0;
assign is_min[101] = (&detect_min[101]) ? 1:0;
assign is_min[102] = (&detect_min[102]) ? 1:0;
assign is_min[103] = (&detect_min[103]) ? 1:0;
assign is_min[104] = (&detect_min[104]) ? 1:0;
assign is_min[105] = (&detect_min[105]) ? 1:0;
assign is_min[106] = (&detect_min[106]) ? 1:0;
assign is_min[107] = (&detect_min[107]) ? 1:0;
assign is_min[108] = (&detect_min[108]) ? 1:0;
assign is_min[109] = (&detect_min[109]) ? 1:0;
assign is_min[110] = (&detect_min[110]) ? 1:0;
assign is_min[111] = (&detect_min[111]) ? 1:0;
assign is_min[112] = (&detect_min[112]) ? 1:0;
assign is_min[113] = (&detect_min[113]) ? 1:0;
assign is_min[114] = (&detect_min[114]) ? 1:0;
assign is_min[115] = (&detect_min[115]) ? 1:0;
assign is_min[116] = (&detect_min[116]) ? 1:0;
assign is_min[117] = (&detect_min[117]) ? 1:0;
assign is_min[118] = (&detect_min[118]) ? 1:0;
assign is_min[119] = (&detect_min[119]) ? 1:0;
assign is_min[120] = (&detect_min[120]) ? 1:0;
assign is_min[121] = (&detect_min[121]) ? 1:0;
assign is_min[122] = (&detect_min[122]) ? 1:0;
assign is_min[123] = (&detect_min[123]) ? 1:0;
assign is_min[124] = (&detect_min[124]) ? 1:0;
assign is_min[125] = (&detect_min[125]) ? 1:0;
assign is_min[126] = (&detect_min[126]) ? 1:0;
assign is_min[127] = (&detect_min[127]) ? 1:0;
assign is_min[128] = (&detect_min[128]) ? 1:0;
assign is_min[129] = (&detect_min[129]) ? 1:0;
assign is_min[130] = (&detect_min[130]) ? 1:0;
assign is_min[131] = (&detect_min[131]) ? 1:0;
assign is_min[132] = (&detect_min[132]) ? 1:0;
assign is_min[133] = (&detect_min[133]) ? 1:0;
assign is_min[134] = (&detect_min[134]) ? 1:0;
assign is_min[135] = (&detect_min[135]) ? 1:0;
assign is_min[136] = (&detect_min[136]) ? 1:0;
assign is_min[137] = (&detect_min[137]) ? 1:0;
assign is_min[138] = (&detect_min[138]) ? 1:0;
assign is_min[139] = (&detect_min[139]) ? 1:0;
assign is_min[140] = (&detect_min[140]) ? 1:0;
assign is_min[141] = (&detect_min[141]) ? 1:0;
assign is_min[142] = (&detect_min[142]) ? 1:0;
assign is_min[143] = (&detect_min[143]) ? 1:0;
assign is_min[144] = (&detect_min[144]) ? 1:0;
assign is_min[145] = (&detect_min[145]) ? 1:0;
assign is_min[146] = (&detect_min[146]) ? 1:0;
assign is_min[147] = (&detect_min[147]) ? 1:0;
assign is_min[148] = (&detect_min[148]) ? 1:0;
assign is_min[149] = (&detect_min[149]) ? 1:0;
assign is_min[150] = (&detect_min[150]) ? 1:0;
assign is_min[151] = (&detect_min[151]) ? 1:0;
assign is_min[152] = (&detect_min[152]) ? 1:0;
assign is_min[153] = (&detect_min[153]) ? 1:0;
assign is_min[154] = (&detect_min[154]) ? 1:0;
assign is_min[155] = (&detect_min[155]) ? 1:0;
assign is_min[156] = (&detect_min[156]) ? 1:0;
assign is_min[157] = (&detect_min[157]) ? 1:0;
assign is_min[158] = (&detect_min[158]) ? 1:0;
assign is_min[159] = (&detect_min[159]) ? 1:0;
assign is_min[160] = (&detect_min[160]) ? 1:0;
assign is_min[161] = (&detect_min[161]) ? 1:0;
assign is_min[162] = (&detect_min[162]) ? 1:0;
assign is_min[163] = (&detect_min[163]) ? 1:0;
assign is_min[164] = (&detect_min[164]) ? 1:0;
assign is_min[165] = (&detect_min[165]) ? 1:0;
assign is_min[166] = (&detect_min[166]) ? 1:0;
assign is_min[167] = (&detect_min[167]) ? 1:0;
assign is_min[168] = (&detect_min[168]) ? 1:0;
assign is_min[169] = (&detect_min[169]) ? 1:0;
assign is_min[170] = (&detect_min[170]) ? 1:0;
assign is_min[171] = (&detect_min[171]) ? 1:0;
assign is_min[172] = (&detect_min[172]) ? 1:0;
assign is_min[173] = (&detect_min[173]) ? 1:0;
assign is_min[174] = (&detect_min[174]) ? 1:0;
assign is_min[175] = (&detect_min[175]) ? 1:0;
assign is_min[176] = (&detect_min[176]) ? 1:0;
assign is_min[177] = (&detect_min[177]) ? 1:0;
assign is_min[178] = (&detect_min[178]) ? 1:0;
assign is_min[179] = (&detect_min[179]) ? 1:0;
assign is_min[180] = (&detect_min[180]) ? 1:0;
assign is_min[181] = (&detect_min[181]) ? 1:0;
assign is_min[182] = (&detect_min[182]) ? 1:0;
assign is_min[183] = (&detect_min[183]) ? 1:0;
assign is_min[184] = (&detect_min[184]) ? 1:0;
assign is_min[185] = (&detect_min[185]) ? 1:0;
assign is_min[186] = (&detect_min[186]) ? 1:0;
assign is_min[187] = (&detect_min[187]) ? 1:0;
assign is_min[188] = (&detect_min[188]) ? 1:0;
assign is_min[189] = (&detect_min[189]) ? 1:0;
assign is_min[190] = (&detect_min[190]) ? 1:0;
assign is_min[191] = (&detect_min[191]) ? 1:0;
assign is_min[192] = (&detect_min[192]) ? 1:0;
assign is_min[193] = (&detect_min[193]) ? 1:0;
assign is_min[194] = (&detect_min[194]) ? 1:0;
assign is_min[195] = (&detect_min[195]) ? 1:0;
assign is_min[196] = (&detect_min[196]) ? 1:0;
assign is_min[197] = (&detect_min[197]) ? 1:0;
assign is_min[198] = (&detect_min[198]) ? 1:0;
assign is_min[199] = (&detect_min[199]) ? 1:0;
assign is_min[200] = (&detect_min[200]) ? 1:0;
assign is_min[201] = (&detect_min[201]) ? 1:0;
assign is_min[202] = (&detect_min[202]) ? 1:0;
assign is_min[203] = (&detect_min[203]) ? 1:0;
assign is_min[204] = (&detect_min[204]) ? 1:0;
assign is_min[205] = (&detect_min[205]) ? 1:0;
assign is_min[206] = (&detect_min[206]) ? 1:0;
assign is_min[207] = (&detect_min[207]) ? 1:0;
assign is_min[208] = (&detect_min[208]) ? 1:0;
assign is_min[209] = (&detect_min[209]) ? 1:0;
assign is_min[210] = (&detect_min[210]) ? 1:0;
assign is_min[211] = (&detect_min[211]) ? 1:0;
assign is_min[212] = (&detect_min[212]) ? 1:0;
assign is_min[213] = (&detect_min[213]) ? 1:0;
assign is_min[214] = (&detect_min[214]) ? 1:0;
assign is_min[215] = (&detect_min[215]) ? 1:0;
assign is_min[216] = (&detect_min[216]) ? 1:0;
assign is_min[217] = (&detect_min[217]) ? 1:0;
assign is_min[218] = (&detect_min[218]) ? 1:0;
assign is_min[219] = (&detect_min[219]) ? 1:0;
assign is_min[220] = (&detect_min[220]) ? 1:0;
assign is_min[221] = (&detect_min[221]) ? 1:0;
assign is_min[222] = (&detect_min[222]) ? 1:0;
assign is_min[223] = (&detect_min[223]) ? 1:0;
assign is_min[224] = (&detect_min[224]) ? 1:0;
assign is_min[225] = (&detect_min[225]) ? 1:0;
assign is_min[226] = (&detect_min[226]) ? 1:0;
assign is_min[227] = (&detect_min[227]) ? 1:0;
assign is_min[228] = (&detect_min[228]) ? 1:0;
assign is_min[229] = (&detect_min[229]) ? 1:0;
assign is_min[230] = (&detect_min[230]) ? 1:0;
assign is_min[231] = (&detect_min[231]) ? 1:0;
assign is_min[232] = (&detect_min[232]) ? 1:0;
assign is_min[233] = (&detect_min[233]) ? 1:0;
assign is_min[234] = (&detect_min[234]) ? 1:0;
assign is_min[235] = (&detect_min[235]) ? 1:0;
assign is_min[236] = (&detect_min[236]) ? 1:0;
assign is_min[237] = (&detect_min[237]) ? 1:0;
assign is_min[238] = (&detect_min[238]) ? 1:0;
assign is_min[239] = (&detect_min[239]) ? 1:0;
assign is_min[240] = (&detect_min[240]) ? 1:0;
assign is_min[241] = (&detect_min[241]) ? 1:0;
assign is_min[242] = (&detect_min[242]) ? 1:0;
assign is_min[243] = (&detect_min[243]) ? 1:0;
assign is_min[244] = (&detect_min[244]) ? 1:0;
assign is_min[245] = (&detect_min[245]) ? 1:0;
assign is_min[246] = (&detect_min[246]) ? 1:0;
assign is_min[247] = (&detect_min[247]) ? 1:0;
assign is_min[248] = (&detect_min[248]) ? 1:0;
assign is_min[249] = (&detect_min[249]) ? 1:0;
assign is_min[250] = (&detect_min[250]) ? 1:0;
assign is_min[251] = (&detect_min[251]) ? 1:0;
assign is_min[252] = (&detect_min[252]) ? 1:0;
assign is_min[253] = (&detect_min[253]) ? 1:0;
assign is_min[254] = (&detect_min[254]) ? 1:0;
assign is_min[255] = (&detect_min[255]) ? 1:0;
assign is_min[256] = (&detect_min[256]) ? 1:0;
assign is_min[257] = (&detect_min[257]) ? 1:0;
assign is_min[258] = (&detect_min[258]) ? 1:0;
assign is_min[259] = (&detect_min[259]) ? 1:0;
assign is_min[260] = (&detect_min[260]) ? 1:0;
assign is_min[261] = (&detect_min[261]) ? 1:0;
assign is_min[262] = (&detect_min[262]) ? 1:0;
assign is_min[263] = (&detect_min[263]) ? 1:0;
assign is_min[264] = (&detect_min[264]) ? 1:0;
assign is_min[265] = (&detect_min[265]) ? 1:0;
assign is_min[266] = (&detect_min[266]) ? 1:0;
assign is_min[267] = (&detect_min[267]) ? 1:0;
assign is_min[268] = (&detect_min[268]) ? 1:0;
assign is_min[269] = (&detect_min[269]) ? 1:0;
assign is_min[270] = (&detect_min[270]) ? 1:0;
assign is_min[271] = (&detect_min[271]) ? 1:0;
assign is_min[272] = (&detect_min[272]) ? 1:0;
assign is_min[273] = (&detect_min[273]) ? 1:0;
assign is_min[274] = (&detect_min[274]) ? 1:0;
assign is_min[275] = (&detect_min[275]) ? 1:0;
assign is_min[276] = (&detect_min[276]) ? 1:0;
assign is_min[277] = (&detect_min[277]) ? 1:0;
assign is_min[278] = (&detect_min[278]) ? 1:0;
assign is_min[279] = (&detect_min[279]) ? 1:0;
assign is_min[280] = (&detect_min[280]) ? 1:0;
assign is_min[281] = (&detect_min[281]) ? 1:0;
assign is_min[282] = (&detect_min[282]) ? 1:0;
assign is_min[283] = (&detect_min[283]) ? 1:0;
assign is_min[284] = (&detect_min[284]) ? 1:0;
assign is_min[285] = (&detect_min[285]) ? 1:0;
assign is_min[286] = (&detect_min[286]) ? 1:0;
assign is_min[287] = (&detect_min[287]) ? 1:0;
assign is_min[288] = (&detect_min[288]) ? 1:0;
assign is_min[289] = (&detect_min[289]) ? 1:0;
assign is_min[290] = (&detect_min[290]) ? 1:0;
assign is_min[291] = (&detect_min[291]) ? 1:0;
assign is_min[292] = (&detect_min[292]) ? 1:0;
assign is_min[293] = (&detect_min[293]) ? 1:0;
assign is_min[294] = (&detect_min[294]) ? 1:0;
assign is_min[295] = (&detect_min[295]) ? 1:0;
assign is_min[296] = (&detect_min[296]) ? 1:0;
assign is_min[297] = (&detect_min[297]) ? 1:0;
assign is_min[298] = (&detect_min[298]) ? 1:0;
assign is_min[299] = (&detect_min[299]) ? 1:0;
assign is_min[300] = (&detect_min[300]) ? 1:0;
assign is_min[301] = (&detect_min[301]) ? 1:0;
assign is_min[302] = (&detect_min[302]) ? 1:0;
assign is_min[303] = (&detect_min[303]) ? 1:0;
assign is_min[304] = (&detect_min[304]) ? 1:0;
assign is_min[305] = (&detect_min[305]) ? 1:0;
assign is_min[306] = (&detect_min[306]) ? 1:0;
assign is_min[307] = (&detect_min[307]) ? 1:0;
assign is_min[308] = (&detect_min[308]) ? 1:0;
assign is_min[309] = (&detect_min[309]) ? 1:0;
assign is_min[310] = (&detect_min[310]) ? 1:0;
assign is_min[311] = (&detect_min[311]) ? 1:0;
assign is_min[312] = (&detect_min[312]) ? 1:0;
assign is_min[313] = (&detect_min[313]) ? 1:0;
assign is_min[314] = (&detect_min[314]) ? 1:0;
assign is_min[315] = (&detect_min[315]) ? 1:0;
assign is_min[316] = (&detect_min[316]) ? 1:0;
assign is_min[317] = (&detect_min[317]) ? 1:0;
assign is_min[318] = (&detect_min[318]) ? 1:0;
assign is_min[319] = (&detect_min[319]) ? 1:0;
assign is_min[320] = (&detect_min[320]) ? 1:0;
assign is_min[321] = (&detect_min[321]) ? 1:0;
assign is_min[322] = (&detect_min[322]) ? 1:0;
assign is_min[323] = (&detect_min[323]) ? 1:0;
assign is_min[324] = (&detect_min[324]) ? 1:0;
assign is_min[325] = (&detect_min[325]) ? 1:0;
assign is_min[326] = (&detect_min[326]) ? 1:0;
assign is_min[327] = (&detect_min[327]) ? 1:0;
assign is_min[328] = (&detect_min[328]) ? 1:0;
assign is_min[329] = (&detect_min[329]) ? 1:0;
assign is_min[330] = (&detect_min[330]) ? 1:0;
assign is_min[331] = (&detect_min[331]) ? 1:0;
assign is_min[332] = (&detect_min[332]) ? 1:0;
assign is_min[333] = (&detect_min[333]) ? 1:0;
assign is_min[334] = (&detect_min[334]) ? 1:0;
assign is_min[335] = (&detect_min[335]) ? 1:0;
assign is_min[336] = (&detect_min[336]) ? 1:0;
assign is_min[337] = (&detect_min[337]) ? 1:0;
assign is_min[338] = (&detect_min[338]) ? 1:0;
assign is_min[339] = (&detect_min[339]) ? 1:0;
assign is_min[340] = (&detect_min[340]) ? 1:0;
assign is_min[341] = (&detect_min[341]) ? 1:0;
assign is_min[342] = (&detect_min[342]) ? 1:0;
assign is_min[343] = (&detect_min[343]) ? 1:0;
assign is_min[344] = (&detect_min[344]) ? 1:0;
assign is_min[345] = (&detect_min[345]) ? 1:0;
assign is_min[346] = (&detect_min[346]) ? 1:0;
assign is_min[347] = (&detect_min[347]) ? 1:0;
assign is_min[348] = (&detect_min[348]) ? 1:0;
assign is_min[349] = (&detect_min[349]) ? 1:0;
assign is_min[350] = (&detect_min[350]) ? 1:0;
assign is_min[351] = (&detect_min[351]) ? 1:0;
assign is_min[352] = (&detect_min[352]) ? 1:0;
assign is_min[353] = (&detect_min[353]) ? 1:0;
assign is_min[354] = (&detect_min[354]) ? 1:0;
assign is_min[355] = (&detect_min[355]) ? 1:0;
assign is_min[356] = (&detect_min[356]) ? 1:0;
assign is_min[357] = (&detect_min[357]) ? 1:0;
assign is_min[358] = (&detect_min[358]) ? 1:0;
assign is_min[359] = (&detect_min[359]) ? 1:0;
assign is_min[360] = (&detect_min[360]) ? 1:0;
assign is_min[361] = (&detect_min[361]) ? 1:0;
assign is_min[362] = (&detect_min[362]) ? 1:0;
assign is_min[363] = (&detect_min[363]) ? 1:0;
assign is_min[364] = (&detect_min[364]) ? 1:0;
assign is_min[365] = (&detect_min[365]) ? 1:0;
assign is_min[366] = (&detect_min[366]) ? 1:0;
assign is_min[367] = (&detect_min[367]) ? 1:0;
assign is_min[368] = (&detect_min[368]) ? 1:0;
assign is_min[369] = (&detect_min[369]) ? 1:0;
assign is_min[370] = (&detect_min[370]) ? 1:0;
assign is_min[371] = (&detect_min[371]) ? 1:0;
assign is_min[372] = (&detect_min[372]) ? 1:0;
assign is_min[373] = (&detect_min[373]) ? 1:0;
assign is_min[374] = (&detect_min[374]) ? 1:0;
assign is_min[375] = (&detect_min[375]) ? 1:0;
assign is_min[376] = (&detect_min[376]) ? 1:0;
assign is_min[377] = (&detect_min[377]) ? 1:0;
assign is_min[378] = (&detect_min[378]) ? 1:0;
assign is_min[379] = (&detect_min[379]) ? 1:0;
assign is_min[380] = (&detect_min[380]) ? 1:0;
assign is_min[381] = (&detect_min[381]) ? 1:0;
assign is_min[382] = (&detect_min[382]) ? 1:0;
assign is_min[383] = (&detect_min[383]) ? 1:0;
assign is_min[384] = (&detect_min[384]) ? 1:0;
assign is_min[385] = (&detect_min[385]) ? 1:0;
assign is_min[386] = (&detect_min[386]) ? 1:0;
assign is_min[387] = (&detect_min[387]) ? 1:0;
assign is_min[388] = (&detect_min[388]) ? 1:0;
assign is_min[389] = (&detect_min[389]) ? 1:0;
assign is_min[390] = (&detect_min[390]) ? 1:0;
assign is_min[391] = (&detect_min[391]) ? 1:0;
assign is_min[392] = (&detect_min[392]) ? 1:0;
assign is_min[393] = (&detect_min[393]) ? 1:0;
assign is_min[394] = (&detect_min[394]) ? 1:0;
assign is_min[395] = (&detect_min[395]) ? 1:0;
assign is_min[396] = (&detect_min[396]) ? 1:0;
assign is_min[397] = (&detect_min[397]) ? 1:0;
assign is_min[398] = (&detect_min[398]) ? 1:0;
assign is_min[399] = (&detect_min[399]) ? 1:0;
assign is_min[400] = (&detect_min[400]) ? 1:0;
assign is_min[401] = (&detect_min[401]) ? 1:0;
assign is_min[402] = (&detect_min[402]) ? 1:0;
assign is_min[403] = (&detect_min[403]) ? 1:0;
assign is_min[404] = (&detect_min[404]) ? 1:0;
assign is_min[405] = (&detect_min[405]) ? 1:0;
assign is_min[406] = (&detect_min[406]) ? 1:0;
assign is_min[407] = (&detect_min[407]) ? 1:0;
assign is_min[408] = (&detect_min[408]) ? 1:0;
assign is_min[409] = (&detect_min[409]) ? 1:0;
assign is_min[410] = (&detect_min[410]) ? 1:0;
assign is_min[411] = (&detect_min[411]) ? 1:0;
assign is_min[412] = (&detect_min[412]) ? 1:0;
assign is_min[413] = (&detect_min[413]) ? 1:0;
assign is_min[414] = (&detect_min[414]) ? 1:0;
assign is_min[415] = (&detect_min[415]) ? 1:0;
assign is_min[416] = (&detect_min[416]) ? 1:0;
assign is_min[417] = (&detect_min[417]) ? 1:0;
assign is_min[418] = (&detect_min[418]) ? 1:0;
assign is_min[419] = (&detect_min[419]) ? 1:0;
assign is_min[420] = (&detect_min[420]) ? 1:0;
assign is_min[421] = (&detect_min[421]) ? 1:0;
assign is_min[422] = (&detect_min[422]) ? 1:0;
assign is_min[423] = (&detect_min[423]) ? 1:0;
assign is_min[424] = (&detect_min[424]) ? 1:0;
assign is_min[425] = (&detect_min[425]) ? 1:0;
assign is_min[426] = (&detect_min[426]) ? 1:0;
assign is_min[427] = (&detect_min[427]) ? 1:0;
assign is_min[428] = (&detect_min[428]) ? 1:0;
assign is_min[429] = (&detect_min[429]) ? 1:0;
assign is_min[430] = (&detect_min[430]) ? 1:0;
assign is_min[431] = (&detect_min[431]) ? 1:0;
assign is_min[432] = (&detect_min[432]) ? 1:0;
assign is_min[433] = (&detect_min[433]) ? 1:0;
assign is_min[434] = (&detect_min[434]) ? 1:0;
assign is_min[435] = (&detect_min[435]) ? 1:0;
assign is_min[436] = (&detect_min[436]) ? 1:0;
assign is_min[437] = (&detect_min[437]) ? 1:0;
assign is_min[438] = (&detect_min[438]) ? 1:0;
assign is_min[439] = (&detect_min[439]) ? 1:0;
assign is_min[440] = (&detect_min[440]) ? 1:0;
assign is_min[441] = (&detect_min[441]) ? 1:0;
assign is_min[442] = (&detect_min[442]) ? 1:0;
assign is_min[443] = (&detect_min[443]) ? 1:0;
assign is_min[444] = (&detect_min[444]) ? 1:0;
assign is_min[445] = (&detect_min[445]) ? 1:0;
assign is_min[446] = (&detect_min[446]) ? 1:0;
assign is_min[447] = (&detect_min[447]) ? 1:0;
assign is_min[448] = (&detect_min[448]) ? 1:0;
assign is_min[449] = (&detect_min[449]) ? 1:0;
assign is_min[450] = (&detect_min[450]) ? 1:0;
assign is_min[451] = (&detect_min[451]) ? 1:0;
assign is_min[452] = (&detect_min[452]) ? 1:0;
assign is_min[453] = (&detect_min[453]) ? 1:0;
assign is_min[454] = (&detect_min[454]) ? 1:0;
assign is_min[455] = (&detect_min[455]) ? 1:0;
assign is_min[456] = (&detect_min[456]) ? 1:0;
assign is_min[457] = (&detect_min[457]) ? 1:0;
assign is_min[458] = (&detect_min[458]) ? 1:0;
assign is_min[459] = (&detect_min[459]) ? 1:0;
assign is_min[460] = (&detect_min[460]) ? 1:0;
assign is_min[461] = (&detect_min[461]) ? 1:0;
assign is_min[462] = (&detect_min[462]) ? 1:0;
assign is_min[463] = (&detect_min[463]) ? 1:0;
assign is_min[464] = (&detect_min[464]) ? 1:0;
assign is_min[465] = (&detect_min[465]) ? 1:0;
assign is_min[466] = (&detect_min[466]) ? 1:0;
assign is_min[467] = (&detect_min[467]) ? 1:0;
assign is_min[468] = (&detect_min[468]) ? 1:0;
assign is_min[469] = (&detect_min[469]) ? 1:0;
assign is_min[470] = (&detect_min[470]) ? 1:0;
assign is_min[471] = (&detect_min[471]) ? 1:0;
assign is_min[472] = (&detect_min[472]) ? 1:0;
assign is_min[473] = (&detect_min[473]) ? 1:0;
assign is_min[474] = (&detect_min[474]) ? 1:0;
assign is_min[475] = (&detect_min[475]) ? 1:0;
assign is_min[476] = (&detect_min[476]) ? 1:0;
assign is_min[477] = (&detect_min[477]) ? 1:0;
assign is_min[478] = (&detect_min[478]) ? 1:0;
assign is_min[479] = (&detect_min[479]) ? 1:0;
assign is_min[480] = (&detect_min[480]) ? 1:0;
assign is_min[481] = (&detect_min[481]) ? 1:0;
assign is_min[482] = (&detect_min[482]) ? 1:0;
assign is_min[483] = (&detect_min[483]) ? 1:0;
assign is_min[484] = (&detect_min[484]) ? 1:0;
assign is_min[485] = (&detect_min[485]) ? 1:0;
assign is_min[486] = (&detect_min[486]) ? 1:0;
assign is_min[487] = (&detect_min[487]) ? 1:0;
assign is_min[488] = (&detect_min[488]) ? 1:0;
assign is_min[489] = (&detect_min[489]) ? 1:0;
assign is_min[490] = (&detect_min[490]) ? 1:0;
assign is_min[491] = (&detect_min[491]) ? 1:0;
assign is_min[492] = (&detect_min[492]) ? 1:0;
assign is_min[493] = (&detect_min[493]) ? 1:0;
assign is_min[494] = (&detect_min[494]) ? 1:0;
assign is_min[495] = (&detect_min[495]) ? 1:0;
assign is_min[496] = (&detect_min[496]) ? 1:0;
assign is_min[497] = (&detect_min[497]) ? 1:0;
assign is_min[498] = (&detect_min[498]) ? 1:0;
assign is_min[499] = (&detect_min[499]) ? 1:0;
assign is_min[500] = (&detect_min[500]) ? 1:0;
assign is_min[501] = (&detect_min[501]) ? 1:0;
assign is_min[502] = (&detect_min[502]) ? 1:0;
assign is_min[503] = (&detect_min[503]) ? 1:0;
assign is_min[504] = (&detect_min[504]) ? 1:0;
assign is_min[505] = (&detect_min[505]) ? 1:0;
assign is_min[506] = (&detect_min[506]) ? 1:0;
assign is_min[507] = (&detect_min[507]) ? 1:0;
assign is_min[508] = (&detect_min[508]) ? 1:0;
assign is_min[509] = (&detect_min[509]) ? 1:0;
assign is_min[510] = (&detect_min[510]) ? 1:0;
assign is_min[511] = (&detect_min[511]) ? 1:0;
assign is_min[512] = (&detect_min[512]) ? 1:0;
assign is_min[513] = (&detect_min[513]) ? 1:0;
assign is_min[514] = (&detect_min[514]) ? 1:0;
assign is_min[515] = (&detect_min[515]) ? 1:0;
assign is_min[516] = (&detect_min[516]) ? 1:0;
assign is_min[517] = (&detect_min[517]) ? 1:0;
assign is_min[518] = (&detect_min[518]) ? 1:0;
assign is_min[519] = (&detect_min[519]) ? 1:0;
assign is_min[520] = (&detect_min[520]) ? 1:0;
assign is_min[521] = (&detect_min[521]) ? 1:0;
assign is_min[522] = (&detect_min[522]) ? 1:0;
assign is_min[523] = (&detect_min[523]) ? 1:0;
assign is_min[524] = (&detect_min[524]) ? 1:0;
assign is_min[525] = (&detect_min[525]) ? 1:0;
assign is_min[526] = (&detect_min[526]) ? 1:0;
assign is_min[527] = (&detect_min[527]) ? 1:0;
assign is_min[528] = (&detect_min[528]) ? 1:0;
assign is_min[529] = (&detect_min[529]) ? 1:0;
assign is_min[530] = (&detect_min[530]) ? 1:0;
assign is_min[531] = (&detect_min[531]) ? 1:0;
assign is_min[532] = (&detect_min[532]) ? 1:0;
assign is_min[533] = (&detect_min[533]) ? 1:0;
assign is_min[534] = (&detect_min[534]) ? 1:0;
assign is_min[535] = (&detect_min[535]) ? 1:0;
assign is_min[536] = (&detect_min[536]) ? 1:0;
assign is_min[537] = (&detect_min[537]) ? 1:0;
assign is_min[538] = (&detect_min[538]) ? 1:0;
assign is_min[539] = (&detect_min[539]) ? 1:0;
assign is_min[540] = (&detect_min[540]) ? 1:0;
assign is_min[541] = (&detect_min[541]) ? 1:0;
assign is_min[542] = (&detect_min[542]) ? 1:0;
assign is_min[543] = (&detect_min[543]) ? 1:0;
assign is_min[544] = (&detect_min[544]) ? 1:0;
assign is_min[545] = (&detect_min[545]) ? 1:0;
assign is_min[546] = (&detect_min[546]) ? 1:0;
assign is_min[547] = (&detect_min[547]) ? 1:0;
assign is_min[548] = (&detect_min[548]) ? 1:0;
assign is_min[549] = (&detect_min[549]) ? 1:0;
assign is_min[550] = (&detect_min[550]) ? 1:0;
assign is_min[551] = (&detect_min[551]) ? 1:0;
assign is_min[552] = (&detect_min[552]) ? 1:0;
assign is_min[553] = (&detect_min[553]) ? 1:0;
assign is_min[554] = (&detect_min[554]) ? 1:0;
assign is_min[555] = (&detect_min[555]) ? 1:0;
assign is_min[556] = (&detect_min[556]) ? 1:0;
assign is_min[557] = (&detect_min[557]) ? 1:0;
assign is_min[558] = (&detect_min[558]) ? 1:0;
assign is_min[559] = (&detect_min[559]) ? 1:0;
assign is_min[560] = (&detect_min[560]) ? 1:0;
assign is_min[561] = (&detect_min[561]) ? 1:0;
assign is_min[562] = (&detect_min[562]) ? 1:0;
assign is_min[563] = (&detect_min[563]) ? 1:0;
assign is_min[564] = (&detect_min[564]) ? 1:0;
assign is_min[565] = (&detect_min[565]) ? 1:0;
assign is_min[566] = (&detect_min[566]) ? 1:0;
assign is_min[567] = (&detect_min[567]) ? 1:0;
assign is_min[568] = (&detect_min[568]) ? 1:0;
assign is_min[569] = (&detect_min[569]) ? 1:0;
assign is_min[570] = (&detect_min[570]) ? 1:0;
assign is_min[571] = (&detect_min[571]) ? 1:0;
assign is_min[572] = (&detect_min[572]) ? 1:0;
assign is_min[573] = (&detect_min[573]) ? 1:0;
assign is_min[574] = (&detect_min[574]) ? 1:0;
assign is_min[575] = (&detect_min[575]) ? 1:0;
assign is_min[576] = (&detect_min[576]) ? 1:0;
assign is_min[577] = (&detect_min[577]) ? 1:0;
assign is_min[578] = (&detect_min[578]) ? 1:0;
assign is_min[579] = (&detect_min[579]) ? 1:0;
assign is_min[580] = (&detect_min[580]) ? 1:0;
assign is_min[581] = (&detect_min[581]) ? 1:0;
assign is_min[582] = (&detect_min[582]) ? 1:0;
assign is_min[583] = (&detect_min[583]) ? 1:0;
assign is_min[584] = (&detect_min[584]) ? 1:0;
assign is_min[585] = (&detect_min[585]) ? 1:0;
assign is_min[586] = (&detect_min[586]) ? 1:0;
assign is_min[587] = (&detect_min[587]) ? 1:0;
assign is_min[588] = (&detect_min[588]) ? 1:0;
assign is_min[589] = (&detect_min[589]) ? 1:0;
assign is_min[590] = (&detect_min[590]) ? 1:0;
assign is_min[591] = (&detect_min[591]) ? 1:0;
assign is_min[592] = (&detect_min[592]) ? 1:0;
assign is_min[593] = (&detect_min[593]) ? 1:0;
assign is_min[594] = (&detect_min[594]) ? 1:0;
assign is_min[595] = (&detect_min[595]) ? 1:0;
assign is_min[596] = (&detect_min[596]) ? 1:0;
assign is_min[597] = (&detect_min[597]) ? 1:0;
assign is_min[598] = (&detect_min[598]) ? 1:0;
assign is_min[599] = (&detect_min[599]) ? 1:0;
assign is_min[600] = (&detect_min[600]) ? 1:0;
assign is_min[601] = (&detect_min[601]) ? 1:0;
assign is_min[602] = (&detect_min[602]) ? 1:0;
assign is_min[603] = (&detect_min[603]) ? 1:0;
assign is_min[604] = (&detect_min[604]) ? 1:0;
assign is_min[605] = (&detect_min[605]) ? 1:0;
assign is_min[606] = (&detect_min[606]) ? 1:0;
assign is_min[607] = (&detect_min[607]) ? 1:0;
assign is_min[608] = (&detect_min[608]) ? 1:0;
assign is_min[609] = (&detect_min[609]) ? 1:0;
assign is_min[610] = (&detect_min[610]) ? 1:0;
assign is_min[611] = (&detect_min[611]) ? 1:0;
assign is_min[612] = (&detect_min[612]) ? 1:0;
assign is_min[613] = (&detect_min[613]) ? 1:0;
assign is_min[614] = (&detect_min[614]) ? 1:0;
assign is_min[615] = (&detect_min[615]) ? 1:0;
assign is_min[616] = (&detect_min[616]) ? 1:0;
assign is_min[617] = (&detect_min[617]) ? 1:0;
assign is_min[618] = (&detect_min[618]) ? 1:0;
assign is_min[619] = (&detect_min[619]) ? 1:0;
assign is_min[620] = (&detect_min[620]) ? 1:0;
assign is_min[621] = (&detect_min[621]) ? 1:0;
assign is_min[622] = (&detect_min[622]) ? 1:0;
assign is_min[623] = (&detect_min[623]) ? 1:0;
assign is_min[624] = (&detect_min[624]) ? 1:0;
assign is_min[625] = (&detect_min[625]) ? 1:0;
assign is_min[626] = (&detect_min[626]) ? 1:0;
assign is_min[627] = (&detect_min[627]) ? 1:0;
assign is_min[628] = (&detect_min[628]) ? 1:0;
assign is_min[629] = (&detect_min[629]) ? 1:0;
assign is_min[630] = (&detect_min[630]) ? 1:0;
assign is_min[631] = (&detect_min[631]) ? 1:0;
assign is_min[632] = (&detect_min[632]) ? 1:0;
assign is_min[633] = (&detect_min[633]) ? 1:0;
assign is_min[634] = (&detect_min[634]) ? 1:0;
assign is_min[635] = (&detect_min[635]) ? 1:0;
assign is_min[636] = (&detect_min[636]) ? 1:0;
assign is_min[637] = (&detect_min[637]) ? 1:0;

assign is_keypoint[0] = is_max[0] | is_min[0];
assign is_keypoint[1] = is_max[1] | is_min[1];
assign is_keypoint[2] = is_max[2] | is_min[2];
assign is_keypoint[3] = is_max[3] | is_min[3];
assign is_keypoint[4] = is_max[4] | is_min[4];
assign is_keypoint[5] = is_max[5] | is_min[5];
assign is_keypoint[6] = is_max[6] | is_min[6];
assign is_keypoint[7] = is_max[7] | is_min[7];
assign is_keypoint[8] = is_max[8] | is_min[8];
assign is_keypoint[9] = is_max[9] | is_min[9];
assign is_keypoint[10] = is_max[10] | is_min[10];
assign is_keypoint[11] = is_max[11] | is_min[11];
assign is_keypoint[12] = is_max[12] | is_min[12];
assign is_keypoint[13] = is_max[13] | is_min[13];
assign is_keypoint[14] = is_max[14] | is_min[14];
assign is_keypoint[15] = is_max[15] | is_min[15];
assign is_keypoint[16] = is_max[16] | is_min[16];
assign is_keypoint[17] = is_max[17] | is_min[17];
assign is_keypoint[18] = is_max[18] | is_min[18];
assign is_keypoint[19] = is_max[19] | is_min[19];
assign is_keypoint[20] = is_max[20] | is_min[20];
assign is_keypoint[21] = is_max[21] | is_min[21];
assign is_keypoint[22] = is_max[22] | is_min[22];
assign is_keypoint[23] = is_max[23] | is_min[23];
assign is_keypoint[24] = is_max[24] | is_min[24];
assign is_keypoint[25] = is_max[25] | is_min[25];
assign is_keypoint[26] = is_max[26] | is_min[26];
assign is_keypoint[27] = is_max[27] | is_min[27];
assign is_keypoint[28] = is_max[28] | is_min[28];
assign is_keypoint[29] = is_max[29] | is_min[29];
assign is_keypoint[30] = is_max[30] | is_min[30];
assign is_keypoint[31] = is_max[31] | is_min[31];
assign is_keypoint[32] = is_max[32] | is_min[32];
assign is_keypoint[33] = is_max[33] | is_min[33];
assign is_keypoint[34] = is_max[34] | is_min[34];
assign is_keypoint[35] = is_max[35] | is_min[35];
assign is_keypoint[36] = is_max[36] | is_min[36];
assign is_keypoint[37] = is_max[37] | is_min[37];
assign is_keypoint[38] = is_max[38] | is_min[38];
assign is_keypoint[39] = is_max[39] | is_min[39];
assign is_keypoint[40] = is_max[40] | is_min[40];
assign is_keypoint[41] = is_max[41] | is_min[41];
assign is_keypoint[42] = is_max[42] | is_min[42];
assign is_keypoint[43] = is_max[43] | is_min[43];
assign is_keypoint[44] = is_max[44] | is_min[44];
assign is_keypoint[45] = is_max[45] | is_min[45];
assign is_keypoint[46] = is_max[46] | is_min[46];
assign is_keypoint[47] = is_max[47] | is_min[47];
assign is_keypoint[48] = is_max[48] | is_min[48];
assign is_keypoint[49] = is_max[49] | is_min[49];
assign is_keypoint[50] = is_max[50] | is_min[50];
assign is_keypoint[51] = is_max[51] | is_min[51];
assign is_keypoint[52] = is_max[52] | is_min[52];
assign is_keypoint[53] = is_max[53] | is_min[53];
assign is_keypoint[54] = is_max[54] | is_min[54];
assign is_keypoint[55] = is_max[55] | is_min[55];
assign is_keypoint[56] = is_max[56] | is_min[56];
assign is_keypoint[57] = is_max[57] | is_min[57];
assign is_keypoint[58] = is_max[58] | is_min[58];
assign is_keypoint[59] = is_max[59] | is_min[59];
assign is_keypoint[60] = is_max[60] | is_min[60];
assign is_keypoint[61] = is_max[61] | is_min[61];
assign is_keypoint[62] = is_max[62] | is_min[62];
assign is_keypoint[63] = is_max[63] | is_min[63];
assign is_keypoint[64] = is_max[64] | is_min[64];
assign is_keypoint[65] = is_max[65] | is_min[65];
assign is_keypoint[66] = is_max[66] | is_min[66];
assign is_keypoint[67] = is_max[67] | is_min[67];
assign is_keypoint[68] = is_max[68] | is_min[68];
assign is_keypoint[69] = is_max[69] | is_min[69];
assign is_keypoint[70] = is_max[70] | is_min[70];
assign is_keypoint[71] = is_max[71] | is_min[71];
assign is_keypoint[72] = is_max[72] | is_min[72];
assign is_keypoint[73] = is_max[73] | is_min[73];
assign is_keypoint[74] = is_max[74] | is_min[74];
assign is_keypoint[75] = is_max[75] | is_min[75];
assign is_keypoint[76] = is_max[76] | is_min[76];
assign is_keypoint[77] = is_max[77] | is_min[77];
assign is_keypoint[78] = is_max[78] | is_min[78];
assign is_keypoint[79] = is_max[79] | is_min[79];
assign is_keypoint[80] = is_max[80] | is_min[80];
assign is_keypoint[81] = is_max[81] | is_min[81];
assign is_keypoint[82] = is_max[82] | is_min[82];
assign is_keypoint[83] = is_max[83] | is_min[83];
assign is_keypoint[84] = is_max[84] | is_min[84];
assign is_keypoint[85] = is_max[85] | is_min[85];
assign is_keypoint[86] = is_max[86] | is_min[86];
assign is_keypoint[87] = is_max[87] | is_min[87];
assign is_keypoint[88] = is_max[88] | is_min[88];
assign is_keypoint[89] = is_max[89] | is_min[89];
assign is_keypoint[90] = is_max[90] | is_min[90];
assign is_keypoint[91] = is_max[91] | is_min[91];
assign is_keypoint[92] = is_max[92] | is_min[92];
assign is_keypoint[93] = is_max[93] | is_min[93];
assign is_keypoint[94] = is_max[94] | is_min[94];
assign is_keypoint[95] = is_max[95] | is_min[95];
assign is_keypoint[96] = is_max[96] | is_min[96];
assign is_keypoint[97] = is_max[97] | is_min[97];
assign is_keypoint[98] = is_max[98] | is_min[98];
assign is_keypoint[99] = is_max[99] | is_min[99];
assign is_keypoint[100] = is_max[100] | is_min[100];
assign is_keypoint[101] = is_max[101] | is_min[101];
assign is_keypoint[102] = is_max[102] | is_min[102];
assign is_keypoint[103] = is_max[103] | is_min[103];
assign is_keypoint[104] = is_max[104] | is_min[104];
assign is_keypoint[105] = is_max[105] | is_min[105];
assign is_keypoint[106] = is_max[106] | is_min[106];
assign is_keypoint[107] = is_max[107] | is_min[107];
assign is_keypoint[108] = is_max[108] | is_min[108];
assign is_keypoint[109] = is_max[109] | is_min[109];
assign is_keypoint[110] = is_max[110] | is_min[110];
assign is_keypoint[111] = is_max[111] | is_min[111];
assign is_keypoint[112] = is_max[112] | is_min[112];
assign is_keypoint[113] = is_max[113] | is_min[113];
assign is_keypoint[114] = is_max[114] | is_min[114];
assign is_keypoint[115] = is_max[115] | is_min[115];
assign is_keypoint[116] = is_max[116] | is_min[116];
assign is_keypoint[117] = is_max[117] | is_min[117];
assign is_keypoint[118] = is_max[118] | is_min[118];
assign is_keypoint[119] = is_max[119] | is_min[119];
assign is_keypoint[120] = is_max[120] | is_min[120];
assign is_keypoint[121] = is_max[121] | is_min[121];
assign is_keypoint[122] = is_max[122] | is_min[122];
assign is_keypoint[123] = is_max[123] | is_min[123];
assign is_keypoint[124] = is_max[124] | is_min[124];
assign is_keypoint[125] = is_max[125] | is_min[125];
assign is_keypoint[126] = is_max[126] | is_min[126];
assign is_keypoint[127] = is_max[127] | is_min[127];
assign is_keypoint[128] = is_max[128] | is_min[128];
assign is_keypoint[129] = is_max[129] | is_min[129];
assign is_keypoint[130] = is_max[130] | is_min[130];
assign is_keypoint[131] = is_max[131] | is_min[131];
assign is_keypoint[132] = is_max[132] | is_min[132];
assign is_keypoint[133] = is_max[133] | is_min[133];
assign is_keypoint[134] = is_max[134] | is_min[134];
assign is_keypoint[135] = is_max[135] | is_min[135];
assign is_keypoint[136] = is_max[136] | is_min[136];
assign is_keypoint[137] = is_max[137] | is_min[137];
assign is_keypoint[138] = is_max[138] | is_min[138];
assign is_keypoint[139] = is_max[139] | is_min[139];
assign is_keypoint[140] = is_max[140] | is_min[140];
assign is_keypoint[141] = is_max[141] | is_min[141];
assign is_keypoint[142] = is_max[142] | is_min[142];
assign is_keypoint[143] = is_max[143] | is_min[143];
assign is_keypoint[144] = is_max[144] | is_min[144];
assign is_keypoint[145] = is_max[145] | is_min[145];
assign is_keypoint[146] = is_max[146] | is_min[146];
assign is_keypoint[147] = is_max[147] | is_min[147];
assign is_keypoint[148] = is_max[148] | is_min[148];
assign is_keypoint[149] = is_max[149] | is_min[149];
assign is_keypoint[150] = is_max[150] | is_min[150];
assign is_keypoint[151] = is_max[151] | is_min[151];
assign is_keypoint[152] = is_max[152] | is_min[152];
assign is_keypoint[153] = is_max[153] | is_min[153];
assign is_keypoint[154] = is_max[154] | is_min[154];
assign is_keypoint[155] = is_max[155] | is_min[155];
assign is_keypoint[156] = is_max[156] | is_min[156];
assign is_keypoint[157] = is_max[157] | is_min[157];
assign is_keypoint[158] = is_max[158] | is_min[158];
assign is_keypoint[159] = is_max[159] | is_min[159];
assign is_keypoint[160] = is_max[160] | is_min[160];
assign is_keypoint[161] = is_max[161] | is_min[161];
assign is_keypoint[162] = is_max[162] | is_min[162];
assign is_keypoint[163] = is_max[163] | is_min[163];
assign is_keypoint[164] = is_max[164] | is_min[164];
assign is_keypoint[165] = is_max[165] | is_min[165];
assign is_keypoint[166] = is_max[166] | is_min[166];
assign is_keypoint[167] = is_max[167] | is_min[167];
assign is_keypoint[168] = is_max[168] | is_min[168];
assign is_keypoint[169] = is_max[169] | is_min[169];
assign is_keypoint[170] = is_max[170] | is_min[170];
assign is_keypoint[171] = is_max[171] | is_min[171];
assign is_keypoint[172] = is_max[172] | is_min[172];
assign is_keypoint[173] = is_max[173] | is_min[173];
assign is_keypoint[174] = is_max[174] | is_min[174];
assign is_keypoint[175] = is_max[175] | is_min[175];
assign is_keypoint[176] = is_max[176] | is_min[176];
assign is_keypoint[177] = is_max[177] | is_min[177];
assign is_keypoint[178] = is_max[178] | is_min[178];
assign is_keypoint[179] = is_max[179] | is_min[179];
assign is_keypoint[180] = is_max[180] | is_min[180];
assign is_keypoint[181] = is_max[181] | is_min[181];
assign is_keypoint[182] = is_max[182] | is_min[182];
assign is_keypoint[183] = is_max[183] | is_min[183];
assign is_keypoint[184] = is_max[184] | is_min[184];
assign is_keypoint[185] = is_max[185] | is_min[185];
assign is_keypoint[186] = is_max[186] | is_min[186];
assign is_keypoint[187] = is_max[187] | is_min[187];
assign is_keypoint[188] = is_max[188] | is_min[188];
assign is_keypoint[189] = is_max[189] | is_min[189];
assign is_keypoint[190] = is_max[190] | is_min[190];
assign is_keypoint[191] = is_max[191] | is_min[191];
assign is_keypoint[192] = is_max[192] | is_min[192];
assign is_keypoint[193] = is_max[193] | is_min[193];
assign is_keypoint[194] = is_max[194] | is_min[194];
assign is_keypoint[195] = is_max[195] | is_min[195];
assign is_keypoint[196] = is_max[196] | is_min[196];
assign is_keypoint[197] = is_max[197] | is_min[197];
assign is_keypoint[198] = is_max[198] | is_min[198];
assign is_keypoint[199] = is_max[199] | is_min[199];
assign is_keypoint[200] = is_max[200] | is_min[200];
assign is_keypoint[201] = is_max[201] | is_min[201];
assign is_keypoint[202] = is_max[202] | is_min[202];
assign is_keypoint[203] = is_max[203] | is_min[203];
assign is_keypoint[204] = is_max[204] | is_min[204];
assign is_keypoint[205] = is_max[205] | is_min[205];
assign is_keypoint[206] = is_max[206] | is_min[206];
assign is_keypoint[207] = is_max[207] | is_min[207];
assign is_keypoint[208] = is_max[208] | is_min[208];
assign is_keypoint[209] = is_max[209] | is_min[209];
assign is_keypoint[210] = is_max[210] | is_min[210];
assign is_keypoint[211] = is_max[211] | is_min[211];
assign is_keypoint[212] = is_max[212] | is_min[212];
assign is_keypoint[213] = is_max[213] | is_min[213];
assign is_keypoint[214] = is_max[214] | is_min[214];
assign is_keypoint[215] = is_max[215] | is_min[215];
assign is_keypoint[216] = is_max[216] | is_min[216];
assign is_keypoint[217] = is_max[217] | is_min[217];
assign is_keypoint[218] = is_max[218] | is_min[218];
assign is_keypoint[219] = is_max[219] | is_min[219];
assign is_keypoint[220] = is_max[220] | is_min[220];
assign is_keypoint[221] = is_max[221] | is_min[221];
assign is_keypoint[222] = is_max[222] | is_min[222];
assign is_keypoint[223] = is_max[223] | is_min[223];
assign is_keypoint[224] = is_max[224] | is_min[224];
assign is_keypoint[225] = is_max[225] | is_min[225];
assign is_keypoint[226] = is_max[226] | is_min[226];
assign is_keypoint[227] = is_max[227] | is_min[227];
assign is_keypoint[228] = is_max[228] | is_min[228];
assign is_keypoint[229] = is_max[229] | is_min[229];
assign is_keypoint[230] = is_max[230] | is_min[230];
assign is_keypoint[231] = is_max[231] | is_min[231];
assign is_keypoint[232] = is_max[232] | is_min[232];
assign is_keypoint[233] = is_max[233] | is_min[233];
assign is_keypoint[234] = is_max[234] | is_min[234];
assign is_keypoint[235] = is_max[235] | is_min[235];
assign is_keypoint[236] = is_max[236] | is_min[236];
assign is_keypoint[237] = is_max[237] | is_min[237];
assign is_keypoint[238] = is_max[238] | is_min[238];
assign is_keypoint[239] = is_max[239] | is_min[239];
assign is_keypoint[240] = is_max[240] | is_min[240];
assign is_keypoint[241] = is_max[241] | is_min[241];
assign is_keypoint[242] = is_max[242] | is_min[242];
assign is_keypoint[243] = is_max[243] | is_min[243];
assign is_keypoint[244] = is_max[244] | is_min[244];
assign is_keypoint[245] = is_max[245] | is_min[245];
assign is_keypoint[246] = is_max[246] | is_min[246];
assign is_keypoint[247] = is_max[247] | is_min[247];
assign is_keypoint[248] = is_max[248] | is_min[248];
assign is_keypoint[249] = is_max[249] | is_min[249];
assign is_keypoint[250] = is_max[250] | is_min[250];
assign is_keypoint[251] = is_max[251] | is_min[251];
assign is_keypoint[252] = is_max[252] | is_min[252];
assign is_keypoint[253] = is_max[253] | is_min[253];
assign is_keypoint[254] = is_max[254] | is_min[254];
assign is_keypoint[255] = is_max[255] | is_min[255];
assign is_keypoint[256] = is_max[256] | is_min[256];
assign is_keypoint[257] = is_max[257] | is_min[257];
assign is_keypoint[258] = is_max[258] | is_min[258];
assign is_keypoint[259] = is_max[259] | is_min[259];
assign is_keypoint[260] = is_max[260] | is_min[260];
assign is_keypoint[261] = is_max[261] | is_min[261];
assign is_keypoint[262] = is_max[262] | is_min[262];
assign is_keypoint[263] = is_max[263] | is_min[263];
assign is_keypoint[264] = is_max[264] | is_min[264];
assign is_keypoint[265] = is_max[265] | is_min[265];
assign is_keypoint[266] = is_max[266] | is_min[266];
assign is_keypoint[267] = is_max[267] | is_min[267];
assign is_keypoint[268] = is_max[268] | is_min[268];
assign is_keypoint[269] = is_max[269] | is_min[269];
assign is_keypoint[270] = is_max[270] | is_min[270];
assign is_keypoint[271] = is_max[271] | is_min[271];
assign is_keypoint[272] = is_max[272] | is_min[272];
assign is_keypoint[273] = is_max[273] | is_min[273];
assign is_keypoint[274] = is_max[274] | is_min[274];
assign is_keypoint[275] = is_max[275] | is_min[275];
assign is_keypoint[276] = is_max[276] | is_min[276];
assign is_keypoint[277] = is_max[277] | is_min[277];
assign is_keypoint[278] = is_max[278] | is_min[278];
assign is_keypoint[279] = is_max[279] | is_min[279];
assign is_keypoint[280] = is_max[280] | is_min[280];
assign is_keypoint[281] = is_max[281] | is_min[281];
assign is_keypoint[282] = is_max[282] | is_min[282];
assign is_keypoint[283] = is_max[283] | is_min[283];
assign is_keypoint[284] = is_max[284] | is_min[284];
assign is_keypoint[285] = is_max[285] | is_min[285];
assign is_keypoint[286] = is_max[286] | is_min[286];
assign is_keypoint[287] = is_max[287] | is_min[287];
assign is_keypoint[288] = is_max[288] | is_min[288];
assign is_keypoint[289] = is_max[289] | is_min[289];
assign is_keypoint[290] = is_max[290] | is_min[290];
assign is_keypoint[291] = is_max[291] | is_min[291];
assign is_keypoint[292] = is_max[292] | is_min[292];
assign is_keypoint[293] = is_max[293] | is_min[293];
assign is_keypoint[294] = is_max[294] | is_min[294];
assign is_keypoint[295] = is_max[295] | is_min[295];
assign is_keypoint[296] = is_max[296] | is_min[296];
assign is_keypoint[297] = is_max[297] | is_min[297];
assign is_keypoint[298] = is_max[298] | is_min[298];
assign is_keypoint[299] = is_max[299] | is_min[299];
assign is_keypoint[300] = is_max[300] | is_min[300];
assign is_keypoint[301] = is_max[301] | is_min[301];
assign is_keypoint[302] = is_max[302] | is_min[302];
assign is_keypoint[303] = is_max[303] | is_min[303];
assign is_keypoint[304] = is_max[304] | is_min[304];
assign is_keypoint[305] = is_max[305] | is_min[305];
assign is_keypoint[306] = is_max[306] | is_min[306];
assign is_keypoint[307] = is_max[307] | is_min[307];
assign is_keypoint[308] = is_max[308] | is_min[308];
assign is_keypoint[309] = is_max[309] | is_min[309];
assign is_keypoint[310] = is_max[310] | is_min[310];
assign is_keypoint[311] = is_max[311] | is_min[311];
assign is_keypoint[312] = is_max[312] | is_min[312];
assign is_keypoint[313] = is_max[313] | is_min[313];
assign is_keypoint[314] = is_max[314] | is_min[314];
assign is_keypoint[315] = is_max[315] | is_min[315];
assign is_keypoint[316] = is_max[316] | is_min[316];
assign is_keypoint[317] = is_max[317] | is_min[317];
assign is_keypoint[318] = is_max[318] | is_min[318];
assign is_keypoint[319] = is_max[319] | is_min[319];
assign is_keypoint[320] = is_max[320] | is_min[320];
assign is_keypoint[321] = is_max[321] | is_min[321];
assign is_keypoint[322] = is_max[322] | is_min[322];
assign is_keypoint[323] = is_max[323] | is_min[323];
assign is_keypoint[324] = is_max[324] | is_min[324];
assign is_keypoint[325] = is_max[325] | is_min[325];
assign is_keypoint[326] = is_max[326] | is_min[326];
assign is_keypoint[327] = is_max[327] | is_min[327];
assign is_keypoint[328] = is_max[328] | is_min[328];
assign is_keypoint[329] = is_max[329] | is_min[329];
assign is_keypoint[330] = is_max[330] | is_min[330];
assign is_keypoint[331] = is_max[331] | is_min[331];
assign is_keypoint[332] = is_max[332] | is_min[332];
assign is_keypoint[333] = is_max[333] | is_min[333];
assign is_keypoint[334] = is_max[334] | is_min[334];
assign is_keypoint[335] = is_max[335] | is_min[335];
assign is_keypoint[336] = is_max[336] | is_min[336];
assign is_keypoint[337] = is_max[337] | is_min[337];
assign is_keypoint[338] = is_max[338] | is_min[338];
assign is_keypoint[339] = is_max[339] | is_min[339];
assign is_keypoint[340] = is_max[340] | is_min[340];
assign is_keypoint[341] = is_max[341] | is_min[341];
assign is_keypoint[342] = is_max[342] | is_min[342];
assign is_keypoint[343] = is_max[343] | is_min[343];
assign is_keypoint[344] = is_max[344] | is_min[344];
assign is_keypoint[345] = is_max[345] | is_min[345];
assign is_keypoint[346] = is_max[346] | is_min[346];
assign is_keypoint[347] = is_max[347] | is_min[347];
assign is_keypoint[348] = is_max[348] | is_min[348];
assign is_keypoint[349] = is_max[349] | is_min[349];
assign is_keypoint[350] = is_max[350] | is_min[350];
assign is_keypoint[351] = is_max[351] | is_min[351];
assign is_keypoint[352] = is_max[352] | is_min[352];
assign is_keypoint[353] = is_max[353] | is_min[353];
assign is_keypoint[354] = is_max[354] | is_min[354];
assign is_keypoint[355] = is_max[355] | is_min[355];
assign is_keypoint[356] = is_max[356] | is_min[356];
assign is_keypoint[357] = is_max[357] | is_min[357];
assign is_keypoint[358] = is_max[358] | is_min[358];
assign is_keypoint[359] = is_max[359] | is_min[359];
assign is_keypoint[360] = is_max[360] | is_min[360];
assign is_keypoint[361] = is_max[361] | is_min[361];
assign is_keypoint[362] = is_max[362] | is_min[362];
assign is_keypoint[363] = is_max[363] | is_min[363];
assign is_keypoint[364] = is_max[364] | is_min[364];
assign is_keypoint[365] = is_max[365] | is_min[365];
assign is_keypoint[366] = is_max[366] | is_min[366];
assign is_keypoint[367] = is_max[367] | is_min[367];
assign is_keypoint[368] = is_max[368] | is_min[368];
assign is_keypoint[369] = is_max[369] | is_min[369];
assign is_keypoint[370] = is_max[370] | is_min[370];
assign is_keypoint[371] = is_max[371] | is_min[371];
assign is_keypoint[372] = is_max[372] | is_min[372];
assign is_keypoint[373] = is_max[373] | is_min[373];
assign is_keypoint[374] = is_max[374] | is_min[374];
assign is_keypoint[375] = is_max[375] | is_min[375];
assign is_keypoint[376] = is_max[376] | is_min[376];
assign is_keypoint[377] = is_max[377] | is_min[377];
assign is_keypoint[378] = is_max[378] | is_min[378];
assign is_keypoint[379] = is_max[379] | is_min[379];
assign is_keypoint[380] = is_max[380] | is_min[380];
assign is_keypoint[381] = is_max[381] | is_min[381];
assign is_keypoint[382] = is_max[382] | is_min[382];
assign is_keypoint[383] = is_max[383] | is_min[383];
assign is_keypoint[384] = is_max[384] | is_min[384];
assign is_keypoint[385] = is_max[385] | is_min[385];
assign is_keypoint[386] = is_max[386] | is_min[386];
assign is_keypoint[387] = is_max[387] | is_min[387];
assign is_keypoint[388] = is_max[388] | is_min[388];
assign is_keypoint[389] = is_max[389] | is_min[389];
assign is_keypoint[390] = is_max[390] | is_min[390];
assign is_keypoint[391] = is_max[391] | is_min[391];
assign is_keypoint[392] = is_max[392] | is_min[392];
assign is_keypoint[393] = is_max[393] | is_min[393];
assign is_keypoint[394] = is_max[394] | is_min[394];
assign is_keypoint[395] = is_max[395] | is_min[395];
assign is_keypoint[396] = is_max[396] | is_min[396];
assign is_keypoint[397] = is_max[397] | is_min[397];
assign is_keypoint[398] = is_max[398] | is_min[398];
assign is_keypoint[399] = is_max[399] | is_min[399];
assign is_keypoint[400] = is_max[400] | is_min[400];
assign is_keypoint[401] = is_max[401] | is_min[401];
assign is_keypoint[402] = is_max[402] | is_min[402];
assign is_keypoint[403] = is_max[403] | is_min[403];
assign is_keypoint[404] = is_max[404] | is_min[404];
assign is_keypoint[405] = is_max[405] | is_min[405];
assign is_keypoint[406] = is_max[406] | is_min[406];
assign is_keypoint[407] = is_max[407] | is_min[407];
assign is_keypoint[408] = is_max[408] | is_min[408];
assign is_keypoint[409] = is_max[409] | is_min[409];
assign is_keypoint[410] = is_max[410] | is_min[410];
assign is_keypoint[411] = is_max[411] | is_min[411];
assign is_keypoint[412] = is_max[412] | is_min[412];
assign is_keypoint[413] = is_max[413] | is_min[413];
assign is_keypoint[414] = is_max[414] | is_min[414];
assign is_keypoint[415] = is_max[415] | is_min[415];
assign is_keypoint[416] = is_max[416] | is_min[416];
assign is_keypoint[417] = is_max[417] | is_min[417];
assign is_keypoint[418] = is_max[418] | is_min[418];
assign is_keypoint[419] = is_max[419] | is_min[419];
assign is_keypoint[420] = is_max[420] | is_min[420];
assign is_keypoint[421] = is_max[421] | is_min[421];
assign is_keypoint[422] = is_max[422] | is_min[422];
assign is_keypoint[423] = is_max[423] | is_min[423];
assign is_keypoint[424] = is_max[424] | is_min[424];
assign is_keypoint[425] = is_max[425] | is_min[425];
assign is_keypoint[426] = is_max[426] | is_min[426];
assign is_keypoint[427] = is_max[427] | is_min[427];
assign is_keypoint[428] = is_max[428] | is_min[428];
assign is_keypoint[429] = is_max[429] | is_min[429];
assign is_keypoint[430] = is_max[430] | is_min[430];
assign is_keypoint[431] = is_max[431] | is_min[431];
assign is_keypoint[432] = is_max[432] | is_min[432];
assign is_keypoint[433] = is_max[433] | is_min[433];
assign is_keypoint[434] = is_max[434] | is_min[434];
assign is_keypoint[435] = is_max[435] | is_min[435];
assign is_keypoint[436] = is_max[436] | is_min[436];
assign is_keypoint[437] = is_max[437] | is_min[437];
assign is_keypoint[438] = is_max[438] | is_min[438];
assign is_keypoint[439] = is_max[439] | is_min[439];
assign is_keypoint[440] = is_max[440] | is_min[440];
assign is_keypoint[441] = is_max[441] | is_min[441];
assign is_keypoint[442] = is_max[442] | is_min[442];
assign is_keypoint[443] = is_max[443] | is_min[443];
assign is_keypoint[444] = is_max[444] | is_min[444];
assign is_keypoint[445] = is_max[445] | is_min[445];
assign is_keypoint[446] = is_max[446] | is_min[446];
assign is_keypoint[447] = is_max[447] | is_min[447];
assign is_keypoint[448] = is_max[448] | is_min[448];
assign is_keypoint[449] = is_max[449] | is_min[449];
assign is_keypoint[450] = is_max[450] | is_min[450];
assign is_keypoint[451] = is_max[451] | is_min[451];
assign is_keypoint[452] = is_max[452] | is_min[452];
assign is_keypoint[453] = is_max[453] | is_min[453];
assign is_keypoint[454] = is_max[454] | is_min[454];
assign is_keypoint[455] = is_max[455] | is_min[455];
assign is_keypoint[456] = is_max[456] | is_min[456];
assign is_keypoint[457] = is_max[457] | is_min[457];
assign is_keypoint[458] = is_max[458] | is_min[458];
assign is_keypoint[459] = is_max[459] | is_min[459];
assign is_keypoint[460] = is_max[460] | is_min[460];
assign is_keypoint[461] = is_max[461] | is_min[461];
assign is_keypoint[462] = is_max[462] | is_min[462];
assign is_keypoint[463] = is_max[463] | is_min[463];
assign is_keypoint[464] = is_max[464] | is_min[464];
assign is_keypoint[465] = is_max[465] | is_min[465];
assign is_keypoint[466] = is_max[466] | is_min[466];
assign is_keypoint[467] = is_max[467] | is_min[467];
assign is_keypoint[468] = is_max[468] | is_min[468];
assign is_keypoint[469] = is_max[469] | is_min[469];
assign is_keypoint[470] = is_max[470] | is_min[470];
assign is_keypoint[471] = is_max[471] | is_min[471];
assign is_keypoint[472] = is_max[472] | is_min[472];
assign is_keypoint[473] = is_max[473] | is_min[473];
assign is_keypoint[474] = is_max[474] | is_min[474];
assign is_keypoint[475] = is_max[475] | is_min[475];
assign is_keypoint[476] = is_max[476] | is_min[476];
assign is_keypoint[477] = is_max[477] | is_min[477];
assign is_keypoint[478] = is_max[478] | is_min[478];
assign is_keypoint[479] = is_max[479] | is_min[479];
assign is_keypoint[480] = is_max[480] | is_min[480];
assign is_keypoint[481] = is_max[481] | is_min[481];
assign is_keypoint[482] = is_max[482] | is_min[482];
assign is_keypoint[483] = is_max[483] | is_min[483];
assign is_keypoint[484] = is_max[484] | is_min[484];
assign is_keypoint[485] = is_max[485] | is_min[485];
assign is_keypoint[486] = is_max[486] | is_min[486];
assign is_keypoint[487] = is_max[487] | is_min[487];
assign is_keypoint[488] = is_max[488] | is_min[488];
assign is_keypoint[489] = is_max[489] | is_min[489];
assign is_keypoint[490] = is_max[490] | is_min[490];
assign is_keypoint[491] = is_max[491] | is_min[491];
assign is_keypoint[492] = is_max[492] | is_min[492];
assign is_keypoint[493] = is_max[493] | is_min[493];
assign is_keypoint[494] = is_max[494] | is_min[494];
assign is_keypoint[495] = is_max[495] | is_min[495];
assign is_keypoint[496] = is_max[496] | is_min[496];
assign is_keypoint[497] = is_max[497] | is_min[497];
assign is_keypoint[498] = is_max[498] | is_min[498];
assign is_keypoint[499] = is_max[499] | is_min[499];
assign is_keypoint[500] = is_max[500] | is_min[500];
assign is_keypoint[501] = is_max[501] | is_min[501];
assign is_keypoint[502] = is_max[502] | is_min[502];
assign is_keypoint[503] = is_max[503] | is_min[503];
assign is_keypoint[504] = is_max[504] | is_min[504];
assign is_keypoint[505] = is_max[505] | is_min[505];
assign is_keypoint[506] = is_max[506] | is_min[506];
assign is_keypoint[507] = is_max[507] | is_min[507];
assign is_keypoint[508] = is_max[508] | is_min[508];
assign is_keypoint[509] = is_max[509] | is_min[509];
assign is_keypoint[510] = is_max[510] | is_min[510];
assign is_keypoint[511] = is_max[511] | is_min[511];
assign is_keypoint[512] = is_max[512] | is_min[512];
assign is_keypoint[513] = is_max[513] | is_min[513];
assign is_keypoint[514] = is_max[514] | is_min[514];
assign is_keypoint[515] = is_max[515] | is_min[515];
assign is_keypoint[516] = is_max[516] | is_min[516];
assign is_keypoint[517] = is_max[517] | is_min[517];
assign is_keypoint[518] = is_max[518] | is_min[518];
assign is_keypoint[519] = is_max[519] | is_min[519];
assign is_keypoint[520] = is_max[520] | is_min[520];
assign is_keypoint[521] = is_max[521] | is_min[521];
assign is_keypoint[522] = is_max[522] | is_min[522];
assign is_keypoint[523] = is_max[523] | is_min[523];
assign is_keypoint[524] = is_max[524] | is_min[524];
assign is_keypoint[525] = is_max[525] | is_min[525];
assign is_keypoint[526] = is_max[526] | is_min[526];
assign is_keypoint[527] = is_max[527] | is_min[527];
assign is_keypoint[528] = is_max[528] | is_min[528];
assign is_keypoint[529] = is_max[529] | is_min[529];
assign is_keypoint[530] = is_max[530] | is_min[530];
assign is_keypoint[531] = is_max[531] | is_min[531];
assign is_keypoint[532] = is_max[532] | is_min[532];
assign is_keypoint[533] = is_max[533] | is_min[533];
assign is_keypoint[534] = is_max[534] | is_min[534];
assign is_keypoint[535] = is_max[535] | is_min[535];
assign is_keypoint[536] = is_max[536] | is_min[536];
assign is_keypoint[537] = is_max[537] | is_min[537];
assign is_keypoint[538] = is_max[538] | is_min[538];
assign is_keypoint[539] = is_max[539] | is_min[539];
assign is_keypoint[540] = is_max[540] | is_min[540];
assign is_keypoint[541] = is_max[541] | is_min[541];
assign is_keypoint[542] = is_max[542] | is_min[542];
assign is_keypoint[543] = is_max[543] | is_min[543];
assign is_keypoint[544] = is_max[544] | is_min[544];
assign is_keypoint[545] = is_max[545] | is_min[545];
assign is_keypoint[546] = is_max[546] | is_min[546];
assign is_keypoint[547] = is_max[547] | is_min[547];
assign is_keypoint[548] = is_max[548] | is_min[548];
assign is_keypoint[549] = is_max[549] | is_min[549];
assign is_keypoint[550] = is_max[550] | is_min[550];
assign is_keypoint[551] = is_max[551] | is_min[551];
assign is_keypoint[552] = is_max[552] | is_min[552];
assign is_keypoint[553] = is_max[553] | is_min[553];
assign is_keypoint[554] = is_max[554] | is_min[554];
assign is_keypoint[555] = is_max[555] | is_min[555];
assign is_keypoint[556] = is_max[556] | is_min[556];
assign is_keypoint[557] = is_max[557] | is_min[557];
assign is_keypoint[558] = is_max[558] | is_min[558];
assign is_keypoint[559] = is_max[559] | is_min[559];
assign is_keypoint[560] = is_max[560] | is_min[560];
assign is_keypoint[561] = is_max[561] | is_min[561];
assign is_keypoint[562] = is_max[562] | is_min[562];
assign is_keypoint[563] = is_max[563] | is_min[563];
assign is_keypoint[564] = is_max[564] | is_min[564];
assign is_keypoint[565] = is_max[565] | is_min[565];
assign is_keypoint[566] = is_max[566] | is_min[566];
assign is_keypoint[567] = is_max[567] | is_min[567];
assign is_keypoint[568] = is_max[568] | is_min[568];
assign is_keypoint[569] = is_max[569] | is_min[569];
assign is_keypoint[570] = is_max[570] | is_min[570];
assign is_keypoint[571] = is_max[571] | is_min[571];
assign is_keypoint[572] = is_max[572] | is_min[572];
assign is_keypoint[573] = is_max[573] | is_min[573];
assign is_keypoint[574] = is_max[574] | is_min[574];
assign is_keypoint[575] = is_max[575] | is_min[575];
assign is_keypoint[576] = is_max[576] | is_min[576];
assign is_keypoint[577] = is_max[577] | is_min[577];
assign is_keypoint[578] = is_max[578] | is_min[578];
assign is_keypoint[579] = is_max[579] | is_min[579];
assign is_keypoint[580] = is_max[580] | is_min[580];
assign is_keypoint[581] = is_max[581] | is_min[581];
assign is_keypoint[582] = is_max[582] | is_min[582];
assign is_keypoint[583] = is_max[583] | is_min[583];
assign is_keypoint[584] = is_max[584] | is_min[584];
assign is_keypoint[585] = is_max[585] | is_min[585];
assign is_keypoint[586] = is_max[586] | is_min[586];
assign is_keypoint[587] = is_max[587] | is_min[587];
assign is_keypoint[588] = is_max[588] | is_min[588];
assign is_keypoint[589] = is_max[589] | is_min[589];
assign is_keypoint[590] = is_max[590] | is_min[590];
assign is_keypoint[591] = is_max[591] | is_min[591];
assign is_keypoint[592] = is_max[592] | is_min[592];
assign is_keypoint[593] = is_max[593] | is_min[593];
assign is_keypoint[594] = is_max[594] | is_min[594];
assign is_keypoint[595] = is_max[595] | is_min[595];
assign is_keypoint[596] = is_max[596] | is_min[596];
assign is_keypoint[597] = is_max[597] | is_min[597];
assign is_keypoint[598] = is_max[598] | is_min[598];
assign is_keypoint[599] = is_max[599] | is_min[599];
assign is_keypoint[600] = is_max[600] | is_min[600];
assign is_keypoint[601] = is_max[601] | is_min[601];
assign is_keypoint[602] = is_max[602] | is_min[602];
assign is_keypoint[603] = is_max[603] | is_min[603];
assign is_keypoint[604] = is_max[604] | is_min[604];
assign is_keypoint[605] = is_max[605] | is_min[605];
assign is_keypoint[606] = is_max[606] | is_min[606];
assign is_keypoint[607] = is_max[607] | is_min[607];
assign is_keypoint[608] = is_max[608] | is_min[608];
assign is_keypoint[609] = is_max[609] | is_min[609];
assign is_keypoint[610] = is_max[610] | is_min[610];
assign is_keypoint[611] = is_max[611] | is_min[611];
assign is_keypoint[612] = is_max[612] | is_min[612];
assign is_keypoint[613] = is_max[613] | is_min[613];
assign is_keypoint[614] = is_max[614] | is_min[614];
assign is_keypoint[615] = is_max[615] | is_min[615];
assign is_keypoint[616] = is_max[616] | is_min[616];
assign is_keypoint[617] = is_max[617] | is_min[617];
assign is_keypoint[618] = is_max[618] | is_min[618];
assign is_keypoint[619] = is_max[619] | is_min[619];
assign is_keypoint[620] = is_max[620] | is_min[620];
assign is_keypoint[621] = is_max[621] | is_min[621];
assign is_keypoint[622] = is_max[622] | is_min[622];
assign is_keypoint[623] = is_max[623] | is_min[623];
assign is_keypoint[624] = is_max[624] | is_min[624];
assign is_keypoint[625] = is_max[625] | is_min[625];
assign is_keypoint[626] = is_max[626] | is_min[626];
assign is_keypoint[627] = is_max[627] | is_min[627];
assign is_keypoint[628] = is_max[628] | is_min[628];
assign is_keypoint[629] = is_max[629] | is_min[629];
assign is_keypoint[630] = is_max[630] | is_min[630];
assign is_keypoint[631] = is_max[631] | is_min[631];
assign is_keypoint[632] = is_max[632] | is_min[632];
assign is_keypoint[633] = is_max[633] | is_min[633];
assign is_keypoint[634] = is_max[634] | is_min[634];
assign is_keypoint[635] = is_max[635] | is_min[635];
assign is_keypoint[636] = is_max[636] | is_min[636];
assign is_keypoint[637] = is_max[637] | is_min[637];

endmodule