`timescale 1ns/10ps
module Gaussian_Blur_5x5_2(
  clk,
  rst_n,
  start,
  done,
  buffer_data_0,
  buffer_data_1,
  buffer_data_2,
  buffer_data_3,
  buffer_data_4,
  blur_mem_we,
  blur_addr,
  blur_din,
  img_addr,
  buffer_we
);


/*SYSTEM*/
input                 clk,
                      rst_n,
                      start;
output reg            done;
output                buffer_we;


/*LINE BUFFER*/
input       [5119:0]  buffer_data_0;
input       [5119:0]  buffer_data_1;
input       [5119:0]  buffer_data_2;
input       [5119:0]  buffer_data_3;
input       [5119:0]  buffer_data_4;

/*Image SRAM Control*/
output reg  [8:0]     img_addr;

/*SRAM Control*/
output reg  [5119:0]  blur_din;
output reg  [8:0]     blur_addr;
output reg            blur_mem_we;

/*Kernel Q0.18 (We take last 6 decimal digits for simplicity (<262144))*/
reg       [159:0]  G_Kernel_5x5[0:2];

/*Module FSM*/
parameter ST_IDLE   = 0,
          ST_READY  = 1,/*Idle 1 state for SRAM to get READY*/
          ST_START  = 2;

reg     [1:0] current_state,
              next_state;

/*Kernel Value*/

always @(posedge clk) begin
  if (!rst_n) begin
    G_Kernel_5x5_1[0][31:0]  <= 32'h07E31AF6; //18'b000001111110001100;//'d030809;         
    G_Kernel_5x5_1[0][63:32] <= 32'h0983EB80; //18'b000010011000001111;//'d037169;         
    G_Kernel_5x5_1[0][95:64] <= 32'h0A212B91; //18'b000010100010000100;//'d039568;        
    G_Kernel_5x5_1[0][127:96] <= 32'h0983EB80; //18'b000010011000001111;//'d037169;         
    G_Kernel_5x5_1[0][159:128] <= 32'h07E31AF6; //18'b000001111110001100;//'d030809;  
    G_Kernel_5x5_1[1][31:0]  <= 32'h0983EB80; //18'b000010011000001111;//'d037169;         
    G_Kernel_5x5_1[1][63:32] <= 32'h0B7AC7A0; //18'b000010110111101011;//'d044842;         
    G_Kernel_5x5_1[1][95:64] <= 32'h0C387DF7; //18'b000011000011100001;//'d047737;        
    G_Kernel_5x5_1[1][127:96] <= 32'h0B7AC7A0; //18'b000010110111101011;//'d044842;         
    G_Kernel_5x5_1[1][159:128] <= 32'h0983EB80; //18'b000010011000001111;//'d037169;   
    G_Kernel_5x5_1[2][31:0]  <= 32'h0A212B91; //18'b000010100010000100;//'d039568;         
    G_Kernel_5x5_1[2][63:32] <= 32'h0C387DF7; //18'b000011000011100001;//'d047737;         
    G_Kernel_5x5_1[2][95:64] <= 32'h0D02737E; //18'b000011010000001001;//'d050818;        
    G_Kernel_5x5_1[2][127:96] <= 32'h0C387DF7; //18'b000011000011100001;//'d047737;         
    G_Kernel_5x5_1[2][159:128] <= 32'h0A212B91; //18'b000010100010000100;//'d039568;          
  end
end


reg   buffer_we_stop;
always @(posedge clk) begin
  if (!rst_n) 
    buffer_we_stop <= 1'b0;    
  else if (img_addr=='d480)
    buffer_we_stop <= 1'b1;
  else
    buffer_we_stop <= 1'b0;
end

assign buffer_we = (start && !(buffer_we_stop || current_state==ST_IDLE)) ? 1:0;

always @(posedge clk) begin
  if (!rst_n) 
    img_addr <= 'd0;    
  else if (start && img_addr<'d480)
    img_addr <= img_addr + 'd1;
  else if (done)
    img_addr <= 'd0;
end

/*Module DONE, inform SYSTEM*/
always @(posedge clk) begin
  if (!rst_n)
    done <= 1'b0;    
  else if (current_state==ST_START && blur_addr=='d480)
    done <= 1'b1;
  else if (current_state==ST_IDLE)
    done <= 1'b0;
end


always @(posedge clk) begin
  if (!rst_n)
    blur_addr <= 'd0;
  else if (blur_mem_we && blur_addr<'d480)
    blur_addr <= blur_addr + 'd1;
  else if (current_state==ST_IDLE)
    blur_addr <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_mem_we <= 1'b0;
  else if (current_state==ST_START && img_addr > 'd3 && blur_addr<'d480)
    blur_mem_we <= 1'b1;
  else if (blur_addr=='d480 || current_state==ST_IDLE)
    blur_mem_we <= 1'b0;
end

reg     ready_start_relay;
always @(posedge clk) begin
  if (!rst_n) 
    ready_start_relay <= 1'b0;
  else if (current_state == ST_READY)
    ready_start_relay <= 1'b1; 
  else if (current_state == ST_IDLE)
    ready_start_relay <= 1'b0;
end

wire  [39:0]  kernel_img_mul_0[0:24];
assign kernel_img_mul_0[0] = buffer_data_4[7:0] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_0[1] = buffer_data_4[15:8] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_0[2] = buffer_data_4[23:16] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_0[5] = buffer_data_3[7:0] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_0[6] = buffer_data_3[15:8] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_0[7] = buffer_data_3[23:16] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_0[10] = buffer_data_2[7:0] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_0[11] = buffer_data_2[15:8] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_0[12] = buffer_data_2[23:16] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_0[15] = buffer_data_1[7:0] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_0[16] = buffer_data_1[15:8] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_0[17] = buffer_data_1[23:16] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_0[20] = buffer_data_0[7:0] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_0[21] = buffer_data_0[15:8] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_0[22] = buffer_data_0[23:16] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_0 = kernel_img_mul_0[0] + kernel_img_mul_0[1] + kernel_img_mul_0[2] + 
                kernel_img_mul_0[5] + kernel_img_mul_0[6] + kernel_img_mul_0[7] + 
                kernel_img_mul_0[10] + kernel_img_mul_0[11] + kernel_img_mul_0[12] + 
                kernel_img_mul_0[15] + kernel_img_mul_0[16] + kernel_img_mul_0[17] + 
                kernel_img_mul_0[20] + kernel_img_mul_0[21] + kernel_img_mul_0[22] + 
                'd0;
always @(posedge clk) begin
  if (!rst_n)
    blur_din[7:0] <= 'd0;
  else if (current_state==ST_START)
    blur_din[7:0] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[7:0] <= 'd0;
end

wire  [39:0]  kernel_img_mul_1[0:24];
assign kernel_img_mul_1[0] = buffer_data_4[7:0] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_1[1] = buffer_data_4[15:8] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_1[2] = buffer_data_4[23:16] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_1[3] = buffer_data_4[31:24] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_1[5] = buffer_data_3[7:0] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_1[6] = buffer_data_3[15:8] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_1[7] = buffer_data_3[23:16] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_1[8] = buffer_data_3[31:24] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_1[10] = buffer_data_2[7:0] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_1[11] = buffer_data_2[15:8] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_1[12] = buffer_data_2[23:16] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_1[13] = buffer_data_2[31:24] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_1[15] = buffer_data_1[7:0] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_1[16] = buffer_data_1[15:8] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_1[17] = buffer_data_1[23:16] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_1[18] = buffer_data_1[31:24] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_1[20] = buffer_data_0[7:0] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_1[21] = buffer_data_0[15:8] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_1[22] = buffer_data_0[23:16] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_1[23] = buffer_data_0[31:24] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_1 = kernel_img_mul_1[0] + kernel_img_mul_1[1] + kernel_img_mul_1[2] + 
                kernel_img_mul_1[3] + kernel_img_mul_1[5] + kernel_img_mul_1[6] + 
                kernel_img_mul_1[7] + kernel_img_mul_1[8] + kernel_img_mul_1[10] + 
                kernel_img_mul_1[11] + kernel_img_mul_1[12] + kernel_img_mul_1[13] + 
                kernel_img_mul_1[15] + kernel_img_mul_1[16] + kernel_img_mul_1[17] + 
                kernel_img_mul_1[18] + kernel_img_mul_1[20] + kernel_img_mul_1[21] + 
                kernel_img_mul_1[22] + kernel_img_mul_1[23] + 'd0;
always @(posedge clk) begin
  if (!rst_n)
    blur_din[15:8] <= 'd0;
  else if (current_state==ST_START)
    blur_din[15:8] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[15:8] <= 'd0;
end

wire  [39:0]  kernel_img_mul_2[0:24];
assign kernel_img_mul_2[0] = buffer_data_4[7:0] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_2[1] = buffer_data_4[15:8] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_2[2] = buffer_data_4[23:16] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_2[3] = buffer_data_4[31:24] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_2[4] = buffer_data_4[39:32] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_2[5] = buffer_data_3[7:0] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_2[6] = buffer_data_3[15:8] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_2[7] = buffer_data_3[23:16] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_2[8] = buffer_data_3[31:24] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_2[9] = buffer_data_3[39:32] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_2[10] = buffer_data_2[7:0] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_2[11] = buffer_data_2[15:8] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_2[12] = buffer_data_2[23:16] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_2[13] = buffer_data_2[31:24] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_2[14] = buffer_data_2[39:32] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_2[15] = buffer_data_1[7:0] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_2[16] = buffer_data_1[15:8] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_2[17] = buffer_data_1[23:16] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_2[18] = buffer_data_1[31:24] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_2[19] = buffer_data_1[39:32] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_2[20] = buffer_data_0[7:0] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_2[21] = buffer_data_0[15:8] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_2[22] = buffer_data_0[23:16] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_2[23] = buffer_data_0[31:24] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_2[24] = buffer_data_0[39:32] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_2 = kernel_img_mul_2[0] + kernel_img_mul_2[1] + kernel_img_mul_2[2] + 
                kernel_img_mul_2[3] + kernel_img_mul_2[4] + kernel_img_mul_2[5] + 
                kernel_img_mul_2[6] + kernel_img_mul_2[7] + kernel_img_mul_2[8] + 
                kernel_img_mul_2[9] + kernel_img_mul_2[10] + kernel_img_mul_2[11] + 
                kernel_img_mul_2[12] + kernel_img_mul_2[13] + kernel_img_mul_2[14] + 
                kernel_img_mul_2[15] + kernel_img_mul_2[16] + kernel_img_mul_2[17] + 
                kernel_img_mul_2[18] + kernel_img_mul_2[19] + kernel_img_mul_2[20] + 
                kernel_img_mul_2[21] + kernel_img_mul_2[22] + kernel_img_mul_2[23] + 
                kernel_img_mul_2[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[23:16] <= 'd0;
  else if (current_state==ST_START)
    blur_din[23:16] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[23:16] <= 'd0;
end

wire  [39:0]  kernel_img_mul_3[0:24];
assign kernel_img_mul_3[0] = buffer_data_4[15:8] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_3[1] = buffer_data_4[23:16] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_3[2] = buffer_data_4[31:24] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_3[3] = buffer_data_4[39:32] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_3[4] = buffer_data_4[47:40] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_3[5] = buffer_data_3[15:8] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_3[6] = buffer_data_3[23:16] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_3[7] = buffer_data_3[31:24] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_3[8] = buffer_data_3[39:32] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_3[9] = buffer_data_3[47:40] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_3[10] = buffer_data_2[15:8] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_3[11] = buffer_data_2[23:16] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_3[12] = buffer_data_2[31:24] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_3[13] = buffer_data_2[39:32] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_3[14] = buffer_data_2[47:40] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_3[15] = buffer_data_1[15:8] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_3[16] = buffer_data_1[23:16] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_3[17] = buffer_data_1[31:24] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_3[18] = buffer_data_1[39:32] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_3[19] = buffer_data_1[47:40] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_3[20] = buffer_data_0[15:8] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_3[21] = buffer_data_0[23:16] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_3[22] = buffer_data_0[31:24] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_3[23] = buffer_data_0[39:32] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_3[24] = buffer_data_0[47:40] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_3 = kernel_img_mul_3[0] + kernel_img_mul_3[1] + kernel_img_mul_3[2] + 
                kernel_img_mul_3[3] + kernel_img_mul_3[4] + kernel_img_mul_3[5] + 
                kernel_img_mul_3[6] + kernel_img_mul_3[7] + kernel_img_mul_3[8] + 
                kernel_img_mul_3[9] + kernel_img_mul_3[10] + kernel_img_mul_3[11] + 
                kernel_img_mul_3[12] + kernel_img_mul_3[13] + kernel_img_mul_3[14] + 
                kernel_img_mul_3[15] + kernel_img_mul_3[16] + kernel_img_mul_3[17] + 
                kernel_img_mul_3[18] + kernel_img_mul_3[19] + kernel_img_mul_3[20] + 
                kernel_img_mul_3[21] + kernel_img_mul_3[22] + kernel_img_mul_3[23] + 
                kernel_img_mul_3[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[31:24] <= 'd0;
  else if (current_state==ST_START)
    blur_din[31:24] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[31:24] <= 'd0;
end

wire  [39:0]  kernel_img_mul_4[0:24];
assign kernel_img_mul_4[0] = buffer_data_4[23:16] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_4[1] = buffer_data_4[31:24] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_4[2] = buffer_data_4[39:32] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_4[3] = buffer_data_4[47:40] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_4[4] = buffer_data_4[55:48] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_4[5] = buffer_data_3[23:16] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_4[6] = buffer_data_3[31:24] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_4[7] = buffer_data_3[39:32] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_4[8] = buffer_data_3[47:40] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_4[9] = buffer_data_3[55:48] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_4[10] = buffer_data_2[23:16] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_4[11] = buffer_data_2[31:24] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_4[12] = buffer_data_2[39:32] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_4[13] = buffer_data_2[47:40] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_4[14] = buffer_data_2[55:48] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_4[15] = buffer_data_1[23:16] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_4[16] = buffer_data_1[31:24] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_4[17] = buffer_data_1[39:32] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_4[18] = buffer_data_1[47:40] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_4[19] = buffer_data_1[55:48] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_4[20] = buffer_data_0[23:16] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_4[21] = buffer_data_0[31:24] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_4[22] = buffer_data_0[39:32] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_4[23] = buffer_data_0[47:40] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_4[24] = buffer_data_0[55:48] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_4 = kernel_img_mul_4[0] + kernel_img_mul_4[1] + kernel_img_mul_4[2] + 
                kernel_img_mul_4[3] + kernel_img_mul_4[4] + kernel_img_mul_4[5] + 
                kernel_img_mul_4[6] + kernel_img_mul_4[7] + kernel_img_mul_4[8] + 
                kernel_img_mul_4[9] + kernel_img_mul_4[10] + kernel_img_mul_4[11] + 
                kernel_img_mul_4[12] + kernel_img_mul_4[13] + kernel_img_mul_4[14] + 
                kernel_img_mul_4[15] + kernel_img_mul_4[16] + kernel_img_mul_4[17] + 
                kernel_img_mul_4[18] + kernel_img_mul_4[19] + kernel_img_mul_4[20] + 
                kernel_img_mul_4[21] + kernel_img_mul_4[22] + kernel_img_mul_4[23] + 
                kernel_img_mul_4[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[39:32] <= 'd0;
  else if (current_state==ST_START)
    blur_din[39:32] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[39:32] <= 'd0;
end

wire  [39:0]  kernel_img_mul_5[0:24];
assign kernel_img_mul_5[0] = buffer_data_4[31:24] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_5[1] = buffer_data_4[39:32] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_5[2] = buffer_data_4[47:40] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_5[3] = buffer_data_4[55:48] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_5[4] = buffer_data_4[63:56] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_5[5] = buffer_data_3[31:24] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_5[6] = buffer_data_3[39:32] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_5[7] = buffer_data_3[47:40] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_5[8] = buffer_data_3[55:48] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_5[9] = buffer_data_3[63:56] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_5[10] = buffer_data_2[31:24] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_5[11] = buffer_data_2[39:32] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_5[12] = buffer_data_2[47:40] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_5[13] = buffer_data_2[55:48] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_5[14] = buffer_data_2[63:56] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_5[15] = buffer_data_1[31:24] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_5[16] = buffer_data_1[39:32] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_5[17] = buffer_data_1[47:40] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_5[18] = buffer_data_1[55:48] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_5[19] = buffer_data_1[63:56] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_5[20] = buffer_data_0[31:24] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_5[21] = buffer_data_0[39:32] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_5[22] = buffer_data_0[47:40] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_5[23] = buffer_data_0[55:48] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_5[24] = buffer_data_0[63:56] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_5 = kernel_img_mul_5[0] + kernel_img_mul_5[1] + kernel_img_mul_5[2] + 
                kernel_img_mul_5[3] + kernel_img_mul_5[4] + kernel_img_mul_5[5] + 
                kernel_img_mul_5[6] + kernel_img_mul_5[7] + kernel_img_mul_5[8] + 
                kernel_img_mul_5[9] + kernel_img_mul_5[10] + kernel_img_mul_5[11] + 
                kernel_img_mul_5[12] + kernel_img_mul_5[13] + kernel_img_mul_5[14] + 
                kernel_img_mul_5[15] + kernel_img_mul_5[16] + kernel_img_mul_5[17] + 
                kernel_img_mul_5[18] + kernel_img_mul_5[19] + kernel_img_mul_5[20] + 
                kernel_img_mul_5[21] + kernel_img_mul_5[22] + kernel_img_mul_5[23] + 
                kernel_img_mul_5[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[47:40] <= 'd0;
  else if (current_state==ST_START)
    blur_din[47:40] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[47:40] <= 'd0;
end

wire  [39:0]  kernel_img_mul_6[0:24];
assign kernel_img_mul_6[0] = buffer_data_4[39:32] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_6[1] = buffer_data_4[47:40] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_6[2] = buffer_data_4[55:48] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_6[3] = buffer_data_4[63:56] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_6[4] = buffer_data_4[71:64] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_6[5] = buffer_data_3[39:32] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_6[6] = buffer_data_3[47:40] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_6[7] = buffer_data_3[55:48] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_6[8] = buffer_data_3[63:56] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_6[9] = buffer_data_3[71:64] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_6[10] = buffer_data_2[39:32] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_6[11] = buffer_data_2[47:40] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_6[12] = buffer_data_2[55:48] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_6[13] = buffer_data_2[63:56] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_6[14] = buffer_data_2[71:64] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_6[15] = buffer_data_1[39:32] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_6[16] = buffer_data_1[47:40] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_6[17] = buffer_data_1[55:48] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_6[18] = buffer_data_1[63:56] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_6[19] = buffer_data_1[71:64] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_6[20] = buffer_data_0[39:32] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_6[21] = buffer_data_0[47:40] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_6[22] = buffer_data_0[55:48] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_6[23] = buffer_data_0[63:56] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_6[24] = buffer_data_0[71:64] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_6 = kernel_img_mul_6[0] + kernel_img_mul_6[1] + kernel_img_mul_6[2] + 
                kernel_img_mul_6[3] + kernel_img_mul_6[4] + kernel_img_mul_6[5] + 
                kernel_img_mul_6[6] + kernel_img_mul_6[7] + kernel_img_mul_6[8] + 
                kernel_img_mul_6[9] + kernel_img_mul_6[10] + kernel_img_mul_6[11] + 
                kernel_img_mul_6[12] + kernel_img_mul_6[13] + kernel_img_mul_6[14] + 
                kernel_img_mul_6[15] + kernel_img_mul_6[16] + kernel_img_mul_6[17] + 
                kernel_img_mul_6[18] + kernel_img_mul_6[19] + kernel_img_mul_6[20] + 
                kernel_img_mul_6[21] + kernel_img_mul_6[22] + kernel_img_mul_6[23] + 
                kernel_img_mul_6[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[55:48] <= 'd0;
  else if (current_state==ST_START)
    blur_din[55:48] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[55:48] <= 'd0;
end

wire  [39:0]  kernel_img_mul_7[0:24];
assign kernel_img_mul_7[0] = buffer_data_4[47:40] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_7[1] = buffer_data_4[55:48] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_7[2] = buffer_data_4[63:56] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_7[3] = buffer_data_4[71:64] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_7[4] = buffer_data_4[79:72] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_7[5] = buffer_data_3[47:40] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_7[6] = buffer_data_3[55:48] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_7[7] = buffer_data_3[63:56] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_7[8] = buffer_data_3[71:64] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_7[9] = buffer_data_3[79:72] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_7[10] = buffer_data_2[47:40] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_7[11] = buffer_data_2[55:48] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_7[12] = buffer_data_2[63:56] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_7[13] = buffer_data_2[71:64] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_7[14] = buffer_data_2[79:72] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_7[15] = buffer_data_1[47:40] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_7[16] = buffer_data_1[55:48] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_7[17] = buffer_data_1[63:56] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_7[18] = buffer_data_1[71:64] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_7[19] = buffer_data_1[79:72] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_7[20] = buffer_data_0[47:40] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_7[21] = buffer_data_0[55:48] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_7[22] = buffer_data_0[63:56] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_7[23] = buffer_data_0[71:64] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_7[24] = buffer_data_0[79:72] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_7 = kernel_img_mul_7[0] + kernel_img_mul_7[1] + kernel_img_mul_7[2] + 
                kernel_img_mul_7[3] + kernel_img_mul_7[4] + kernel_img_mul_7[5] + 
                kernel_img_mul_7[6] + kernel_img_mul_7[7] + kernel_img_mul_7[8] + 
                kernel_img_mul_7[9] + kernel_img_mul_7[10] + kernel_img_mul_7[11] + 
                kernel_img_mul_7[12] + kernel_img_mul_7[13] + kernel_img_mul_7[14] + 
                kernel_img_mul_7[15] + kernel_img_mul_7[16] + kernel_img_mul_7[17] + 
                kernel_img_mul_7[18] + kernel_img_mul_7[19] + kernel_img_mul_7[20] + 
                kernel_img_mul_7[21] + kernel_img_mul_7[22] + kernel_img_mul_7[23] + 
                kernel_img_mul_7[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[63:56] <= 'd0;
  else if (current_state==ST_START)
    blur_din[63:56] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[63:56] <= 'd0;
end

wire  [39:0]  kernel_img_mul_8[0:24];
assign kernel_img_mul_8[0] = buffer_data_4[55:48] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_8[1] = buffer_data_4[63:56] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_8[2] = buffer_data_4[71:64] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_8[3] = buffer_data_4[79:72] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_8[4] = buffer_data_4[87:80] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_8[5] = buffer_data_3[55:48] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_8[6] = buffer_data_3[63:56] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_8[7] = buffer_data_3[71:64] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_8[8] = buffer_data_3[79:72] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_8[9] = buffer_data_3[87:80] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_8[10] = buffer_data_2[55:48] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_8[11] = buffer_data_2[63:56] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_8[12] = buffer_data_2[71:64] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_8[13] = buffer_data_2[79:72] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_8[14] = buffer_data_2[87:80] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_8[15] = buffer_data_1[55:48] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_8[16] = buffer_data_1[63:56] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_8[17] = buffer_data_1[71:64] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_8[18] = buffer_data_1[79:72] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_8[19] = buffer_data_1[87:80] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_8[20] = buffer_data_0[55:48] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_8[21] = buffer_data_0[63:56] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_8[22] = buffer_data_0[71:64] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_8[23] = buffer_data_0[79:72] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_8[24] = buffer_data_0[87:80] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_8 = kernel_img_mul_8[0] + kernel_img_mul_8[1] + kernel_img_mul_8[2] + 
                kernel_img_mul_8[3] + kernel_img_mul_8[4] + kernel_img_mul_8[5] + 
                kernel_img_mul_8[6] + kernel_img_mul_8[7] + kernel_img_mul_8[8] + 
                kernel_img_mul_8[9] + kernel_img_mul_8[10] + kernel_img_mul_8[11] + 
                kernel_img_mul_8[12] + kernel_img_mul_8[13] + kernel_img_mul_8[14] + 
                kernel_img_mul_8[15] + kernel_img_mul_8[16] + kernel_img_mul_8[17] + 
                kernel_img_mul_8[18] + kernel_img_mul_8[19] + kernel_img_mul_8[20] + 
                kernel_img_mul_8[21] + kernel_img_mul_8[22] + kernel_img_mul_8[23] + 
                kernel_img_mul_8[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[71:64] <= 'd0;
  else if (current_state==ST_START)
    blur_din[71:64] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[71:64] <= 'd0;
end

wire  [39:0]  kernel_img_mul_9[0:24];
assign kernel_img_mul_9[0] = buffer_data_4[63:56] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_9[1] = buffer_data_4[71:64] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_9[2] = buffer_data_4[79:72] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_9[3] = buffer_data_4[87:80] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_9[4] = buffer_data_4[95:88] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_9[5] = buffer_data_3[63:56] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_9[6] = buffer_data_3[71:64] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_9[7] = buffer_data_3[79:72] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_9[8] = buffer_data_3[87:80] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_9[9] = buffer_data_3[95:88] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_9[10] = buffer_data_2[63:56] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_9[11] = buffer_data_2[71:64] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_9[12] = buffer_data_2[79:72] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_9[13] = buffer_data_2[87:80] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_9[14] = buffer_data_2[95:88] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_9[15] = buffer_data_1[63:56] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_9[16] = buffer_data_1[71:64] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_9[17] = buffer_data_1[79:72] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_9[18] = buffer_data_1[87:80] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_9[19] = buffer_data_1[95:88] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_9[20] = buffer_data_0[63:56] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_9[21] = buffer_data_0[71:64] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_9[22] = buffer_data_0[79:72] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_9[23] = buffer_data_0[87:80] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_9[24] = buffer_data_0[95:88] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_9 = kernel_img_mul_9[0] + kernel_img_mul_9[1] + kernel_img_mul_9[2] + 
                kernel_img_mul_9[3] + kernel_img_mul_9[4] + kernel_img_mul_9[5] + 
                kernel_img_mul_9[6] + kernel_img_mul_9[7] + kernel_img_mul_9[8] + 
                kernel_img_mul_9[9] + kernel_img_mul_9[10] + kernel_img_mul_9[11] + 
                kernel_img_mul_9[12] + kernel_img_mul_9[13] + kernel_img_mul_9[14] + 
                kernel_img_mul_9[15] + kernel_img_mul_9[16] + kernel_img_mul_9[17] + 
                kernel_img_mul_9[18] + kernel_img_mul_9[19] + kernel_img_mul_9[20] + 
                kernel_img_mul_9[21] + kernel_img_mul_9[22] + kernel_img_mul_9[23] + 
                kernel_img_mul_9[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[79:72] <= 'd0;
  else if (current_state==ST_START)
    blur_din[79:72] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[79:72] <= 'd0;
end

wire  [39:0]  kernel_img_mul_10[0:24];
assign kernel_img_mul_10[0] = buffer_data_4[71:64] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_10[1] = buffer_data_4[79:72] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_10[2] = buffer_data_4[87:80] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_10[3] = buffer_data_4[95:88] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_10[4] = buffer_data_4[103:96] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_10[5] = buffer_data_3[71:64] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_10[6] = buffer_data_3[79:72] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_10[7] = buffer_data_3[87:80] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_10[8] = buffer_data_3[95:88] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_10[9] = buffer_data_3[103:96] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_10[10] = buffer_data_2[71:64] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_10[11] = buffer_data_2[79:72] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_10[12] = buffer_data_2[87:80] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_10[13] = buffer_data_2[95:88] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_10[14] = buffer_data_2[103:96] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_10[15] = buffer_data_1[71:64] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_10[16] = buffer_data_1[79:72] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_10[17] = buffer_data_1[87:80] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_10[18] = buffer_data_1[95:88] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_10[19] = buffer_data_1[103:96] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_10[20] = buffer_data_0[71:64] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_10[21] = buffer_data_0[79:72] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_10[22] = buffer_data_0[87:80] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_10[23] = buffer_data_0[95:88] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_10[24] = buffer_data_0[103:96] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_10 = kernel_img_mul_10[0] + kernel_img_mul_10[1] + kernel_img_mul_10[2] + 
                kernel_img_mul_10[3] + kernel_img_mul_10[4] + kernel_img_mul_10[5] + 
                kernel_img_mul_10[6] + kernel_img_mul_10[7] + kernel_img_mul_10[8] + 
                kernel_img_mul_10[9] + kernel_img_mul_10[10] + kernel_img_mul_10[11] + 
                kernel_img_mul_10[12] + kernel_img_mul_10[13] + kernel_img_mul_10[14] + 
                kernel_img_mul_10[15] + kernel_img_mul_10[16] + kernel_img_mul_10[17] + 
                kernel_img_mul_10[18] + kernel_img_mul_10[19] + kernel_img_mul_10[20] + 
                kernel_img_mul_10[21] + kernel_img_mul_10[22] + kernel_img_mul_10[23] + 
                kernel_img_mul_10[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[87:80] <= 'd0;
  else if (current_state==ST_START)
    blur_din[87:80] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[87:80] <= 'd0;
end

wire  [39:0]  kernel_img_mul_11[0:24];
assign kernel_img_mul_11[0] = buffer_data_4[79:72] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_11[1] = buffer_data_4[87:80] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_11[2] = buffer_data_4[95:88] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_11[3] = buffer_data_4[103:96] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_11[4] = buffer_data_4[111:104] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_11[5] = buffer_data_3[79:72] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_11[6] = buffer_data_3[87:80] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_11[7] = buffer_data_3[95:88] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_11[8] = buffer_data_3[103:96] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_11[9] = buffer_data_3[111:104] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_11[10] = buffer_data_2[79:72] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_11[11] = buffer_data_2[87:80] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_11[12] = buffer_data_2[95:88] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_11[13] = buffer_data_2[103:96] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_11[14] = buffer_data_2[111:104] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_11[15] = buffer_data_1[79:72] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_11[16] = buffer_data_1[87:80] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_11[17] = buffer_data_1[95:88] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_11[18] = buffer_data_1[103:96] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_11[19] = buffer_data_1[111:104] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_11[20] = buffer_data_0[79:72] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_11[21] = buffer_data_0[87:80] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_11[22] = buffer_data_0[95:88] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_11[23] = buffer_data_0[103:96] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_11[24] = buffer_data_0[111:104] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_11 = kernel_img_mul_11[0] + kernel_img_mul_11[1] + kernel_img_mul_11[2] + 
                kernel_img_mul_11[3] + kernel_img_mul_11[4] + kernel_img_mul_11[5] + 
                kernel_img_mul_11[6] + kernel_img_mul_11[7] + kernel_img_mul_11[8] + 
                kernel_img_mul_11[9] + kernel_img_mul_11[10] + kernel_img_mul_11[11] + 
                kernel_img_mul_11[12] + kernel_img_mul_11[13] + kernel_img_mul_11[14] + 
                kernel_img_mul_11[15] + kernel_img_mul_11[16] + kernel_img_mul_11[17] + 
                kernel_img_mul_11[18] + kernel_img_mul_11[19] + kernel_img_mul_11[20] + 
                kernel_img_mul_11[21] + kernel_img_mul_11[22] + kernel_img_mul_11[23] + 
                kernel_img_mul_11[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[95:88] <= 'd0;
  else if (current_state==ST_START)
    blur_din[95:88] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[95:88] <= 'd0;
end

wire  [39:0]  kernel_img_mul_12[0:24];
assign kernel_img_mul_12[0] = buffer_data_4[87:80] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_12[1] = buffer_data_4[95:88] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_12[2] = buffer_data_4[103:96] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_12[3] = buffer_data_4[111:104] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_12[4] = buffer_data_4[119:112] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_12[5] = buffer_data_3[87:80] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_12[6] = buffer_data_3[95:88] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_12[7] = buffer_data_3[103:96] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_12[8] = buffer_data_3[111:104] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_12[9] = buffer_data_3[119:112] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_12[10] = buffer_data_2[87:80] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_12[11] = buffer_data_2[95:88] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_12[12] = buffer_data_2[103:96] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_12[13] = buffer_data_2[111:104] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_12[14] = buffer_data_2[119:112] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_12[15] = buffer_data_1[87:80] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_12[16] = buffer_data_1[95:88] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_12[17] = buffer_data_1[103:96] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_12[18] = buffer_data_1[111:104] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_12[19] = buffer_data_1[119:112] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_12[20] = buffer_data_0[87:80] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_12[21] = buffer_data_0[95:88] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_12[22] = buffer_data_0[103:96] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_12[23] = buffer_data_0[111:104] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_12[24] = buffer_data_0[119:112] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_12 = kernel_img_mul_12[0] + kernel_img_mul_12[1] + kernel_img_mul_12[2] + 
                kernel_img_mul_12[3] + kernel_img_mul_12[4] + kernel_img_mul_12[5] + 
                kernel_img_mul_12[6] + kernel_img_mul_12[7] + kernel_img_mul_12[8] + 
                kernel_img_mul_12[9] + kernel_img_mul_12[10] + kernel_img_mul_12[11] + 
                kernel_img_mul_12[12] + kernel_img_mul_12[13] + kernel_img_mul_12[14] + 
                kernel_img_mul_12[15] + kernel_img_mul_12[16] + kernel_img_mul_12[17] + 
                kernel_img_mul_12[18] + kernel_img_mul_12[19] + kernel_img_mul_12[20] + 
                kernel_img_mul_12[21] + kernel_img_mul_12[22] + kernel_img_mul_12[23] + 
                kernel_img_mul_12[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[103:96] <= 'd0;
  else if (current_state==ST_START)
    blur_din[103:96] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[103:96] <= 'd0;
end

wire  [39:0]  kernel_img_mul_13[0:24];
assign kernel_img_mul_13[0] = buffer_data_4[95:88] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_13[1] = buffer_data_4[103:96] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_13[2] = buffer_data_4[111:104] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_13[3] = buffer_data_4[119:112] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_13[4] = buffer_data_4[127:120] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_13[5] = buffer_data_3[95:88] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_13[6] = buffer_data_3[103:96] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_13[7] = buffer_data_3[111:104] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_13[8] = buffer_data_3[119:112] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_13[9] = buffer_data_3[127:120] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_13[10] = buffer_data_2[95:88] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_13[11] = buffer_data_2[103:96] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_13[12] = buffer_data_2[111:104] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_13[13] = buffer_data_2[119:112] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_13[14] = buffer_data_2[127:120] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_13[15] = buffer_data_1[95:88] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_13[16] = buffer_data_1[103:96] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_13[17] = buffer_data_1[111:104] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_13[18] = buffer_data_1[119:112] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_13[19] = buffer_data_1[127:120] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_13[20] = buffer_data_0[95:88] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_13[21] = buffer_data_0[103:96] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_13[22] = buffer_data_0[111:104] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_13[23] = buffer_data_0[119:112] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_13[24] = buffer_data_0[127:120] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_13 = kernel_img_mul_13[0] + kernel_img_mul_13[1] + kernel_img_mul_13[2] + 
                kernel_img_mul_13[3] + kernel_img_mul_13[4] + kernel_img_mul_13[5] + 
                kernel_img_mul_13[6] + kernel_img_mul_13[7] + kernel_img_mul_13[8] + 
                kernel_img_mul_13[9] + kernel_img_mul_13[10] + kernel_img_mul_13[11] + 
                kernel_img_mul_13[12] + kernel_img_mul_13[13] + kernel_img_mul_13[14] + 
                kernel_img_mul_13[15] + kernel_img_mul_13[16] + kernel_img_mul_13[17] + 
                kernel_img_mul_13[18] + kernel_img_mul_13[19] + kernel_img_mul_13[20] + 
                kernel_img_mul_13[21] + kernel_img_mul_13[22] + kernel_img_mul_13[23] + 
                kernel_img_mul_13[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[111:104] <= 'd0;
  else if (current_state==ST_START)
    blur_din[111:104] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[111:104] <= 'd0;
end

wire  [39:0]  kernel_img_mul_14[0:24];
assign kernel_img_mul_14[0] = buffer_data_4[103:96] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_14[1] = buffer_data_4[111:104] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_14[2] = buffer_data_4[119:112] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_14[3] = buffer_data_4[127:120] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_14[4] = buffer_data_4[135:128] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_14[5] = buffer_data_3[103:96] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_14[6] = buffer_data_3[111:104] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_14[7] = buffer_data_3[119:112] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_14[8] = buffer_data_3[127:120] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_14[9] = buffer_data_3[135:128] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_14[10] = buffer_data_2[103:96] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_14[11] = buffer_data_2[111:104] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_14[12] = buffer_data_2[119:112] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_14[13] = buffer_data_2[127:120] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_14[14] = buffer_data_2[135:128] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_14[15] = buffer_data_1[103:96] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_14[16] = buffer_data_1[111:104] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_14[17] = buffer_data_1[119:112] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_14[18] = buffer_data_1[127:120] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_14[19] = buffer_data_1[135:128] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_14[20] = buffer_data_0[103:96] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_14[21] = buffer_data_0[111:104] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_14[22] = buffer_data_0[119:112] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_14[23] = buffer_data_0[127:120] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_14[24] = buffer_data_0[135:128] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_14 = kernel_img_mul_14[0] + kernel_img_mul_14[1] + kernel_img_mul_14[2] + 
                kernel_img_mul_14[3] + kernel_img_mul_14[4] + kernel_img_mul_14[5] + 
                kernel_img_mul_14[6] + kernel_img_mul_14[7] + kernel_img_mul_14[8] + 
                kernel_img_mul_14[9] + kernel_img_mul_14[10] + kernel_img_mul_14[11] + 
                kernel_img_mul_14[12] + kernel_img_mul_14[13] + kernel_img_mul_14[14] + 
                kernel_img_mul_14[15] + kernel_img_mul_14[16] + kernel_img_mul_14[17] + 
                kernel_img_mul_14[18] + kernel_img_mul_14[19] + kernel_img_mul_14[20] + 
                kernel_img_mul_14[21] + kernel_img_mul_14[22] + kernel_img_mul_14[23] + 
                kernel_img_mul_14[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[119:112] <= 'd0;
  else if (current_state==ST_START)
    blur_din[119:112] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[119:112] <= 'd0;
end

wire  [39:0]  kernel_img_mul_15[0:24];
assign kernel_img_mul_15[0] = buffer_data_4[111:104] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_15[1] = buffer_data_4[119:112] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_15[2] = buffer_data_4[127:120] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_15[3] = buffer_data_4[135:128] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_15[4] = buffer_data_4[143:136] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_15[5] = buffer_data_3[111:104] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_15[6] = buffer_data_3[119:112] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_15[7] = buffer_data_3[127:120] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_15[8] = buffer_data_3[135:128] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_15[9] = buffer_data_3[143:136] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_15[10] = buffer_data_2[111:104] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_15[11] = buffer_data_2[119:112] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_15[12] = buffer_data_2[127:120] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_15[13] = buffer_data_2[135:128] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_15[14] = buffer_data_2[143:136] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_15[15] = buffer_data_1[111:104] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_15[16] = buffer_data_1[119:112] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_15[17] = buffer_data_1[127:120] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_15[18] = buffer_data_1[135:128] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_15[19] = buffer_data_1[143:136] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_15[20] = buffer_data_0[111:104] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_15[21] = buffer_data_0[119:112] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_15[22] = buffer_data_0[127:120] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_15[23] = buffer_data_0[135:128] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_15[24] = buffer_data_0[143:136] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_15 = kernel_img_mul_15[0] + kernel_img_mul_15[1] + kernel_img_mul_15[2] + 
                kernel_img_mul_15[3] + kernel_img_mul_15[4] + kernel_img_mul_15[5] + 
                kernel_img_mul_15[6] + kernel_img_mul_15[7] + kernel_img_mul_15[8] + 
                kernel_img_mul_15[9] + kernel_img_mul_15[10] + kernel_img_mul_15[11] + 
                kernel_img_mul_15[12] + kernel_img_mul_15[13] + kernel_img_mul_15[14] + 
                kernel_img_mul_15[15] + kernel_img_mul_15[16] + kernel_img_mul_15[17] + 
                kernel_img_mul_15[18] + kernel_img_mul_15[19] + kernel_img_mul_15[20] + 
                kernel_img_mul_15[21] + kernel_img_mul_15[22] + kernel_img_mul_15[23] + 
                kernel_img_mul_15[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[127:120] <= 'd0;
  else if (current_state==ST_START)
    blur_din[127:120] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[127:120] <= 'd0;
end

wire  [39:0]  kernel_img_mul_16[0:24];
assign kernel_img_mul_16[0] = buffer_data_4[119:112] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_16[1] = buffer_data_4[127:120] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_16[2] = buffer_data_4[135:128] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_16[3] = buffer_data_4[143:136] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_16[4] = buffer_data_4[151:144] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_16[5] = buffer_data_3[119:112] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_16[6] = buffer_data_3[127:120] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_16[7] = buffer_data_3[135:128] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_16[8] = buffer_data_3[143:136] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_16[9] = buffer_data_3[151:144] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_16[10] = buffer_data_2[119:112] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_16[11] = buffer_data_2[127:120] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_16[12] = buffer_data_2[135:128] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_16[13] = buffer_data_2[143:136] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_16[14] = buffer_data_2[151:144] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_16[15] = buffer_data_1[119:112] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_16[16] = buffer_data_1[127:120] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_16[17] = buffer_data_1[135:128] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_16[18] = buffer_data_1[143:136] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_16[19] = buffer_data_1[151:144] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_16[20] = buffer_data_0[119:112] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_16[21] = buffer_data_0[127:120] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_16[22] = buffer_data_0[135:128] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_16[23] = buffer_data_0[143:136] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_16[24] = buffer_data_0[151:144] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_16 = kernel_img_mul_16[0] + kernel_img_mul_16[1] + kernel_img_mul_16[2] + 
                kernel_img_mul_16[3] + kernel_img_mul_16[4] + kernel_img_mul_16[5] + 
                kernel_img_mul_16[6] + kernel_img_mul_16[7] + kernel_img_mul_16[8] + 
                kernel_img_mul_16[9] + kernel_img_mul_16[10] + kernel_img_mul_16[11] + 
                kernel_img_mul_16[12] + kernel_img_mul_16[13] + kernel_img_mul_16[14] + 
                kernel_img_mul_16[15] + kernel_img_mul_16[16] + kernel_img_mul_16[17] + 
                kernel_img_mul_16[18] + kernel_img_mul_16[19] + kernel_img_mul_16[20] + 
                kernel_img_mul_16[21] + kernel_img_mul_16[22] + kernel_img_mul_16[23] + 
                kernel_img_mul_16[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[135:128] <= 'd0;
  else if (current_state==ST_START)
    blur_din[135:128] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[135:128] <= 'd0;
end

wire  [39:0]  kernel_img_mul_17[0:24];
assign kernel_img_mul_17[0] = buffer_data_4[127:120] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_17[1] = buffer_data_4[135:128] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_17[2] = buffer_data_4[143:136] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_17[3] = buffer_data_4[151:144] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_17[4] = buffer_data_4[159:152] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_17[5] = buffer_data_3[127:120] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_17[6] = buffer_data_3[135:128] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_17[7] = buffer_data_3[143:136] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_17[8] = buffer_data_3[151:144] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_17[9] = buffer_data_3[159:152] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_17[10] = buffer_data_2[127:120] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_17[11] = buffer_data_2[135:128] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_17[12] = buffer_data_2[143:136] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_17[13] = buffer_data_2[151:144] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_17[14] = buffer_data_2[159:152] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_17[15] = buffer_data_1[127:120] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_17[16] = buffer_data_1[135:128] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_17[17] = buffer_data_1[143:136] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_17[18] = buffer_data_1[151:144] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_17[19] = buffer_data_1[159:152] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_17[20] = buffer_data_0[127:120] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_17[21] = buffer_data_0[135:128] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_17[22] = buffer_data_0[143:136] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_17[23] = buffer_data_0[151:144] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_17[24] = buffer_data_0[159:152] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_17 = kernel_img_mul_17[0] + kernel_img_mul_17[1] + kernel_img_mul_17[2] + 
                kernel_img_mul_17[3] + kernel_img_mul_17[4] + kernel_img_mul_17[5] + 
                kernel_img_mul_17[6] + kernel_img_mul_17[7] + kernel_img_mul_17[8] + 
                kernel_img_mul_17[9] + kernel_img_mul_17[10] + kernel_img_mul_17[11] + 
                kernel_img_mul_17[12] + kernel_img_mul_17[13] + kernel_img_mul_17[14] + 
                kernel_img_mul_17[15] + kernel_img_mul_17[16] + kernel_img_mul_17[17] + 
                kernel_img_mul_17[18] + kernel_img_mul_17[19] + kernel_img_mul_17[20] + 
                kernel_img_mul_17[21] + kernel_img_mul_17[22] + kernel_img_mul_17[23] + 
                kernel_img_mul_17[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[143:136] <= 'd0;
  else if (current_state==ST_START)
    blur_din[143:136] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[143:136] <= 'd0;
end

wire  [39:0]  kernel_img_mul_18[0:24];
assign kernel_img_mul_18[0] = buffer_data_4[135:128] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_18[1] = buffer_data_4[143:136] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_18[2] = buffer_data_4[151:144] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_18[3] = buffer_data_4[159:152] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_18[4] = buffer_data_4[167:160] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_18[5] = buffer_data_3[135:128] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_18[6] = buffer_data_3[143:136] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_18[7] = buffer_data_3[151:144] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_18[8] = buffer_data_3[159:152] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_18[9] = buffer_data_3[167:160] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_18[10] = buffer_data_2[135:128] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_18[11] = buffer_data_2[143:136] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_18[12] = buffer_data_2[151:144] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_18[13] = buffer_data_2[159:152] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_18[14] = buffer_data_2[167:160] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_18[15] = buffer_data_1[135:128] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_18[16] = buffer_data_1[143:136] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_18[17] = buffer_data_1[151:144] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_18[18] = buffer_data_1[159:152] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_18[19] = buffer_data_1[167:160] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_18[20] = buffer_data_0[135:128] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_18[21] = buffer_data_0[143:136] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_18[22] = buffer_data_0[151:144] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_18[23] = buffer_data_0[159:152] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_18[24] = buffer_data_0[167:160] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_18 = kernel_img_mul_18[0] + kernel_img_mul_18[1] + kernel_img_mul_18[2] + 
                kernel_img_mul_18[3] + kernel_img_mul_18[4] + kernel_img_mul_18[5] + 
                kernel_img_mul_18[6] + kernel_img_mul_18[7] + kernel_img_mul_18[8] + 
                kernel_img_mul_18[9] + kernel_img_mul_18[10] + kernel_img_mul_18[11] + 
                kernel_img_mul_18[12] + kernel_img_mul_18[13] + kernel_img_mul_18[14] + 
                kernel_img_mul_18[15] + kernel_img_mul_18[16] + kernel_img_mul_18[17] + 
                kernel_img_mul_18[18] + kernel_img_mul_18[19] + kernel_img_mul_18[20] + 
                kernel_img_mul_18[21] + kernel_img_mul_18[22] + kernel_img_mul_18[23] + 
                kernel_img_mul_18[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[151:144] <= 'd0;
  else if (current_state==ST_START)
    blur_din[151:144] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[151:144] <= 'd0;
end

wire  [39:0]  kernel_img_mul_19[0:24];
assign kernel_img_mul_19[0] = buffer_data_4[143:136] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_19[1] = buffer_data_4[151:144] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_19[2] = buffer_data_4[159:152] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_19[3] = buffer_data_4[167:160] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_19[4] = buffer_data_4[175:168] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_19[5] = buffer_data_3[143:136] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_19[6] = buffer_data_3[151:144] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_19[7] = buffer_data_3[159:152] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_19[8] = buffer_data_3[167:160] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_19[9] = buffer_data_3[175:168] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_19[10] = buffer_data_2[143:136] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_19[11] = buffer_data_2[151:144] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_19[12] = buffer_data_2[159:152] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_19[13] = buffer_data_2[167:160] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_19[14] = buffer_data_2[175:168] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_19[15] = buffer_data_1[143:136] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_19[16] = buffer_data_1[151:144] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_19[17] = buffer_data_1[159:152] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_19[18] = buffer_data_1[167:160] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_19[19] = buffer_data_1[175:168] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_19[20] = buffer_data_0[143:136] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_19[21] = buffer_data_0[151:144] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_19[22] = buffer_data_0[159:152] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_19[23] = buffer_data_0[167:160] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_19[24] = buffer_data_0[175:168] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_19 = kernel_img_mul_19[0] + kernel_img_mul_19[1] + kernel_img_mul_19[2] + 
                kernel_img_mul_19[3] + kernel_img_mul_19[4] + kernel_img_mul_19[5] + 
                kernel_img_mul_19[6] + kernel_img_mul_19[7] + kernel_img_mul_19[8] + 
                kernel_img_mul_19[9] + kernel_img_mul_19[10] + kernel_img_mul_19[11] + 
                kernel_img_mul_19[12] + kernel_img_mul_19[13] + kernel_img_mul_19[14] + 
                kernel_img_mul_19[15] + kernel_img_mul_19[16] + kernel_img_mul_19[17] + 
                kernel_img_mul_19[18] + kernel_img_mul_19[19] + kernel_img_mul_19[20] + 
                kernel_img_mul_19[21] + kernel_img_mul_19[22] + kernel_img_mul_19[23] + 
                kernel_img_mul_19[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[159:152] <= 'd0;
  else if (current_state==ST_START)
    blur_din[159:152] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[159:152] <= 'd0;
end

wire  [39:0]  kernel_img_mul_20[0:24];
assign kernel_img_mul_20[0] = buffer_data_4[151:144] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_20[1] = buffer_data_4[159:152] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_20[2] = buffer_data_4[167:160] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_20[3] = buffer_data_4[175:168] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_20[4] = buffer_data_4[183:176] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_20[5] = buffer_data_3[151:144] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_20[6] = buffer_data_3[159:152] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_20[7] = buffer_data_3[167:160] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_20[8] = buffer_data_3[175:168] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_20[9] = buffer_data_3[183:176] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_20[10] = buffer_data_2[151:144] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_20[11] = buffer_data_2[159:152] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_20[12] = buffer_data_2[167:160] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_20[13] = buffer_data_2[175:168] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_20[14] = buffer_data_2[183:176] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_20[15] = buffer_data_1[151:144] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_20[16] = buffer_data_1[159:152] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_20[17] = buffer_data_1[167:160] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_20[18] = buffer_data_1[175:168] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_20[19] = buffer_data_1[183:176] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_20[20] = buffer_data_0[151:144] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_20[21] = buffer_data_0[159:152] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_20[22] = buffer_data_0[167:160] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_20[23] = buffer_data_0[175:168] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_20[24] = buffer_data_0[183:176] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_20 = kernel_img_mul_20[0] + kernel_img_mul_20[1] + kernel_img_mul_20[2] + 
                kernel_img_mul_20[3] + kernel_img_mul_20[4] + kernel_img_mul_20[5] + 
                kernel_img_mul_20[6] + kernel_img_mul_20[7] + kernel_img_mul_20[8] + 
                kernel_img_mul_20[9] + kernel_img_mul_20[10] + kernel_img_mul_20[11] + 
                kernel_img_mul_20[12] + kernel_img_mul_20[13] + kernel_img_mul_20[14] + 
                kernel_img_mul_20[15] + kernel_img_mul_20[16] + kernel_img_mul_20[17] + 
                kernel_img_mul_20[18] + kernel_img_mul_20[19] + kernel_img_mul_20[20] + 
                kernel_img_mul_20[21] + kernel_img_mul_20[22] + kernel_img_mul_20[23] + 
                kernel_img_mul_20[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[167:160] <= 'd0;
  else if (current_state==ST_START)
    blur_din[167:160] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[167:160] <= 'd0;
end

wire  [39:0]  kernel_img_mul_21[0:24];
assign kernel_img_mul_21[0] = buffer_data_4[159:152] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_21[1] = buffer_data_4[167:160] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_21[2] = buffer_data_4[175:168] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_21[3] = buffer_data_4[183:176] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_21[4] = buffer_data_4[191:184] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_21[5] = buffer_data_3[159:152] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_21[6] = buffer_data_3[167:160] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_21[7] = buffer_data_3[175:168] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_21[8] = buffer_data_3[183:176] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_21[9] = buffer_data_3[191:184] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_21[10] = buffer_data_2[159:152] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_21[11] = buffer_data_2[167:160] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_21[12] = buffer_data_2[175:168] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_21[13] = buffer_data_2[183:176] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_21[14] = buffer_data_2[191:184] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_21[15] = buffer_data_1[159:152] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_21[16] = buffer_data_1[167:160] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_21[17] = buffer_data_1[175:168] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_21[18] = buffer_data_1[183:176] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_21[19] = buffer_data_1[191:184] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_21[20] = buffer_data_0[159:152] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_21[21] = buffer_data_0[167:160] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_21[22] = buffer_data_0[175:168] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_21[23] = buffer_data_0[183:176] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_21[24] = buffer_data_0[191:184] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_21 = kernel_img_mul_21[0] + kernel_img_mul_21[1] + kernel_img_mul_21[2] + 
                kernel_img_mul_21[3] + kernel_img_mul_21[4] + kernel_img_mul_21[5] + 
                kernel_img_mul_21[6] + kernel_img_mul_21[7] + kernel_img_mul_21[8] + 
                kernel_img_mul_21[9] + kernel_img_mul_21[10] + kernel_img_mul_21[11] + 
                kernel_img_mul_21[12] + kernel_img_mul_21[13] + kernel_img_mul_21[14] + 
                kernel_img_mul_21[15] + kernel_img_mul_21[16] + kernel_img_mul_21[17] + 
                kernel_img_mul_21[18] + kernel_img_mul_21[19] + kernel_img_mul_21[20] + 
                kernel_img_mul_21[21] + kernel_img_mul_21[22] + kernel_img_mul_21[23] + 
                kernel_img_mul_21[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[175:168] <= 'd0;
  else if (current_state==ST_START)
    blur_din[175:168] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[175:168] <= 'd0;
end

wire  [39:0]  kernel_img_mul_22[0:24];
assign kernel_img_mul_22[0] = buffer_data_4[167:160] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_22[1] = buffer_data_4[175:168] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_22[2] = buffer_data_4[183:176] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_22[3] = buffer_data_4[191:184] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_22[4] = buffer_data_4[199:192] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_22[5] = buffer_data_3[167:160] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_22[6] = buffer_data_3[175:168] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_22[7] = buffer_data_3[183:176] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_22[8] = buffer_data_3[191:184] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_22[9] = buffer_data_3[199:192] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_22[10] = buffer_data_2[167:160] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_22[11] = buffer_data_2[175:168] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_22[12] = buffer_data_2[183:176] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_22[13] = buffer_data_2[191:184] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_22[14] = buffer_data_2[199:192] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_22[15] = buffer_data_1[167:160] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_22[16] = buffer_data_1[175:168] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_22[17] = buffer_data_1[183:176] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_22[18] = buffer_data_1[191:184] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_22[19] = buffer_data_1[199:192] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_22[20] = buffer_data_0[167:160] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_22[21] = buffer_data_0[175:168] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_22[22] = buffer_data_0[183:176] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_22[23] = buffer_data_0[191:184] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_22[24] = buffer_data_0[199:192] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_22 = kernel_img_mul_22[0] + kernel_img_mul_22[1] + kernel_img_mul_22[2] + 
                kernel_img_mul_22[3] + kernel_img_mul_22[4] + kernel_img_mul_22[5] + 
                kernel_img_mul_22[6] + kernel_img_mul_22[7] + kernel_img_mul_22[8] + 
                kernel_img_mul_22[9] + kernel_img_mul_22[10] + kernel_img_mul_22[11] + 
                kernel_img_mul_22[12] + kernel_img_mul_22[13] + kernel_img_mul_22[14] + 
                kernel_img_mul_22[15] + kernel_img_mul_22[16] + kernel_img_mul_22[17] + 
                kernel_img_mul_22[18] + kernel_img_mul_22[19] + kernel_img_mul_22[20] + 
                kernel_img_mul_22[21] + kernel_img_mul_22[22] + kernel_img_mul_22[23] + 
                kernel_img_mul_22[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[183:176] <= 'd0;
  else if (current_state==ST_START)
    blur_din[183:176] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[183:176] <= 'd0;
end

wire  [39:0]  kernel_img_mul_23[0:24];
assign kernel_img_mul_23[0] = buffer_data_4[175:168] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_23[1] = buffer_data_4[183:176] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_23[2] = buffer_data_4[191:184] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_23[3] = buffer_data_4[199:192] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_23[4] = buffer_data_4[207:200] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_23[5] = buffer_data_3[175:168] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_23[6] = buffer_data_3[183:176] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_23[7] = buffer_data_3[191:184] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_23[8] = buffer_data_3[199:192] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_23[9] = buffer_data_3[207:200] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_23[10] = buffer_data_2[175:168] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_23[11] = buffer_data_2[183:176] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_23[12] = buffer_data_2[191:184] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_23[13] = buffer_data_2[199:192] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_23[14] = buffer_data_2[207:200] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_23[15] = buffer_data_1[175:168] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_23[16] = buffer_data_1[183:176] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_23[17] = buffer_data_1[191:184] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_23[18] = buffer_data_1[199:192] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_23[19] = buffer_data_1[207:200] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_23[20] = buffer_data_0[175:168] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_23[21] = buffer_data_0[183:176] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_23[22] = buffer_data_0[191:184] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_23[23] = buffer_data_0[199:192] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_23[24] = buffer_data_0[207:200] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_23 = kernel_img_mul_23[0] + kernel_img_mul_23[1] + kernel_img_mul_23[2] + 
                kernel_img_mul_23[3] + kernel_img_mul_23[4] + kernel_img_mul_23[5] + 
                kernel_img_mul_23[6] + kernel_img_mul_23[7] + kernel_img_mul_23[8] + 
                kernel_img_mul_23[9] + kernel_img_mul_23[10] + kernel_img_mul_23[11] + 
                kernel_img_mul_23[12] + kernel_img_mul_23[13] + kernel_img_mul_23[14] + 
                kernel_img_mul_23[15] + kernel_img_mul_23[16] + kernel_img_mul_23[17] + 
                kernel_img_mul_23[18] + kernel_img_mul_23[19] + kernel_img_mul_23[20] + 
                kernel_img_mul_23[21] + kernel_img_mul_23[22] + kernel_img_mul_23[23] + 
                kernel_img_mul_23[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[191:184] <= 'd0;
  else if (current_state==ST_START)
    blur_din[191:184] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[191:184] <= 'd0;
end

wire  [39:0]  kernel_img_mul_24[0:24];
assign kernel_img_mul_24[0] = buffer_data_4[183:176] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_24[1] = buffer_data_4[191:184] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_24[2] = buffer_data_4[199:192] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_24[3] = buffer_data_4[207:200] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_24[4] = buffer_data_4[215:208] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_24[5] = buffer_data_3[183:176] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_24[6] = buffer_data_3[191:184] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_24[7] = buffer_data_3[199:192] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_24[8] = buffer_data_3[207:200] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_24[9] = buffer_data_3[215:208] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_24[10] = buffer_data_2[183:176] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_24[11] = buffer_data_2[191:184] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_24[12] = buffer_data_2[199:192] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_24[13] = buffer_data_2[207:200] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_24[14] = buffer_data_2[215:208] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_24[15] = buffer_data_1[183:176] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_24[16] = buffer_data_1[191:184] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_24[17] = buffer_data_1[199:192] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_24[18] = buffer_data_1[207:200] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_24[19] = buffer_data_1[215:208] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_24[20] = buffer_data_0[183:176] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_24[21] = buffer_data_0[191:184] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_24[22] = buffer_data_0[199:192] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_24[23] = buffer_data_0[207:200] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_24[24] = buffer_data_0[215:208] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_24 = kernel_img_mul_24[0] + kernel_img_mul_24[1] + kernel_img_mul_24[2] + 
                kernel_img_mul_24[3] + kernel_img_mul_24[4] + kernel_img_mul_24[5] + 
                kernel_img_mul_24[6] + kernel_img_mul_24[7] + kernel_img_mul_24[8] + 
                kernel_img_mul_24[9] + kernel_img_mul_24[10] + kernel_img_mul_24[11] + 
                kernel_img_mul_24[12] + kernel_img_mul_24[13] + kernel_img_mul_24[14] + 
                kernel_img_mul_24[15] + kernel_img_mul_24[16] + kernel_img_mul_24[17] + 
                kernel_img_mul_24[18] + kernel_img_mul_24[19] + kernel_img_mul_24[20] + 
                kernel_img_mul_24[21] + kernel_img_mul_24[22] + kernel_img_mul_24[23] + 
                kernel_img_mul_24[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[199:192] <= 'd0;
  else if (current_state==ST_START)
    blur_din[199:192] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[199:192] <= 'd0;
end

wire  [39:0]  kernel_img_mul_25[0:24];
assign kernel_img_mul_25[0] = buffer_data_4[191:184] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_25[1] = buffer_data_4[199:192] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_25[2] = buffer_data_4[207:200] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_25[3] = buffer_data_4[215:208] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_25[4] = buffer_data_4[223:216] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_25[5] = buffer_data_3[191:184] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_25[6] = buffer_data_3[199:192] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_25[7] = buffer_data_3[207:200] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_25[8] = buffer_data_3[215:208] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_25[9] = buffer_data_3[223:216] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_25[10] = buffer_data_2[191:184] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_25[11] = buffer_data_2[199:192] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_25[12] = buffer_data_2[207:200] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_25[13] = buffer_data_2[215:208] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_25[14] = buffer_data_2[223:216] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_25[15] = buffer_data_1[191:184] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_25[16] = buffer_data_1[199:192] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_25[17] = buffer_data_1[207:200] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_25[18] = buffer_data_1[215:208] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_25[19] = buffer_data_1[223:216] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_25[20] = buffer_data_0[191:184] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_25[21] = buffer_data_0[199:192] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_25[22] = buffer_data_0[207:200] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_25[23] = buffer_data_0[215:208] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_25[24] = buffer_data_0[223:216] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_25 = kernel_img_mul_25[0] + kernel_img_mul_25[1] + kernel_img_mul_25[2] + 
                kernel_img_mul_25[3] + kernel_img_mul_25[4] + kernel_img_mul_25[5] + 
                kernel_img_mul_25[6] + kernel_img_mul_25[7] + kernel_img_mul_25[8] + 
                kernel_img_mul_25[9] + kernel_img_mul_25[10] + kernel_img_mul_25[11] + 
                kernel_img_mul_25[12] + kernel_img_mul_25[13] + kernel_img_mul_25[14] + 
                kernel_img_mul_25[15] + kernel_img_mul_25[16] + kernel_img_mul_25[17] + 
                kernel_img_mul_25[18] + kernel_img_mul_25[19] + kernel_img_mul_25[20] + 
                kernel_img_mul_25[21] + kernel_img_mul_25[22] + kernel_img_mul_25[23] + 
                kernel_img_mul_25[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[207:200] <= 'd0;
  else if (current_state==ST_START)
    blur_din[207:200] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[207:200] <= 'd0;
end

wire  [39:0]  kernel_img_mul_26[0:24];
assign kernel_img_mul_26[0] = buffer_data_4[199:192] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_26[1] = buffer_data_4[207:200] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_26[2] = buffer_data_4[215:208] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_26[3] = buffer_data_4[223:216] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_26[4] = buffer_data_4[231:224] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_26[5] = buffer_data_3[199:192] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_26[6] = buffer_data_3[207:200] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_26[7] = buffer_data_3[215:208] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_26[8] = buffer_data_3[223:216] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_26[9] = buffer_data_3[231:224] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_26[10] = buffer_data_2[199:192] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_26[11] = buffer_data_2[207:200] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_26[12] = buffer_data_2[215:208] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_26[13] = buffer_data_2[223:216] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_26[14] = buffer_data_2[231:224] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_26[15] = buffer_data_1[199:192] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_26[16] = buffer_data_1[207:200] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_26[17] = buffer_data_1[215:208] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_26[18] = buffer_data_1[223:216] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_26[19] = buffer_data_1[231:224] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_26[20] = buffer_data_0[199:192] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_26[21] = buffer_data_0[207:200] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_26[22] = buffer_data_0[215:208] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_26[23] = buffer_data_0[223:216] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_26[24] = buffer_data_0[231:224] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_26 = kernel_img_mul_26[0] + kernel_img_mul_26[1] + kernel_img_mul_26[2] + 
                kernel_img_mul_26[3] + kernel_img_mul_26[4] + kernel_img_mul_26[5] + 
                kernel_img_mul_26[6] + kernel_img_mul_26[7] + kernel_img_mul_26[8] + 
                kernel_img_mul_26[9] + kernel_img_mul_26[10] + kernel_img_mul_26[11] + 
                kernel_img_mul_26[12] + kernel_img_mul_26[13] + kernel_img_mul_26[14] + 
                kernel_img_mul_26[15] + kernel_img_mul_26[16] + kernel_img_mul_26[17] + 
                kernel_img_mul_26[18] + kernel_img_mul_26[19] + kernel_img_mul_26[20] + 
                kernel_img_mul_26[21] + kernel_img_mul_26[22] + kernel_img_mul_26[23] + 
                kernel_img_mul_26[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[215:208] <= 'd0;
  else if (current_state==ST_START)
    blur_din[215:208] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[215:208] <= 'd0;
end

wire  [39:0]  kernel_img_mul_27[0:24];
assign kernel_img_mul_27[0] = buffer_data_4[207:200] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_27[1] = buffer_data_4[215:208] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_27[2] = buffer_data_4[223:216] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_27[3] = buffer_data_4[231:224] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_27[4] = buffer_data_4[239:232] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_27[5] = buffer_data_3[207:200] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_27[6] = buffer_data_3[215:208] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_27[7] = buffer_data_3[223:216] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_27[8] = buffer_data_3[231:224] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_27[9] = buffer_data_3[239:232] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_27[10] = buffer_data_2[207:200] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_27[11] = buffer_data_2[215:208] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_27[12] = buffer_data_2[223:216] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_27[13] = buffer_data_2[231:224] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_27[14] = buffer_data_2[239:232] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_27[15] = buffer_data_1[207:200] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_27[16] = buffer_data_1[215:208] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_27[17] = buffer_data_1[223:216] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_27[18] = buffer_data_1[231:224] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_27[19] = buffer_data_1[239:232] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_27[20] = buffer_data_0[207:200] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_27[21] = buffer_data_0[215:208] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_27[22] = buffer_data_0[223:216] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_27[23] = buffer_data_0[231:224] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_27[24] = buffer_data_0[239:232] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_27 = kernel_img_mul_27[0] + kernel_img_mul_27[1] + kernel_img_mul_27[2] + 
                kernel_img_mul_27[3] + kernel_img_mul_27[4] + kernel_img_mul_27[5] + 
                kernel_img_mul_27[6] + kernel_img_mul_27[7] + kernel_img_mul_27[8] + 
                kernel_img_mul_27[9] + kernel_img_mul_27[10] + kernel_img_mul_27[11] + 
                kernel_img_mul_27[12] + kernel_img_mul_27[13] + kernel_img_mul_27[14] + 
                kernel_img_mul_27[15] + kernel_img_mul_27[16] + kernel_img_mul_27[17] + 
                kernel_img_mul_27[18] + kernel_img_mul_27[19] + kernel_img_mul_27[20] + 
                kernel_img_mul_27[21] + kernel_img_mul_27[22] + kernel_img_mul_27[23] + 
                kernel_img_mul_27[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[223:216] <= 'd0;
  else if (current_state==ST_START)
    blur_din[223:216] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[223:216] <= 'd0;
end

wire  [39:0]  kernel_img_mul_28[0:24];
assign kernel_img_mul_28[0] = buffer_data_4[215:208] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_28[1] = buffer_data_4[223:216] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_28[2] = buffer_data_4[231:224] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_28[3] = buffer_data_4[239:232] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_28[4] = buffer_data_4[247:240] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_28[5] = buffer_data_3[215:208] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_28[6] = buffer_data_3[223:216] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_28[7] = buffer_data_3[231:224] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_28[8] = buffer_data_3[239:232] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_28[9] = buffer_data_3[247:240] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_28[10] = buffer_data_2[215:208] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_28[11] = buffer_data_2[223:216] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_28[12] = buffer_data_2[231:224] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_28[13] = buffer_data_2[239:232] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_28[14] = buffer_data_2[247:240] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_28[15] = buffer_data_1[215:208] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_28[16] = buffer_data_1[223:216] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_28[17] = buffer_data_1[231:224] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_28[18] = buffer_data_1[239:232] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_28[19] = buffer_data_1[247:240] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_28[20] = buffer_data_0[215:208] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_28[21] = buffer_data_0[223:216] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_28[22] = buffer_data_0[231:224] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_28[23] = buffer_data_0[239:232] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_28[24] = buffer_data_0[247:240] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_28 = kernel_img_mul_28[0] + kernel_img_mul_28[1] + kernel_img_mul_28[2] + 
                kernel_img_mul_28[3] + kernel_img_mul_28[4] + kernel_img_mul_28[5] + 
                kernel_img_mul_28[6] + kernel_img_mul_28[7] + kernel_img_mul_28[8] + 
                kernel_img_mul_28[9] + kernel_img_mul_28[10] + kernel_img_mul_28[11] + 
                kernel_img_mul_28[12] + kernel_img_mul_28[13] + kernel_img_mul_28[14] + 
                kernel_img_mul_28[15] + kernel_img_mul_28[16] + kernel_img_mul_28[17] + 
                kernel_img_mul_28[18] + kernel_img_mul_28[19] + kernel_img_mul_28[20] + 
                kernel_img_mul_28[21] + kernel_img_mul_28[22] + kernel_img_mul_28[23] + 
                kernel_img_mul_28[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[231:224] <= 'd0;
  else if (current_state==ST_START)
    blur_din[231:224] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[231:224] <= 'd0;
end

wire  [39:0]  kernel_img_mul_29[0:24];
assign kernel_img_mul_29[0] = buffer_data_4[223:216] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_29[1] = buffer_data_4[231:224] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_29[2] = buffer_data_4[239:232] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_29[3] = buffer_data_4[247:240] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_29[4] = buffer_data_4[255:248] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_29[5] = buffer_data_3[223:216] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_29[6] = buffer_data_3[231:224] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_29[7] = buffer_data_3[239:232] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_29[8] = buffer_data_3[247:240] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_29[9] = buffer_data_3[255:248] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_29[10] = buffer_data_2[223:216] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_29[11] = buffer_data_2[231:224] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_29[12] = buffer_data_2[239:232] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_29[13] = buffer_data_2[247:240] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_29[14] = buffer_data_2[255:248] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_29[15] = buffer_data_1[223:216] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_29[16] = buffer_data_1[231:224] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_29[17] = buffer_data_1[239:232] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_29[18] = buffer_data_1[247:240] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_29[19] = buffer_data_1[255:248] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_29[20] = buffer_data_0[223:216] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_29[21] = buffer_data_0[231:224] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_29[22] = buffer_data_0[239:232] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_29[23] = buffer_data_0[247:240] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_29[24] = buffer_data_0[255:248] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_29 = kernel_img_mul_29[0] + kernel_img_mul_29[1] + kernel_img_mul_29[2] + 
                kernel_img_mul_29[3] + kernel_img_mul_29[4] + kernel_img_mul_29[5] + 
                kernel_img_mul_29[6] + kernel_img_mul_29[7] + kernel_img_mul_29[8] + 
                kernel_img_mul_29[9] + kernel_img_mul_29[10] + kernel_img_mul_29[11] + 
                kernel_img_mul_29[12] + kernel_img_mul_29[13] + kernel_img_mul_29[14] + 
                kernel_img_mul_29[15] + kernel_img_mul_29[16] + kernel_img_mul_29[17] + 
                kernel_img_mul_29[18] + kernel_img_mul_29[19] + kernel_img_mul_29[20] + 
                kernel_img_mul_29[21] + kernel_img_mul_29[22] + kernel_img_mul_29[23] + 
                kernel_img_mul_29[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[239:232] <= 'd0;
  else if (current_state==ST_START)
    blur_din[239:232] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[239:232] <= 'd0;
end

wire  [39:0]  kernel_img_mul_30[0:24];
assign kernel_img_mul_30[0] = buffer_data_4[231:224] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_30[1] = buffer_data_4[239:232] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_30[2] = buffer_data_4[247:240] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_30[3] = buffer_data_4[255:248] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_30[4] = buffer_data_4[263:256] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_30[5] = buffer_data_3[231:224] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_30[6] = buffer_data_3[239:232] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_30[7] = buffer_data_3[247:240] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_30[8] = buffer_data_3[255:248] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_30[9] = buffer_data_3[263:256] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_30[10] = buffer_data_2[231:224] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_30[11] = buffer_data_2[239:232] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_30[12] = buffer_data_2[247:240] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_30[13] = buffer_data_2[255:248] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_30[14] = buffer_data_2[263:256] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_30[15] = buffer_data_1[231:224] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_30[16] = buffer_data_1[239:232] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_30[17] = buffer_data_1[247:240] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_30[18] = buffer_data_1[255:248] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_30[19] = buffer_data_1[263:256] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_30[20] = buffer_data_0[231:224] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_30[21] = buffer_data_0[239:232] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_30[22] = buffer_data_0[247:240] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_30[23] = buffer_data_0[255:248] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_30[24] = buffer_data_0[263:256] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_30 = kernel_img_mul_30[0] + kernel_img_mul_30[1] + kernel_img_mul_30[2] + 
                kernel_img_mul_30[3] + kernel_img_mul_30[4] + kernel_img_mul_30[5] + 
                kernel_img_mul_30[6] + kernel_img_mul_30[7] + kernel_img_mul_30[8] + 
                kernel_img_mul_30[9] + kernel_img_mul_30[10] + kernel_img_mul_30[11] + 
                kernel_img_mul_30[12] + kernel_img_mul_30[13] + kernel_img_mul_30[14] + 
                kernel_img_mul_30[15] + kernel_img_mul_30[16] + kernel_img_mul_30[17] + 
                kernel_img_mul_30[18] + kernel_img_mul_30[19] + kernel_img_mul_30[20] + 
                kernel_img_mul_30[21] + kernel_img_mul_30[22] + kernel_img_mul_30[23] + 
                kernel_img_mul_30[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[247:240] <= 'd0;
  else if (current_state==ST_START)
    blur_din[247:240] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[247:240] <= 'd0;
end

wire  [39:0]  kernel_img_mul_31[0:24];
assign kernel_img_mul_31[0] = buffer_data_4[239:232] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_31[1] = buffer_data_4[247:240] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_31[2] = buffer_data_4[255:248] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_31[3] = buffer_data_4[263:256] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_31[4] = buffer_data_4[271:264] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_31[5] = buffer_data_3[239:232] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_31[6] = buffer_data_3[247:240] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_31[7] = buffer_data_3[255:248] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_31[8] = buffer_data_3[263:256] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_31[9] = buffer_data_3[271:264] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_31[10] = buffer_data_2[239:232] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_31[11] = buffer_data_2[247:240] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_31[12] = buffer_data_2[255:248] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_31[13] = buffer_data_2[263:256] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_31[14] = buffer_data_2[271:264] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_31[15] = buffer_data_1[239:232] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_31[16] = buffer_data_1[247:240] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_31[17] = buffer_data_1[255:248] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_31[18] = buffer_data_1[263:256] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_31[19] = buffer_data_1[271:264] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_31[20] = buffer_data_0[239:232] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_31[21] = buffer_data_0[247:240] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_31[22] = buffer_data_0[255:248] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_31[23] = buffer_data_0[263:256] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_31[24] = buffer_data_0[271:264] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_31 = kernel_img_mul_31[0] + kernel_img_mul_31[1] + kernel_img_mul_31[2] + 
                kernel_img_mul_31[3] + kernel_img_mul_31[4] + kernel_img_mul_31[5] + 
                kernel_img_mul_31[6] + kernel_img_mul_31[7] + kernel_img_mul_31[8] + 
                kernel_img_mul_31[9] + kernel_img_mul_31[10] + kernel_img_mul_31[11] + 
                kernel_img_mul_31[12] + kernel_img_mul_31[13] + kernel_img_mul_31[14] + 
                kernel_img_mul_31[15] + kernel_img_mul_31[16] + kernel_img_mul_31[17] + 
                kernel_img_mul_31[18] + kernel_img_mul_31[19] + kernel_img_mul_31[20] + 
                kernel_img_mul_31[21] + kernel_img_mul_31[22] + kernel_img_mul_31[23] + 
                kernel_img_mul_31[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[255:248] <= 'd0;
  else if (current_state==ST_START)
    blur_din[255:248] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[255:248] <= 'd0;
end

wire  [39:0]  kernel_img_mul_32[0:24];
assign kernel_img_mul_32[0] = buffer_data_4[247:240] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_32[1] = buffer_data_4[255:248] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_32[2] = buffer_data_4[263:256] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_32[3] = buffer_data_4[271:264] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_32[4] = buffer_data_4[279:272] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_32[5] = buffer_data_3[247:240] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_32[6] = buffer_data_3[255:248] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_32[7] = buffer_data_3[263:256] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_32[8] = buffer_data_3[271:264] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_32[9] = buffer_data_3[279:272] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_32[10] = buffer_data_2[247:240] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_32[11] = buffer_data_2[255:248] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_32[12] = buffer_data_2[263:256] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_32[13] = buffer_data_2[271:264] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_32[14] = buffer_data_2[279:272] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_32[15] = buffer_data_1[247:240] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_32[16] = buffer_data_1[255:248] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_32[17] = buffer_data_1[263:256] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_32[18] = buffer_data_1[271:264] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_32[19] = buffer_data_1[279:272] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_32[20] = buffer_data_0[247:240] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_32[21] = buffer_data_0[255:248] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_32[22] = buffer_data_0[263:256] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_32[23] = buffer_data_0[271:264] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_32[24] = buffer_data_0[279:272] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_32 = kernel_img_mul_32[0] + kernel_img_mul_32[1] + kernel_img_mul_32[2] + 
                kernel_img_mul_32[3] + kernel_img_mul_32[4] + kernel_img_mul_32[5] + 
                kernel_img_mul_32[6] + kernel_img_mul_32[7] + kernel_img_mul_32[8] + 
                kernel_img_mul_32[9] + kernel_img_mul_32[10] + kernel_img_mul_32[11] + 
                kernel_img_mul_32[12] + kernel_img_mul_32[13] + kernel_img_mul_32[14] + 
                kernel_img_mul_32[15] + kernel_img_mul_32[16] + kernel_img_mul_32[17] + 
                kernel_img_mul_32[18] + kernel_img_mul_32[19] + kernel_img_mul_32[20] + 
                kernel_img_mul_32[21] + kernel_img_mul_32[22] + kernel_img_mul_32[23] + 
                kernel_img_mul_32[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[263:256] <= 'd0;
  else if (current_state==ST_START)
    blur_din[263:256] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[263:256] <= 'd0;
end

wire  [39:0]  kernel_img_mul_33[0:24];
assign kernel_img_mul_33[0] = buffer_data_4[255:248] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_33[1] = buffer_data_4[263:256] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_33[2] = buffer_data_4[271:264] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_33[3] = buffer_data_4[279:272] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_33[4] = buffer_data_4[287:280] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_33[5] = buffer_data_3[255:248] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_33[6] = buffer_data_3[263:256] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_33[7] = buffer_data_3[271:264] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_33[8] = buffer_data_3[279:272] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_33[9] = buffer_data_3[287:280] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_33[10] = buffer_data_2[255:248] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_33[11] = buffer_data_2[263:256] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_33[12] = buffer_data_2[271:264] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_33[13] = buffer_data_2[279:272] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_33[14] = buffer_data_2[287:280] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_33[15] = buffer_data_1[255:248] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_33[16] = buffer_data_1[263:256] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_33[17] = buffer_data_1[271:264] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_33[18] = buffer_data_1[279:272] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_33[19] = buffer_data_1[287:280] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_33[20] = buffer_data_0[255:248] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_33[21] = buffer_data_0[263:256] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_33[22] = buffer_data_0[271:264] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_33[23] = buffer_data_0[279:272] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_33[24] = buffer_data_0[287:280] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_33 = kernel_img_mul_33[0] + kernel_img_mul_33[1] + kernel_img_mul_33[2] + 
                kernel_img_mul_33[3] + kernel_img_mul_33[4] + kernel_img_mul_33[5] + 
                kernel_img_mul_33[6] + kernel_img_mul_33[7] + kernel_img_mul_33[8] + 
                kernel_img_mul_33[9] + kernel_img_mul_33[10] + kernel_img_mul_33[11] + 
                kernel_img_mul_33[12] + kernel_img_mul_33[13] + kernel_img_mul_33[14] + 
                kernel_img_mul_33[15] + kernel_img_mul_33[16] + kernel_img_mul_33[17] + 
                kernel_img_mul_33[18] + kernel_img_mul_33[19] + kernel_img_mul_33[20] + 
                kernel_img_mul_33[21] + kernel_img_mul_33[22] + kernel_img_mul_33[23] + 
                kernel_img_mul_33[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[271:264] <= 'd0;
  else if (current_state==ST_START)
    blur_din[271:264] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[271:264] <= 'd0;
end

wire  [39:0]  kernel_img_mul_34[0:24];
assign kernel_img_mul_34[0] = buffer_data_4[263:256] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_34[1] = buffer_data_4[271:264] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_34[2] = buffer_data_4[279:272] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_34[3] = buffer_data_4[287:280] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_34[4] = buffer_data_4[295:288] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_34[5] = buffer_data_3[263:256] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_34[6] = buffer_data_3[271:264] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_34[7] = buffer_data_3[279:272] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_34[8] = buffer_data_3[287:280] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_34[9] = buffer_data_3[295:288] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_34[10] = buffer_data_2[263:256] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_34[11] = buffer_data_2[271:264] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_34[12] = buffer_data_2[279:272] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_34[13] = buffer_data_2[287:280] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_34[14] = buffer_data_2[295:288] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_34[15] = buffer_data_1[263:256] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_34[16] = buffer_data_1[271:264] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_34[17] = buffer_data_1[279:272] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_34[18] = buffer_data_1[287:280] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_34[19] = buffer_data_1[295:288] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_34[20] = buffer_data_0[263:256] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_34[21] = buffer_data_0[271:264] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_34[22] = buffer_data_0[279:272] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_34[23] = buffer_data_0[287:280] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_34[24] = buffer_data_0[295:288] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_34 = kernel_img_mul_34[0] + kernel_img_mul_34[1] + kernel_img_mul_34[2] + 
                kernel_img_mul_34[3] + kernel_img_mul_34[4] + kernel_img_mul_34[5] + 
                kernel_img_mul_34[6] + kernel_img_mul_34[7] + kernel_img_mul_34[8] + 
                kernel_img_mul_34[9] + kernel_img_mul_34[10] + kernel_img_mul_34[11] + 
                kernel_img_mul_34[12] + kernel_img_mul_34[13] + kernel_img_mul_34[14] + 
                kernel_img_mul_34[15] + kernel_img_mul_34[16] + kernel_img_mul_34[17] + 
                kernel_img_mul_34[18] + kernel_img_mul_34[19] + kernel_img_mul_34[20] + 
                kernel_img_mul_34[21] + kernel_img_mul_34[22] + kernel_img_mul_34[23] + 
                kernel_img_mul_34[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[279:272] <= 'd0;
  else if (current_state==ST_START)
    blur_din[279:272] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[279:272] <= 'd0;
end

wire  [39:0]  kernel_img_mul_35[0:24];
assign kernel_img_mul_35[0] = buffer_data_4[271:264] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_35[1] = buffer_data_4[279:272] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_35[2] = buffer_data_4[287:280] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_35[3] = buffer_data_4[295:288] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_35[4] = buffer_data_4[303:296] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_35[5] = buffer_data_3[271:264] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_35[6] = buffer_data_3[279:272] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_35[7] = buffer_data_3[287:280] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_35[8] = buffer_data_3[295:288] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_35[9] = buffer_data_3[303:296] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_35[10] = buffer_data_2[271:264] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_35[11] = buffer_data_2[279:272] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_35[12] = buffer_data_2[287:280] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_35[13] = buffer_data_2[295:288] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_35[14] = buffer_data_2[303:296] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_35[15] = buffer_data_1[271:264] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_35[16] = buffer_data_1[279:272] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_35[17] = buffer_data_1[287:280] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_35[18] = buffer_data_1[295:288] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_35[19] = buffer_data_1[303:296] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_35[20] = buffer_data_0[271:264] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_35[21] = buffer_data_0[279:272] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_35[22] = buffer_data_0[287:280] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_35[23] = buffer_data_0[295:288] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_35[24] = buffer_data_0[303:296] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_35 = kernel_img_mul_35[0] + kernel_img_mul_35[1] + kernel_img_mul_35[2] + 
                kernel_img_mul_35[3] + kernel_img_mul_35[4] + kernel_img_mul_35[5] + 
                kernel_img_mul_35[6] + kernel_img_mul_35[7] + kernel_img_mul_35[8] + 
                kernel_img_mul_35[9] + kernel_img_mul_35[10] + kernel_img_mul_35[11] + 
                kernel_img_mul_35[12] + kernel_img_mul_35[13] + kernel_img_mul_35[14] + 
                kernel_img_mul_35[15] + kernel_img_mul_35[16] + kernel_img_mul_35[17] + 
                kernel_img_mul_35[18] + kernel_img_mul_35[19] + kernel_img_mul_35[20] + 
                kernel_img_mul_35[21] + kernel_img_mul_35[22] + kernel_img_mul_35[23] + 
                kernel_img_mul_35[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[287:280] <= 'd0;
  else if (current_state==ST_START)
    blur_din[287:280] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[287:280] <= 'd0;
end

wire  [39:0]  kernel_img_mul_36[0:24];
assign kernel_img_mul_36[0] = buffer_data_4[279:272] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_36[1] = buffer_data_4[287:280] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_36[2] = buffer_data_4[295:288] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_36[3] = buffer_data_4[303:296] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_36[4] = buffer_data_4[311:304] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_36[5] = buffer_data_3[279:272] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_36[6] = buffer_data_3[287:280] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_36[7] = buffer_data_3[295:288] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_36[8] = buffer_data_3[303:296] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_36[9] = buffer_data_3[311:304] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_36[10] = buffer_data_2[279:272] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_36[11] = buffer_data_2[287:280] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_36[12] = buffer_data_2[295:288] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_36[13] = buffer_data_2[303:296] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_36[14] = buffer_data_2[311:304] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_36[15] = buffer_data_1[279:272] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_36[16] = buffer_data_1[287:280] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_36[17] = buffer_data_1[295:288] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_36[18] = buffer_data_1[303:296] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_36[19] = buffer_data_1[311:304] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_36[20] = buffer_data_0[279:272] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_36[21] = buffer_data_0[287:280] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_36[22] = buffer_data_0[295:288] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_36[23] = buffer_data_0[303:296] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_36[24] = buffer_data_0[311:304] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_36 = kernel_img_mul_36[0] + kernel_img_mul_36[1] + kernel_img_mul_36[2] + 
                kernel_img_mul_36[3] + kernel_img_mul_36[4] + kernel_img_mul_36[5] + 
                kernel_img_mul_36[6] + kernel_img_mul_36[7] + kernel_img_mul_36[8] + 
                kernel_img_mul_36[9] + kernel_img_mul_36[10] + kernel_img_mul_36[11] + 
                kernel_img_mul_36[12] + kernel_img_mul_36[13] + kernel_img_mul_36[14] + 
                kernel_img_mul_36[15] + kernel_img_mul_36[16] + kernel_img_mul_36[17] + 
                kernel_img_mul_36[18] + kernel_img_mul_36[19] + kernel_img_mul_36[20] + 
                kernel_img_mul_36[21] + kernel_img_mul_36[22] + kernel_img_mul_36[23] + 
                kernel_img_mul_36[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[295:288] <= 'd0;
  else if (current_state==ST_START)
    blur_din[295:288] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[295:288] <= 'd0;
end

wire  [39:0]  kernel_img_mul_37[0:24];
assign kernel_img_mul_37[0] = buffer_data_4[287:280] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_37[1] = buffer_data_4[295:288] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_37[2] = buffer_data_4[303:296] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_37[3] = buffer_data_4[311:304] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_37[4] = buffer_data_4[319:312] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_37[5] = buffer_data_3[287:280] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_37[6] = buffer_data_3[295:288] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_37[7] = buffer_data_3[303:296] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_37[8] = buffer_data_3[311:304] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_37[9] = buffer_data_3[319:312] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_37[10] = buffer_data_2[287:280] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_37[11] = buffer_data_2[295:288] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_37[12] = buffer_data_2[303:296] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_37[13] = buffer_data_2[311:304] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_37[14] = buffer_data_2[319:312] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_37[15] = buffer_data_1[287:280] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_37[16] = buffer_data_1[295:288] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_37[17] = buffer_data_1[303:296] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_37[18] = buffer_data_1[311:304] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_37[19] = buffer_data_1[319:312] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_37[20] = buffer_data_0[287:280] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_37[21] = buffer_data_0[295:288] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_37[22] = buffer_data_0[303:296] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_37[23] = buffer_data_0[311:304] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_37[24] = buffer_data_0[319:312] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_37 = kernel_img_mul_37[0] + kernel_img_mul_37[1] + kernel_img_mul_37[2] + 
                kernel_img_mul_37[3] + kernel_img_mul_37[4] + kernel_img_mul_37[5] + 
                kernel_img_mul_37[6] + kernel_img_mul_37[7] + kernel_img_mul_37[8] + 
                kernel_img_mul_37[9] + kernel_img_mul_37[10] + kernel_img_mul_37[11] + 
                kernel_img_mul_37[12] + kernel_img_mul_37[13] + kernel_img_mul_37[14] + 
                kernel_img_mul_37[15] + kernel_img_mul_37[16] + kernel_img_mul_37[17] + 
                kernel_img_mul_37[18] + kernel_img_mul_37[19] + kernel_img_mul_37[20] + 
                kernel_img_mul_37[21] + kernel_img_mul_37[22] + kernel_img_mul_37[23] + 
                kernel_img_mul_37[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[303:296] <= 'd0;
  else if (current_state==ST_START)
    blur_din[303:296] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[303:296] <= 'd0;
end

wire  [39:0]  kernel_img_mul_38[0:24];
assign kernel_img_mul_38[0] = buffer_data_4[295:288] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_38[1] = buffer_data_4[303:296] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_38[2] = buffer_data_4[311:304] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_38[3] = buffer_data_4[319:312] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_38[4] = buffer_data_4[327:320] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_38[5] = buffer_data_3[295:288] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_38[6] = buffer_data_3[303:296] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_38[7] = buffer_data_3[311:304] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_38[8] = buffer_data_3[319:312] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_38[9] = buffer_data_3[327:320] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_38[10] = buffer_data_2[295:288] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_38[11] = buffer_data_2[303:296] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_38[12] = buffer_data_2[311:304] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_38[13] = buffer_data_2[319:312] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_38[14] = buffer_data_2[327:320] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_38[15] = buffer_data_1[295:288] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_38[16] = buffer_data_1[303:296] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_38[17] = buffer_data_1[311:304] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_38[18] = buffer_data_1[319:312] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_38[19] = buffer_data_1[327:320] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_38[20] = buffer_data_0[295:288] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_38[21] = buffer_data_0[303:296] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_38[22] = buffer_data_0[311:304] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_38[23] = buffer_data_0[319:312] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_38[24] = buffer_data_0[327:320] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_38 = kernel_img_mul_38[0] + kernel_img_mul_38[1] + kernel_img_mul_38[2] + 
                kernel_img_mul_38[3] + kernel_img_mul_38[4] + kernel_img_mul_38[5] + 
                kernel_img_mul_38[6] + kernel_img_mul_38[7] + kernel_img_mul_38[8] + 
                kernel_img_mul_38[9] + kernel_img_mul_38[10] + kernel_img_mul_38[11] + 
                kernel_img_mul_38[12] + kernel_img_mul_38[13] + kernel_img_mul_38[14] + 
                kernel_img_mul_38[15] + kernel_img_mul_38[16] + kernel_img_mul_38[17] + 
                kernel_img_mul_38[18] + kernel_img_mul_38[19] + kernel_img_mul_38[20] + 
                kernel_img_mul_38[21] + kernel_img_mul_38[22] + kernel_img_mul_38[23] + 
                kernel_img_mul_38[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[311:304] <= 'd0;
  else if (current_state==ST_START)
    blur_din[311:304] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[311:304] <= 'd0;
end

wire  [39:0]  kernel_img_mul_39[0:24];
assign kernel_img_mul_39[0] = buffer_data_4[303:296] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_39[1] = buffer_data_4[311:304] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_39[2] = buffer_data_4[319:312] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_39[3] = buffer_data_4[327:320] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_39[4] = buffer_data_4[335:328] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_39[5] = buffer_data_3[303:296] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_39[6] = buffer_data_3[311:304] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_39[7] = buffer_data_3[319:312] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_39[8] = buffer_data_3[327:320] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_39[9] = buffer_data_3[335:328] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_39[10] = buffer_data_2[303:296] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_39[11] = buffer_data_2[311:304] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_39[12] = buffer_data_2[319:312] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_39[13] = buffer_data_2[327:320] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_39[14] = buffer_data_2[335:328] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_39[15] = buffer_data_1[303:296] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_39[16] = buffer_data_1[311:304] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_39[17] = buffer_data_1[319:312] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_39[18] = buffer_data_1[327:320] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_39[19] = buffer_data_1[335:328] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_39[20] = buffer_data_0[303:296] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_39[21] = buffer_data_0[311:304] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_39[22] = buffer_data_0[319:312] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_39[23] = buffer_data_0[327:320] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_39[24] = buffer_data_0[335:328] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_39 = kernel_img_mul_39[0] + kernel_img_mul_39[1] + kernel_img_mul_39[2] + 
                kernel_img_mul_39[3] + kernel_img_mul_39[4] + kernel_img_mul_39[5] + 
                kernel_img_mul_39[6] + kernel_img_mul_39[7] + kernel_img_mul_39[8] + 
                kernel_img_mul_39[9] + kernel_img_mul_39[10] + kernel_img_mul_39[11] + 
                kernel_img_mul_39[12] + kernel_img_mul_39[13] + kernel_img_mul_39[14] + 
                kernel_img_mul_39[15] + kernel_img_mul_39[16] + kernel_img_mul_39[17] + 
                kernel_img_mul_39[18] + kernel_img_mul_39[19] + kernel_img_mul_39[20] + 
                kernel_img_mul_39[21] + kernel_img_mul_39[22] + kernel_img_mul_39[23] + 
                kernel_img_mul_39[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[319:312] <= 'd0;
  else if (current_state==ST_START)
    blur_din[319:312] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[319:312] <= 'd0;
end

wire  [39:0]  kernel_img_mul_40[0:24];
assign kernel_img_mul_40[0] = buffer_data_4[311:304] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_40[1] = buffer_data_4[319:312] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_40[2] = buffer_data_4[327:320] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_40[3] = buffer_data_4[335:328] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_40[4] = buffer_data_4[343:336] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_40[5] = buffer_data_3[311:304] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_40[6] = buffer_data_3[319:312] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_40[7] = buffer_data_3[327:320] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_40[8] = buffer_data_3[335:328] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_40[9] = buffer_data_3[343:336] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_40[10] = buffer_data_2[311:304] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_40[11] = buffer_data_2[319:312] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_40[12] = buffer_data_2[327:320] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_40[13] = buffer_data_2[335:328] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_40[14] = buffer_data_2[343:336] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_40[15] = buffer_data_1[311:304] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_40[16] = buffer_data_1[319:312] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_40[17] = buffer_data_1[327:320] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_40[18] = buffer_data_1[335:328] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_40[19] = buffer_data_1[343:336] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_40[20] = buffer_data_0[311:304] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_40[21] = buffer_data_0[319:312] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_40[22] = buffer_data_0[327:320] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_40[23] = buffer_data_0[335:328] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_40[24] = buffer_data_0[343:336] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_40 = kernel_img_mul_40[0] + kernel_img_mul_40[1] + kernel_img_mul_40[2] + 
                kernel_img_mul_40[3] + kernel_img_mul_40[4] + kernel_img_mul_40[5] + 
                kernel_img_mul_40[6] + kernel_img_mul_40[7] + kernel_img_mul_40[8] + 
                kernel_img_mul_40[9] + kernel_img_mul_40[10] + kernel_img_mul_40[11] + 
                kernel_img_mul_40[12] + kernel_img_mul_40[13] + kernel_img_mul_40[14] + 
                kernel_img_mul_40[15] + kernel_img_mul_40[16] + kernel_img_mul_40[17] + 
                kernel_img_mul_40[18] + kernel_img_mul_40[19] + kernel_img_mul_40[20] + 
                kernel_img_mul_40[21] + kernel_img_mul_40[22] + kernel_img_mul_40[23] + 
                kernel_img_mul_40[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[327:320] <= 'd0;
  else if (current_state==ST_START)
    blur_din[327:320] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[327:320] <= 'd0;
end

wire  [39:0]  kernel_img_mul_41[0:24];
assign kernel_img_mul_41[0] = buffer_data_4[319:312] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_41[1] = buffer_data_4[327:320] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_41[2] = buffer_data_4[335:328] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_41[3] = buffer_data_4[343:336] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_41[4] = buffer_data_4[351:344] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_41[5] = buffer_data_3[319:312] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_41[6] = buffer_data_3[327:320] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_41[7] = buffer_data_3[335:328] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_41[8] = buffer_data_3[343:336] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_41[9] = buffer_data_3[351:344] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_41[10] = buffer_data_2[319:312] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_41[11] = buffer_data_2[327:320] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_41[12] = buffer_data_2[335:328] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_41[13] = buffer_data_2[343:336] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_41[14] = buffer_data_2[351:344] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_41[15] = buffer_data_1[319:312] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_41[16] = buffer_data_1[327:320] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_41[17] = buffer_data_1[335:328] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_41[18] = buffer_data_1[343:336] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_41[19] = buffer_data_1[351:344] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_41[20] = buffer_data_0[319:312] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_41[21] = buffer_data_0[327:320] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_41[22] = buffer_data_0[335:328] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_41[23] = buffer_data_0[343:336] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_41[24] = buffer_data_0[351:344] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_41 = kernel_img_mul_41[0] + kernel_img_mul_41[1] + kernel_img_mul_41[2] + 
                kernel_img_mul_41[3] + kernel_img_mul_41[4] + kernel_img_mul_41[5] + 
                kernel_img_mul_41[6] + kernel_img_mul_41[7] + kernel_img_mul_41[8] + 
                kernel_img_mul_41[9] + kernel_img_mul_41[10] + kernel_img_mul_41[11] + 
                kernel_img_mul_41[12] + kernel_img_mul_41[13] + kernel_img_mul_41[14] + 
                kernel_img_mul_41[15] + kernel_img_mul_41[16] + kernel_img_mul_41[17] + 
                kernel_img_mul_41[18] + kernel_img_mul_41[19] + kernel_img_mul_41[20] + 
                kernel_img_mul_41[21] + kernel_img_mul_41[22] + kernel_img_mul_41[23] + 
                kernel_img_mul_41[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[335:328] <= 'd0;
  else if (current_state==ST_START)
    blur_din[335:328] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[335:328] <= 'd0;
end

wire  [39:0]  kernel_img_mul_42[0:24];
assign kernel_img_mul_42[0] = buffer_data_4[327:320] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_42[1] = buffer_data_4[335:328] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_42[2] = buffer_data_4[343:336] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_42[3] = buffer_data_4[351:344] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_42[4] = buffer_data_4[359:352] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_42[5] = buffer_data_3[327:320] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_42[6] = buffer_data_3[335:328] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_42[7] = buffer_data_3[343:336] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_42[8] = buffer_data_3[351:344] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_42[9] = buffer_data_3[359:352] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_42[10] = buffer_data_2[327:320] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_42[11] = buffer_data_2[335:328] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_42[12] = buffer_data_2[343:336] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_42[13] = buffer_data_2[351:344] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_42[14] = buffer_data_2[359:352] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_42[15] = buffer_data_1[327:320] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_42[16] = buffer_data_1[335:328] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_42[17] = buffer_data_1[343:336] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_42[18] = buffer_data_1[351:344] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_42[19] = buffer_data_1[359:352] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_42[20] = buffer_data_0[327:320] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_42[21] = buffer_data_0[335:328] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_42[22] = buffer_data_0[343:336] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_42[23] = buffer_data_0[351:344] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_42[24] = buffer_data_0[359:352] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_42 = kernel_img_mul_42[0] + kernel_img_mul_42[1] + kernel_img_mul_42[2] + 
                kernel_img_mul_42[3] + kernel_img_mul_42[4] + kernel_img_mul_42[5] + 
                kernel_img_mul_42[6] + kernel_img_mul_42[7] + kernel_img_mul_42[8] + 
                kernel_img_mul_42[9] + kernel_img_mul_42[10] + kernel_img_mul_42[11] + 
                kernel_img_mul_42[12] + kernel_img_mul_42[13] + kernel_img_mul_42[14] + 
                kernel_img_mul_42[15] + kernel_img_mul_42[16] + kernel_img_mul_42[17] + 
                kernel_img_mul_42[18] + kernel_img_mul_42[19] + kernel_img_mul_42[20] + 
                kernel_img_mul_42[21] + kernel_img_mul_42[22] + kernel_img_mul_42[23] + 
                kernel_img_mul_42[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[343:336] <= 'd0;
  else if (current_state==ST_START)
    blur_din[343:336] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[343:336] <= 'd0;
end

wire  [39:0]  kernel_img_mul_43[0:24];
assign kernel_img_mul_43[0] = buffer_data_4[335:328] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_43[1] = buffer_data_4[343:336] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_43[2] = buffer_data_4[351:344] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_43[3] = buffer_data_4[359:352] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_43[4] = buffer_data_4[367:360] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_43[5] = buffer_data_3[335:328] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_43[6] = buffer_data_3[343:336] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_43[7] = buffer_data_3[351:344] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_43[8] = buffer_data_3[359:352] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_43[9] = buffer_data_3[367:360] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_43[10] = buffer_data_2[335:328] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_43[11] = buffer_data_2[343:336] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_43[12] = buffer_data_2[351:344] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_43[13] = buffer_data_2[359:352] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_43[14] = buffer_data_2[367:360] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_43[15] = buffer_data_1[335:328] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_43[16] = buffer_data_1[343:336] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_43[17] = buffer_data_1[351:344] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_43[18] = buffer_data_1[359:352] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_43[19] = buffer_data_1[367:360] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_43[20] = buffer_data_0[335:328] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_43[21] = buffer_data_0[343:336] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_43[22] = buffer_data_0[351:344] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_43[23] = buffer_data_0[359:352] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_43[24] = buffer_data_0[367:360] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_43 = kernel_img_mul_43[0] + kernel_img_mul_43[1] + kernel_img_mul_43[2] + 
                kernel_img_mul_43[3] + kernel_img_mul_43[4] + kernel_img_mul_43[5] + 
                kernel_img_mul_43[6] + kernel_img_mul_43[7] + kernel_img_mul_43[8] + 
                kernel_img_mul_43[9] + kernel_img_mul_43[10] + kernel_img_mul_43[11] + 
                kernel_img_mul_43[12] + kernel_img_mul_43[13] + kernel_img_mul_43[14] + 
                kernel_img_mul_43[15] + kernel_img_mul_43[16] + kernel_img_mul_43[17] + 
                kernel_img_mul_43[18] + kernel_img_mul_43[19] + kernel_img_mul_43[20] + 
                kernel_img_mul_43[21] + kernel_img_mul_43[22] + kernel_img_mul_43[23] + 
                kernel_img_mul_43[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[351:344] <= 'd0;
  else if (current_state==ST_START)
    blur_din[351:344] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[351:344] <= 'd0;
end

wire  [39:0]  kernel_img_mul_44[0:24];
assign kernel_img_mul_44[0] = buffer_data_4[343:336] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_44[1] = buffer_data_4[351:344] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_44[2] = buffer_data_4[359:352] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_44[3] = buffer_data_4[367:360] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_44[4] = buffer_data_4[375:368] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_44[5] = buffer_data_3[343:336] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_44[6] = buffer_data_3[351:344] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_44[7] = buffer_data_3[359:352] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_44[8] = buffer_data_3[367:360] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_44[9] = buffer_data_3[375:368] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_44[10] = buffer_data_2[343:336] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_44[11] = buffer_data_2[351:344] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_44[12] = buffer_data_2[359:352] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_44[13] = buffer_data_2[367:360] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_44[14] = buffer_data_2[375:368] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_44[15] = buffer_data_1[343:336] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_44[16] = buffer_data_1[351:344] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_44[17] = buffer_data_1[359:352] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_44[18] = buffer_data_1[367:360] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_44[19] = buffer_data_1[375:368] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_44[20] = buffer_data_0[343:336] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_44[21] = buffer_data_0[351:344] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_44[22] = buffer_data_0[359:352] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_44[23] = buffer_data_0[367:360] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_44[24] = buffer_data_0[375:368] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_44 = kernel_img_mul_44[0] + kernel_img_mul_44[1] + kernel_img_mul_44[2] + 
                kernel_img_mul_44[3] + kernel_img_mul_44[4] + kernel_img_mul_44[5] + 
                kernel_img_mul_44[6] + kernel_img_mul_44[7] + kernel_img_mul_44[8] + 
                kernel_img_mul_44[9] + kernel_img_mul_44[10] + kernel_img_mul_44[11] + 
                kernel_img_mul_44[12] + kernel_img_mul_44[13] + kernel_img_mul_44[14] + 
                kernel_img_mul_44[15] + kernel_img_mul_44[16] + kernel_img_mul_44[17] + 
                kernel_img_mul_44[18] + kernel_img_mul_44[19] + kernel_img_mul_44[20] + 
                kernel_img_mul_44[21] + kernel_img_mul_44[22] + kernel_img_mul_44[23] + 
                kernel_img_mul_44[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[359:352] <= 'd0;
  else if (current_state==ST_START)
    blur_din[359:352] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[359:352] <= 'd0;
end

wire  [39:0]  kernel_img_mul_45[0:24];
assign kernel_img_mul_45[0] = buffer_data_4[351:344] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_45[1] = buffer_data_4[359:352] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_45[2] = buffer_data_4[367:360] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_45[3] = buffer_data_4[375:368] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_45[4] = buffer_data_4[383:376] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_45[5] = buffer_data_3[351:344] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_45[6] = buffer_data_3[359:352] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_45[7] = buffer_data_3[367:360] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_45[8] = buffer_data_3[375:368] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_45[9] = buffer_data_3[383:376] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_45[10] = buffer_data_2[351:344] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_45[11] = buffer_data_2[359:352] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_45[12] = buffer_data_2[367:360] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_45[13] = buffer_data_2[375:368] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_45[14] = buffer_data_2[383:376] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_45[15] = buffer_data_1[351:344] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_45[16] = buffer_data_1[359:352] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_45[17] = buffer_data_1[367:360] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_45[18] = buffer_data_1[375:368] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_45[19] = buffer_data_1[383:376] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_45[20] = buffer_data_0[351:344] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_45[21] = buffer_data_0[359:352] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_45[22] = buffer_data_0[367:360] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_45[23] = buffer_data_0[375:368] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_45[24] = buffer_data_0[383:376] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_45 = kernel_img_mul_45[0] + kernel_img_mul_45[1] + kernel_img_mul_45[2] + 
                kernel_img_mul_45[3] + kernel_img_mul_45[4] + kernel_img_mul_45[5] + 
                kernel_img_mul_45[6] + kernel_img_mul_45[7] + kernel_img_mul_45[8] + 
                kernel_img_mul_45[9] + kernel_img_mul_45[10] + kernel_img_mul_45[11] + 
                kernel_img_mul_45[12] + kernel_img_mul_45[13] + kernel_img_mul_45[14] + 
                kernel_img_mul_45[15] + kernel_img_mul_45[16] + kernel_img_mul_45[17] + 
                kernel_img_mul_45[18] + kernel_img_mul_45[19] + kernel_img_mul_45[20] + 
                kernel_img_mul_45[21] + kernel_img_mul_45[22] + kernel_img_mul_45[23] + 
                kernel_img_mul_45[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[367:360] <= 'd0;
  else if (current_state==ST_START)
    blur_din[367:360] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[367:360] <= 'd0;
end

wire  [39:0]  kernel_img_mul_46[0:24];
assign kernel_img_mul_46[0] = buffer_data_4[359:352] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_46[1] = buffer_data_4[367:360] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_46[2] = buffer_data_4[375:368] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_46[3] = buffer_data_4[383:376] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_46[4] = buffer_data_4[391:384] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_46[5] = buffer_data_3[359:352] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_46[6] = buffer_data_3[367:360] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_46[7] = buffer_data_3[375:368] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_46[8] = buffer_data_3[383:376] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_46[9] = buffer_data_3[391:384] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_46[10] = buffer_data_2[359:352] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_46[11] = buffer_data_2[367:360] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_46[12] = buffer_data_2[375:368] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_46[13] = buffer_data_2[383:376] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_46[14] = buffer_data_2[391:384] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_46[15] = buffer_data_1[359:352] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_46[16] = buffer_data_1[367:360] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_46[17] = buffer_data_1[375:368] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_46[18] = buffer_data_1[383:376] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_46[19] = buffer_data_1[391:384] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_46[20] = buffer_data_0[359:352] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_46[21] = buffer_data_0[367:360] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_46[22] = buffer_data_0[375:368] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_46[23] = buffer_data_0[383:376] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_46[24] = buffer_data_0[391:384] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_46 = kernel_img_mul_46[0] + kernel_img_mul_46[1] + kernel_img_mul_46[2] + 
                kernel_img_mul_46[3] + kernel_img_mul_46[4] + kernel_img_mul_46[5] + 
                kernel_img_mul_46[6] + kernel_img_mul_46[7] + kernel_img_mul_46[8] + 
                kernel_img_mul_46[9] + kernel_img_mul_46[10] + kernel_img_mul_46[11] + 
                kernel_img_mul_46[12] + kernel_img_mul_46[13] + kernel_img_mul_46[14] + 
                kernel_img_mul_46[15] + kernel_img_mul_46[16] + kernel_img_mul_46[17] + 
                kernel_img_mul_46[18] + kernel_img_mul_46[19] + kernel_img_mul_46[20] + 
                kernel_img_mul_46[21] + kernel_img_mul_46[22] + kernel_img_mul_46[23] + 
                kernel_img_mul_46[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[375:368] <= 'd0;
  else if (current_state==ST_START)
    blur_din[375:368] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[375:368] <= 'd0;
end

wire  [39:0]  kernel_img_mul_47[0:24];
assign kernel_img_mul_47[0] = buffer_data_4[367:360] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_47[1] = buffer_data_4[375:368] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_47[2] = buffer_data_4[383:376] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_47[3] = buffer_data_4[391:384] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_47[4] = buffer_data_4[399:392] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_47[5] = buffer_data_3[367:360] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_47[6] = buffer_data_3[375:368] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_47[7] = buffer_data_3[383:376] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_47[8] = buffer_data_3[391:384] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_47[9] = buffer_data_3[399:392] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_47[10] = buffer_data_2[367:360] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_47[11] = buffer_data_2[375:368] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_47[12] = buffer_data_2[383:376] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_47[13] = buffer_data_2[391:384] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_47[14] = buffer_data_2[399:392] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_47[15] = buffer_data_1[367:360] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_47[16] = buffer_data_1[375:368] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_47[17] = buffer_data_1[383:376] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_47[18] = buffer_data_1[391:384] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_47[19] = buffer_data_1[399:392] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_47[20] = buffer_data_0[367:360] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_47[21] = buffer_data_0[375:368] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_47[22] = buffer_data_0[383:376] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_47[23] = buffer_data_0[391:384] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_47[24] = buffer_data_0[399:392] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_47 = kernel_img_mul_47[0] + kernel_img_mul_47[1] + kernel_img_mul_47[2] + 
                kernel_img_mul_47[3] + kernel_img_mul_47[4] + kernel_img_mul_47[5] + 
                kernel_img_mul_47[6] + kernel_img_mul_47[7] + kernel_img_mul_47[8] + 
                kernel_img_mul_47[9] + kernel_img_mul_47[10] + kernel_img_mul_47[11] + 
                kernel_img_mul_47[12] + kernel_img_mul_47[13] + kernel_img_mul_47[14] + 
                kernel_img_mul_47[15] + kernel_img_mul_47[16] + kernel_img_mul_47[17] + 
                kernel_img_mul_47[18] + kernel_img_mul_47[19] + kernel_img_mul_47[20] + 
                kernel_img_mul_47[21] + kernel_img_mul_47[22] + kernel_img_mul_47[23] + 
                kernel_img_mul_47[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[383:376] <= 'd0;
  else if (current_state==ST_START)
    blur_din[383:376] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[383:376] <= 'd0;
end

wire  [39:0]  kernel_img_mul_48[0:24];
assign kernel_img_mul_48[0] = buffer_data_4[375:368] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_48[1] = buffer_data_4[383:376] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_48[2] = buffer_data_4[391:384] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_48[3] = buffer_data_4[399:392] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_48[4] = buffer_data_4[407:400] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_48[5] = buffer_data_3[375:368] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_48[6] = buffer_data_3[383:376] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_48[7] = buffer_data_3[391:384] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_48[8] = buffer_data_3[399:392] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_48[9] = buffer_data_3[407:400] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_48[10] = buffer_data_2[375:368] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_48[11] = buffer_data_2[383:376] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_48[12] = buffer_data_2[391:384] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_48[13] = buffer_data_2[399:392] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_48[14] = buffer_data_2[407:400] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_48[15] = buffer_data_1[375:368] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_48[16] = buffer_data_1[383:376] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_48[17] = buffer_data_1[391:384] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_48[18] = buffer_data_1[399:392] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_48[19] = buffer_data_1[407:400] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_48[20] = buffer_data_0[375:368] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_48[21] = buffer_data_0[383:376] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_48[22] = buffer_data_0[391:384] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_48[23] = buffer_data_0[399:392] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_48[24] = buffer_data_0[407:400] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_48 = kernel_img_mul_48[0] + kernel_img_mul_48[1] + kernel_img_mul_48[2] + 
                kernel_img_mul_48[3] + kernel_img_mul_48[4] + kernel_img_mul_48[5] + 
                kernel_img_mul_48[6] + kernel_img_mul_48[7] + kernel_img_mul_48[8] + 
                kernel_img_mul_48[9] + kernel_img_mul_48[10] + kernel_img_mul_48[11] + 
                kernel_img_mul_48[12] + kernel_img_mul_48[13] + kernel_img_mul_48[14] + 
                kernel_img_mul_48[15] + kernel_img_mul_48[16] + kernel_img_mul_48[17] + 
                kernel_img_mul_48[18] + kernel_img_mul_48[19] + kernel_img_mul_48[20] + 
                kernel_img_mul_48[21] + kernel_img_mul_48[22] + kernel_img_mul_48[23] + 
                kernel_img_mul_48[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[391:384] <= 'd0;
  else if (current_state==ST_START)
    blur_din[391:384] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[391:384] <= 'd0;
end

wire  [39:0]  kernel_img_mul_49[0:24];
assign kernel_img_mul_49[0] = buffer_data_4[383:376] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_49[1] = buffer_data_4[391:384] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_49[2] = buffer_data_4[399:392] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_49[3] = buffer_data_4[407:400] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_49[4] = buffer_data_4[415:408] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_49[5] = buffer_data_3[383:376] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_49[6] = buffer_data_3[391:384] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_49[7] = buffer_data_3[399:392] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_49[8] = buffer_data_3[407:400] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_49[9] = buffer_data_3[415:408] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_49[10] = buffer_data_2[383:376] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_49[11] = buffer_data_2[391:384] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_49[12] = buffer_data_2[399:392] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_49[13] = buffer_data_2[407:400] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_49[14] = buffer_data_2[415:408] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_49[15] = buffer_data_1[383:376] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_49[16] = buffer_data_1[391:384] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_49[17] = buffer_data_1[399:392] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_49[18] = buffer_data_1[407:400] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_49[19] = buffer_data_1[415:408] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_49[20] = buffer_data_0[383:376] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_49[21] = buffer_data_0[391:384] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_49[22] = buffer_data_0[399:392] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_49[23] = buffer_data_0[407:400] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_49[24] = buffer_data_0[415:408] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_49 = kernel_img_mul_49[0] + kernel_img_mul_49[1] + kernel_img_mul_49[2] + 
                kernel_img_mul_49[3] + kernel_img_mul_49[4] + kernel_img_mul_49[5] + 
                kernel_img_mul_49[6] + kernel_img_mul_49[7] + kernel_img_mul_49[8] + 
                kernel_img_mul_49[9] + kernel_img_mul_49[10] + kernel_img_mul_49[11] + 
                kernel_img_mul_49[12] + kernel_img_mul_49[13] + kernel_img_mul_49[14] + 
                kernel_img_mul_49[15] + kernel_img_mul_49[16] + kernel_img_mul_49[17] + 
                kernel_img_mul_49[18] + kernel_img_mul_49[19] + kernel_img_mul_49[20] + 
                kernel_img_mul_49[21] + kernel_img_mul_49[22] + kernel_img_mul_49[23] + 
                kernel_img_mul_49[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[399:392] <= 'd0;
  else if (current_state==ST_START)
    blur_din[399:392] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[399:392] <= 'd0;
end

wire  [39:0]  kernel_img_mul_50[0:24];
assign kernel_img_mul_50[0] = buffer_data_4[391:384] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_50[1] = buffer_data_4[399:392] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_50[2] = buffer_data_4[407:400] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_50[3] = buffer_data_4[415:408] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_50[4] = buffer_data_4[423:416] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_50[5] = buffer_data_3[391:384] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_50[6] = buffer_data_3[399:392] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_50[7] = buffer_data_3[407:400] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_50[8] = buffer_data_3[415:408] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_50[9] = buffer_data_3[423:416] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_50[10] = buffer_data_2[391:384] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_50[11] = buffer_data_2[399:392] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_50[12] = buffer_data_2[407:400] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_50[13] = buffer_data_2[415:408] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_50[14] = buffer_data_2[423:416] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_50[15] = buffer_data_1[391:384] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_50[16] = buffer_data_1[399:392] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_50[17] = buffer_data_1[407:400] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_50[18] = buffer_data_1[415:408] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_50[19] = buffer_data_1[423:416] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_50[20] = buffer_data_0[391:384] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_50[21] = buffer_data_0[399:392] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_50[22] = buffer_data_0[407:400] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_50[23] = buffer_data_0[415:408] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_50[24] = buffer_data_0[423:416] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_50 = kernel_img_mul_50[0] + kernel_img_mul_50[1] + kernel_img_mul_50[2] + 
                kernel_img_mul_50[3] + kernel_img_mul_50[4] + kernel_img_mul_50[5] + 
                kernel_img_mul_50[6] + kernel_img_mul_50[7] + kernel_img_mul_50[8] + 
                kernel_img_mul_50[9] + kernel_img_mul_50[10] + kernel_img_mul_50[11] + 
                kernel_img_mul_50[12] + kernel_img_mul_50[13] + kernel_img_mul_50[14] + 
                kernel_img_mul_50[15] + kernel_img_mul_50[16] + kernel_img_mul_50[17] + 
                kernel_img_mul_50[18] + kernel_img_mul_50[19] + kernel_img_mul_50[20] + 
                kernel_img_mul_50[21] + kernel_img_mul_50[22] + kernel_img_mul_50[23] + 
                kernel_img_mul_50[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[407:400] <= 'd0;
  else if (current_state==ST_START)
    blur_din[407:400] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[407:400] <= 'd0;
end

wire  [39:0]  kernel_img_mul_51[0:24];
assign kernel_img_mul_51[0] = buffer_data_4[399:392] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_51[1] = buffer_data_4[407:400] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_51[2] = buffer_data_4[415:408] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_51[3] = buffer_data_4[423:416] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_51[4] = buffer_data_4[431:424] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_51[5] = buffer_data_3[399:392] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_51[6] = buffer_data_3[407:400] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_51[7] = buffer_data_3[415:408] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_51[8] = buffer_data_3[423:416] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_51[9] = buffer_data_3[431:424] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_51[10] = buffer_data_2[399:392] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_51[11] = buffer_data_2[407:400] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_51[12] = buffer_data_2[415:408] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_51[13] = buffer_data_2[423:416] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_51[14] = buffer_data_2[431:424] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_51[15] = buffer_data_1[399:392] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_51[16] = buffer_data_1[407:400] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_51[17] = buffer_data_1[415:408] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_51[18] = buffer_data_1[423:416] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_51[19] = buffer_data_1[431:424] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_51[20] = buffer_data_0[399:392] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_51[21] = buffer_data_0[407:400] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_51[22] = buffer_data_0[415:408] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_51[23] = buffer_data_0[423:416] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_51[24] = buffer_data_0[431:424] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_51 = kernel_img_mul_51[0] + kernel_img_mul_51[1] + kernel_img_mul_51[2] + 
                kernel_img_mul_51[3] + kernel_img_mul_51[4] + kernel_img_mul_51[5] + 
                kernel_img_mul_51[6] + kernel_img_mul_51[7] + kernel_img_mul_51[8] + 
                kernel_img_mul_51[9] + kernel_img_mul_51[10] + kernel_img_mul_51[11] + 
                kernel_img_mul_51[12] + kernel_img_mul_51[13] + kernel_img_mul_51[14] + 
                kernel_img_mul_51[15] + kernel_img_mul_51[16] + kernel_img_mul_51[17] + 
                kernel_img_mul_51[18] + kernel_img_mul_51[19] + kernel_img_mul_51[20] + 
                kernel_img_mul_51[21] + kernel_img_mul_51[22] + kernel_img_mul_51[23] + 
                kernel_img_mul_51[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[415:408] <= 'd0;
  else if (current_state==ST_START)
    blur_din[415:408] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[415:408] <= 'd0;
end

wire  [39:0]  kernel_img_mul_52[0:24];
assign kernel_img_mul_52[0] = buffer_data_4[407:400] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_52[1] = buffer_data_4[415:408] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_52[2] = buffer_data_4[423:416] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_52[3] = buffer_data_4[431:424] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_52[4] = buffer_data_4[439:432] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_52[5] = buffer_data_3[407:400] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_52[6] = buffer_data_3[415:408] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_52[7] = buffer_data_3[423:416] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_52[8] = buffer_data_3[431:424] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_52[9] = buffer_data_3[439:432] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_52[10] = buffer_data_2[407:400] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_52[11] = buffer_data_2[415:408] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_52[12] = buffer_data_2[423:416] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_52[13] = buffer_data_2[431:424] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_52[14] = buffer_data_2[439:432] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_52[15] = buffer_data_1[407:400] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_52[16] = buffer_data_1[415:408] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_52[17] = buffer_data_1[423:416] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_52[18] = buffer_data_1[431:424] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_52[19] = buffer_data_1[439:432] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_52[20] = buffer_data_0[407:400] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_52[21] = buffer_data_0[415:408] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_52[22] = buffer_data_0[423:416] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_52[23] = buffer_data_0[431:424] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_52[24] = buffer_data_0[439:432] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_52 = kernel_img_mul_52[0] + kernel_img_mul_52[1] + kernel_img_mul_52[2] + 
                kernel_img_mul_52[3] + kernel_img_mul_52[4] + kernel_img_mul_52[5] + 
                kernel_img_mul_52[6] + kernel_img_mul_52[7] + kernel_img_mul_52[8] + 
                kernel_img_mul_52[9] + kernel_img_mul_52[10] + kernel_img_mul_52[11] + 
                kernel_img_mul_52[12] + kernel_img_mul_52[13] + kernel_img_mul_52[14] + 
                kernel_img_mul_52[15] + kernel_img_mul_52[16] + kernel_img_mul_52[17] + 
                kernel_img_mul_52[18] + kernel_img_mul_52[19] + kernel_img_mul_52[20] + 
                kernel_img_mul_52[21] + kernel_img_mul_52[22] + kernel_img_mul_52[23] + 
                kernel_img_mul_52[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[423:416] <= 'd0;
  else if (current_state==ST_START)
    blur_din[423:416] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[423:416] <= 'd0;
end

wire  [39:0]  kernel_img_mul_53[0:24];
assign kernel_img_mul_53[0] = buffer_data_4[415:408] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_53[1] = buffer_data_4[423:416] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_53[2] = buffer_data_4[431:424] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_53[3] = buffer_data_4[439:432] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_53[4] = buffer_data_4[447:440] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_53[5] = buffer_data_3[415:408] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_53[6] = buffer_data_3[423:416] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_53[7] = buffer_data_3[431:424] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_53[8] = buffer_data_3[439:432] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_53[9] = buffer_data_3[447:440] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_53[10] = buffer_data_2[415:408] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_53[11] = buffer_data_2[423:416] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_53[12] = buffer_data_2[431:424] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_53[13] = buffer_data_2[439:432] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_53[14] = buffer_data_2[447:440] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_53[15] = buffer_data_1[415:408] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_53[16] = buffer_data_1[423:416] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_53[17] = buffer_data_1[431:424] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_53[18] = buffer_data_1[439:432] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_53[19] = buffer_data_1[447:440] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_53[20] = buffer_data_0[415:408] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_53[21] = buffer_data_0[423:416] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_53[22] = buffer_data_0[431:424] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_53[23] = buffer_data_0[439:432] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_53[24] = buffer_data_0[447:440] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_53 = kernel_img_mul_53[0] + kernel_img_mul_53[1] + kernel_img_mul_53[2] + 
                kernel_img_mul_53[3] + kernel_img_mul_53[4] + kernel_img_mul_53[5] + 
                kernel_img_mul_53[6] + kernel_img_mul_53[7] + kernel_img_mul_53[8] + 
                kernel_img_mul_53[9] + kernel_img_mul_53[10] + kernel_img_mul_53[11] + 
                kernel_img_mul_53[12] + kernel_img_mul_53[13] + kernel_img_mul_53[14] + 
                kernel_img_mul_53[15] + kernel_img_mul_53[16] + kernel_img_mul_53[17] + 
                kernel_img_mul_53[18] + kernel_img_mul_53[19] + kernel_img_mul_53[20] + 
                kernel_img_mul_53[21] + kernel_img_mul_53[22] + kernel_img_mul_53[23] + 
                kernel_img_mul_53[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[431:424] <= 'd0;
  else if (current_state==ST_START)
    blur_din[431:424] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[431:424] <= 'd0;
end

wire  [39:0]  kernel_img_mul_54[0:24];
assign kernel_img_mul_54[0] = buffer_data_4[423:416] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_54[1] = buffer_data_4[431:424] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_54[2] = buffer_data_4[439:432] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_54[3] = buffer_data_4[447:440] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_54[4] = buffer_data_4[455:448] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_54[5] = buffer_data_3[423:416] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_54[6] = buffer_data_3[431:424] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_54[7] = buffer_data_3[439:432] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_54[8] = buffer_data_3[447:440] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_54[9] = buffer_data_3[455:448] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_54[10] = buffer_data_2[423:416] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_54[11] = buffer_data_2[431:424] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_54[12] = buffer_data_2[439:432] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_54[13] = buffer_data_2[447:440] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_54[14] = buffer_data_2[455:448] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_54[15] = buffer_data_1[423:416] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_54[16] = buffer_data_1[431:424] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_54[17] = buffer_data_1[439:432] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_54[18] = buffer_data_1[447:440] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_54[19] = buffer_data_1[455:448] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_54[20] = buffer_data_0[423:416] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_54[21] = buffer_data_0[431:424] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_54[22] = buffer_data_0[439:432] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_54[23] = buffer_data_0[447:440] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_54[24] = buffer_data_0[455:448] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_54 = kernel_img_mul_54[0] + kernel_img_mul_54[1] + kernel_img_mul_54[2] + 
                kernel_img_mul_54[3] + kernel_img_mul_54[4] + kernel_img_mul_54[5] + 
                kernel_img_mul_54[6] + kernel_img_mul_54[7] + kernel_img_mul_54[8] + 
                kernel_img_mul_54[9] + kernel_img_mul_54[10] + kernel_img_mul_54[11] + 
                kernel_img_mul_54[12] + kernel_img_mul_54[13] + kernel_img_mul_54[14] + 
                kernel_img_mul_54[15] + kernel_img_mul_54[16] + kernel_img_mul_54[17] + 
                kernel_img_mul_54[18] + kernel_img_mul_54[19] + kernel_img_mul_54[20] + 
                kernel_img_mul_54[21] + kernel_img_mul_54[22] + kernel_img_mul_54[23] + 
                kernel_img_mul_54[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[439:432] <= 'd0;
  else if (current_state==ST_START)
    blur_din[439:432] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[439:432] <= 'd0;
end

wire  [39:0]  kernel_img_mul_55[0:24];
assign kernel_img_mul_55[0] = buffer_data_4[431:424] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_55[1] = buffer_data_4[439:432] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_55[2] = buffer_data_4[447:440] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_55[3] = buffer_data_4[455:448] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_55[4] = buffer_data_4[463:456] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_55[5] = buffer_data_3[431:424] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_55[6] = buffer_data_3[439:432] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_55[7] = buffer_data_3[447:440] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_55[8] = buffer_data_3[455:448] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_55[9] = buffer_data_3[463:456] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_55[10] = buffer_data_2[431:424] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_55[11] = buffer_data_2[439:432] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_55[12] = buffer_data_2[447:440] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_55[13] = buffer_data_2[455:448] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_55[14] = buffer_data_2[463:456] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_55[15] = buffer_data_1[431:424] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_55[16] = buffer_data_1[439:432] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_55[17] = buffer_data_1[447:440] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_55[18] = buffer_data_1[455:448] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_55[19] = buffer_data_1[463:456] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_55[20] = buffer_data_0[431:424] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_55[21] = buffer_data_0[439:432] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_55[22] = buffer_data_0[447:440] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_55[23] = buffer_data_0[455:448] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_55[24] = buffer_data_0[463:456] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_55 = kernel_img_mul_55[0] + kernel_img_mul_55[1] + kernel_img_mul_55[2] + 
                kernel_img_mul_55[3] + kernel_img_mul_55[4] + kernel_img_mul_55[5] + 
                kernel_img_mul_55[6] + kernel_img_mul_55[7] + kernel_img_mul_55[8] + 
                kernel_img_mul_55[9] + kernel_img_mul_55[10] + kernel_img_mul_55[11] + 
                kernel_img_mul_55[12] + kernel_img_mul_55[13] + kernel_img_mul_55[14] + 
                kernel_img_mul_55[15] + kernel_img_mul_55[16] + kernel_img_mul_55[17] + 
                kernel_img_mul_55[18] + kernel_img_mul_55[19] + kernel_img_mul_55[20] + 
                kernel_img_mul_55[21] + kernel_img_mul_55[22] + kernel_img_mul_55[23] + 
                kernel_img_mul_55[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[447:440] <= 'd0;
  else if (current_state==ST_START)
    blur_din[447:440] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[447:440] <= 'd0;
end

wire  [39:0]  kernel_img_mul_56[0:24];
assign kernel_img_mul_56[0] = buffer_data_4[439:432] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_56[1] = buffer_data_4[447:440] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_56[2] = buffer_data_4[455:448] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_56[3] = buffer_data_4[463:456] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_56[4] = buffer_data_4[471:464] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_56[5] = buffer_data_3[439:432] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_56[6] = buffer_data_3[447:440] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_56[7] = buffer_data_3[455:448] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_56[8] = buffer_data_3[463:456] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_56[9] = buffer_data_3[471:464] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_56[10] = buffer_data_2[439:432] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_56[11] = buffer_data_2[447:440] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_56[12] = buffer_data_2[455:448] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_56[13] = buffer_data_2[463:456] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_56[14] = buffer_data_2[471:464] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_56[15] = buffer_data_1[439:432] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_56[16] = buffer_data_1[447:440] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_56[17] = buffer_data_1[455:448] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_56[18] = buffer_data_1[463:456] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_56[19] = buffer_data_1[471:464] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_56[20] = buffer_data_0[439:432] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_56[21] = buffer_data_0[447:440] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_56[22] = buffer_data_0[455:448] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_56[23] = buffer_data_0[463:456] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_56[24] = buffer_data_0[471:464] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_56 = kernel_img_mul_56[0] + kernel_img_mul_56[1] + kernel_img_mul_56[2] + 
                kernel_img_mul_56[3] + kernel_img_mul_56[4] + kernel_img_mul_56[5] + 
                kernel_img_mul_56[6] + kernel_img_mul_56[7] + kernel_img_mul_56[8] + 
                kernel_img_mul_56[9] + kernel_img_mul_56[10] + kernel_img_mul_56[11] + 
                kernel_img_mul_56[12] + kernel_img_mul_56[13] + kernel_img_mul_56[14] + 
                kernel_img_mul_56[15] + kernel_img_mul_56[16] + kernel_img_mul_56[17] + 
                kernel_img_mul_56[18] + kernel_img_mul_56[19] + kernel_img_mul_56[20] + 
                kernel_img_mul_56[21] + kernel_img_mul_56[22] + kernel_img_mul_56[23] + 
                kernel_img_mul_56[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[455:448] <= 'd0;
  else if (current_state==ST_START)
    blur_din[455:448] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[455:448] <= 'd0;
end

wire  [39:0]  kernel_img_mul_57[0:24];
assign kernel_img_mul_57[0] = buffer_data_4[447:440] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_57[1] = buffer_data_4[455:448] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_57[2] = buffer_data_4[463:456] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_57[3] = buffer_data_4[471:464] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_57[4] = buffer_data_4[479:472] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_57[5] = buffer_data_3[447:440] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_57[6] = buffer_data_3[455:448] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_57[7] = buffer_data_3[463:456] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_57[8] = buffer_data_3[471:464] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_57[9] = buffer_data_3[479:472] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_57[10] = buffer_data_2[447:440] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_57[11] = buffer_data_2[455:448] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_57[12] = buffer_data_2[463:456] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_57[13] = buffer_data_2[471:464] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_57[14] = buffer_data_2[479:472] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_57[15] = buffer_data_1[447:440] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_57[16] = buffer_data_1[455:448] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_57[17] = buffer_data_1[463:456] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_57[18] = buffer_data_1[471:464] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_57[19] = buffer_data_1[479:472] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_57[20] = buffer_data_0[447:440] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_57[21] = buffer_data_0[455:448] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_57[22] = buffer_data_0[463:456] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_57[23] = buffer_data_0[471:464] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_57[24] = buffer_data_0[479:472] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_57 = kernel_img_mul_57[0] + kernel_img_mul_57[1] + kernel_img_mul_57[2] + 
                kernel_img_mul_57[3] + kernel_img_mul_57[4] + kernel_img_mul_57[5] + 
                kernel_img_mul_57[6] + kernel_img_mul_57[7] + kernel_img_mul_57[8] + 
                kernel_img_mul_57[9] + kernel_img_mul_57[10] + kernel_img_mul_57[11] + 
                kernel_img_mul_57[12] + kernel_img_mul_57[13] + kernel_img_mul_57[14] + 
                kernel_img_mul_57[15] + kernel_img_mul_57[16] + kernel_img_mul_57[17] + 
                kernel_img_mul_57[18] + kernel_img_mul_57[19] + kernel_img_mul_57[20] + 
                kernel_img_mul_57[21] + kernel_img_mul_57[22] + kernel_img_mul_57[23] + 
                kernel_img_mul_57[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[463:456] <= 'd0;
  else if (current_state==ST_START)
    blur_din[463:456] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[463:456] <= 'd0;
end

wire  [39:0]  kernel_img_mul_58[0:24];
assign kernel_img_mul_58[0] = buffer_data_4[455:448] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_58[1] = buffer_data_4[463:456] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_58[2] = buffer_data_4[471:464] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_58[3] = buffer_data_4[479:472] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_58[4] = buffer_data_4[487:480] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_58[5] = buffer_data_3[455:448] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_58[6] = buffer_data_3[463:456] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_58[7] = buffer_data_3[471:464] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_58[8] = buffer_data_3[479:472] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_58[9] = buffer_data_3[487:480] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_58[10] = buffer_data_2[455:448] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_58[11] = buffer_data_2[463:456] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_58[12] = buffer_data_2[471:464] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_58[13] = buffer_data_2[479:472] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_58[14] = buffer_data_2[487:480] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_58[15] = buffer_data_1[455:448] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_58[16] = buffer_data_1[463:456] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_58[17] = buffer_data_1[471:464] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_58[18] = buffer_data_1[479:472] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_58[19] = buffer_data_1[487:480] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_58[20] = buffer_data_0[455:448] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_58[21] = buffer_data_0[463:456] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_58[22] = buffer_data_0[471:464] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_58[23] = buffer_data_0[479:472] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_58[24] = buffer_data_0[487:480] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_58 = kernel_img_mul_58[0] + kernel_img_mul_58[1] + kernel_img_mul_58[2] + 
                kernel_img_mul_58[3] + kernel_img_mul_58[4] + kernel_img_mul_58[5] + 
                kernel_img_mul_58[6] + kernel_img_mul_58[7] + kernel_img_mul_58[8] + 
                kernel_img_mul_58[9] + kernel_img_mul_58[10] + kernel_img_mul_58[11] + 
                kernel_img_mul_58[12] + kernel_img_mul_58[13] + kernel_img_mul_58[14] + 
                kernel_img_mul_58[15] + kernel_img_mul_58[16] + kernel_img_mul_58[17] + 
                kernel_img_mul_58[18] + kernel_img_mul_58[19] + kernel_img_mul_58[20] + 
                kernel_img_mul_58[21] + kernel_img_mul_58[22] + kernel_img_mul_58[23] + 
                kernel_img_mul_58[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[471:464] <= 'd0;
  else if (current_state==ST_START)
    blur_din[471:464] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[471:464] <= 'd0;
end

wire  [39:0]  kernel_img_mul_59[0:24];
assign kernel_img_mul_59[0] = buffer_data_4[463:456] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_59[1] = buffer_data_4[471:464] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_59[2] = buffer_data_4[479:472] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_59[3] = buffer_data_4[487:480] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_59[4] = buffer_data_4[495:488] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_59[5] = buffer_data_3[463:456] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_59[6] = buffer_data_3[471:464] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_59[7] = buffer_data_3[479:472] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_59[8] = buffer_data_3[487:480] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_59[9] = buffer_data_3[495:488] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_59[10] = buffer_data_2[463:456] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_59[11] = buffer_data_2[471:464] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_59[12] = buffer_data_2[479:472] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_59[13] = buffer_data_2[487:480] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_59[14] = buffer_data_2[495:488] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_59[15] = buffer_data_1[463:456] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_59[16] = buffer_data_1[471:464] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_59[17] = buffer_data_1[479:472] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_59[18] = buffer_data_1[487:480] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_59[19] = buffer_data_1[495:488] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_59[20] = buffer_data_0[463:456] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_59[21] = buffer_data_0[471:464] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_59[22] = buffer_data_0[479:472] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_59[23] = buffer_data_0[487:480] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_59[24] = buffer_data_0[495:488] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_59 = kernel_img_mul_59[0] + kernel_img_mul_59[1] + kernel_img_mul_59[2] + 
                kernel_img_mul_59[3] + kernel_img_mul_59[4] + kernel_img_mul_59[5] + 
                kernel_img_mul_59[6] + kernel_img_mul_59[7] + kernel_img_mul_59[8] + 
                kernel_img_mul_59[9] + kernel_img_mul_59[10] + kernel_img_mul_59[11] + 
                kernel_img_mul_59[12] + kernel_img_mul_59[13] + kernel_img_mul_59[14] + 
                kernel_img_mul_59[15] + kernel_img_mul_59[16] + kernel_img_mul_59[17] + 
                kernel_img_mul_59[18] + kernel_img_mul_59[19] + kernel_img_mul_59[20] + 
                kernel_img_mul_59[21] + kernel_img_mul_59[22] + kernel_img_mul_59[23] + 
                kernel_img_mul_59[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[479:472] <= 'd0;
  else if (current_state==ST_START)
    blur_din[479:472] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[479:472] <= 'd0;
end

wire  [39:0]  kernel_img_mul_60[0:24];
assign kernel_img_mul_60[0] = buffer_data_4[471:464] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_60[1] = buffer_data_4[479:472] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_60[2] = buffer_data_4[487:480] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_60[3] = buffer_data_4[495:488] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_60[4] = buffer_data_4[503:496] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_60[5] = buffer_data_3[471:464] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_60[6] = buffer_data_3[479:472] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_60[7] = buffer_data_3[487:480] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_60[8] = buffer_data_3[495:488] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_60[9] = buffer_data_3[503:496] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_60[10] = buffer_data_2[471:464] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_60[11] = buffer_data_2[479:472] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_60[12] = buffer_data_2[487:480] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_60[13] = buffer_data_2[495:488] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_60[14] = buffer_data_2[503:496] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_60[15] = buffer_data_1[471:464] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_60[16] = buffer_data_1[479:472] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_60[17] = buffer_data_1[487:480] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_60[18] = buffer_data_1[495:488] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_60[19] = buffer_data_1[503:496] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_60[20] = buffer_data_0[471:464] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_60[21] = buffer_data_0[479:472] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_60[22] = buffer_data_0[487:480] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_60[23] = buffer_data_0[495:488] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_60[24] = buffer_data_0[503:496] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_60 = kernel_img_mul_60[0] + kernel_img_mul_60[1] + kernel_img_mul_60[2] + 
                kernel_img_mul_60[3] + kernel_img_mul_60[4] + kernel_img_mul_60[5] + 
                kernel_img_mul_60[6] + kernel_img_mul_60[7] + kernel_img_mul_60[8] + 
                kernel_img_mul_60[9] + kernel_img_mul_60[10] + kernel_img_mul_60[11] + 
                kernel_img_mul_60[12] + kernel_img_mul_60[13] + kernel_img_mul_60[14] + 
                kernel_img_mul_60[15] + kernel_img_mul_60[16] + kernel_img_mul_60[17] + 
                kernel_img_mul_60[18] + kernel_img_mul_60[19] + kernel_img_mul_60[20] + 
                kernel_img_mul_60[21] + kernel_img_mul_60[22] + kernel_img_mul_60[23] + 
                kernel_img_mul_60[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[487:480] <= 'd0;
  else if (current_state==ST_START)
    blur_din[487:480] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[487:480] <= 'd0;
end

wire  [39:0]  kernel_img_mul_61[0:24];
assign kernel_img_mul_61[0] = buffer_data_4[479:472] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_61[1] = buffer_data_4[487:480] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_61[2] = buffer_data_4[495:488] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_61[3] = buffer_data_4[503:496] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_61[4] = buffer_data_4[511:504] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_61[5] = buffer_data_3[479:472] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_61[6] = buffer_data_3[487:480] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_61[7] = buffer_data_3[495:488] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_61[8] = buffer_data_3[503:496] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_61[9] = buffer_data_3[511:504] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_61[10] = buffer_data_2[479:472] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_61[11] = buffer_data_2[487:480] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_61[12] = buffer_data_2[495:488] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_61[13] = buffer_data_2[503:496] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_61[14] = buffer_data_2[511:504] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_61[15] = buffer_data_1[479:472] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_61[16] = buffer_data_1[487:480] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_61[17] = buffer_data_1[495:488] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_61[18] = buffer_data_1[503:496] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_61[19] = buffer_data_1[511:504] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_61[20] = buffer_data_0[479:472] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_61[21] = buffer_data_0[487:480] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_61[22] = buffer_data_0[495:488] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_61[23] = buffer_data_0[503:496] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_61[24] = buffer_data_0[511:504] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_61 = kernel_img_mul_61[0] + kernel_img_mul_61[1] + kernel_img_mul_61[2] + 
                kernel_img_mul_61[3] + kernel_img_mul_61[4] + kernel_img_mul_61[5] + 
                kernel_img_mul_61[6] + kernel_img_mul_61[7] + kernel_img_mul_61[8] + 
                kernel_img_mul_61[9] + kernel_img_mul_61[10] + kernel_img_mul_61[11] + 
                kernel_img_mul_61[12] + kernel_img_mul_61[13] + kernel_img_mul_61[14] + 
                kernel_img_mul_61[15] + kernel_img_mul_61[16] + kernel_img_mul_61[17] + 
                kernel_img_mul_61[18] + kernel_img_mul_61[19] + kernel_img_mul_61[20] + 
                kernel_img_mul_61[21] + kernel_img_mul_61[22] + kernel_img_mul_61[23] + 
                kernel_img_mul_61[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[495:488] <= 'd0;
  else if (current_state==ST_START)
    blur_din[495:488] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[495:488] <= 'd0;
end

wire  [39:0]  kernel_img_mul_62[0:24];
assign kernel_img_mul_62[0] = buffer_data_4[487:480] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_62[1] = buffer_data_4[495:488] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_62[2] = buffer_data_4[503:496] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_62[3] = buffer_data_4[511:504] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_62[4] = buffer_data_4[519:512] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_62[5] = buffer_data_3[487:480] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_62[6] = buffer_data_3[495:488] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_62[7] = buffer_data_3[503:496] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_62[8] = buffer_data_3[511:504] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_62[9] = buffer_data_3[519:512] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_62[10] = buffer_data_2[487:480] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_62[11] = buffer_data_2[495:488] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_62[12] = buffer_data_2[503:496] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_62[13] = buffer_data_2[511:504] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_62[14] = buffer_data_2[519:512] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_62[15] = buffer_data_1[487:480] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_62[16] = buffer_data_1[495:488] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_62[17] = buffer_data_1[503:496] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_62[18] = buffer_data_1[511:504] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_62[19] = buffer_data_1[519:512] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_62[20] = buffer_data_0[487:480] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_62[21] = buffer_data_0[495:488] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_62[22] = buffer_data_0[503:496] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_62[23] = buffer_data_0[511:504] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_62[24] = buffer_data_0[519:512] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_62 = kernel_img_mul_62[0] + kernel_img_mul_62[1] + kernel_img_mul_62[2] + 
                kernel_img_mul_62[3] + kernel_img_mul_62[4] + kernel_img_mul_62[5] + 
                kernel_img_mul_62[6] + kernel_img_mul_62[7] + kernel_img_mul_62[8] + 
                kernel_img_mul_62[9] + kernel_img_mul_62[10] + kernel_img_mul_62[11] + 
                kernel_img_mul_62[12] + kernel_img_mul_62[13] + kernel_img_mul_62[14] + 
                kernel_img_mul_62[15] + kernel_img_mul_62[16] + kernel_img_mul_62[17] + 
                kernel_img_mul_62[18] + kernel_img_mul_62[19] + kernel_img_mul_62[20] + 
                kernel_img_mul_62[21] + kernel_img_mul_62[22] + kernel_img_mul_62[23] + 
                kernel_img_mul_62[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[503:496] <= 'd0;
  else if (current_state==ST_START)
    blur_din[503:496] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[503:496] <= 'd0;
end

wire  [39:0]  kernel_img_mul_63[0:24];
assign kernel_img_mul_63[0] = buffer_data_4[495:488] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_63[1] = buffer_data_4[503:496] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_63[2] = buffer_data_4[511:504] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_63[3] = buffer_data_4[519:512] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_63[4] = buffer_data_4[527:520] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_63[5] = buffer_data_3[495:488] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_63[6] = buffer_data_3[503:496] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_63[7] = buffer_data_3[511:504] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_63[8] = buffer_data_3[519:512] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_63[9] = buffer_data_3[527:520] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_63[10] = buffer_data_2[495:488] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_63[11] = buffer_data_2[503:496] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_63[12] = buffer_data_2[511:504] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_63[13] = buffer_data_2[519:512] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_63[14] = buffer_data_2[527:520] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_63[15] = buffer_data_1[495:488] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_63[16] = buffer_data_1[503:496] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_63[17] = buffer_data_1[511:504] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_63[18] = buffer_data_1[519:512] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_63[19] = buffer_data_1[527:520] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_63[20] = buffer_data_0[495:488] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_63[21] = buffer_data_0[503:496] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_63[22] = buffer_data_0[511:504] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_63[23] = buffer_data_0[519:512] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_63[24] = buffer_data_0[527:520] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_63 = kernel_img_mul_63[0] + kernel_img_mul_63[1] + kernel_img_mul_63[2] + 
                kernel_img_mul_63[3] + kernel_img_mul_63[4] + kernel_img_mul_63[5] + 
                kernel_img_mul_63[6] + kernel_img_mul_63[7] + kernel_img_mul_63[8] + 
                kernel_img_mul_63[9] + kernel_img_mul_63[10] + kernel_img_mul_63[11] + 
                kernel_img_mul_63[12] + kernel_img_mul_63[13] + kernel_img_mul_63[14] + 
                kernel_img_mul_63[15] + kernel_img_mul_63[16] + kernel_img_mul_63[17] + 
                kernel_img_mul_63[18] + kernel_img_mul_63[19] + kernel_img_mul_63[20] + 
                kernel_img_mul_63[21] + kernel_img_mul_63[22] + kernel_img_mul_63[23] + 
                kernel_img_mul_63[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[511:504] <= 'd0;
  else if (current_state==ST_START)
    blur_din[511:504] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[511:504] <= 'd0;
end

wire  [39:0]  kernel_img_mul_64[0:24];
assign kernel_img_mul_64[0] = buffer_data_4[503:496] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_64[1] = buffer_data_4[511:504] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_64[2] = buffer_data_4[519:512] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_64[3] = buffer_data_4[527:520] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_64[4] = buffer_data_4[535:528] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_64[5] = buffer_data_3[503:496] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_64[6] = buffer_data_3[511:504] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_64[7] = buffer_data_3[519:512] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_64[8] = buffer_data_3[527:520] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_64[9] = buffer_data_3[535:528] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_64[10] = buffer_data_2[503:496] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_64[11] = buffer_data_2[511:504] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_64[12] = buffer_data_2[519:512] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_64[13] = buffer_data_2[527:520] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_64[14] = buffer_data_2[535:528] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_64[15] = buffer_data_1[503:496] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_64[16] = buffer_data_1[511:504] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_64[17] = buffer_data_1[519:512] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_64[18] = buffer_data_1[527:520] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_64[19] = buffer_data_1[535:528] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_64[20] = buffer_data_0[503:496] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_64[21] = buffer_data_0[511:504] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_64[22] = buffer_data_0[519:512] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_64[23] = buffer_data_0[527:520] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_64[24] = buffer_data_0[535:528] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_64 = kernel_img_mul_64[0] + kernel_img_mul_64[1] + kernel_img_mul_64[2] + 
                kernel_img_mul_64[3] + kernel_img_mul_64[4] + kernel_img_mul_64[5] + 
                kernel_img_mul_64[6] + kernel_img_mul_64[7] + kernel_img_mul_64[8] + 
                kernel_img_mul_64[9] + kernel_img_mul_64[10] + kernel_img_mul_64[11] + 
                kernel_img_mul_64[12] + kernel_img_mul_64[13] + kernel_img_mul_64[14] + 
                kernel_img_mul_64[15] + kernel_img_mul_64[16] + kernel_img_mul_64[17] + 
                kernel_img_mul_64[18] + kernel_img_mul_64[19] + kernel_img_mul_64[20] + 
                kernel_img_mul_64[21] + kernel_img_mul_64[22] + kernel_img_mul_64[23] + 
                kernel_img_mul_64[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[519:512] <= 'd0;
  else if (current_state==ST_START)
    blur_din[519:512] <= kernel_img_sum_64[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[519:512] <= 'd0;
end

wire  [39:0]  kernel_img_mul_65[0:24];
assign kernel_img_mul_65[0] = buffer_data_4[511:504] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_65[1] = buffer_data_4[519:512] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_65[2] = buffer_data_4[527:520] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_65[3] = buffer_data_4[535:528] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_65[4] = buffer_data_4[543:536] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_65[5] = buffer_data_3[511:504] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_65[6] = buffer_data_3[519:512] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_65[7] = buffer_data_3[527:520] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_65[8] = buffer_data_3[535:528] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_65[9] = buffer_data_3[543:536] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_65[10] = buffer_data_2[511:504] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_65[11] = buffer_data_2[519:512] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_65[12] = buffer_data_2[527:520] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_65[13] = buffer_data_2[535:528] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_65[14] = buffer_data_2[543:536] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_65[15] = buffer_data_1[511:504] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_65[16] = buffer_data_1[519:512] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_65[17] = buffer_data_1[527:520] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_65[18] = buffer_data_1[535:528] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_65[19] = buffer_data_1[543:536] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_65[20] = buffer_data_0[511:504] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_65[21] = buffer_data_0[519:512] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_65[22] = buffer_data_0[527:520] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_65[23] = buffer_data_0[535:528] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_65[24] = buffer_data_0[543:536] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_65 = kernel_img_mul_65[0] + kernel_img_mul_65[1] + kernel_img_mul_65[2] + 
                kernel_img_mul_65[3] + kernel_img_mul_65[4] + kernel_img_mul_65[5] + 
                kernel_img_mul_65[6] + kernel_img_mul_65[7] + kernel_img_mul_65[8] + 
                kernel_img_mul_65[9] + kernel_img_mul_65[10] + kernel_img_mul_65[11] + 
                kernel_img_mul_65[12] + kernel_img_mul_65[13] + kernel_img_mul_65[14] + 
                kernel_img_mul_65[15] + kernel_img_mul_65[16] + kernel_img_mul_65[17] + 
                kernel_img_mul_65[18] + kernel_img_mul_65[19] + kernel_img_mul_65[20] + 
                kernel_img_mul_65[21] + kernel_img_mul_65[22] + kernel_img_mul_65[23] + 
                kernel_img_mul_65[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[527:520] <= 'd0;
  else if (current_state==ST_START)
    blur_din[527:520] <= kernel_img_sum_65[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[527:520] <= 'd0;
end

wire  [39:0]  kernel_img_mul_66[0:24];
assign kernel_img_mul_66[0] = buffer_data_4[519:512] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_66[1] = buffer_data_4[527:520] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_66[2] = buffer_data_4[535:528] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_66[3] = buffer_data_4[543:536] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_66[4] = buffer_data_4[551:544] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_66[5] = buffer_data_3[519:512] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_66[6] = buffer_data_3[527:520] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_66[7] = buffer_data_3[535:528] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_66[8] = buffer_data_3[543:536] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_66[9] = buffer_data_3[551:544] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_66[10] = buffer_data_2[519:512] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_66[11] = buffer_data_2[527:520] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_66[12] = buffer_data_2[535:528] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_66[13] = buffer_data_2[543:536] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_66[14] = buffer_data_2[551:544] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_66[15] = buffer_data_1[519:512] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_66[16] = buffer_data_1[527:520] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_66[17] = buffer_data_1[535:528] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_66[18] = buffer_data_1[543:536] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_66[19] = buffer_data_1[551:544] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_66[20] = buffer_data_0[519:512] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_66[21] = buffer_data_0[527:520] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_66[22] = buffer_data_0[535:528] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_66[23] = buffer_data_0[543:536] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_66[24] = buffer_data_0[551:544] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_66 = kernel_img_mul_66[0] + kernel_img_mul_66[1] + kernel_img_mul_66[2] + 
                kernel_img_mul_66[3] + kernel_img_mul_66[4] + kernel_img_mul_66[5] + 
                kernel_img_mul_66[6] + kernel_img_mul_66[7] + kernel_img_mul_66[8] + 
                kernel_img_mul_66[9] + kernel_img_mul_66[10] + kernel_img_mul_66[11] + 
                kernel_img_mul_66[12] + kernel_img_mul_66[13] + kernel_img_mul_66[14] + 
                kernel_img_mul_66[15] + kernel_img_mul_66[16] + kernel_img_mul_66[17] + 
                kernel_img_mul_66[18] + kernel_img_mul_66[19] + kernel_img_mul_66[20] + 
                kernel_img_mul_66[21] + kernel_img_mul_66[22] + kernel_img_mul_66[23] + 
                kernel_img_mul_66[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[535:528] <= 'd0;
  else if (current_state==ST_START)
    blur_din[535:528] <= kernel_img_sum_66[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[535:528] <= 'd0;
end

wire  [39:0]  kernel_img_mul_67[0:24];
assign kernel_img_mul_67[0] = buffer_data_4[527:520] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_67[1] = buffer_data_4[535:528] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_67[2] = buffer_data_4[543:536] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_67[3] = buffer_data_4[551:544] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_67[4] = buffer_data_4[559:552] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_67[5] = buffer_data_3[527:520] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_67[6] = buffer_data_3[535:528] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_67[7] = buffer_data_3[543:536] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_67[8] = buffer_data_3[551:544] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_67[9] = buffer_data_3[559:552] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_67[10] = buffer_data_2[527:520] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_67[11] = buffer_data_2[535:528] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_67[12] = buffer_data_2[543:536] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_67[13] = buffer_data_2[551:544] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_67[14] = buffer_data_2[559:552] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_67[15] = buffer_data_1[527:520] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_67[16] = buffer_data_1[535:528] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_67[17] = buffer_data_1[543:536] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_67[18] = buffer_data_1[551:544] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_67[19] = buffer_data_1[559:552] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_67[20] = buffer_data_0[527:520] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_67[21] = buffer_data_0[535:528] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_67[22] = buffer_data_0[543:536] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_67[23] = buffer_data_0[551:544] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_67[24] = buffer_data_0[559:552] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_67 = kernel_img_mul_67[0] + kernel_img_mul_67[1] + kernel_img_mul_67[2] + 
                kernel_img_mul_67[3] + kernel_img_mul_67[4] + kernel_img_mul_67[5] + 
                kernel_img_mul_67[6] + kernel_img_mul_67[7] + kernel_img_mul_67[8] + 
                kernel_img_mul_67[9] + kernel_img_mul_67[10] + kernel_img_mul_67[11] + 
                kernel_img_mul_67[12] + kernel_img_mul_67[13] + kernel_img_mul_67[14] + 
                kernel_img_mul_67[15] + kernel_img_mul_67[16] + kernel_img_mul_67[17] + 
                kernel_img_mul_67[18] + kernel_img_mul_67[19] + kernel_img_mul_67[20] + 
                kernel_img_mul_67[21] + kernel_img_mul_67[22] + kernel_img_mul_67[23] + 
                kernel_img_mul_67[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[543:536] <= 'd0;
  else if (current_state==ST_START)
    blur_din[543:536] <= kernel_img_sum_67[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[543:536] <= 'd0;
end

wire  [39:0]  kernel_img_mul_68[0:24];
assign kernel_img_mul_68[0] = buffer_data_4[535:528] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_68[1] = buffer_data_4[543:536] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_68[2] = buffer_data_4[551:544] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_68[3] = buffer_data_4[559:552] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_68[4] = buffer_data_4[567:560] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_68[5] = buffer_data_3[535:528] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_68[6] = buffer_data_3[543:536] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_68[7] = buffer_data_3[551:544] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_68[8] = buffer_data_3[559:552] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_68[9] = buffer_data_3[567:560] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_68[10] = buffer_data_2[535:528] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_68[11] = buffer_data_2[543:536] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_68[12] = buffer_data_2[551:544] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_68[13] = buffer_data_2[559:552] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_68[14] = buffer_data_2[567:560] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_68[15] = buffer_data_1[535:528] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_68[16] = buffer_data_1[543:536] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_68[17] = buffer_data_1[551:544] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_68[18] = buffer_data_1[559:552] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_68[19] = buffer_data_1[567:560] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_68[20] = buffer_data_0[535:528] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_68[21] = buffer_data_0[543:536] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_68[22] = buffer_data_0[551:544] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_68[23] = buffer_data_0[559:552] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_68[24] = buffer_data_0[567:560] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_68 = kernel_img_mul_68[0] + kernel_img_mul_68[1] + kernel_img_mul_68[2] + 
                kernel_img_mul_68[3] + kernel_img_mul_68[4] + kernel_img_mul_68[5] + 
                kernel_img_mul_68[6] + kernel_img_mul_68[7] + kernel_img_mul_68[8] + 
                kernel_img_mul_68[9] + kernel_img_mul_68[10] + kernel_img_mul_68[11] + 
                kernel_img_mul_68[12] + kernel_img_mul_68[13] + kernel_img_mul_68[14] + 
                kernel_img_mul_68[15] + kernel_img_mul_68[16] + kernel_img_mul_68[17] + 
                kernel_img_mul_68[18] + kernel_img_mul_68[19] + kernel_img_mul_68[20] + 
                kernel_img_mul_68[21] + kernel_img_mul_68[22] + kernel_img_mul_68[23] + 
                kernel_img_mul_68[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[551:544] <= 'd0;
  else if (current_state==ST_START)
    blur_din[551:544] <= kernel_img_sum_68[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[551:544] <= 'd0;
end

wire  [39:0]  kernel_img_mul_69[0:24];
assign kernel_img_mul_69[0] = buffer_data_4[543:536] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_69[1] = buffer_data_4[551:544] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_69[2] = buffer_data_4[559:552] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_69[3] = buffer_data_4[567:560] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_69[4] = buffer_data_4[575:568] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_69[5] = buffer_data_3[543:536] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_69[6] = buffer_data_3[551:544] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_69[7] = buffer_data_3[559:552] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_69[8] = buffer_data_3[567:560] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_69[9] = buffer_data_3[575:568] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_69[10] = buffer_data_2[543:536] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_69[11] = buffer_data_2[551:544] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_69[12] = buffer_data_2[559:552] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_69[13] = buffer_data_2[567:560] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_69[14] = buffer_data_2[575:568] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_69[15] = buffer_data_1[543:536] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_69[16] = buffer_data_1[551:544] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_69[17] = buffer_data_1[559:552] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_69[18] = buffer_data_1[567:560] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_69[19] = buffer_data_1[575:568] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_69[20] = buffer_data_0[543:536] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_69[21] = buffer_data_0[551:544] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_69[22] = buffer_data_0[559:552] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_69[23] = buffer_data_0[567:560] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_69[24] = buffer_data_0[575:568] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_69 = kernel_img_mul_69[0] + kernel_img_mul_69[1] + kernel_img_mul_69[2] + 
                kernel_img_mul_69[3] + kernel_img_mul_69[4] + kernel_img_mul_69[5] + 
                kernel_img_mul_69[6] + kernel_img_mul_69[7] + kernel_img_mul_69[8] + 
                kernel_img_mul_69[9] + kernel_img_mul_69[10] + kernel_img_mul_69[11] + 
                kernel_img_mul_69[12] + kernel_img_mul_69[13] + kernel_img_mul_69[14] + 
                kernel_img_mul_69[15] + kernel_img_mul_69[16] + kernel_img_mul_69[17] + 
                kernel_img_mul_69[18] + kernel_img_mul_69[19] + kernel_img_mul_69[20] + 
                kernel_img_mul_69[21] + kernel_img_mul_69[22] + kernel_img_mul_69[23] + 
                kernel_img_mul_69[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[559:552] <= 'd0;
  else if (current_state==ST_START)
    blur_din[559:552] <= kernel_img_sum_69[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[559:552] <= 'd0;
end

wire  [39:0]  kernel_img_mul_70[0:24];
assign kernel_img_mul_70[0] = buffer_data_4[551:544] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_70[1] = buffer_data_4[559:552] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_70[2] = buffer_data_4[567:560] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_70[3] = buffer_data_4[575:568] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_70[4] = buffer_data_4[583:576] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_70[5] = buffer_data_3[551:544] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_70[6] = buffer_data_3[559:552] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_70[7] = buffer_data_3[567:560] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_70[8] = buffer_data_3[575:568] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_70[9] = buffer_data_3[583:576] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_70[10] = buffer_data_2[551:544] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_70[11] = buffer_data_2[559:552] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_70[12] = buffer_data_2[567:560] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_70[13] = buffer_data_2[575:568] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_70[14] = buffer_data_2[583:576] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_70[15] = buffer_data_1[551:544] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_70[16] = buffer_data_1[559:552] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_70[17] = buffer_data_1[567:560] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_70[18] = buffer_data_1[575:568] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_70[19] = buffer_data_1[583:576] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_70[20] = buffer_data_0[551:544] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_70[21] = buffer_data_0[559:552] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_70[22] = buffer_data_0[567:560] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_70[23] = buffer_data_0[575:568] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_70[24] = buffer_data_0[583:576] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_70 = kernel_img_mul_70[0] + kernel_img_mul_70[1] + kernel_img_mul_70[2] + 
                kernel_img_mul_70[3] + kernel_img_mul_70[4] + kernel_img_mul_70[5] + 
                kernel_img_mul_70[6] + kernel_img_mul_70[7] + kernel_img_mul_70[8] + 
                kernel_img_mul_70[9] + kernel_img_mul_70[10] + kernel_img_mul_70[11] + 
                kernel_img_mul_70[12] + kernel_img_mul_70[13] + kernel_img_mul_70[14] + 
                kernel_img_mul_70[15] + kernel_img_mul_70[16] + kernel_img_mul_70[17] + 
                kernel_img_mul_70[18] + kernel_img_mul_70[19] + kernel_img_mul_70[20] + 
                kernel_img_mul_70[21] + kernel_img_mul_70[22] + kernel_img_mul_70[23] + 
                kernel_img_mul_70[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[567:560] <= 'd0;
  else if (current_state==ST_START)
    blur_din[567:560] <= kernel_img_sum_70[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[567:560] <= 'd0;
end

wire  [39:0]  kernel_img_mul_71[0:24];
assign kernel_img_mul_71[0] = buffer_data_4[559:552] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_71[1] = buffer_data_4[567:560] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_71[2] = buffer_data_4[575:568] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_71[3] = buffer_data_4[583:576] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_71[4] = buffer_data_4[591:584] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_71[5] = buffer_data_3[559:552] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_71[6] = buffer_data_3[567:560] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_71[7] = buffer_data_3[575:568] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_71[8] = buffer_data_3[583:576] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_71[9] = buffer_data_3[591:584] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_71[10] = buffer_data_2[559:552] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_71[11] = buffer_data_2[567:560] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_71[12] = buffer_data_2[575:568] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_71[13] = buffer_data_2[583:576] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_71[14] = buffer_data_2[591:584] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_71[15] = buffer_data_1[559:552] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_71[16] = buffer_data_1[567:560] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_71[17] = buffer_data_1[575:568] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_71[18] = buffer_data_1[583:576] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_71[19] = buffer_data_1[591:584] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_71[20] = buffer_data_0[559:552] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_71[21] = buffer_data_0[567:560] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_71[22] = buffer_data_0[575:568] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_71[23] = buffer_data_0[583:576] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_71[24] = buffer_data_0[591:584] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_71 = kernel_img_mul_71[0] + kernel_img_mul_71[1] + kernel_img_mul_71[2] + 
                kernel_img_mul_71[3] + kernel_img_mul_71[4] + kernel_img_mul_71[5] + 
                kernel_img_mul_71[6] + kernel_img_mul_71[7] + kernel_img_mul_71[8] + 
                kernel_img_mul_71[9] + kernel_img_mul_71[10] + kernel_img_mul_71[11] + 
                kernel_img_mul_71[12] + kernel_img_mul_71[13] + kernel_img_mul_71[14] + 
                kernel_img_mul_71[15] + kernel_img_mul_71[16] + kernel_img_mul_71[17] + 
                kernel_img_mul_71[18] + kernel_img_mul_71[19] + kernel_img_mul_71[20] + 
                kernel_img_mul_71[21] + kernel_img_mul_71[22] + kernel_img_mul_71[23] + 
                kernel_img_mul_71[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[575:568] <= 'd0;
  else if (current_state==ST_START)
    blur_din[575:568] <= kernel_img_sum_71[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[575:568] <= 'd0;
end

wire  [39:0]  kernel_img_mul_72[0:24];
assign kernel_img_mul_72[0] = buffer_data_4[567:560] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_72[1] = buffer_data_4[575:568] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_72[2] = buffer_data_4[583:576] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_72[3] = buffer_data_4[591:584] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_72[4] = buffer_data_4[599:592] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_72[5] = buffer_data_3[567:560] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_72[6] = buffer_data_3[575:568] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_72[7] = buffer_data_3[583:576] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_72[8] = buffer_data_3[591:584] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_72[9] = buffer_data_3[599:592] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_72[10] = buffer_data_2[567:560] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_72[11] = buffer_data_2[575:568] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_72[12] = buffer_data_2[583:576] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_72[13] = buffer_data_2[591:584] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_72[14] = buffer_data_2[599:592] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_72[15] = buffer_data_1[567:560] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_72[16] = buffer_data_1[575:568] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_72[17] = buffer_data_1[583:576] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_72[18] = buffer_data_1[591:584] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_72[19] = buffer_data_1[599:592] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_72[20] = buffer_data_0[567:560] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_72[21] = buffer_data_0[575:568] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_72[22] = buffer_data_0[583:576] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_72[23] = buffer_data_0[591:584] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_72[24] = buffer_data_0[599:592] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_72 = kernel_img_mul_72[0] + kernel_img_mul_72[1] + kernel_img_mul_72[2] + 
                kernel_img_mul_72[3] + kernel_img_mul_72[4] + kernel_img_mul_72[5] + 
                kernel_img_mul_72[6] + kernel_img_mul_72[7] + kernel_img_mul_72[8] + 
                kernel_img_mul_72[9] + kernel_img_mul_72[10] + kernel_img_mul_72[11] + 
                kernel_img_mul_72[12] + kernel_img_mul_72[13] + kernel_img_mul_72[14] + 
                kernel_img_mul_72[15] + kernel_img_mul_72[16] + kernel_img_mul_72[17] + 
                kernel_img_mul_72[18] + kernel_img_mul_72[19] + kernel_img_mul_72[20] + 
                kernel_img_mul_72[21] + kernel_img_mul_72[22] + kernel_img_mul_72[23] + 
                kernel_img_mul_72[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[583:576] <= 'd0;
  else if (current_state==ST_START)
    blur_din[583:576] <= kernel_img_sum_72[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[583:576] <= 'd0;
end

wire  [39:0]  kernel_img_mul_73[0:24];
assign kernel_img_mul_73[0] = buffer_data_4[575:568] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_73[1] = buffer_data_4[583:576] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_73[2] = buffer_data_4[591:584] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_73[3] = buffer_data_4[599:592] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_73[4] = buffer_data_4[607:600] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_73[5] = buffer_data_3[575:568] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_73[6] = buffer_data_3[583:576] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_73[7] = buffer_data_3[591:584] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_73[8] = buffer_data_3[599:592] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_73[9] = buffer_data_3[607:600] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_73[10] = buffer_data_2[575:568] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_73[11] = buffer_data_2[583:576] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_73[12] = buffer_data_2[591:584] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_73[13] = buffer_data_2[599:592] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_73[14] = buffer_data_2[607:600] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_73[15] = buffer_data_1[575:568] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_73[16] = buffer_data_1[583:576] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_73[17] = buffer_data_1[591:584] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_73[18] = buffer_data_1[599:592] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_73[19] = buffer_data_1[607:600] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_73[20] = buffer_data_0[575:568] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_73[21] = buffer_data_0[583:576] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_73[22] = buffer_data_0[591:584] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_73[23] = buffer_data_0[599:592] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_73[24] = buffer_data_0[607:600] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_73 = kernel_img_mul_73[0] + kernel_img_mul_73[1] + kernel_img_mul_73[2] + 
                kernel_img_mul_73[3] + kernel_img_mul_73[4] + kernel_img_mul_73[5] + 
                kernel_img_mul_73[6] + kernel_img_mul_73[7] + kernel_img_mul_73[8] + 
                kernel_img_mul_73[9] + kernel_img_mul_73[10] + kernel_img_mul_73[11] + 
                kernel_img_mul_73[12] + kernel_img_mul_73[13] + kernel_img_mul_73[14] + 
                kernel_img_mul_73[15] + kernel_img_mul_73[16] + kernel_img_mul_73[17] + 
                kernel_img_mul_73[18] + kernel_img_mul_73[19] + kernel_img_mul_73[20] + 
                kernel_img_mul_73[21] + kernel_img_mul_73[22] + kernel_img_mul_73[23] + 
                kernel_img_mul_73[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[591:584] <= 'd0;
  else if (current_state==ST_START)
    blur_din[591:584] <= kernel_img_sum_73[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[591:584] <= 'd0;
end

wire  [39:0]  kernel_img_mul_74[0:24];
assign kernel_img_mul_74[0] = buffer_data_4[583:576] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_74[1] = buffer_data_4[591:584] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_74[2] = buffer_data_4[599:592] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_74[3] = buffer_data_4[607:600] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_74[4] = buffer_data_4[615:608] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_74[5] = buffer_data_3[583:576] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_74[6] = buffer_data_3[591:584] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_74[7] = buffer_data_3[599:592] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_74[8] = buffer_data_3[607:600] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_74[9] = buffer_data_3[615:608] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_74[10] = buffer_data_2[583:576] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_74[11] = buffer_data_2[591:584] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_74[12] = buffer_data_2[599:592] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_74[13] = buffer_data_2[607:600] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_74[14] = buffer_data_2[615:608] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_74[15] = buffer_data_1[583:576] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_74[16] = buffer_data_1[591:584] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_74[17] = buffer_data_1[599:592] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_74[18] = buffer_data_1[607:600] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_74[19] = buffer_data_1[615:608] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_74[20] = buffer_data_0[583:576] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_74[21] = buffer_data_0[591:584] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_74[22] = buffer_data_0[599:592] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_74[23] = buffer_data_0[607:600] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_74[24] = buffer_data_0[615:608] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_74 = kernel_img_mul_74[0] + kernel_img_mul_74[1] + kernel_img_mul_74[2] + 
                kernel_img_mul_74[3] + kernel_img_mul_74[4] + kernel_img_mul_74[5] + 
                kernel_img_mul_74[6] + kernel_img_mul_74[7] + kernel_img_mul_74[8] + 
                kernel_img_mul_74[9] + kernel_img_mul_74[10] + kernel_img_mul_74[11] + 
                kernel_img_mul_74[12] + kernel_img_mul_74[13] + kernel_img_mul_74[14] + 
                kernel_img_mul_74[15] + kernel_img_mul_74[16] + kernel_img_mul_74[17] + 
                kernel_img_mul_74[18] + kernel_img_mul_74[19] + kernel_img_mul_74[20] + 
                kernel_img_mul_74[21] + kernel_img_mul_74[22] + kernel_img_mul_74[23] + 
                kernel_img_mul_74[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[599:592] <= 'd0;
  else if (current_state==ST_START)
    blur_din[599:592] <= kernel_img_sum_74[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[599:592] <= 'd0;
end

wire  [39:0]  kernel_img_mul_75[0:24];
assign kernel_img_mul_75[0] = buffer_data_4[591:584] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_75[1] = buffer_data_4[599:592] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_75[2] = buffer_data_4[607:600] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_75[3] = buffer_data_4[615:608] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_75[4] = buffer_data_4[623:616] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_75[5] = buffer_data_3[591:584] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_75[6] = buffer_data_3[599:592] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_75[7] = buffer_data_3[607:600] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_75[8] = buffer_data_3[615:608] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_75[9] = buffer_data_3[623:616] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_75[10] = buffer_data_2[591:584] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_75[11] = buffer_data_2[599:592] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_75[12] = buffer_data_2[607:600] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_75[13] = buffer_data_2[615:608] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_75[14] = buffer_data_2[623:616] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_75[15] = buffer_data_1[591:584] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_75[16] = buffer_data_1[599:592] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_75[17] = buffer_data_1[607:600] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_75[18] = buffer_data_1[615:608] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_75[19] = buffer_data_1[623:616] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_75[20] = buffer_data_0[591:584] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_75[21] = buffer_data_0[599:592] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_75[22] = buffer_data_0[607:600] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_75[23] = buffer_data_0[615:608] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_75[24] = buffer_data_0[623:616] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_75 = kernel_img_mul_75[0] + kernel_img_mul_75[1] + kernel_img_mul_75[2] + 
                kernel_img_mul_75[3] + kernel_img_mul_75[4] + kernel_img_mul_75[5] + 
                kernel_img_mul_75[6] + kernel_img_mul_75[7] + kernel_img_mul_75[8] + 
                kernel_img_mul_75[9] + kernel_img_mul_75[10] + kernel_img_mul_75[11] + 
                kernel_img_mul_75[12] + kernel_img_mul_75[13] + kernel_img_mul_75[14] + 
                kernel_img_mul_75[15] + kernel_img_mul_75[16] + kernel_img_mul_75[17] + 
                kernel_img_mul_75[18] + kernel_img_mul_75[19] + kernel_img_mul_75[20] + 
                kernel_img_mul_75[21] + kernel_img_mul_75[22] + kernel_img_mul_75[23] + 
                kernel_img_mul_75[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[607:600] <= 'd0;
  else if (current_state==ST_START)
    blur_din[607:600] <= kernel_img_sum_75[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[607:600] <= 'd0;
end

wire  [39:0]  kernel_img_mul_76[0:24];
assign kernel_img_mul_76[0] = buffer_data_4[599:592] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_76[1] = buffer_data_4[607:600] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_76[2] = buffer_data_4[615:608] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_76[3] = buffer_data_4[623:616] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_76[4] = buffer_data_4[631:624] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_76[5] = buffer_data_3[599:592] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_76[6] = buffer_data_3[607:600] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_76[7] = buffer_data_3[615:608] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_76[8] = buffer_data_3[623:616] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_76[9] = buffer_data_3[631:624] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_76[10] = buffer_data_2[599:592] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_76[11] = buffer_data_2[607:600] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_76[12] = buffer_data_2[615:608] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_76[13] = buffer_data_2[623:616] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_76[14] = buffer_data_2[631:624] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_76[15] = buffer_data_1[599:592] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_76[16] = buffer_data_1[607:600] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_76[17] = buffer_data_1[615:608] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_76[18] = buffer_data_1[623:616] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_76[19] = buffer_data_1[631:624] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_76[20] = buffer_data_0[599:592] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_76[21] = buffer_data_0[607:600] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_76[22] = buffer_data_0[615:608] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_76[23] = buffer_data_0[623:616] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_76[24] = buffer_data_0[631:624] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_76 = kernel_img_mul_76[0] + kernel_img_mul_76[1] + kernel_img_mul_76[2] + 
                kernel_img_mul_76[3] + kernel_img_mul_76[4] + kernel_img_mul_76[5] + 
                kernel_img_mul_76[6] + kernel_img_mul_76[7] + kernel_img_mul_76[8] + 
                kernel_img_mul_76[9] + kernel_img_mul_76[10] + kernel_img_mul_76[11] + 
                kernel_img_mul_76[12] + kernel_img_mul_76[13] + kernel_img_mul_76[14] + 
                kernel_img_mul_76[15] + kernel_img_mul_76[16] + kernel_img_mul_76[17] + 
                kernel_img_mul_76[18] + kernel_img_mul_76[19] + kernel_img_mul_76[20] + 
                kernel_img_mul_76[21] + kernel_img_mul_76[22] + kernel_img_mul_76[23] + 
                kernel_img_mul_76[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[615:608] <= 'd0;
  else if (current_state==ST_START)
    blur_din[615:608] <= kernel_img_sum_76[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[615:608] <= 'd0;
end

wire  [39:0]  kernel_img_mul_77[0:24];
assign kernel_img_mul_77[0] = buffer_data_4[607:600] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_77[1] = buffer_data_4[615:608] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_77[2] = buffer_data_4[623:616] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_77[3] = buffer_data_4[631:624] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_77[4] = buffer_data_4[639:632] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_77[5] = buffer_data_3[607:600] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_77[6] = buffer_data_3[615:608] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_77[7] = buffer_data_3[623:616] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_77[8] = buffer_data_3[631:624] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_77[9] = buffer_data_3[639:632] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_77[10] = buffer_data_2[607:600] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_77[11] = buffer_data_2[615:608] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_77[12] = buffer_data_2[623:616] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_77[13] = buffer_data_2[631:624] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_77[14] = buffer_data_2[639:632] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_77[15] = buffer_data_1[607:600] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_77[16] = buffer_data_1[615:608] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_77[17] = buffer_data_1[623:616] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_77[18] = buffer_data_1[631:624] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_77[19] = buffer_data_1[639:632] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_77[20] = buffer_data_0[607:600] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_77[21] = buffer_data_0[615:608] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_77[22] = buffer_data_0[623:616] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_77[23] = buffer_data_0[631:624] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_77[24] = buffer_data_0[639:632] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_77 = kernel_img_mul_77[0] + kernel_img_mul_77[1] + kernel_img_mul_77[2] + 
                kernel_img_mul_77[3] + kernel_img_mul_77[4] + kernel_img_mul_77[5] + 
                kernel_img_mul_77[6] + kernel_img_mul_77[7] + kernel_img_mul_77[8] + 
                kernel_img_mul_77[9] + kernel_img_mul_77[10] + kernel_img_mul_77[11] + 
                kernel_img_mul_77[12] + kernel_img_mul_77[13] + kernel_img_mul_77[14] + 
                kernel_img_mul_77[15] + kernel_img_mul_77[16] + kernel_img_mul_77[17] + 
                kernel_img_mul_77[18] + kernel_img_mul_77[19] + kernel_img_mul_77[20] + 
                kernel_img_mul_77[21] + kernel_img_mul_77[22] + kernel_img_mul_77[23] + 
                kernel_img_mul_77[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[623:616] <= 'd0;
  else if (current_state==ST_START)
    blur_din[623:616] <= kernel_img_sum_77[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[623:616] <= 'd0;
end

wire  [39:0]  kernel_img_mul_78[0:24];
assign kernel_img_mul_78[0] = buffer_data_4[615:608] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_78[1] = buffer_data_4[623:616] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_78[2] = buffer_data_4[631:624] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_78[3] = buffer_data_4[639:632] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_78[4] = buffer_data_4[647:640] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_78[5] = buffer_data_3[615:608] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_78[6] = buffer_data_3[623:616] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_78[7] = buffer_data_3[631:624] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_78[8] = buffer_data_3[639:632] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_78[9] = buffer_data_3[647:640] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_78[10] = buffer_data_2[615:608] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_78[11] = buffer_data_2[623:616] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_78[12] = buffer_data_2[631:624] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_78[13] = buffer_data_2[639:632] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_78[14] = buffer_data_2[647:640] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_78[15] = buffer_data_1[615:608] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_78[16] = buffer_data_1[623:616] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_78[17] = buffer_data_1[631:624] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_78[18] = buffer_data_1[639:632] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_78[19] = buffer_data_1[647:640] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_78[20] = buffer_data_0[615:608] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_78[21] = buffer_data_0[623:616] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_78[22] = buffer_data_0[631:624] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_78[23] = buffer_data_0[639:632] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_78[24] = buffer_data_0[647:640] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_78 = kernel_img_mul_78[0] + kernel_img_mul_78[1] + kernel_img_mul_78[2] + 
                kernel_img_mul_78[3] + kernel_img_mul_78[4] + kernel_img_mul_78[5] + 
                kernel_img_mul_78[6] + kernel_img_mul_78[7] + kernel_img_mul_78[8] + 
                kernel_img_mul_78[9] + kernel_img_mul_78[10] + kernel_img_mul_78[11] + 
                kernel_img_mul_78[12] + kernel_img_mul_78[13] + kernel_img_mul_78[14] + 
                kernel_img_mul_78[15] + kernel_img_mul_78[16] + kernel_img_mul_78[17] + 
                kernel_img_mul_78[18] + kernel_img_mul_78[19] + kernel_img_mul_78[20] + 
                kernel_img_mul_78[21] + kernel_img_mul_78[22] + kernel_img_mul_78[23] + 
                kernel_img_mul_78[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[631:624] <= 'd0;
  else if (current_state==ST_START)
    blur_din[631:624] <= kernel_img_sum_78[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[631:624] <= 'd0;
end

wire  [39:0]  kernel_img_mul_79[0:24];
assign kernel_img_mul_79[0] = buffer_data_4[623:616] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_79[1] = buffer_data_4[631:624] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_79[2] = buffer_data_4[639:632] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_79[3] = buffer_data_4[647:640] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_79[4] = buffer_data_4[655:648] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_79[5] = buffer_data_3[623:616] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_79[6] = buffer_data_3[631:624] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_79[7] = buffer_data_3[639:632] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_79[8] = buffer_data_3[647:640] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_79[9] = buffer_data_3[655:648] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_79[10] = buffer_data_2[623:616] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_79[11] = buffer_data_2[631:624] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_79[12] = buffer_data_2[639:632] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_79[13] = buffer_data_2[647:640] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_79[14] = buffer_data_2[655:648] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_79[15] = buffer_data_1[623:616] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_79[16] = buffer_data_1[631:624] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_79[17] = buffer_data_1[639:632] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_79[18] = buffer_data_1[647:640] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_79[19] = buffer_data_1[655:648] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_79[20] = buffer_data_0[623:616] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_79[21] = buffer_data_0[631:624] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_79[22] = buffer_data_0[639:632] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_79[23] = buffer_data_0[647:640] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_79[24] = buffer_data_0[655:648] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_79 = kernel_img_mul_79[0] + kernel_img_mul_79[1] + kernel_img_mul_79[2] + 
                kernel_img_mul_79[3] + kernel_img_mul_79[4] + kernel_img_mul_79[5] + 
                kernel_img_mul_79[6] + kernel_img_mul_79[7] + kernel_img_mul_79[8] + 
                kernel_img_mul_79[9] + kernel_img_mul_79[10] + kernel_img_mul_79[11] + 
                kernel_img_mul_79[12] + kernel_img_mul_79[13] + kernel_img_mul_79[14] + 
                kernel_img_mul_79[15] + kernel_img_mul_79[16] + kernel_img_mul_79[17] + 
                kernel_img_mul_79[18] + kernel_img_mul_79[19] + kernel_img_mul_79[20] + 
                kernel_img_mul_79[21] + kernel_img_mul_79[22] + kernel_img_mul_79[23] + 
                kernel_img_mul_79[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[639:632] <= 'd0;
  else if (current_state==ST_START)
    blur_din[639:632] <= kernel_img_sum_79[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[639:632] <= 'd0;
end

wire  [39:0]  kernel_img_mul_80[0:24];
assign kernel_img_mul_80[0] = buffer_data_4[631:624] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_80[1] = buffer_data_4[639:632] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_80[2] = buffer_data_4[647:640] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_80[3] = buffer_data_4[655:648] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_80[4] = buffer_data_4[663:656] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_80[5] = buffer_data_3[631:624] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_80[6] = buffer_data_3[639:632] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_80[7] = buffer_data_3[647:640] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_80[8] = buffer_data_3[655:648] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_80[9] = buffer_data_3[663:656] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_80[10] = buffer_data_2[631:624] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_80[11] = buffer_data_2[639:632] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_80[12] = buffer_data_2[647:640] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_80[13] = buffer_data_2[655:648] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_80[14] = buffer_data_2[663:656] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_80[15] = buffer_data_1[631:624] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_80[16] = buffer_data_1[639:632] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_80[17] = buffer_data_1[647:640] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_80[18] = buffer_data_1[655:648] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_80[19] = buffer_data_1[663:656] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_80[20] = buffer_data_0[631:624] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_80[21] = buffer_data_0[639:632] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_80[22] = buffer_data_0[647:640] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_80[23] = buffer_data_0[655:648] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_80[24] = buffer_data_0[663:656] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_80 = kernel_img_mul_80[0] + kernel_img_mul_80[1] + kernel_img_mul_80[2] + 
                kernel_img_mul_80[3] + kernel_img_mul_80[4] + kernel_img_mul_80[5] + 
                kernel_img_mul_80[6] + kernel_img_mul_80[7] + kernel_img_mul_80[8] + 
                kernel_img_mul_80[9] + kernel_img_mul_80[10] + kernel_img_mul_80[11] + 
                kernel_img_mul_80[12] + kernel_img_mul_80[13] + kernel_img_mul_80[14] + 
                kernel_img_mul_80[15] + kernel_img_mul_80[16] + kernel_img_mul_80[17] + 
                kernel_img_mul_80[18] + kernel_img_mul_80[19] + kernel_img_mul_80[20] + 
                kernel_img_mul_80[21] + kernel_img_mul_80[22] + kernel_img_mul_80[23] + 
                kernel_img_mul_80[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[647:640] <= 'd0;
  else if (current_state==ST_START)
    blur_din[647:640] <= kernel_img_sum_80[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[647:640] <= 'd0;
end

wire  [39:0]  kernel_img_mul_81[0:24];
assign kernel_img_mul_81[0] = buffer_data_4[639:632] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_81[1] = buffer_data_4[647:640] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_81[2] = buffer_data_4[655:648] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_81[3] = buffer_data_4[663:656] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_81[4] = buffer_data_4[671:664] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_81[5] = buffer_data_3[639:632] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_81[6] = buffer_data_3[647:640] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_81[7] = buffer_data_3[655:648] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_81[8] = buffer_data_3[663:656] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_81[9] = buffer_data_3[671:664] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_81[10] = buffer_data_2[639:632] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_81[11] = buffer_data_2[647:640] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_81[12] = buffer_data_2[655:648] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_81[13] = buffer_data_2[663:656] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_81[14] = buffer_data_2[671:664] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_81[15] = buffer_data_1[639:632] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_81[16] = buffer_data_1[647:640] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_81[17] = buffer_data_1[655:648] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_81[18] = buffer_data_1[663:656] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_81[19] = buffer_data_1[671:664] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_81[20] = buffer_data_0[639:632] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_81[21] = buffer_data_0[647:640] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_81[22] = buffer_data_0[655:648] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_81[23] = buffer_data_0[663:656] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_81[24] = buffer_data_0[671:664] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_81 = kernel_img_mul_81[0] + kernel_img_mul_81[1] + kernel_img_mul_81[2] + 
                kernel_img_mul_81[3] + kernel_img_mul_81[4] + kernel_img_mul_81[5] + 
                kernel_img_mul_81[6] + kernel_img_mul_81[7] + kernel_img_mul_81[8] + 
                kernel_img_mul_81[9] + kernel_img_mul_81[10] + kernel_img_mul_81[11] + 
                kernel_img_mul_81[12] + kernel_img_mul_81[13] + kernel_img_mul_81[14] + 
                kernel_img_mul_81[15] + kernel_img_mul_81[16] + kernel_img_mul_81[17] + 
                kernel_img_mul_81[18] + kernel_img_mul_81[19] + kernel_img_mul_81[20] + 
                kernel_img_mul_81[21] + kernel_img_mul_81[22] + kernel_img_mul_81[23] + 
                kernel_img_mul_81[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[655:648] <= 'd0;
  else if (current_state==ST_START)
    blur_din[655:648] <= kernel_img_sum_81[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[655:648] <= 'd0;
end

wire  [39:0]  kernel_img_mul_82[0:24];
assign kernel_img_mul_82[0] = buffer_data_4[647:640] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_82[1] = buffer_data_4[655:648] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_82[2] = buffer_data_4[663:656] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_82[3] = buffer_data_4[671:664] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_82[4] = buffer_data_4[679:672] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_82[5] = buffer_data_3[647:640] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_82[6] = buffer_data_3[655:648] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_82[7] = buffer_data_3[663:656] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_82[8] = buffer_data_3[671:664] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_82[9] = buffer_data_3[679:672] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_82[10] = buffer_data_2[647:640] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_82[11] = buffer_data_2[655:648] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_82[12] = buffer_data_2[663:656] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_82[13] = buffer_data_2[671:664] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_82[14] = buffer_data_2[679:672] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_82[15] = buffer_data_1[647:640] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_82[16] = buffer_data_1[655:648] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_82[17] = buffer_data_1[663:656] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_82[18] = buffer_data_1[671:664] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_82[19] = buffer_data_1[679:672] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_82[20] = buffer_data_0[647:640] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_82[21] = buffer_data_0[655:648] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_82[22] = buffer_data_0[663:656] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_82[23] = buffer_data_0[671:664] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_82[24] = buffer_data_0[679:672] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_82 = kernel_img_mul_82[0] + kernel_img_mul_82[1] + kernel_img_mul_82[2] + 
                kernel_img_mul_82[3] + kernel_img_mul_82[4] + kernel_img_mul_82[5] + 
                kernel_img_mul_82[6] + kernel_img_mul_82[7] + kernel_img_mul_82[8] + 
                kernel_img_mul_82[9] + kernel_img_mul_82[10] + kernel_img_mul_82[11] + 
                kernel_img_mul_82[12] + kernel_img_mul_82[13] + kernel_img_mul_82[14] + 
                kernel_img_mul_82[15] + kernel_img_mul_82[16] + kernel_img_mul_82[17] + 
                kernel_img_mul_82[18] + kernel_img_mul_82[19] + kernel_img_mul_82[20] + 
                kernel_img_mul_82[21] + kernel_img_mul_82[22] + kernel_img_mul_82[23] + 
                kernel_img_mul_82[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[663:656] <= 'd0;
  else if (current_state==ST_START)
    blur_din[663:656] <= kernel_img_sum_82[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[663:656] <= 'd0;
end

wire  [39:0]  kernel_img_mul_83[0:24];
assign kernel_img_mul_83[0] = buffer_data_4[655:648] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_83[1] = buffer_data_4[663:656] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_83[2] = buffer_data_4[671:664] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_83[3] = buffer_data_4[679:672] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_83[4] = buffer_data_4[687:680] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_83[5] = buffer_data_3[655:648] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_83[6] = buffer_data_3[663:656] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_83[7] = buffer_data_3[671:664] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_83[8] = buffer_data_3[679:672] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_83[9] = buffer_data_3[687:680] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_83[10] = buffer_data_2[655:648] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_83[11] = buffer_data_2[663:656] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_83[12] = buffer_data_2[671:664] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_83[13] = buffer_data_2[679:672] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_83[14] = buffer_data_2[687:680] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_83[15] = buffer_data_1[655:648] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_83[16] = buffer_data_1[663:656] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_83[17] = buffer_data_1[671:664] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_83[18] = buffer_data_1[679:672] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_83[19] = buffer_data_1[687:680] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_83[20] = buffer_data_0[655:648] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_83[21] = buffer_data_0[663:656] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_83[22] = buffer_data_0[671:664] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_83[23] = buffer_data_0[679:672] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_83[24] = buffer_data_0[687:680] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_83 = kernel_img_mul_83[0] + kernel_img_mul_83[1] + kernel_img_mul_83[2] + 
                kernel_img_mul_83[3] + kernel_img_mul_83[4] + kernel_img_mul_83[5] + 
                kernel_img_mul_83[6] + kernel_img_mul_83[7] + kernel_img_mul_83[8] + 
                kernel_img_mul_83[9] + kernel_img_mul_83[10] + kernel_img_mul_83[11] + 
                kernel_img_mul_83[12] + kernel_img_mul_83[13] + kernel_img_mul_83[14] + 
                kernel_img_mul_83[15] + kernel_img_mul_83[16] + kernel_img_mul_83[17] + 
                kernel_img_mul_83[18] + kernel_img_mul_83[19] + kernel_img_mul_83[20] + 
                kernel_img_mul_83[21] + kernel_img_mul_83[22] + kernel_img_mul_83[23] + 
                kernel_img_mul_83[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[671:664] <= 'd0;
  else if (current_state==ST_START)
    blur_din[671:664] <= kernel_img_sum_83[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[671:664] <= 'd0;
end

wire  [39:0]  kernel_img_mul_84[0:24];
assign kernel_img_mul_84[0] = buffer_data_4[663:656] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_84[1] = buffer_data_4[671:664] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_84[2] = buffer_data_4[679:672] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_84[3] = buffer_data_4[687:680] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_84[4] = buffer_data_4[695:688] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_84[5] = buffer_data_3[663:656] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_84[6] = buffer_data_3[671:664] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_84[7] = buffer_data_3[679:672] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_84[8] = buffer_data_3[687:680] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_84[9] = buffer_data_3[695:688] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_84[10] = buffer_data_2[663:656] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_84[11] = buffer_data_2[671:664] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_84[12] = buffer_data_2[679:672] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_84[13] = buffer_data_2[687:680] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_84[14] = buffer_data_2[695:688] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_84[15] = buffer_data_1[663:656] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_84[16] = buffer_data_1[671:664] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_84[17] = buffer_data_1[679:672] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_84[18] = buffer_data_1[687:680] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_84[19] = buffer_data_1[695:688] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_84[20] = buffer_data_0[663:656] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_84[21] = buffer_data_0[671:664] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_84[22] = buffer_data_0[679:672] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_84[23] = buffer_data_0[687:680] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_84[24] = buffer_data_0[695:688] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_84 = kernel_img_mul_84[0] + kernel_img_mul_84[1] + kernel_img_mul_84[2] + 
                kernel_img_mul_84[3] + kernel_img_mul_84[4] + kernel_img_mul_84[5] + 
                kernel_img_mul_84[6] + kernel_img_mul_84[7] + kernel_img_mul_84[8] + 
                kernel_img_mul_84[9] + kernel_img_mul_84[10] + kernel_img_mul_84[11] + 
                kernel_img_mul_84[12] + kernel_img_mul_84[13] + kernel_img_mul_84[14] + 
                kernel_img_mul_84[15] + kernel_img_mul_84[16] + kernel_img_mul_84[17] + 
                kernel_img_mul_84[18] + kernel_img_mul_84[19] + kernel_img_mul_84[20] + 
                kernel_img_mul_84[21] + kernel_img_mul_84[22] + kernel_img_mul_84[23] + 
                kernel_img_mul_84[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[679:672] <= 'd0;
  else if (current_state==ST_START)
    blur_din[679:672] <= kernel_img_sum_84[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[679:672] <= 'd0;
end

wire  [39:0]  kernel_img_mul_85[0:24];
assign kernel_img_mul_85[0] = buffer_data_4[671:664] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_85[1] = buffer_data_4[679:672] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_85[2] = buffer_data_4[687:680] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_85[3] = buffer_data_4[695:688] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_85[4] = buffer_data_4[703:696] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_85[5] = buffer_data_3[671:664] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_85[6] = buffer_data_3[679:672] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_85[7] = buffer_data_3[687:680] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_85[8] = buffer_data_3[695:688] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_85[9] = buffer_data_3[703:696] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_85[10] = buffer_data_2[671:664] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_85[11] = buffer_data_2[679:672] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_85[12] = buffer_data_2[687:680] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_85[13] = buffer_data_2[695:688] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_85[14] = buffer_data_2[703:696] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_85[15] = buffer_data_1[671:664] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_85[16] = buffer_data_1[679:672] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_85[17] = buffer_data_1[687:680] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_85[18] = buffer_data_1[695:688] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_85[19] = buffer_data_1[703:696] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_85[20] = buffer_data_0[671:664] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_85[21] = buffer_data_0[679:672] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_85[22] = buffer_data_0[687:680] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_85[23] = buffer_data_0[695:688] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_85[24] = buffer_data_0[703:696] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_85 = kernel_img_mul_85[0] + kernel_img_mul_85[1] + kernel_img_mul_85[2] + 
                kernel_img_mul_85[3] + kernel_img_mul_85[4] + kernel_img_mul_85[5] + 
                kernel_img_mul_85[6] + kernel_img_mul_85[7] + kernel_img_mul_85[8] + 
                kernel_img_mul_85[9] + kernel_img_mul_85[10] + kernel_img_mul_85[11] + 
                kernel_img_mul_85[12] + kernel_img_mul_85[13] + kernel_img_mul_85[14] + 
                kernel_img_mul_85[15] + kernel_img_mul_85[16] + kernel_img_mul_85[17] + 
                kernel_img_mul_85[18] + kernel_img_mul_85[19] + kernel_img_mul_85[20] + 
                kernel_img_mul_85[21] + kernel_img_mul_85[22] + kernel_img_mul_85[23] + 
                kernel_img_mul_85[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[687:680] <= 'd0;
  else if (current_state==ST_START)
    blur_din[687:680] <= kernel_img_sum_85[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[687:680] <= 'd0;
end

wire  [39:0]  kernel_img_mul_86[0:24];
assign kernel_img_mul_86[0] = buffer_data_4[679:672] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_86[1] = buffer_data_4[687:680] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_86[2] = buffer_data_4[695:688] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_86[3] = buffer_data_4[703:696] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_86[4] = buffer_data_4[711:704] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_86[5] = buffer_data_3[679:672] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_86[6] = buffer_data_3[687:680] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_86[7] = buffer_data_3[695:688] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_86[8] = buffer_data_3[703:696] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_86[9] = buffer_data_3[711:704] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_86[10] = buffer_data_2[679:672] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_86[11] = buffer_data_2[687:680] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_86[12] = buffer_data_2[695:688] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_86[13] = buffer_data_2[703:696] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_86[14] = buffer_data_2[711:704] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_86[15] = buffer_data_1[679:672] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_86[16] = buffer_data_1[687:680] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_86[17] = buffer_data_1[695:688] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_86[18] = buffer_data_1[703:696] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_86[19] = buffer_data_1[711:704] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_86[20] = buffer_data_0[679:672] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_86[21] = buffer_data_0[687:680] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_86[22] = buffer_data_0[695:688] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_86[23] = buffer_data_0[703:696] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_86[24] = buffer_data_0[711:704] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_86 = kernel_img_mul_86[0] + kernel_img_mul_86[1] + kernel_img_mul_86[2] + 
                kernel_img_mul_86[3] + kernel_img_mul_86[4] + kernel_img_mul_86[5] + 
                kernel_img_mul_86[6] + kernel_img_mul_86[7] + kernel_img_mul_86[8] + 
                kernel_img_mul_86[9] + kernel_img_mul_86[10] + kernel_img_mul_86[11] + 
                kernel_img_mul_86[12] + kernel_img_mul_86[13] + kernel_img_mul_86[14] + 
                kernel_img_mul_86[15] + kernel_img_mul_86[16] + kernel_img_mul_86[17] + 
                kernel_img_mul_86[18] + kernel_img_mul_86[19] + kernel_img_mul_86[20] + 
                kernel_img_mul_86[21] + kernel_img_mul_86[22] + kernel_img_mul_86[23] + 
                kernel_img_mul_86[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[695:688] <= 'd0;
  else if (current_state==ST_START)
    blur_din[695:688] <= kernel_img_sum_86[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[695:688] <= 'd0;
end

wire  [39:0]  kernel_img_mul_87[0:24];
assign kernel_img_mul_87[0] = buffer_data_4[687:680] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_87[1] = buffer_data_4[695:688] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_87[2] = buffer_data_4[703:696] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_87[3] = buffer_data_4[711:704] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_87[4] = buffer_data_4[719:712] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_87[5] = buffer_data_3[687:680] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_87[6] = buffer_data_3[695:688] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_87[7] = buffer_data_3[703:696] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_87[8] = buffer_data_3[711:704] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_87[9] = buffer_data_3[719:712] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_87[10] = buffer_data_2[687:680] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_87[11] = buffer_data_2[695:688] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_87[12] = buffer_data_2[703:696] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_87[13] = buffer_data_2[711:704] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_87[14] = buffer_data_2[719:712] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_87[15] = buffer_data_1[687:680] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_87[16] = buffer_data_1[695:688] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_87[17] = buffer_data_1[703:696] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_87[18] = buffer_data_1[711:704] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_87[19] = buffer_data_1[719:712] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_87[20] = buffer_data_0[687:680] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_87[21] = buffer_data_0[695:688] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_87[22] = buffer_data_0[703:696] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_87[23] = buffer_data_0[711:704] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_87[24] = buffer_data_0[719:712] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_87 = kernel_img_mul_87[0] + kernel_img_mul_87[1] + kernel_img_mul_87[2] + 
                kernel_img_mul_87[3] + kernel_img_mul_87[4] + kernel_img_mul_87[5] + 
                kernel_img_mul_87[6] + kernel_img_mul_87[7] + kernel_img_mul_87[8] + 
                kernel_img_mul_87[9] + kernel_img_mul_87[10] + kernel_img_mul_87[11] + 
                kernel_img_mul_87[12] + kernel_img_mul_87[13] + kernel_img_mul_87[14] + 
                kernel_img_mul_87[15] + kernel_img_mul_87[16] + kernel_img_mul_87[17] + 
                kernel_img_mul_87[18] + kernel_img_mul_87[19] + kernel_img_mul_87[20] + 
                kernel_img_mul_87[21] + kernel_img_mul_87[22] + kernel_img_mul_87[23] + 
                kernel_img_mul_87[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[703:696] <= 'd0;
  else if (current_state==ST_START)
    blur_din[703:696] <= kernel_img_sum_87[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[703:696] <= 'd0;
end

wire  [39:0]  kernel_img_mul_88[0:24];
assign kernel_img_mul_88[0] = buffer_data_4[695:688] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_88[1] = buffer_data_4[703:696] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_88[2] = buffer_data_4[711:704] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_88[3] = buffer_data_4[719:712] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_88[4] = buffer_data_4[727:720] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_88[5] = buffer_data_3[695:688] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_88[6] = buffer_data_3[703:696] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_88[7] = buffer_data_3[711:704] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_88[8] = buffer_data_3[719:712] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_88[9] = buffer_data_3[727:720] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_88[10] = buffer_data_2[695:688] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_88[11] = buffer_data_2[703:696] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_88[12] = buffer_data_2[711:704] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_88[13] = buffer_data_2[719:712] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_88[14] = buffer_data_2[727:720] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_88[15] = buffer_data_1[695:688] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_88[16] = buffer_data_1[703:696] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_88[17] = buffer_data_1[711:704] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_88[18] = buffer_data_1[719:712] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_88[19] = buffer_data_1[727:720] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_88[20] = buffer_data_0[695:688] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_88[21] = buffer_data_0[703:696] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_88[22] = buffer_data_0[711:704] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_88[23] = buffer_data_0[719:712] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_88[24] = buffer_data_0[727:720] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_88 = kernel_img_mul_88[0] + kernel_img_mul_88[1] + kernel_img_mul_88[2] + 
                kernel_img_mul_88[3] + kernel_img_mul_88[4] + kernel_img_mul_88[5] + 
                kernel_img_mul_88[6] + kernel_img_mul_88[7] + kernel_img_mul_88[8] + 
                kernel_img_mul_88[9] + kernel_img_mul_88[10] + kernel_img_mul_88[11] + 
                kernel_img_mul_88[12] + kernel_img_mul_88[13] + kernel_img_mul_88[14] + 
                kernel_img_mul_88[15] + kernel_img_mul_88[16] + kernel_img_mul_88[17] + 
                kernel_img_mul_88[18] + kernel_img_mul_88[19] + kernel_img_mul_88[20] + 
                kernel_img_mul_88[21] + kernel_img_mul_88[22] + kernel_img_mul_88[23] + 
                kernel_img_mul_88[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[711:704] <= 'd0;
  else if (current_state==ST_START)
    blur_din[711:704] <= kernel_img_sum_88[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[711:704] <= 'd0;
end

wire  [39:0]  kernel_img_mul_89[0:24];
assign kernel_img_mul_89[0] = buffer_data_4[703:696] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_89[1] = buffer_data_4[711:704] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_89[2] = buffer_data_4[719:712] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_89[3] = buffer_data_4[727:720] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_89[4] = buffer_data_4[735:728] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_89[5] = buffer_data_3[703:696] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_89[6] = buffer_data_3[711:704] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_89[7] = buffer_data_3[719:712] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_89[8] = buffer_data_3[727:720] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_89[9] = buffer_data_3[735:728] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_89[10] = buffer_data_2[703:696] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_89[11] = buffer_data_2[711:704] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_89[12] = buffer_data_2[719:712] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_89[13] = buffer_data_2[727:720] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_89[14] = buffer_data_2[735:728] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_89[15] = buffer_data_1[703:696] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_89[16] = buffer_data_1[711:704] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_89[17] = buffer_data_1[719:712] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_89[18] = buffer_data_1[727:720] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_89[19] = buffer_data_1[735:728] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_89[20] = buffer_data_0[703:696] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_89[21] = buffer_data_0[711:704] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_89[22] = buffer_data_0[719:712] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_89[23] = buffer_data_0[727:720] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_89[24] = buffer_data_0[735:728] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_89 = kernel_img_mul_89[0] + kernel_img_mul_89[1] + kernel_img_mul_89[2] + 
                kernel_img_mul_89[3] + kernel_img_mul_89[4] + kernel_img_mul_89[5] + 
                kernel_img_mul_89[6] + kernel_img_mul_89[7] + kernel_img_mul_89[8] + 
                kernel_img_mul_89[9] + kernel_img_mul_89[10] + kernel_img_mul_89[11] + 
                kernel_img_mul_89[12] + kernel_img_mul_89[13] + kernel_img_mul_89[14] + 
                kernel_img_mul_89[15] + kernel_img_mul_89[16] + kernel_img_mul_89[17] + 
                kernel_img_mul_89[18] + kernel_img_mul_89[19] + kernel_img_mul_89[20] + 
                kernel_img_mul_89[21] + kernel_img_mul_89[22] + kernel_img_mul_89[23] + 
                kernel_img_mul_89[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[719:712] <= 'd0;
  else if (current_state==ST_START)
    blur_din[719:712] <= kernel_img_sum_89[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[719:712] <= 'd0;
end

wire  [39:0]  kernel_img_mul_90[0:24];
assign kernel_img_mul_90[0] = buffer_data_4[711:704] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_90[1] = buffer_data_4[719:712] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_90[2] = buffer_data_4[727:720] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_90[3] = buffer_data_4[735:728] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_90[4] = buffer_data_4[743:736] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_90[5] = buffer_data_3[711:704] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_90[6] = buffer_data_3[719:712] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_90[7] = buffer_data_3[727:720] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_90[8] = buffer_data_3[735:728] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_90[9] = buffer_data_3[743:736] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_90[10] = buffer_data_2[711:704] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_90[11] = buffer_data_2[719:712] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_90[12] = buffer_data_2[727:720] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_90[13] = buffer_data_2[735:728] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_90[14] = buffer_data_2[743:736] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_90[15] = buffer_data_1[711:704] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_90[16] = buffer_data_1[719:712] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_90[17] = buffer_data_1[727:720] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_90[18] = buffer_data_1[735:728] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_90[19] = buffer_data_1[743:736] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_90[20] = buffer_data_0[711:704] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_90[21] = buffer_data_0[719:712] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_90[22] = buffer_data_0[727:720] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_90[23] = buffer_data_0[735:728] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_90[24] = buffer_data_0[743:736] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_90 = kernel_img_mul_90[0] + kernel_img_mul_90[1] + kernel_img_mul_90[2] + 
                kernel_img_mul_90[3] + kernel_img_mul_90[4] + kernel_img_mul_90[5] + 
                kernel_img_mul_90[6] + kernel_img_mul_90[7] + kernel_img_mul_90[8] + 
                kernel_img_mul_90[9] + kernel_img_mul_90[10] + kernel_img_mul_90[11] + 
                kernel_img_mul_90[12] + kernel_img_mul_90[13] + kernel_img_mul_90[14] + 
                kernel_img_mul_90[15] + kernel_img_mul_90[16] + kernel_img_mul_90[17] + 
                kernel_img_mul_90[18] + kernel_img_mul_90[19] + kernel_img_mul_90[20] + 
                kernel_img_mul_90[21] + kernel_img_mul_90[22] + kernel_img_mul_90[23] + 
                kernel_img_mul_90[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[727:720] <= 'd0;
  else if (current_state==ST_START)
    blur_din[727:720] <= kernel_img_sum_90[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[727:720] <= 'd0;
end

wire  [39:0]  kernel_img_mul_91[0:24];
assign kernel_img_mul_91[0] = buffer_data_4[719:712] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_91[1] = buffer_data_4[727:720] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_91[2] = buffer_data_4[735:728] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_91[3] = buffer_data_4[743:736] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_91[4] = buffer_data_4[751:744] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_91[5] = buffer_data_3[719:712] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_91[6] = buffer_data_3[727:720] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_91[7] = buffer_data_3[735:728] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_91[8] = buffer_data_3[743:736] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_91[9] = buffer_data_3[751:744] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_91[10] = buffer_data_2[719:712] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_91[11] = buffer_data_2[727:720] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_91[12] = buffer_data_2[735:728] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_91[13] = buffer_data_2[743:736] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_91[14] = buffer_data_2[751:744] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_91[15] = buffer_data_1[719:712] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_91[16] = buffer_data_1[727:720] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_91[17] = buffer_data_1[735:728] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_91[18] = buffer_data_1[743:736] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_91[19] = buffer_data_1[751:744] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_91[20] = buffer_data_0[719:712] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_91[21] = buffer_data_0[727:720] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_91[22] = buffer_data_0[735:728] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_91[23] = buffer_data_0[743:736] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_91[24] = buffer_data_0[751:744] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_91 = kernel_img_mul_91[0] + kernel_img_mul_91[1] + kernel_img_mul_91[2] + 
                kernel_img_mul_91[3] + kernel_img_mul_91[4] + kernel_img_mul_91[5] + 
                kernel_img_mul_91[6] + kernel_img_mul_91[7] + kernel_img_mul_91[8] + 
                kernel_img_mul_91[9] + kernel_img_mul_91[10] + kernel_img_mul_91[11] + 
                kernel_img_mul_91[12] + kernel_img_mul_91[13] + kernel_img_mul_91[14] + 
                kernel_img_mul_91[15] + kernel_img_mul_91[16] + kernel_img_mul_91[17] + 
                kernel_img_mul_91[18] + kernel_img_mul_91[19] + kernel_img_mul_91[20] + 
                kernel_img_mul_91[21] + kernel_img_mul_91[22] + kernel_img_mul_91[23] + 
                kernel_img_mul_91[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[735:728] <= 'd0;
  else if (current_state==ST_START)
    blur_din[735:728] <= kernel_img_sum_91[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[735:728] <= 'd0;
end

wire  [39:0]  kernel_img_mul_92[0:24];
assign kernel_img_mul_92[0] = buffer_data_4[727:720] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_92[1] = buffer_data_4[735:728] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_92[2] = buffer_data_4[743:736] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_92[3] = buffer_data_4[751:744] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_92[4] = buffer_data_4[759:752] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_92[5] = buffer_data_3[727:720] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_92[6] = buffer_data_3[735:728] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_92[7] = buffer_data_3[743:736] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_92[8] = buffer_data_3[751:744] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_92[9] = buffer_data_3[759:752] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_92[10] = buffer_data_2[727:720] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_92[11] = buffer_data_2[735:728] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_92[12] = buffer_data_2[743:736] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_92[13] = buffer_data_2[751:744] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_92[14] = buffer_data_2[759:752] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_92[15] = buffer_data_1[727:720] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_92[16] = buffer_data_1[735:728] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_92[17] = buffer_data_1[743:736] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_92[18] = buffer_data_1[751:744] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_92[19] = buffer_data_1[759:752] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_92[20] = buffer_data_0[727:720] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_92[21] = buffer_data_0[735:728] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_92[22] = buffer_data_0[743:736] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_92[23] = buffer_data_0[751:744] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_92[24] = buffer_data_0[759:752] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_92 = kernel_img_mul_92[0] + kernel_img_mul_92[1] + kernel_img_mul_92[2] + 
                kernel_img_mul_92[3] + kernel_img_mul_92[4] + kernel_img_mul_92[5] + 
                kernel_img_mul_92[6] + kernel_img_mul_92[7] + kernel_img_mul_92[8] + 
                kernel_img_mul_92[9] + kernel_img_mul_92[10] + kernel_img_mul_92[11] + 
                kernel_img_mul_92[12] + kernel_img_mul_92[13] + kernel_img_mul_92[14] + 
                kernel_img_mul_92[15] + kernel_img_mul_92[16] + kernel_img_mul_92[17] + 
                kernel_img_mul_92[18] + kernel_img_mul_92[19] + kernel_img_mul_92[20] + 
                kernel_img_mul_92[21] + kernel_img_mul_92[22] + kernel_img_mul_92[23] + 
                kernel_img_mul_92[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[743:736] <= 'd0;
  else if (current_state==ST_START)
    blur_din[743:736] <= kernel_img_sum_92[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[743:736] <= 'd0;
end

wire  [39:0]  kernel_img_mul_93[0:24];
assign kernel_img_mul_93[0] = buffer_data_4[735:728] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_93[1] = buffer_data_4[743:736] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_93[2] = buffer_data_4[751:744] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_93[3] = buffer_data_4[759:752] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_93[4] = buffer_data_4[767:760] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_93[5] = buffer_data_3[735:728] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_93[6] = buffer_data_3[743:736] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_93[7] = buffer_data_3[751:744] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_93[8] = buffer_data_3[759:752] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_93[9] = buffer_data_3[767:760] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_93[10] = buffer_data_2[735:728] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_93[11] = buffer_data_2[743:736] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_93[12] = buffer_data_2[751:744] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_93[13] = buffer_data_2[759:752] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_93[14] = buffer_data_2[767:760] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_93[15] = buffer_data_1[735:728] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_93[16] = buffer_data_1[743:736] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_93[17] = buffer_data_1[751:744] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_93[18] = buffer_data_1[759:752] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_93[19] = buffer_data_1[767:760] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_93[20] = buffer_data_0[735:728] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_93[21] = buffer_data_0[743:736] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_93[22] = buffer_data_0[751:744] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_93[23] = buffer_data_0[759:752] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_93[24] = buffer_data_0[767:760] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_93 = kernel_img_mul_93[0] + kernel_img_mul_93[1] + kernel_img_mul_93[2] + 
                kernel_img_mul_93[3] + kernel_img_mul_93[4] + kernel_img_mul_93[5] + 
                kernel_img_mul_93[6] + kernel_img_mul_93[7] + kernel_img_mul_93[8] + 
                kernel_img_mul_93[9] + kernel_img_mul_93[10] + kernel_img_mul_93[11] + 
                kernel_img_mul_93[12] + kernel_img_mul_93[13] + kernel_img_mul_93[14] + 
                kernel_img_mul_93[15] + kernel_img_mul_93[16] + kernel_img_mul_93[17] + 
                kernel_img_mul_93[18] + kernel_img_mul_93[19] + kernel_img_mul_93[20] + 
                kernel_img_mul_93[21] + kernel_img_mul_93[22] + kernel_img_mul_93[23] + 
                kernel_img_mul_93[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[751:744] <= 'd0;
  else if (current_state==ST_START)
    blur_din[751:744] <= kernel_img_sum_93[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[751:744] <= 'd0;
end

wire  [39:0]  kernel_img_mul_94[0:24];
assign kernel_img_mul_94[0] = buffer_data_4[743:736] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_94[1] = buffer_data_4[751:744] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_94[2] = buffer_data_4[759:752] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_94[3] = buffer_data_4[767:760] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_94[4] = buffer_data_4[775:768] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_94[5] = buffer_data_3[743:736] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_94[6] = buffer_data_3[751:744] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_94[7] = buffer_data_3[759:752] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_94[8] = buffer_data_3[767:760] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_94[9] = buffer_data_3[775:768] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_94[10] = buffer_data_2[743:736] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_94[11] = buffer_data_2[751:744] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_94[12] = buffer_data_2[759:752] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_94[13] = buffer_data_2[767:760] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_94[14] = buffer_data_2[775:768] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_94[15] = buffer_data_1[743:736] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_94[16] = buffer_data_1[751:744] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_94[17] = buffer_data_1[759:752] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_94[18] = buffer_data_1[767:760] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_94[19] = buffer_data_1[775:768] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_94[20] = buffer_data_0[743:736] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_94[21] = buffer_data_0[751:744] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_94[22] = buffer_data_0[759:752] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_94[23] = buffer_data_0[767:760] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_94[24] = buffer_data_0[775:768] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_94 = kernel_img_mul_94[0] + kernel_img_mul_94[1] + kernel_img_mul_94[2] + 
                kernel_img_mul_94[3] + kernel_img_mul_94[4] + kernel_img_mul_94[5] + 
                kernel_img_mul_94[6] + kernel_img_mul_94[7] + kernel_img_mul_94[8] + 
                kernel_img_mul_94[9] + kernel_img_mul_94[10] + kernel_img_mul_94[11] + 
                kernel_img_mul_94[12] + kernel_img_mul_94[13] + kernel_img_mul_94[14] + 
                kernel_img_mul_94[15] + kernel_img_mul_94[16] + kernel_img_mul_94[17] + 
                kernel_img_mul_94[18] + kernel_img_mul_94[19] + kernel_img_mul_94[20] + 
                kernel_img_mul_94[21] + kernel_img_mul_94[22] + kernel_img_mul_94[23] + 
                kernel_img_mul_94[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[759:752] <= 'd0;
  else if (current_state==ST_START)
    blur_din[759:752] <= kernel_img_sum_94[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[759:752] <= 'd0;
end

wire  [39:0]  kernel_img_mul_95[0:24];
assign kernel_img_mul_95[0] = buffer_data_4[751:744] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_95[1] = buffer_data_4[759:752] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_95[2] = buffer_data_4[767:760] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_95[3] = buffer_data_4[775:768] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_95[4] = buffer_data_4[783:776] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_95[5] = buffer_data_3[751:744] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_95[6] = buffer_data_3[759:752] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_95[7] = buffer_data_3[767:760] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_95[8] = buffer_data_3[775:768] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_95[9] = buffer_data_3[783:776] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_95[10] = buffer_data_2[751:744] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_95[11] = buffer_data_2[759:752] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_95[12] = buffer_data_2[767:760] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_95[13] = buffer_data_2[775:768] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_95[14] = buffer_data_2[783:776] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_95[15] = buffer_data_1[751:744] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_95[16] = buffer_data_1[759:752] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_95[17] = buffer_data_1[767:760] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_95[18] = buffer_data_1[775:768] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_95[19] = buffer_data_1[783:776] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_95[20] = buffer_data_0[751:744] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_95[21] = buffer_data_0[759:752] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_95[22] = buffer_data_0[767:760] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_95[23] = buffer_data_0[775:768] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_95[24] = buffer_data_0[783:776] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_95 = kernel_img_mul_95[0] + kernel_img_mul_95[1] + kernel_img_mul_95[2] + 
                kernel_img_mul_95[3] + kernel_img_mul_95[4] + kernel_img_mul_95[5] + 
                kernel_img_mul_95[6] + kernel_img_mul_95[7] + kernel_img_mul_95[8] + 
                kernel_img_mul_95[9] + kernel_img_mul_95[10] + kernel_img_mul_95[11] + 
                kernel_img_mul_95[12] + kernel_img_mul_95[13] + kernel_img_mul_95[14] + 
                kernel_img_mul_95[15] + kernel_img_mul_95[16] + kernel_img_mul_95[17] + 
                kernel_img_mul_95[18] + kernel_img_mul_95[19] + kernel_img_mul_95[20] + 
                kernel_img_mul_95[21] + kernel_img_mul_95[22] + kernel_img_mul_95[23] + 
                kernel_img_mul_95[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[767:760] <= 'd0;
  else if (current_state==ST_START)
    blur_din[767:760] <= kernel_img_sum_95[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[767:760] <= 'd0;
end

wire  [39:0]  kernel_img_mul_96[0:24];
assign kernel_img_mul_96[0] = buffer_data_4[759:752] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_96[1] = buffer_data_4[767:760] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_96[2] = buffer_data_4[775:768] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_96[3] = buffer_data_4[783:776] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_96[4] = buffer_data_4[791:784] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_96[5] = buffer_data_3[759:752] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_96[6] = buffer_data_3[767:760] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_96[7] = buffer_data_3[775:768] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_96[8] = buffer_data_3[783:776] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_96[9] = buffer_data_3[791:784] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_96[10] = buffer_data_2[759:752] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_96[11] = buffer_data_2[767:760] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_96[12] = buffer_data_2[775:768] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_96[13] = buffer_data_2[783:776] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_96[14] = buffer_data_2[791:784] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_96[15] = buffer_data_1[759:752] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_96[16] = buffer_data_1[767:760] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_96[17] = buffer_data_1[775:768] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_96[18] = buffer_data_1[783:776] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_96[19] = buffer_data_1[791:784] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_96[20] = buffer_data_0[759:752] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_96[21] = buffer_data_0[767:760] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_96[22] = buffer_data_0[775:768] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_96[23] = buffer_data_0[783:776] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_96[24] = buffer_data_0[791:784] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_96 = kernel_img_mul_96[0] + kernel_img_mul_96[1] + kernel_img_mul_96[2] + 
                kernel_img_mul_96[3] + kernel_img_mul_96[4] + kernel_img_mul_96[5] + 
                kernel_img_mul_96[6] + kernel_img_mul_96[7] + kernel_img_mul_96[8] + 
                kernel_img_mul_96[9] + kernel_img_mul_96[10] + kernel_img_mul_96[11] + 
                kernel_img_mul_96[12] + kernel_img_mul_96[13] + kernel_img_mul_96[14] + 
                kernel_img_mul_96[15] + kernel_img_mul_96[16] + kernel_img_mul_96[17] + 
                kernel_img_mul_96[18] + kernel_img_mul_96[19] + kernel_img_mul_96[20] + 
                kernel_img_mul_96[21] + kernel_img_mul_96[22] + kernel_img_mul_96[23] + 
                kernel_img_mul_96[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[775:768] <= 'd0;
  else if (current_state==ST_START)
    blur_din[775:768] <= kernel_img_sum_96[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[775:768] <= 'd0;
end

wire  [39:0]  kernel_img_mul_97[0:24];
assign kernel_img_mul_97[0] = buffer_data_4[767:760] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_97[1] = buffer_data_4[775:768] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_97[2] = buffer_data_4[783:776] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_97[3] = buffer_data_4[791:784] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_97[4] = buffer_data_4[799:792] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_97[5] = buffer_data_3[767:760] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_97[6] = buffer_data_3[775:768] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_97[7] = buffer_data_3[783:776] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_97[8] = buffer_data_3[791:784] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_97[9] = buffer_data_3[799:792] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_97[10] = buffer_data_2[767:760] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_97[11] = buffer_data_2[775:768] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_97[12] = buffer_data_2[783:776] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_97[13] = buffer_data_2[791:784] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_97[14] = buffer_data_2[799:792] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_97[15] = buffer_data_1[767:760] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_97[16] = buffer_data_1[775:768] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_97[17] = buffer_data_1[783:776] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_97[18] = buffer_data_1[791:784] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_97[19] = buffer_data_1[799:792] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_97[20] = buffer_data_0[767:760] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_97[21] = buffer_data_0[775:768] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_97[22] = buffer_data_0[783:776] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_97[23] = buffer_data_0[791:784] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_97[24] = buffer_data_0[799:792] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_97 = kernel_img_mul_97[0] + kernel_img_mul_97[1] + kernel_img_mul_97[2] + 
                kernel_img_mul_97[3] + kernel_img_mul_97[4] + kernel_img_mul_97[5] + 
                kernel_img_mul_97[6] + kernel_img_mul_97[7] + kernel_img_mul_97[8] + 
                kernel_img_mul_97[9] + kernel_img_mul_97[10] + kernel_img_mul_97[11] + 
                kernel_img_mul_97[12] + kernel_img_mul_97[13] + kernel_img_mul_97[14] + 
                kernel_img_mul_97[15] + kernel_img_mul_97[16] + kernel_img_mul_97[17] + 
                kernel_img_mul_97[18] + kernel_img_mul_97[19] + kernel_img_mul_97[20] + 
                kernel_img_mul_97[21] + kernel_img_mul_97[22] + kernel_img_mul_97[23] + 
                kernel_img_mul_97[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[783:776] <= 'd0;
  else if (current_state==ST_START)
    blur_din[783:776] <= kernel_img_sum_97[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[783:776] <= 'd0;
end

wire  [39:0]  kernel_img_mul_98[0:24];
assign kernel_img_mul_98[0] = buffer_data_4[775:768] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_98[1] = buffer_data_4[783:776] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_98[2] = buffer_data_4[791:784] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_98[3] = buffer_data_4[799:792] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_98[4] = buffer_data_4[807:800] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_98[5] = buffer_data_3[775:768] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_98[6] = buffer_data_3[783:776] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_98[7] = buffer_data_3[791:784] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_98[8] = buffer_data_3[799:792] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_98[9] = buffer_data_3[807:800] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_98[10] = buffer_data_2[775:768] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_98[11] = buffer_data_2[783:776] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_98[12] = buffer_data_2[791:784] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_98[13] = buffer_data_2[799:792] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_98[14] = buffer_data_2[807:800] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_98[15] = buffer_data_1[775:768] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_98[16] = buffer_data_1[783:776] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_98[17] = buffer_data_1[791:784] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_98[18] = buffer_data_1[799:792] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_98[19] = buffer_data_1[807:800] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_98[20] = buffer_data_0[775:768] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_98[21] = buffer_data_0[783:776] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_98[22] = buffer_data_0[791:784] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_98[23] = buffer_data_0[799:792] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_98[24] = buffer_data_0[807:800] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_98 = kernel_img_mul_98[0] + kernel_img_mul_98[1] + kernel_img_mul_98[2] + 
                kernel_img_mul_98[3] + kernel_img_mul_98[4] + kernel_img_mul_98[5] + 
                kernel_img_mul_98[6] + kernel_img_mul_98[7] + kernel_img_mul_98[8] + 
                kernel_img_mul_98[9] + kernel_img_mul_98[10] + kernel_img_mul_98[11] + 
                kernel_img_mul_98[12] + kernel_img_mul_98[13] + kernel_img_mul_98[14] + 
                kernel_img_mul_98[15] + kernel_img_mul_98[16] + kernel_img_mul_98[17] + 
                kernel_img_mul_98[18] + kernel_img_mul_98[19] + kernel_img_mul_98[20] + 
                kernel_img_mul_98[21] + kernel_img_mul_98[22] + kernel_img_mul_98[23] + 
                kernel_img_mul_98[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[791:784] <= 'd0;
  else if (current_state==ST_START)
    blur_din[791:784] <= kernel_img_sum_98[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[791:784] <= 'd0;
end

wire  [39:0]  kernel_img_mul_99[0:24];
assign kernel_img_mul_99[0] = buffer_data_4[783:776] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_99[1] = buffer_data_4[791:784] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_99[2] = buffer_data_4[799:792] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_99[3] = buffer_data_4[807:800] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_99[4] = buffer_data_4[815:808] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_99[5] = buffer_data_3[783:776] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_99[6] = buffer_data_3[791:784] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_99[7] = buffer_data_3[799:792] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_99[8] = buffer_data_3[807:800] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_99[9] = buffer_data_3[815:808] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_99[10] = buffer_data_2[783:776] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_99[11] = buffer_data_2[791:784] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_99[12] = buffer_data_2[799:792] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_99[13] = buffer_data_2[807:800] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_99[14] = buffer_data_2[815:808] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_99[15] = buffer_data_1[783:776] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_99[16] = buffer_data_1[791:784] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_99[17] = buffer_data_1[799:792] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_99[18] = buffer_data_1[807:800] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_99[19] = buffer_data_1[815:808] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_99[20] = buffer_data_0[783:776] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_99[21] = buffer_data_0[791:784] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_99[22] = buffer_data_0[799:792] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_99[23] = buffer_data_0[807:800] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_99[24] = buffer_data_0[815:808] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_99 = kernel_img_mul_99[0] + kernel_img_mul_99[1] + kernel_img_mul_99[2] + 
                kernel_img_mul_99[3] + kernel_img_mul_99[4] + kernel_img_mul_99[5] + 
                kernel_img_mul_99[6] + kernel_img_mul_99[7] + kernel_img_mul_99[8] + 
                kernel_img_mul_99[9] + kernel_img_mul_99[10] + kernel_img_mul_99[11] + 
                kernel_img_mul_99[12] + kernel_img_mul_99[13] + kernel_img_mul_99[14] + 
                kernel_img_mul_99[15] + kernel_img_mul_99[16] + kernel_img_mul_99[17] + 
                kernel_img_mul_99[18] + kernel_img_mul_99[19] + kernel_img_mul_99[20] + 
                kernel_img_mul_99[21] + kernel_img_mul_99[22] + kernel_img_mul_99[23] + 
                kernel_img_mul_99[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[799:792] <= 'd0;
  else if (current_state==ST_START)
    blur_din[799:792] <= kernel_img_sum_99[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[799:792] <= 'd0;
end

wire  [39:0]  kernel_img_mul_100[0:24];
assign kernel_img_mul_100[0] = buffer_data_4[791:784] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_100[1] = buffer_data_4[799:792] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_100[2] = buffer_data_4[807:800] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_100[3] = buffer_data_4[815:808] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_100[4] = buffer_data_4[823:816] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_100[5] = buffer_data_3[791:784] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_100[6] = buffer_data_3[799:792] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_100[7] = buffer_data_3[807:800] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_100[8] = buffer_data_3[815:808] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_100[9] = buffer_data_3[823:816] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_100[10] = buffer_data_2[791:784] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_100[11] = buffer_data_2[799:792] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_100[12] = buffer_data_2[807:800] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_100[13] = buffer_data_2[815:808] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_100[14] = buffer_data_2[823:816] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_100[15] = buffer_data_1[791:784] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_100[16] = buffer_data_1[799:792] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_100[17] = buffer_data_1[807:800] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_100[18] = buffer_data_1[815:808] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_100[19] = buffer_data_1[823:816] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_100[20] = buffer_data_0[791:784] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_100[21] = buffer_data_0[799:792] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_100[22] = buffer_data_0[807:800] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_100[23] = buffer_data_0[815:808] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_100[24] = buffer_data_0[823:816] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_100 = kernel_img_mul_100[0] + kernel_img_mul_100[1] + kernel_img_mul_100[2] + 
                kernel_img_mul_100[3] + kernel_img_mul_100[4] + kernel_img_mul_100[5] + 
                kernel_img_mul_100[6] + kernel_img_mul_100[7] + kernel_img_mul_100[8] + 
                kernel_img_mul_100[9] + kernel_img_mul_100[10] + kernel_img_mul_100[11] + 
                kernel_img_mul_100[12] + kernel_img_mul_100[13] + kernel_img_mul_100[14] + 
                kernel_img_mul_100[15] + kernel_img_mul_100[16] + kernel_img_mul_100[17] + 
                kernel_img_mul_100[18] + kernel_img_mul_100[19] + kernel_img_mul_100[20] + 
                kernel_img_mul_100[21] + kernel_img_mul_100[22] + kernel_img_mul_100[23] + 
                kernel_img_mul_100[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[807:800] <= 'd0;
  else if (current_state==ST_START)
    blur_din[807:800] <= kernel_img_sum_100[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[807:800] <= 'd0;
end

wire  [39:0]  kernel_img_mul_101[0:24];
assign kernel_img_mul_101[0] = buffer_data_4[799:792] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_101[1] = buffer_data_4[807:800] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_101[2] = buffer_data_4[815:808] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_101[3] = buffer_data_4[823:816] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_101[4] = buffer_data_4[831:824] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_101[5] = buffer_data_3[799:792] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_101[6] = buffer_data_3[807:800] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_101[7] = buffer_data_3[815:808] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_101[8] = buffer_data_3[823:816] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_101[9] = buffer_data_3[831:824] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_101[10] = buffer_data_2[799:792] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_101[11] = buffer_data_2[807:800] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_101[12] = buffer_data_2[815:808] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_101[13] = buffer_data_2[823:816] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_101[14] = buffer_data_2[831:824] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_101[15] = buffer_data_1[799:792] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_101[16] = buffer_data_1[807:800] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_101[17] = buffer_data_1[815:808] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_101[18] = buffer_data_1[823:816] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_101[19] = buffer_data_1[831:824] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_101[20] = buffer_data_0[799:792] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_101[21] = buffer_data_0[807:800] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_101[22] = buffer_data_0[815:808] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_101[23] = buffer_data_0[823:816] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_101[24] = buffer_data_0[831:824] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_101 = kernel_img_mul_101[0] + kernel_img_mul_101[1] + kernel_img_mul_101[2] + 
                kernel_img_mul_101[3] + kernel_img_mul_101[4] + kernel_img_mul_101[5] + 
                kernel_img_mul_101[6] + kernel_img_mul_101[7] + kernel_img_mul_101[8] + 
                kernel_img_mul_101[9] + kernel_img_mul_101[10] + kernel_img_mul_101[11] + 
                kernel_img_mul_101[12] + kernel_img_mul_101[13] + kernel_img_mul_101[14] + 
                kernel_img_mul_101[15] + kernel_img_mul_101[16] + kernel_img_mul_101[17] + 
                kernel_img_mul_101[18] + kernel_img_mul_101[19] + kernel_img_mul_101[20] + 
                kernel_img_mul_101[21] + kernel_img_mul_101[22] + kernel_img_mul_101[23] + 
                kernel_img_mul_101[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[815:808] <= 'd0;
  else if (current_state==ST_START)
    blur_din[815:808] <= kernel_img_sum_101[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[815:808] <= 'd0;
end

wire  [39:0]  kernel_img_mul_102[0:24];
assign kernel_img_mul_102[0] = buffer_data_4[807:800] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_102[1] = buffer_data_4[815:808] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_102[2] = buffer_data_4[823:816] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_102[3] = buffer_data_4[831:824] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_102[4] = buffer_data_4[839:832] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_102[5] = buffer_data_3[807:800] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_102[6] = buffer_data_3[815:808] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_102[7] = buffer_data_3[823:816] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_102[8] = buffer_data_3[831:824] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_102[9] = buffer_data_3[839:832] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_102[10] = buffer_data_2[807:800] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_102[11] = buffer_data_2[815:808] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_102[12] = buffer_data_2[823:816] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_102[13] = buffer_data_2[831:824] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_102[14] = buffer_data_2[839:832] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_102[15] = buffer_data_1[807:800] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_102[16] = buffer_data_1[815:808] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_102[17] = buffer_data_1[823:816] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_102[18] = buffer_data_1[831:824] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_102[19] = buffer_data_1[839:832] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_102[20] = buffer_data_0[807:800] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_102[21] = buffer_data_0[815:808] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_102[22] = buffer_data_0[823:816] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_102[23] = buffer_data_0[831:824] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_102[24] = buffer_data_0[839:832] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_102 = kernel_img_mul_102[0] + kernel_img_mul_102[1] + kernel_img_mul_102[2] + 
                kernel_img_mul_102[3] + kernel_img_mul_102[4] + kernel_img_mul_102[5] + 
                kernel_img_mul_102[6] + kernel_img_mul_102[7] + kernel_img_mul_102[8] + 
                kernel_img_mul_102[9] + kernel_img_mul_102[10] + kernel_img_mul_102[11] + 
                kernel_img_mul_102[12] + kernel_img_mul_102[13] + kernel_img_mul_102[14] + 
                kernel_img_mul_102[15] + kernel_img_mul_102[16] + kernel_img_mul_102[17] + 
                kernel_img_mul_102[18] + kernel_img_mul_102[19] + kernel_img_mul_102[20] + 
                kernel_img_mul_102[21] + kernel_img_mul_102[22] + kernel_img_mul_102[23] + 
                kernel_img_mul_102[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[823:816] <= 'd0;
  else if (current_state==ST_START)
    blur_din[823:816] <= kernel_img_sum_102[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[823:816] <= 'd0;
end

wire  [39:0]  kernel_img_mul_103[0:24];
assign kernel_img_mul_103[0] = buffer_data_4[815:808] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_103[1] = buffer_data_4[823:816] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_103[2] = buffer_data_4[831:824] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_103[3] = buffer_data_4[839:832] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_103[4] = buffer_data_4[847:840] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_103[5] = buffer_data_3[815:808] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_103[6] = buffer_data_3[823:816] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_103[7] = buffer_data_3[831:824] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_103[8] = buffer_data_3[839:832] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_103[9] = buffer_data_3[847:840] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_103[10] = buffer_data_2[815:808] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_103[11] = buffer_data_2[823:816] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_103[12] = buffer_data_2[831:824] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_103[13] = buffer_data_2[839:832] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_103[14] = buffer_data_2[847:840] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_103[15] = buffer_data_1[815:808] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_103[16] = buffer_data_1[823:816] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_103[17] = buffer_data_1[831:824] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_103[18] = buffer_data_1[839:832] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_103[19] = buffer_data_1[847:840] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_103[20] = buffer_data_0[815:808] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_103[21] = buffer_data_0[823:816] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_103[22] = buffer_data_0[831:824] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_103[23] = buffer_data_0[839:832] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_103[24] = buffer_data_0[847:840] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_103 = kernel_img_mul_103[0] + kernel_img_mul_103[1] + kernel_img_mul_103[2] + 
                kernel_img_mul_103[3] + kernel_img_mul_103[4] + kernel_img_mul_103[5] + 
                kernel_img_mul_103[6] + kernel_img_mul_103[7] + kernel_img_mul_103[8] + 
                kernel_img_mul_103[9] + kernel_img_mul_103[10] + kernel_img_mul_103[11] + 
                kernel_img_mul_103[12] + kernel_img_mul_103[13] + kernel_img_mul_103[14] + 
                kernel_img_mul_103[15] + kernel_img_mul_103[16] + kernel_img_mul_103[17] + 
                kernel_img_mul_103[18] + kernel_img_mul_103[19] + kernel_img_mul_103[20] + 
                kernel_img_mul_103[21] + kernel_img_mul_103[22] + kernel_img_mul_103[23] + 
                kernel_img_mul_103[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[831:824] <= 'd0;
  else if (current_state==ST_START)
    blur_din[831:824] <= kernel_img_sum_103[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[831:824] <= 'd0;
end

wire  [39:0]  kernel_img_mul_104[0:24];
assign kernel_img_mul_104[0] = buffer_data_4[823:816] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_104[1] = buffer_data_4[831:824] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_104[2] = buffer_data_4[839:832] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_104[3] = buffer_data_4[847:840] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_104[4] = buffer_data_4[855:848] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_104[5] = buffer_data_3[823:816] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_104[6] = buffer_data_3[831:824] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_104[7] = buffer_data_3[839:832] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_104[8] = buffer_data_3[847:840] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_104[9] = buffer_data_3[855:848] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_104[10] = buffer_data_2[823:816] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_104[11] = buffer_data_2[831:824] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_104[12] = buffer_data_2[839:832] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_104[13] = buffer_data_2[847:840] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_104[14] = buffer_data_2[855:848] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_104[15] = buffer_data_1[823:816] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_104[16] = buffer_data_1[831:824] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_104[17] = buffer_data_1[839:832] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_104[18] = buffer_data_1[847:840] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_104[19] = buffer_data_1[855:848] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_104[20] = buffer_data_0[823:816] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_104[21] = buffer_data_0[831:824] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_104[22] = buffer_data_0[839:832] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_104[23] = buffer_data_0[847:840] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_104[24] = buffer_data_0[855:848] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_104 = kernel_img_mul_104[0] + kernel_img_mul_104[1] + kernel_img_mul_104[2] + 
                kernel_img_mul_104[3] + kernel_img_mul_104[4] + kernel_img_mul_104[5] + 
                kernel_img_mul_104[6] + kernel_img_mul_104[7] + kernel_img_mul_104[8] + 
                kernel_img_mul_104[9] + kernel_img_mul_104[10] + kernel_img_mul_104[11] + 
                kernel_img_mul_104[12] + kernel_img_mul_104[13] + kernel_img_mul_104[14] + 
                kernel_img_mul_104[15] + kernel_img_mul_104[16] + kernel_img_mul_104[17] + 
                kernel_img_mul_104[18] + kernel_img_mul_104[19] + kernel_img_mul_104[20] + 
                kernel_img_mul_104[21] + kernel_img_mul_104[22] + kernel_img_mul_104[23] + 
                kernel_img_mul_104[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[839:832] <= 'd0;
  else if (current_state==ST_START)
    blur_din[839:832] <= kernel_img_sum_104[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[839:832] <= 'd0;
end

wire  [39:0]  kernel_img_mul_105[0:24];
assign kernel_img_mul_105[0] = buffer_data_4[831:824] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_105[1] = buffer_data_4[839:832] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_105[2] = buffer_data_4[847:840] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_105[3] = buffer_data_4[855:848] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_105[4] = buffer_data_4[863:856] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_105[5] = buffer_data_3[831:824] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_105[6] = buffer_data_3[839:832] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_105[7] = buffer_data_3[847:840] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_105[8] = buffer_data_3[855:848] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_105[9] = buffer_data_3[863:856] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_105[10] = buffer_data_2[831:824] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_105[11] = buffer_data_2[839:832] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_105[12] = buffer_data_2[847:840] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_105[13] = buffer_data_2[855:848] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_105[14] = buffer_data_2[863:856] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_105[15] = buffer_data_1[831:824] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_105[16] = buffer_data_1[839:832] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_105[17] = buffer_data_1[847:840] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_105[18] = buffer_data_1[855:848] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_105[19] = buffer_data_1[863:856] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_105[20] = buffer_data_0[831:824] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_105[21] = buffer_data_0[839:832] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_105[22] = buffer_data_0[847:840] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_105[23] = buffer_data_0[855:848] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_105[24] = buffer_data_0[863:856] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_105 = kernel_img_mul_105[0] + kernel_img_mul_105[1] + kernel_img_mul_105[2] + 
                kernel_img_mul_105[3] + kernel_img_mul_105[4] + kernel_img_mul_105[5] + 
                kernel_img_mul_105[6] + kernel_img_mul_105[7] + kernel_img_mul_105[8] + 
                kernel_img_mul_105[9] + kernel_img_mul_105[10] + kernel_img_mul_105[11] + 
                kernel_img_mul_105[12] + kernel_img_mul_105[13] + kernel_img_mul_105[14] + 
                kernel_img_mul_105[15] + kernel_img_mul_105[16] + kernel_img_mul_105[17] + 
                kernel_img_mul_105[18] + kernel_img_mul_105[19] + kernel_img_mul_105[20] + 
                kernel_img_mul_105[21] + kernel_img_mul_105[22] + kernel_img_mul_105[23] + 
                kernel_img_mul_105[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[847:840] <= 'd0;
  else if (current_state==ST_START)
    blur_din[847:840] <= kernel_img_sum_105[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[847:840] <= 'd0;
end

wire  [39:0]  kernel_img_mul_106[0:24];
assign kernel_img_mul_106[0] = buffer_data_4[839:832] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_106[1] = buffer_data_4[847:840] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_106[2] = buffer_data_4[855:848] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_106[3] = buffer_data_4[863:856] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_106[4] = buffer_data_4[871:864] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_106[5] = buffer_data_3[839:832] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_106[6] = buffer_data_3[847:840] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_106[7] = buffer_data_3[855:848] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_106[8] = buffer_data_3[863:856] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_106[9] = buffer_data_3[871:864] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_106[10] = buffer_data_2[839:832] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_106[11] = buffer_data_2[847:840] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_106[12] = buffer_data_2[855:848] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_106[13] = buffer_data_2[863:856] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_106[14] = buffer_data_2[871:864] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_106[15] = buffer_data_1[839:832] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_106[16] = buffer_data_1[847:840] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_106[17] = buffer_data_1[855:848] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_106[18] = buffer_data_1[863:856] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_106[19] = buffer_data_1[871:864] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_106[20] = buffer_data_0[839:832] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_106[21] = buffer_data_0[847:840] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_106[22] = buffer_data_0[855:848] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_106[23] = buffer_data_0[863:856] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_106[24] = buffer_data_0[871:864] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_106 = kernel_img_mul_106[0] + kernel_img_mul_106[1] + kernel_img_mul_106[2] + 
                kernel_img_mul_106[3] + kernel_img_mul_106[4] + kernel_img_mul_106[5] + 
                kernel_img_mul_106[6] + kernel_img_mul_106[7] + kernel_img_mul_106[8] + 
                kernel_img_mul_106[9] + kernel_img_mul_106[10] + kernel_img_mul_106[11] + 
                kernel_img_mul_106[12] + kernel_img_mul_106[13] + kernel_img_mul_106[14] + 
                kernel_img_mul_106[15] + kernel_img_mul_106[16] + kernel_img_mul_106[17] + 
                kernel_img_mul_106[18] + kernel_img_mul_106[19] + kernel_img_mul_106[20] + 
                kernel_img_mul_106[21] + kernel_img_mul_106[22] + kernel_img_mul_106[23] + 
                kernel_img_mul_106[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[855:848] <= 'd0;
  else if (current_state==ST_START)
    blur_din[855:848] <= kernel_img_sum_106[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[855:848] <= 'd0;
end

wire  [39:0]  kernel_img_mul_107[0:24];
assign kernel_img_mul_107[0] = buffer_data_4[847:840] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_107[1] = buffer_data_4[855:848] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_107[2] = buffer_data_4[863:856] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_107[3] = buffer_data_4[871:864] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_107[4] = buffer_data_4[879:872] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_107[5] = buffer_data_3[847:840] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_107[6] = buffer_data_3[855:848] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_107[7] = buffer_data_3[863:856] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_107[8] = buffer_data_3[871:864] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_107[9] = buffer_data_3[879:872] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_107[10] = buffer_data_2[847:840] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_107[11] = buffer_data_2[855:848] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_107[12] = buffer_data_2[863:856] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_107[13] = buffer_data_2[871:864] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_107[14] = buffer_data_2[879:872] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_107[15] = buffer_data_1[847:840] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_107[16] = buffer_data_1[855:848] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_107[17] = buffer_data_1[863:856] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_107[18] = buffer_data_1[871:864] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_107[19] = buffer_data_1[879:872] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_107[20] = buffer_data_0[847:840] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_107[21] = buffer_data_0[855:848] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_107[22] = buffer_data_0[863:856] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_107[23] = buffer_data_0[871:864] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_107[24] = buffer_data_0[879:872] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_107 = kernel_img_mul_107[0] + kernel_img_mul_107[1] + kernel_img_mul_107[2] + 
                kernel_img_mul_107[3] + kernel_img_mul_107[4] + kernel_img_mul_107[5] + 
                kernel_img_mul_107[6] + kernel_img_mul_107[7] + kernel_img_mul_107[8] + 
                kernel_img_mul_107[9] + kernel_img_mul_107[10] + kernel_img_mul_107[11] + 
                kernel_img_mul_107[12] + kernel_img_mul_107[13] + kernel_img_mul_107[14] + 
                kernel_img_mul_107[15] + kernel_img_mul_107[16] + kernel_img_mul_107[17] + 
                kernel_img_mul_107[18] + kernel_img_mul_107[19] + kernel_img_mul_107[20] + 
                kernel_img_mul_107[21] + kernel_img_mul_107[22] + kernel_img_mul_107[23] + 
                kernel_img_mul_107[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[863:856] <= 'd0;
  else if (current_state==ST_START)
    blur_din[863:856] <= kernel_img_sum_107[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[863:856] <= 'd0;
end

wire  [39:0]  kernel_img_mul_108[0:24];
assign kernel_img_mul_108[0] = buffer_data_4[855:848] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_108[1] = buffer_data_4[863:856] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_108[2] = buffer_data_4[871:864] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_108[3] = buffer_data_4[879:872] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_108[4] = buffer_data_4[887:880] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_108[5] = buffer_data_3[855:848] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_108[6] = buffer_data_3[863:856] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_108[7] = buffer_data_3[871:864] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_108[8] = buffer_data_3[879:872] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_108[9] = buffer_data_3[887:880] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_108[10] = buffer_data_2[855:848] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_108[11] = buffer_data_2[863:856] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_108[12] = buffer_data_2[871:864] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_108[13] = buffer_data_2[879:872] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_108[14] = buffer_data_2[887:880] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_108[15] = buffer_data_1[855:848] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_108[16] = buffer_data_1[863:856] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_108[17] = buffer_data_1[871:864] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_108[18] = buffer_data_1[879:872] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_108[19] = buffer_data_1[887:880] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_108[20] = buffer_data_0[855:848] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_108[21] = buffer_data_0[863:856] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_108[22] = buffer_data_0[871:864] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_108[23] = buffer_data_0[879:872] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_108[24] = buffer_data_0[887:880] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_108 = kernel_img_mul_108[0] + kernel_img_mul_108[1] + kernel_img_mul_108[2] + 
                kernel_img_mul_108[3] + kernel_img_mul_108[4] + kernel_img_mul_108[5] + 
                kernel_img_mul_108[6] + kernel_img_mul_108[7] + kernel_img_mul_108[8] + 
                kernel_img_mul_108[9] + kernel_img_mul_108[10] + kernel_img_mul_108[11] + 
                kernel_img_mul_108[12] + kernel_img_mul_108[13] + kernel_img_mul_108[14] + 
                kernel_img_mul_108[15] + kernel_img_mul_108[16] + kernel_img_mul_108[17] + 
                kernel_img_mul_108[18] + kernel_img_mul_108[19] + kernel_img_mul_108[20] + 
                kernel_img_mul_108[21] + kernel_img_mul_108[22] + kernel_img_mul_108[23] + 
                kernel_img_mul_108[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[871:864] <= 'd0;
  else if (current_state==ST_START)
    blur_din[871:864] <= kernel_img_sum_108[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[871:864] <= 'd0;
end

wire  [39:0]  kernel_img_mul_109[0:24];
assign kernel_img_mul_109[0] = buffer_data_4[863:856] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_109[1] = buffer_data_4[871:864] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_109[2] = buffer_data_4[879:872] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_109[3] = buffer_data_4[887:880] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_109[4] = buffer_data_4[895:888] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_109[5] = buffer_data_3[863:856] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_109[6] = buffer_data_3[871:864] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_109[7] = buffer_data_3[879:872] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_109[8] = buffer_data_3[887:880] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_109[9] = buffer_data_3[895:888] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_109[10] = buffer_data_2[863:856] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_109[11] = buffer_data_2[871:864] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_109[12] = buffer_data_2[879:872] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_109[13] = buffer_data_2[887:880] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_109[14] = buffer_data_2[895:888] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_109[15] = buffer_data_1[863:856] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_109[16] = buffer_data_1[871:864] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_109[17] = buffer_data_1[879:872] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_109[18] = buffer_data_1[887:880] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_109[19] = buffer_data_1[895:888] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_109[20] = buffer_data_0[863:856] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_109[21] = buffer_data_0[871:864] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_109[22] = buffer_data_0[879:872] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_109[23] = buffer_data_0[887:880] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_109[24] = buffer_data_0[895:888] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_109 = kernel_img_mul_109[0] + kernel_img_mul_109[1] + kernel_img_mul_109[2] + 
                kernel_img_mul_109[3] + kernel_img_mul_109[4] + kernel_img_mul_109[5] + 
                kernel_img_mul_109[6] + kernel_img_mul_109[7] + kernel_img_mul_109[8] + 
                kernel_img_mul_109[9] + kernel_img_mul_109[10] + kernel_img_mul_109[11] + 
                kernel_img_mul_109[12] + kernel_img_mul_109[13] + kernel_img_mul_109[14] + 
                kernel_img_mul_109[15] + kernel_img_mul_109[16] + kernel_img_mul_109[17] + 
                kernel_img_mul_109[18] + kernel_img_mul_109[19] + kernel_img_mul_109[20] + 
                kernel_img_mul_109[21] + kernel_img_mul_109[22] + kernel_img_mul_109[23] + 
                kernel_img_mul_109[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[879:872] <= 'd0;
  else if (current_state==ST_START)
    blur_din[879:872] <= kernel_img_sum_109[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[879:872] <= 'd0;
end

wire  [39:0]  kernel_img_mul_110[0:24];
assign kernel_img_mul_110[0] = buffer_data_4[871:864] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_110[1] = buffer_data_4[879:872] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_110[2] = buffer_data_4[887:880] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_110[3] = buffer_data_4[895:888] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_110[4] = buffer_data_4[903:896] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_110[5] = buffer_data_3[871:864] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_110[6] = buffer_data_3[879:872] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_110[7] = buffer_data_3[887:880] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_110[8] = buffer_data_3[895:888] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_110[9] = buffer_data_3[903:896] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_110[10] = buffer_data_2[871:864] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_110[11] = buffer_data_2[879:872] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_110[12] = buffer_data_2[887:880] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_110[13] = buffer_data_2[895:888] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_110[14] = buffer_data_2[903:896] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_110[15] = buffer_data_1[871:864] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_110[16] = buffer_data_1[879:872] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_110[17] = buffer_data_1[887:880] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_110[18] = buffer_data_1[895:888] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_110[19] = buffer_data_1[903:896] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_110[20] = buffer_data_0[871:864] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_110[21] = buffer_data_0[879:872] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_110[22] = buffer_data_0[887:880] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_110[23] = buffer_data_0[895:888] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_110[24] = buffer_data_0[903:896] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_110 = kernel_img_mul_110[0] + kernel_img_mul_110[1] + kernel_img_mul_110[2] + 
                kernel_img_mul_110[3] + kernel_img_mul_110[4] + kernel_img_mul_110[5] + 
                kernel_img_mul_110[6] + kernel_img_mul_110[7] + kernel_img_mul_110[8] + 
                kernel_img_mul_110[9] + kernel_img_mul_110[10] + kernel_img_mul_110[11] + 
                kernel_img_mul_110[12] + kernel_img_mul_110[13] + kernel_img_mul_110[14] + 
                kernel_img_mul_110[15] + kernel_img_mul_110[16] + kernel_img_mul_110[17] + 
                kernel_img_mul_110[18] + kernel_img_mul_110[19] + kernel_img_mul_110[20] + 
                kernel_img_mul_110[21] + kernel_img_mul_110[22] + kernel_img_mul_110[23] + 
                kernel_img_mul_110[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[887:880] <= 'd0;
  else if (current_state==ST_START)
    blur_din[887:880] <= kernel_img_sum_110[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[887:880] <= 'd0;
end

wire  [39:0]  kernel_img_mul_111[0:24];
assign kernel_img_mul_111[0] = buffer_data_4[879:872] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_111[1] = buffer_data_4[887:880] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_111[2] = buffer_data_4[895:888] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_111[3] = buffer_data_4[903:896] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_111[4] = buffer_data_4[911:904] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_111[5] = buffer_data_3[879:872] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_111[6] = buffer_data_3[887:880] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_111[7] = buffer_data_3[895:888] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_111[8] = buffer_data_3[903:896] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_111[9] = buffer_data_3[911:904] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_111[10] = buffer_data_2[879:872] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_111[11] = buffer_data_2[887:880] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_111[12] = buffer_data_2[895:888] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_111[13] = buffer_data_2[903:896] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_111[14] = buffer_data_2[911:904] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_111[15] = buffer_data_1[879:872] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_111[16] = buffer_data_1[887:880] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_111[17] = buffer_data_1[895:888] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_111[18] = buffer_data_1[903:896] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_111[19] = buffer_data_1[911:904] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_111[20] = buffer_data_0[879:872] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_111[21] = buffer_data_0[887:880] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_111[22] = buffer_data_0[895:888] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_111[23] = buffer_data_0[903:896] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_111[24] = buffer_data_0[911:904] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_111 = kernel_img_mul_111[0] + kernel_img_mul_111[1] + kernel_img_mul_111[2] + 
                kernel_img_mul_111[3] + kernel_img_mul_111[4] + kernel_img_mul_111[5] + 
                kernel_img_mul_111[6] + kernel_img_mul_111[7] + kernel_img_mul_111[8] + 
                kernel_img_mul_111[9] + kernel_img_mul_111[10] + kernel_img_mul_111[11] + 
                kernel_img_mul_111[12] + kernel_img_mul_111[13] + kernel_img_mul_111[14] + 
                kernel_img_mul_111[15] + kernel_img_mul_111[16] + kernel_img_mul_111[17] + 
                kernel_img_mul_111[18] + kernel_img_mul_111[19] + kernel_img_mul_111[20] + 
                kernel_img_mul_111[21] + kernel_img_mul_111[22] + kernel_img_mul_111[23] + 
                kernel_img_mul_111[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[895:888] <= 'd0;
  else if (current_state==ST_START)
    blur_din[895:888] <= kernel_img_sum_111[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[895:888] <= 'd0;
end

wire  [39:0]  kernel_img_mul_112[0:24];
assign kernel_img_mul_112[0] = buffer_data_4[887:880] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_112[1] = buffer_data_4[895:888] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_112[2] = buffer_data_4[903:896] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_112[3] = buffer_data_4[911:904] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_112[4] = buffer_data_4[919:912] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_112[5] = buffer_data_3[887:880] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_112[6] = buffer_data_3[895:888] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_112[7] = buffer_data_3[903:896] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_112[8] = buffer_data_3[911:904] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_112[9] = buffer_data_3[919:912] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_112[10] = buffer_data_2[887:880] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_112[11] = buffer_data_2[895:888] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_112[12] = buffer_data_2[903:896] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_112[13] = buffer_data_2[911:904] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_112[14] = buffer_data_2[919:912] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_112[15] = buffer_data_1[887:880] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_112[16] = buffer_data_1[895:888] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_112[17] = buffer_data_1[903:896] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_112[18] = buffer_data_1[911:904] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_112[19] = buffer_data_1[919:912] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_112[20] = buffer_data_0[887:880] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_112[21] = buffer_data_0[895:888] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_112[22] = buffer_data_0[903:896] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_112[23] = buffer_data_0[911:904] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_112[24] = buffer_data_0[919:912] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_112 = kernel_img_mul_112[0] + kernel_img_mul_112[1] + kernel_img_mul_112[2] + 
                kernel_img_mul_112[3] + kernel_img_mul_112[4] + kernel_img_mul_112[5] + 
                kernel_img_mul_112[6] + kernel_img_mul_112[7] + kernel_img_mul_112[8] + 
                kernel_img_mul_112[9] + kernel_img_mul_112[10] + kernel_img_mul_112[11] + 
                kernel_img_mul_112[12] + kernel_img_mul_112[13] + kernel_img_mul_112[14] + 
                kernel_img_mul_112[15] + kernel_img_mul_112[16] + kernel_img_mul_112[17] + 
                kernel_img_mul_112[18] + kernel_img_mul_112[19] + kernel_img_mul_112[20] + 
                kernel_img_mul_112[21] + kernel_img_mul_112[22] + kernel_img_mul_112[23] + 
                kernel_img_mul_112[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[903:896] <= 'd0;
  else if (current_state==ST_START)
    blur_din[903:896] <= kernel_img_sum_112[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[903:896] <= 'd0;
end

wire  [39:0]  kernel_img_mul_113[0:24];
assign kernel_img_mul_113[0] = buffer_data_4[895:888] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_113[1] = buffer_data_4[903:896] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_113[2] = buffer_data_4[911:904] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_113[3] = buffer_data_4[919:912] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_113[4] = buffer_data_4[927:920] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_113[5] = buffer_data_3[895:888] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_113[6] = buffer_data_3[903:896] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_113[7] = buffer_data_3[911:904] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_113[8] = buffer_data_3[919:912] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_113[9] = buffer_data_3[927:920] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_113[10] = buffer_data_2[895:888] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_113[11] = buffer_data_2[903:896] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_113[12] = buffer_data_2[911:904] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_113[13] = buffer_data_2[919:912] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_113[14] = buffer_data_2[927:920] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_113[15] = buffer_data_1[895:888] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_113[16] = buffer_data_1[903:896] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_113[17] = buffer_data_1[911:904] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_113[18] = buffer_data_1[919:912] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_113[19] = buffer_data_1[927:920] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_113[20] = buffer_data_0[895:888] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_113[21] = buffer_data_0[903:896] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_113[22] = buffer_data_0[911:904] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_113[23] = buffer_data_0[919:912] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_113[24] = buffer_data_0[927:920] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_113 = kernel_img_mul_113[0] + kernel_img_mul_113[1] + kernel_img_mul_113[2] + 
                kernel_img_mul_113[3] + kernel_img_mul_113[4] + kernel_img_mul_113[5] + 
                kernel_img_mul_113[6] + kernel_img_mul_113[7] + kernel_img_mul_113[8] + 
                kernel_img_mul_113[9] + kernel_img_mul_113[10] + kernel_img_mul_113[11] + 
                kernel_img_mul_113[12] + kernel_img_mul_113[13] + kernel_img_mul_113[14] + 
                kernel_img_mul_113[15] + kernel_img_mul_113[16] + kernel_img_mul_113[17] + 
                kernel_img_mul_113[18] + kernel_img_mul_113[19] + kernel_img_mul_113[20] + 
                kernel_img_mul_113[21] + kernel_img_mul_113[22] + kernel_img_mul_113[23] + 
                kernel_img_mul_113[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[911:904] <= 'd0;
  else if (current_state==ST_START)
    blur_din[911:904] <= kernel_img_sum_113[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[911:904] <= 'd0;
end

wire  [39:0]  kernel_img_mul_114[0:24];
assign kernel_img_mul_114[0] = buffer_data_4[903:896] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_114[1] = buffer_data_4[911:904] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_114[2] = buffer_data_4[919:912] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_114[3] = buffer_data_4[927:920] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_114[4] = buffer_data_4[935:928] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_114[5] = buffer_data_3[903:896] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_114[6] = buffer_data_3[911:904] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_114[7] = buffer_data_3[919:912] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_114[8] = buffer_data_3[927:920] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_114[9] = buffer_data_3[935:928] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_114[10] = buffer_data_2[903:896] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_114[11] = buffer_data_2[911:904] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_114[12] = buffer_data_2[919:912] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_114[13] = buffer_data_2[927:920] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_114[14] = buffer_data_2[935:928] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_114[15] = buffer_data_1[903:896] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_114[16] = buffer_data_1[911:904] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_114[17] = buffer_data_1[919:912] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_114[18] = buffer_data_1[927:920] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_114[19] = buffer_data_1[935:928] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_114[20] = buffer_data_0[903:896] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_114[21] = buffer_data_0[911:904] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_114[22] = buffer_data_0[919:912] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_114[23] = buffer_data_0[927:920] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_114[24] = buffer_data_0[935:928] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_114 = kernel_img_mul_114[0] + kernel_img_mul_114[1] + kernel_img_mul_114[2] + 
                kernel_img_mul_114[3] + kernel_img_mul_114[4] + kernel_img_mul_114[5] + 
                kernel_img_mul_114[6] + kernel_img_mul_114[7] + kernel_img_mul_114[8] + 
                kernel_img_mul_114[9] + kernel_img_mul_114[10] + kernel_img_mul_114[11] + 
                kernel_img_mul_114[12] + kernel_img_mul_114[13] + kernel_img_mul_114[14] + 
                kernel_img_mul_114[15] + kernel_img_mul_114[16] + kernel_img_mul_114[17] + 
                kernel_img_mul_114[18] + kernel_img_mul_114[19] + kernel_img_mul_114[20] + 
                kernel_img_mul_114[21] + kernel_img_mul_114[22] + kernel_img_mul_114[23] + 
                kernel_img_mul_114[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[919:912] <= 'd0;
  else if (current_state==ST_START)
    blur_din[919:912] <= kernel_img_sum_114[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[919:912] <= 'd0;
end

wire  [39:0]  kernel_img_mul_115[0:24];
assign kernel_img_mul_115[0] = buffer_data_4[911:904] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_115[1] = buffer_data_4[919:912] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_115[2] = buffer_data_4[927:920] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_115[3] = buffer_data_4[935:928] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_115[4] = buffer_data_4[943:936] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_115[5] = buffer_data_3[911:904] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_115[6] = buffer_data_3[919:912] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_115[7] = buffer_data_3[927:920] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_115[8] = buffer_data_3[935:928] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_115[9] = buffer_data_3[943:936] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_115[10] = buffer_data_2[911:904] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_115[11] = buffer_data_2[919:912] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_115[12] = buffer_data_2[927:920] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_115[13] = buffer_data_2[935:928] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_115[14] = buffer_data_2[943:936] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_115[15] = buffer_data_1[911:904] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_115[16] = buffer_data_1[919:912] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_115[17] = buffer_data_1[927:920] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_115[18] = buffer_data_1[935:928] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_115[19] = buffer_data_1[943:936] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_115[20] = buffer_data_0[911:904] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_115[21] = buffer_data_0[919:912] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_115[22] = buffer_data_0[927:920] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_115[23] = buffer_data_0[935:928] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_115[24] = buffer_data_0[943:936] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_115 = kernel_img_mul_115[0] + kernel_img_mul_115[1] + kernel_img_mul_115[2] + 
                kernel_img_mul_115[3] + kernel_img_mul_115[4] + kernel_img_mul_115[5] + 
                kernel_img_mul_115[6] + kernel_img_mul_115[7] + kernel_img_mul_115[8] + 
                kernel_img_mul_115[9] + kernel_img_mul_115[10] + kernel_img_mul_115[11] + 
                kernel_img_mul_115[12] + kernel_img_mul_115[13] + kernel_img_mul_115[14] + 
                kernel_img_mul_115[15] + kernel_img_mul_115[16] + kernel_img_mul_115[17] + 
                kernel_img_mul_115[18] + kernel_img_mul_115[19] + kernel_img_mul_115[20] + 
                kernel_img_mul_115[21] + kernel_img_mul_115[22] + kernel_img_mul_115[23] + 
                kernel_img_mul_115[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[927:920] <= 'd0;
  else if (current_state==ST_START)
    blur_din[927:920] <= kernel_img_sum_115[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[927:920] <= 'd0;
end

wire  [39:0]  kernel_img_mul_116[0:24];
assign kernel_img_mul_116[0] = buffer_data_4[919:912] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_116[1] = buffer_data_4[927:920] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_116[2] = buffer_data_4[935:928] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_116[3] = buffer_data_4[943:936] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_116[4] = buffer_data_4[951:944] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_116[5] = buffer_data_3[919:912] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_116[6] = buffer_data_3[927:920] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_116[7] = buffer_data_3[935:928] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_116[8] = buffer_data_3[943:936] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_116[9] = buffer_data_3[951:944] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_116[10] = buffer_data_2[919:912] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_116[11] = buffer_data_2[927:920] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_116[12] = buffer_data_2[935:928] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_116[13] = buffer_data_2[943:936] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_116[14] = buffer_data_2[951:944] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_116[15] = buffer_data_1[919:912] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_116[16] = buffer_data_1[927:920] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_116[17] = buffer_data_1[935:928] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_116[18] = buffer_data_1[943:936] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_116[19] = buffer_data_1[951:944] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_116[20] = buffer_data_0[919:912] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_116[21] = buffer_data_0[927:920] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_116[22] = buffer_data_0[935:928] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_116[23] = buffer_data_0[943:936] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_116[24] = buffer_data_0[951:944] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_116 = kernel_img_mul_116[0] + kernel_img_mul_116[1] + kernel_img_mul_116[2] + 
                kernel_img_mul_116[3] + kernel_img_mul_116[4] + kernel_img_mul_116[5] + 
                kernel_img_mul_116[6] + kernel_img_mul_116[7] + kernel_img_mul_116[8] + 
                kernel_img_mul_116[9] + kernel_img_mul_116[10] + kernel_img_mul_116[11] + 
                kernel_img_mul_116[12] + kernel_img_mul_116[13] + kernel_img_mul_116[14] + 
                kernel_img_mul_116[15] + kernel_img_mul_116[16] + kernel_img_mul_116[17] + 
                kernel_img_mul_116[18] + kernel_img_mul_116[19] + kernel_img_mul_116[20] + 
                kernel_img_mul_116[21] + kernel_img_mul_116[22] + kernel_img_mul_116[23] + 
                kernel_img_mul_116[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[935:928] <= 'd0;
  else if (current_state==ST_START)
    blur_din[935:928] <= kernel_img_sum_116[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[935:928] <= 'd0;
end

wire  [39:0]  kernel_img_mul_117[0:24];
assign kernel_img_mul_117[0] = buffer_data_4[927:920] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_117[1] = buffer_data_4[935:928] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_117[2] = buffer_data_4[943:936] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_117[3] = buffer_data_4[951:944] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_117[4] = buffer_data_4[959:952] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_117[5] = buffer_data_3[927:920] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_117[6] = buffer_data_3[935:928] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_117[7] = buffer_data_3[943:936] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_117[8] = buffer_data_3[951:944] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_117[9] = buffer_data_3[959:952] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_117[10] = buffer_data_2[927:920] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_117[11] = buffer_data_2[935:928] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_117[12] = buffer_data_2[943:936] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_117[13] = buffer_data_2[951:944] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_117[14] = buffer_data_2[959:952] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_117[15] = buffer_data_1[927:920] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_117[16] = buffer_data_1[935:928] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_117[17] = buffer_data_1[943:936] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_117[18] = buffer_data_1[951:944] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_117[19] = buffer_data_1[959:952] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_117[20] = buffer_data_0[927:920] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_117[21] = buffer_data_0[935:928] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_117[22] = buffer_data_0[943:936] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_117[23] = buffer_data_0[951:944] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_117[24] = buffer_data_0[959:952] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_117 = kernel_img_mul_117[0] + kernel_img_mul_117[1] + kernel_img_mul_117[2] + 
                kernel_img_mul_117[3] + kernel_img_mul_117[4] + kernel_img_mul_117[5] + 
                kernel_img_mul_117[6] + kernel_img_mul_117[7] + kernel_img_mul_117[8] + 
                kernel_img_mul_117[9] + kernel_img_mul_117[10] + kernel_img_mul_117[11] + 
                kernel_img_mul_117[12] + kernel_img_mul_117[13] + kernel_img_mul_117[14] + 
                kernel_img_mul_117[15] + kernel_img_mul_117[16] + kernel_img_mul_117[17] + 
                kernel_img_mul_117[18] + kernel_img_mul_117[19] + kernel_img_mul_117[20] + 
                kernel_img_mul_117[21] + kernel_img_mul_117[22] + kernel_img_mul_117[23] + 
                kernel_img_mul_117[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[943:936] <= 'd0;
  else if (current_state==ST_START)
    blur_din[943:936] <= kernel_img_sum_117[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[943:936] <= 'd0;
end

wire  [39:0]  kernel_img_mul_118[0:24];
assign kernel_img_mul_118[0] = buffer_data_4[935:928] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_118[1] = buffer_data_4[943:936] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_118[2] = buffer_data_4[951:944] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_118[3] = buffer_data_4[959:952] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_118[4] = buffer_data_4[967:960] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_118[5] = buffer_data_3[935:928] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_118[6] = buffer_data_3[943:936] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_118[7] = buffer_data_3[951:944] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_118[8] = buffer_data_3[959:952] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_118[9] = buffer_data_3[967:960] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_118[10] = buffer_data_2[935:928] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_118[11] = buffer_data_2[943:936] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_118[12] = buffer_data_2[951:944] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_118[13] = buffer_data_2[959:952] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_118[14] = buffer_data_2[967:960] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_118[15] = buffer_data_1[935:928] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_118[16] = buffer_data_1[943:936] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_118[17] = buffer_data_1[951:944] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_118[18] = buffer_data_1[959:952] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_118[19] = buffer_data_1[967:960] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_118[20] = buffer_data_0[935:928] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_118[21] = buffer_data_0[943:936] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_118[22] = buffer_data_0[951:944] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_118[23] = buffer_data_0[959:952] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_118[24] = buffer_data_0[967:960] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_118 = kernel_img_mul_118[0] + kernel_img_mul_118[1] + kernel_img_mul_118[2] + 
                kernel_img_mul_118[3] + kernel_img_mul_118[4] + kernel_img_mul_118[5] + 
                kernel_img_mul_118[6] + kernel_img_mul_118[7] + kernel_img_mul_118[8] + 
                kernel_img_mul_118[9] + kernel_img_mul_118[10] + kernel_img_mul_118[11] + 
                kernel_img_mul_118[12] + kernel_img_mul_118[13] + kernel_img_mul_118[14] + 
                kernel_img_mul_118[15] + kernel_img_mul_118[16] + kernel_img_mul_118[17] + 
                kernel_img_mul_118[18] + kernel_img_mul_118[19] + kernel_img_mul_118[20] + 
                kernel_img_mul_118[21] + kernel_img_mul_118[22] + kernel_img_mul_118[23] + 
                kernel_img_mul_118[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[951:944] <= 'd0;
  else if (current_state==ST_START)
    blur_din[951:944] <= kernel_img_sum_118[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[951:944] <= 'd0;
end

wire  [39:0]  kernel_img_mul_119[0:24];
assign kernel_img_mul_119[0] = buffer_data_4[943:936] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_119[1] = buffer_data_4[951:944] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_119[2] = buffer_data_4[959:952] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_119[3] = buffer_data_4[967:960] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_119[4] = buffer_data_4[975:968] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_119[5] = buffer_data_3[943:936] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_119[6] = buffer_data_3[951:944] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_119[7] = buffer_data_3[959:952] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_119[8] = buffer_data_3[967:960] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_119[9] = buffer_data_3[975:968] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_119[10] = buffer_data_2[943:936] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_119[11] = buffer_data_2[951:944] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_119[12] = buffer_data_2[959:952] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_119[13] = buffer_data_2[967:960] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_119[14] = buffer_data_2[975:968] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_119[15] = buffer_data_1[943:936] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_119[16] = buffer_data_1[951:944] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_119[17] = buffer_data_1[959:952] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_119[18] = buffer_data_1[967:960] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_119[19] = buffer_data_1[975:968] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_119[20] = buffer_data_0[943:936] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_119[21] = buffer_data_0[951:944] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_119[22] = buffer_data_0[959:952] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_119[23] = buffer_data_0[967:960] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_119[24] = buffer_data_0[975:968] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_119 = kernel_img_mul_119[0] + kernel_img_mul_119[1] + kernel_img_mul_119[2] + 
                kernel_img_mul_119[3] + kernel_img_mul_119[4] + kernel_img_mul_119[5] + 
                kernel_img_mul_119[6] + kernel_img_mul_119[7] + kernel_img_mul_119[8] + 
                kernel_img_mul_119[9] + kernel_img_mul_119[10] + kernel_img_mul_119[11] + 
                kernel_img_mul_119[12] + kernel_img_mul_119[13] + kernel_img_mul_119[14] + 
                kernel_img_mul_119[15] + kernel_img_mul_119[16] + kernel_img_mul_119[17] + 
                kernel_img_mul_119[18] + kernel_img_mul_119[19] + kernel_img_mul_119[20] + 
                kernel_img_mul_119[21] + kernel_img_mul_119[22] + kernel_img_mul_119[23] + 
                kernel_img_mul_119[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[959:952] <= 'd0;
  else if (current_state==ST_START)
    blur_din[959:952] <= kernel_img_sum_119[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[959:952] <= 'd0;
end

wire  [39:0]  kernel_img_mul_120[0:24];
assign kernel_img_mul_120[0] = buffer_data_4[951:944] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_120[1] = buffer_data_4[959:952] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_120[2] = buffer_data_4[967:960] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_120[3] = buffer_data_4[975:968] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_120[4] = buffer_data_4[983:976] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_120[5] = buffer_data_3[951:944] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_120[6] = buffer_data_3[959:952] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_120[7] = buffer_data_3[967:960] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_120[8] = buffer_data_3[975:968] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_120[9] = buffer_data_3[983:976] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_120[10] = buffer_data_2[951:944] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_120[11] = buffer_data_2[959:952] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_120[12] = buffer_data_2[967:960] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_120[13] = buffer_data_2[975:968] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_120[14] = buffer_data_2[983:976] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_120[15] = buffer_data_1[951:944] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_120[16] = buffer_data_1[959:952] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_120[17] = buffer_data_1[967:960] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_120[18] = buffer_data_1[975:968] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_120[19] = buffer_data_1[983:976] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_120[20] = buffer_data_0[951:944] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_120[21] = buffer_data_0[959:952] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_120[22] = buffer_data_0[967:960] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_120[23] = buffer_data_0[975:968] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_120[24] = buffer_data_0[983:976] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_120 = kernel_img_mul_120[0] + kernel_img_mul_120[1] + kernel_img_mul_120[2] + 
                kernel_img_mul_120[3] + kernel_img_mul_120[4] + kernel_img_mul_120[5] + 
                kernel_img_mul_120[6] + kernel_img_mul_120[7] + kernel_img_mul_120[8] + 
                kernel_img_mul_120[9] + kernel_img_mul_120[10] + kernel_img_mul_120[11] + 
                kernel_img_mul_120[12] + kernel_img_mul_120[13] + kernel_img_mul_120[14] + 
                kernel_img_mul_120[15] + kernel_img_mul_120[16] + kernel_img_mul_120[17] + 
                kernel_img_mul_120[18] + kernel_img_mul_120[19] + kernel_img_mul_120[20] + 
                kernel_img_mul_120[21] + kernel_img_mul_120[22] + kernel_img_mul_120[23] + 
                kernel_img_mul_120[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[967:960] <= 'd0;
  else if (current_state==ST_START)
    blur_din[967:960] <= kernel_img_sum_120[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[967:960] <= 'd0;
end

wire  [39:0]  kernel_img_mul_121[0:24];
assign kernel_img_mul_121[0] = buffer_data_4[959:952] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_121[1] = buffer_data_4[967:960] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_121[2] = buffer_data_4[975:968] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_121[3] = buffer_data_4[983:976] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_121[4] = buffer_data_4[991:984] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_121[5] = buffer_data_3[959:952] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_121[6] = buffer_data_3[967:960] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_121[7] = buffer_data_3[975:968] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_121[8] = buffer_data_3[983:976] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_121[9] = buffer_data_3[991:984] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_121[10] = buffer_data_2[959:952] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_121[11] = buffer_data_2[967:960] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_121[12] = buffer_data_2[975:968] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_121[13] = buffer_data_2[983:976] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_121[14] = buffer_data_2[991:984] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_121[15] = buffer_data_1[959:952] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_121[16] = buffer_data_1[967:960] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_121[17] = buffer_data_1[975:968] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_121[18] = buffer_data_1[983:976] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_121[19] = buffer_data_1[991:984] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_121[20] = buffer_data_0[959:952] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_121[21] = buffer_data_0[967:960] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_121[22] = buffer_data_0[975:968] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_121[23] = buffer_data_0[983:976] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_121[24] = buffer_data_0[991:984] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_121 = kernel_img_mul_121[0] + kernel_img_mul_121[1] + kernel_img_mul_121[2] + 
                kernel_img_mul_121[3] + kernel_img_mul_121[4] + kernel_img_mul_121[5] + 
                kernel_img_mul_121[6] + kernel_img_mul_121[7] + kernel_img_mul_121[8] + 
                kernel_img_mul_121[9] + kernel_img_mul_121[10] + kernel_img_mul_121[11] + 
                kernel_img_mul_121[12] + kernel_img_mul_121[13] + kernel_img_mul_121[14] + 
                kernel_img_mul_121[15] + kernel_img_mul_121[16] + kernel_img_mul_121[17] + 
                kernel_img_mul_121[18] + kernel_img_mul_121[19] + kernel_img_mul_121[20] + 
                kernel_img_mul_121[21] + kernel_img_mul_121[22] + kernel_img_mul_121[23] + 
                kernel_img_mul_121[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[975:968] <= 'd0;
  else if (current_state==ST_START)
    blur_din[975:968] <= kernel_img_sum_121[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[975:968] <= 'd0;
end

wire  [39:0]  kernel_img_mul_122[0:24];
assign kernel_img_mul_122[0] = buffer_data_4[967:960] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_122[1] = buffer_data_4[975:968] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_122[2] = buffer_data_4[983:976] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_122[3] = buffer_data_4[991:984] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_122[4] = buffer_data_4[999:992] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_122[5] = buffer_data_3[967:960] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_122[6] = buffer_data_3[975:968] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_122[7] = buffer_data_3[983:976] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_122[8] = buffer_data_3[991:984] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_122[9] = buffer_data_3[999:992] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_122[10] = buffer_data_2[967:960] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_122[11] = buffer_data_2[975:968] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_122[12] = buffer_data_2[983:976] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_122[13] = buffer_data_2[991:984] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_122[14] = buffer_data_2[999:992] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_122[15] = buffer_data_1[967:960] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_122[16] = buffer_data_1[975:968] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_122[17] = buffer_data_1[983:976] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_122[18] = buffer_data_1[991:984] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_122[19] = buffer_data_1[999:992] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_122[20] = buffer_data_0[967:960] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_122[21] = buffer_data_0[975:968] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_122[22] = buffer_data_0[983:976] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_122[23] = buffer_data_0[991:984] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_122[24] = buffer_data_0[999:992] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_122 = kernel_img_mul_122[0] + kernel_img_mul_122[1] + kernel_img_mul_122[2] + 
                kernel_img_mul_122[3] + kernel_img_mul_122[4] + kernel_img_mul_122[5] + 
                kernel_img_mul_122[6] + kernel_img_mul_122[7] + kernel_img_mul_122[8] + 
                kernel_img_mul_122[9] + kernel_img_mul_122[10] + kernel_img_mul_122[11] + 
                kernel_img_mul_122[12] + kernel_img_mul_122[13] + kernel_img_mul_122[14] + 
                kernel_img_mul_122[15] + kernel_img_mul_122[16] + kernel_img_mul_122[17] + 
                kernel_img_mul_122[18] + kernel_img_mul_122[19] + kernel_img_mul_122[20] + 
                kernel_img_mul_122[21] + kernel_img_mul_122[22] + kernel_img_mul_122[23] + 
                kernel_img_mul_122[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[983:976] <= 'd0;
  else if (current_state==ST_START)
    blur_din[983:976] <= kernel_img_sum_122[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[983:976] <= 'd0;
end

wire  [39:0]  kernel_img_mul_123[0:24];
assign kernel_img_mul_123[0] = buffer_data_4[975:968] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_123[1] = buffer_data_4[983:976] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_123[2] = buffer_data_4[991:984] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_123[3] = buffer_data_4[999:992] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_123[4] = buffer_data_4[1007:1000] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_123[5] = buffer_data_3[975:968] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_123[6] = buffer_data_3[983:976] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_123[7] = buffer_data_3[991:984] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_123[8] = buffer_data_3[999:992] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_123[9] = buffer_data_3[1007:1000] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_123[10] = buffer_data_2[975:968] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_123[11] = buffer_data_2[983:976] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_123[12] = buffer_data_2[991:984] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_123[13] = buffer_data_2[999:992] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_123[14] = buffer_data_2[1007:1000] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_123[15] = buffer_data_1[975:968] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_123[16] = buffer_data_1[983:976] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_123[17] = buffer_data_1[991:984] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_123[18] = buffer_data_1[999:992] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_123[19] = buffer_data_1[1007:1000] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_123[20] = buffer_data_0[975:968] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_123[21] = buffer_data_0[983:976] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_123[22] = buffer_data_0[991:984] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_123[23] = buffer_data_0[999:992] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_123[24] = buffer_data_0[1007:1000] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_123 = kernel_img_mul_123[0] + kernel_img_mul_123[1] + kernel_img_mul_123[2] + 
                kernel_img_mul_123[3] + kernel_img_mul_123[4] + kernel_img_mul_123[5] + 
                kernel_img_mul_123[6] + kernel_img_mul_123[7] + kernel_img_mul_123[8] + 
                kernel_img_mul_123[9] + kernel_img_mul_123[10] + kernel_img_mul_123[11] + 
                kernel_img_mul_123[12] + kernel_img_mul_123[13] + kernel_img_mul_123[14] + 
                kernel_img_mul_123[15] + kernel_img_mul_123[16] + kernel_img_mul_123[17] + 
                kernel_img_mul_123[18] + kernel_img_mul_123[19] + kernel_img_mul_123[20] + 
                kernel_img_mul_123[21] + kernel_img_mul_123[22] + kernel_img_mul_123[23] + 
                kernel_img_mul_123[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[991:984] <= 'd0;
  else if (current_state==ST_START)
    blur_din[991:984] <= kernel_img_sum_123[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[991:984] <= 'd0;
end

wire  [39:0]  kernel_img_mul_124[0:24];
assign kernel_img_mul_124[0] = buffer_data_4[983:976] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_124[1] = buffer_data_4[991:984] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_124[2] = buffer_data_4[999:992] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_124[3] = buffer_data_4[1007:1000] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_124[4] = buffer_data_4[1015:1008] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_124[5] = buffer_data_3[983:976] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_124[6] = buffer_data_3[991:984] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_124[7] = buffer_data_3[999:992] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_124[8] = buffer_data_3[1007:1000] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_124[9] = buffer_data_3[1015:1008] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_124[10] = buffer_data_2[983:976] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_124[11] = buffer_data_2[991:984] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_124[12] = buffer_data_2[999:992] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_124[13] = buffer_data_2[1007:1000] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_124[14] = buffer_data_2[1015:1008] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_124[15] = buffer_data_1[983:976] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_124[16] = buffer_data_1[991:984] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_124[17] = buffer_data_1[999:992] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_124[18] = buffer_data_1[1007:1000] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_124[19] = buffer_data_1[1015:1008] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_124[20] = buffer_data_0[983:976] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_124[21] = buffer_data_0[991:984] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_124[22] = buffer_data_0[999:992] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_124[23] = buffer_data_0[1007:1000] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_124[24] = buffer_data_0[1015:1008] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_124 = kernel_img_mul_124[0] + kernel_img_mul_124[1] + kernel_img_mul_124[2] + 
                kernel_img_mul_124[3] + kernel_img_mul_124[4] + kernel_img_mul_124[5] + 
                kernel_img_mul_124[6] + kernel_img_mul_124[7] + kernel_img_mul_124[8] + 
                kernel_img_mul_124[9] + kernel_img_mul_124[10] + kernel_img_mul_124[11] + 
                kernel_img_mul_124[12] + kernel_img_mul_124[13] + kernel_img_mul_124[14] + 
                kernel_img_mul_124[15] + kernel_img_mul_124[16] + kernel_img_mul_124[17] + 
                kernel_img_mul_124[18] + kernel_img_mul_124[19] + kernel_img_mul_124[20] + 
                kernel_img_mul_124[21] + kernel_img_mul_124[22] + kernel_img_mul_124[23] + 
                kernel_img_mul_124[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[999:992] <= 'd0;
  else if (current_state==ST_START)
    blur_din[999:992] <= kernel_img_sum_124[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[999:992] <= 'd0;
end

wire  [39:0]  kernel_img_mul_125[0:24];
assign kernel_img_mul_125[0] = buffer_data_4[991:984] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_125[1] = buffer_data_4[999:992] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_125[2] = buffer_data_4[1007:1000] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_125[3] = buffer_data_4[1015:1008] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_125[4] = buffer_data_4[1023:1016] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_125[5] = buffer_data_3[991:984] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_125[6] = buffer_data_3[999:992] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_125[7] = buffer_data_3[1007:1000] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_125[8] = buffer_data_3[1015:1008] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_125[9] = buffer_data_3[1023:1016] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_125[10] = buffer_data_2[991:984] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_125[11] = buffer_data_2[999:992] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_125[12] = buffer_data_2[1007:1000] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_125[13] = buffer_data_2[1015:1008] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_125[14] = buffer_data_2[1023:1016] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_125[15] = buffer_data_1[991:984] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_125[16] = buffer_data_1[999:992] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_125[17] = buffer_data_1[1007:1000] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_125[18] = buffer_data_1[1015:1008] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_125[19] = buffer_data_1[1023:1016] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_125[20] = buffer_data_0[991:984] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_125[21] = buffer_data_0[999:992] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_125[22] = buffer_data_0[1007:1000] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_125[23] = buffer_data_0[1015:1008] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_125[24] = buffer_data_0[1023:1016] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_125 = kernel_img_mul_125[0] + kernel_img_mul_125[1] + kernel_img_mul_125[2] + 
                kernel_img_mul_125[3] + kernel_img_mul_125[4] + kernel_img_mul_125[5] + 
                kernel_img_mul_125[6] + kernel_img_mul_125[7] + kernel_img_mul_125[8] + 
                kernel_img_mul_125[9] + kernel_img_mul_125[10] + kernel_img_mul_125[11] + 
                kernel_img_mul_125[12] + kernel_img_mul_125[13] + kernel_img_mul_125[14] + 
                kernel_img_mul_125[15] + kernel_img_mul_125[16] + kernel_img_mul_125[17] + 
                kernel_img_mul_125[18] + kernel_img_mul_125[19] + kernel_img_mul_125[20] + 
                kernel_img_mul_125[21] + kernel_img_mul_125[22] + kernel_img_mul_125[23] + 
                kernel_img_mul_125[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1007:1000] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1007:1000] <= kernel_img_sum_125[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1007:1000] <= 'd0;
end

wire  [39:0]  kernel_img_mul_126[0:24];
assign kernel_img_mul_126[0] = buffer_data_4[999:992] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_126[1] = buffer_data_4[1007:1000] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_126[2] = buffer_data_4[1015:1008] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_126[3] = buffer_data_4[1023:1016] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_126[4] = buffer_data_4[1031:1024] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_126[5] = buffer_data_3[999:992] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_126[6] = buffer_data_3[1007:1000] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_126[7] = buffer_data_3[1015:1008] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_126[8] = buffer_data_3[1023:1016] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_126[9] = buffer_data_3[1031:1024] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_126[10] = buffer_data_2[999:992] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_126[11] = buffer_data_2[1007:1000] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_126[12] = buffer_data_2[1015:1008] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_126[13] = buffer_data_2[1023:1016] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_126[14] = buffer_data_2[1031:1024] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_126[15] = buffer_data_1[999:992] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_126[16] = buffer_data_1[1007:1000] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_126[17] = buffer_data_1[1015:1008] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_126[18] = buffer_data_1[1023:1016] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_126[19] = buffer_data_1[1031:1024] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_126[20] = buffer_data_0[999:992] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_126[21] = buffer_data_0[1007:1000] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_126[22] = buffer_data_0[1015:1008] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_126[23] = buffer_data_0[1023:1016] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_126[24] = buffer_data_0[1031:1024] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_126 = kernel_img_mul_126[0] + kernel_img_mul_126[1] + kernel_img_mul_126[2] + 
                kernel_img_mul_126[3] + kernel_img_mul_126[4] + kernel_img_mul_126[5] + 
                kernel_img_mul_126[6] + kernel_img_mul_126[7] + kernel_img_mul_126[8] + 
                kernel_img_mul_126[9] + kernel_img_mul_126[10] + kernel_img_mul_126[11] + 
                kernel_img_mul_126[12] + kernel_img_mul_126[13] + kernel_img_mul_126[14] + 
                kernel_img_mul_126[15] + kernel_img_mul_126[16] + kernel_img_mul_126[17] + 
                kernel_img_mul_126[18] + kernel_img_mul_126[19] + kernel_img_mul_126[20] + 
                kernel_img_mul_126[21] + kernel_img_mul_126[22] + kernel_img_mul_126[23] + 
                kernel_img_mul_126[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1015:1008] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1015:1008] <= kernel_img_sum_126[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1015:1008] <= 'd0;
end

wire  [39:0]  kernel_img_mul_127[0:24];
assign kernel_img_mul_127[0] = buffer_data_4[1007:1000] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_127[1] = buffer_data_4[1015:1008] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_127[2] = buffer_data_4[1023:1016] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_127[3] = buffer_data_4[1031:1024] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_127[4] = buffer_data_4[1039:1032] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_127[5] = buffer_data_3[1007:1000] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_127[6] = buffer_data_3[1015:1008] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_127[7] = buffer_data_3[1023:1016] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_127[8] = buffer_data_3[1031:1024] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_127[9] = buffer_data_3[1039:1032] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_127[10] = buffer_data_2[1007:1000] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_127[11] = buffer_data_2[1015:1008] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_127[12] = buffer_data_2[1023:1016] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_127[13] = buffer_data_2[1031:1024] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_127[14] = buffer_data_2[1039:1032] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_127[15] = buffer_data_1[1007:1000] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_127[16] = buffer_data_1[1015:1008] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_127[17] = buffer_data_1[1023:1016] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_127[18] = buffer_data_1[1031:1024] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_127[19] = buffer_data_1[1039:1032] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_127[20] = buffer_data_0[1007:1000] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_127[21] = buffer_data_0[1015:1008] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_127[22] = buffer_data_0[1023:1016] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_127[23] = buffer_data_0[1031:1024] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_127[24] = buffer_data_0[1039:1032] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_127 = kernel_img_mul_127[0] + kernel_img_mul_127[1] + kernel_img_mul_127[2] + 
                kernel_img_mul_127[3] + kernel_img_mul_127[4] + kernel_img_mul_127[5] + 
                kernel_img_mul_127[6] + kernel_img_mul_127[7] + kernel_img_mul_127[8] + 
                kernel_img_mul_127[9] + kernel_img_mul_127[10] + kernel_img_mul_127[11] + 
                kernel_img_mul_127[12] + kernel_img_mul_127[13] + kernel_img_mul_127[14] + 
                kernel_img_mul_127[15] + kernel_img_mul_127[16] + kernel_img_mul_127[17] + 
                kernel_img_mul_127[18] + kernel_img_mul_127[19] + kernel_img_mul_127[20] + 
                kernel_img_mul_127[21] + kernel_img_mul_127[22] + kernel_img_mul_127[23] + 
                kernel_img_mul_127[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1023:1016] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1023:1016] <= kernel_img_sum_127[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1023:1016] <= 'd0;
end

wire  [39:0]  kernel_img_mul_128[0:24];
assign kernel_img_mul_128[0] = buffer_data_4[1015:1008] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_128[1] = buffer_data_4[1023:1016] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_128[2] = buffer_data_4[1031:1024] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_128[3] = buffer_data_4[1039:1032] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_128[4] = buffer_data_4[1047:1040] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_128[5] = buffer_data_3[1015:1008] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_128[6] = buffer_data_3[1023:1016] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_128[7] = buffer_data_3[1031:1024] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_128[8] = buffer_data_3[1039:1032] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_128[9] = buffer_data_3[1047:1040] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_128[10] = buffer_data_2[1015:1008] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_128[11] = buffer_data_2[1023:1016] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_128[12] = buffer_data_2[1031:1024] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_128[13] = buffer_data_2[1039:1032] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_128[14] = buffer_data_2[1047:1040] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_128[15] = buffer_data_1[1015:1008] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_128[16] = buffer_data_1[1023:1016] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_128[17] = buffer_data_1[1031:1024] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_128[18] = buffer_data_1[1039:1032] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_128[19] = buffer_data_1[1047:1040] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_128[20] = buffer_data_0[1015:1008] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_128[21] = buffer_data_0[1023:1016] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_128[22] = buffer_data_0[1031:1024] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_128[23] = buffer_data_0[1039:1032] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_128[24] = buffer_data_0[1047:1040] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_128 = kernel_img_mul_128[0] + kernel_img_mul_128[1] + kernel_img_mul_128[2] + 
                kernel_img_mul_128[3] + kernel_img_mul_128[4] + kernel_img_mul_128[5] + 
                kernel_img_mul_128[6] + kernel_img_mul_128[7] + kernel_img_mul_128[8] + 
                kernel_img_mul_128[9] + kernel_img_mul_128[10] + kernel_img_mul_128[11] + 
                kernel_img_mul_128[12] + kernel_img_mul_128[13] + kernel_img_mul_128[14] + 
                kernel_img_mul_128[15] + kernel_img_mul_128[16] + kernel_img_mul_128[17] + 
                kernel_img_mul_128[18] + kernel_img_mul_128[19] + kernel_img_mul_128[20] + 
                kernel_img_mul_128[21] + kernel_img_mul_128[22] + kernel_img_mul_128[23] + 
                kernel_img_mul_128[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1031:1024] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1031:1024] <= kernel_img_sum_128[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1031:1024] <= 'd0;
end

wire  [39:0]  kernel_img_mul_129[0:24];
assign kernel_img_mul_129[0] = buffer_data_4[1023:1016] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_129[1] = buffer_data_4[1031:1024] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_129[2] = buffer_data_4[1039:1032] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_129[3] = buffer_data_4[1047:1040] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_129[4] = buffer_data_4[1055:1048] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_129[5] = buffer_data_3[1023:1016] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_129[6] = buffer_data_3[1031:1024] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_129[7] = buffer_data_3[1039:1032] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_129[8] = buffer_data_3[1047:1040] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_129[9] = buffer_data_3[1055:1048] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_129[10] = buffer_data_2[1023:1016] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_129[11] = buffer_data_2[1031:1024] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_129[12] = buffer_data_2[1039:1032] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_129[13] = buffer_data_2[1047:1040] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_129[14] = buffer_data_2[1055:1048] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_129[15] = buffer_data_1[1023:1016] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_129[16] = buffer_data_1[1031:1024] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_129[17] = buffer_data_1[1039:1032] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_129[18] = buffer_data_1[1047:1040] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_129[19] = buffer_data_1[1055:1048] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_129[20] = buffer_data_0[1023:1016] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_129[21] = buffer_data_0[1031:1024] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_129[22] = buffer_data_0[1039:1032] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_129[23] = buffer_data_0[1047:1040] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_129[24] = buffer_data_0[1055:1048] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_129 = kernel_img_mul_129[0] + kernel_img_mul_129[1] + kernel_img_mul_129[2] + 
                kernel_img_mul_129[3] + kernel_img_mul_129[4] + kernel_img_mul_129[5] + 
                kernel_img_mul_129[6] + kernel_img_mul_129[7] + kernel_img_mul_129[8] + 
                kernel_img_mul_129[9] + kernel_img_mul_129[10] + kernel_img_mul_129[11] + 
                kernel_img_mul_129[12] + kernel_img_mul_129[13] + kernel_img_mul_129[14] + 
                kernel_img_mul_129[15] + kernel_img_mul_129[16] + kernel_img_mul_129[17] + 
                kernel_img_mul_129[18] + kernel_img_mul_129[19] + kernel_img_mul_129[20] + 
                kernel_img_mul_129[21] + kernel_img_mul_129[22] + kernel_img_mul_129[23] + 
                kernel_img_mul_129[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1039:1032] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1039:1032] <= kernel_img_sum_129[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1039:1032] <= 'd0;
end

wire  [39:0]  kernel_img_mul_130[0:24];
assign kernel_img_mul_130[0] = buffer_data_4[1031:1024] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_130[1] = buffer_data_4[1039:1032] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_130[2] = buffer_data_4[1047:1040] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_130[3] = buffer_data_4[1055:1048] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_130[4] = buffer_data_4[1063:1056] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_130[5] = buffer_data_3[1031:1024] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_130[6] = buffer_data_3[1039:1032] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_130[7] = buffer_data_3[1047:1040] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_130[8] = buffer_data_3[1055:1048] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_130[9] = buffer_data_3[1063:1056] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_130[10] = buffer_data_2[1031:1024] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_130[11] = buffer_data_2[1039:1032] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_130[12] = buffer_data_2[1047:1040] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_130[13] = buffer_data_2[1055:1048] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_130[14] = buffer_data_2[1063:1056] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_130[15] = buffer_data_1[1031:1024] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_130[16] = buffer_data_1[1039:1032] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_130[17] = buffer_data_1[1047:1040] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_130[18] = buffer_data_1[1055:1048] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_130[19] = buffer_data_1[1063:1056] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_130[20] = buffer_data_0[1031:1024] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_130[21] = buffer_data_0[1039:1032] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_130[22] = buffer_data_0[1047:1040] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_130[23] = buffer_data_0[1055:1048] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_130[24] = buffer_data_0[1063:1056] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_130 = kernel_img_mul_130[0] + kernel_img_mul_130[1] + kernel_img_mul_130[2] + 
                kernel_img_mul_130[3] + kernel_img_mul_130[4] + kernel_img_mul_130[5] + 
                kernel_img_mul_130[6] + kernel_img_mul_130[7] + kernel_img_mul_130[8] + 
                kernel_img_mul_130[9] + kernel_img_mul_130[10] + kernel_img_mul_130[11] + 
                kernel_img_mul_130[12] + kernel_img_mul_130[13] + kernel_img_mul_130[14] + 
                kernel_img_mul_130[15] + kernel_img_mul_130[16] + kernel_img_mul_130[17] + 
                kernel_img_mul_130[18] + kernel_img_mul_130[19] + kernel_img_mul_130[20] + 
                kernel_img_mul_130[21] + kernel_img_mul_130[22] + kernel_img_mul_130[23] + 
                kernel_img_mul_130[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1047:1040] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1047:1040] <= kernel_img_sum_130[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1047:1040] <= 'd0;
end

wire  [39:0]  kernel_img_mul_131[0:24];
assign kernel_img_mul_131[0] = buffer_data_4[1039:1032] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_131[1] = buffer_data_4[1047:1040] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_131[2] = buffer_data_4[1055:1048] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_131[3] = buffer_data_4[1063:1056] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_131[4] = buffer_data_4[1071:1064] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_131[5] = buffer_data_3[1039:1032] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_131[6] = buffer_data_3[1047:1040] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_131[7] = buffer_data_3[1055:1048] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_131[8] = buffer_data_3[1063:1056] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_131[9] = buffer_data_3[1071:1064] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_131[10] = buffer_data_2[1039:1032] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_131[11] = buffer_data_2[1047:1040] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_131[12] = buffer_data_2[1055:1048] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_131[13] = buffer_data_2[1063:1056] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_131[14] = buffer_data_2[1071:1064] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_131[15] = buffer_data_1[1039:1032] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_131[16] = buffer_data_1[1047:1040] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_131[17] = buffer_data_1[1055:1048] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_131[18] = buffer_data_1[1063:1056] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_131[19] = buffer_data_1[1071:1064] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_131[20] = buffer_data_0[1039:1032] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_131[21] = buffer_data_0[1047:1040] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_131[22] = buffer_data_0[1055:1048] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_131[23] = buffer_data_0[1063:1056] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_131[24] = buffer_data_0[1071:1064] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_131 = kernel_img_mul_131[0] + kernel_img_mul_131[1] + kernel_img_mul_131[2] + 
                kernel_img_mul_131[3] + kernel_img_mul_131[4] + kernel_img_mul_131[5] + 
                kernel_img_mul_131[6] + kernel_img_mul_131[7] + kernel_img_mul_131[8] + 
                kernel_img_mul_131[9] + kernel_img_mul_131[10] + kernel_img_mul_131[11] + 
                kernel_img_mul_131[12] + kernel_img_mul_131[13] + kernel_img_mul_131[14] + 
                kernel_img_mul_131[15] + kernel_img_mul_131[16] + kernel_img_mul_131[17] + 
                kernel_img_mul_131[18] + kernel_img_mul_131[19] + kernel_img_mul_131[20] + 
                kernel_img_mul_131[21] + kernel_img_mul_131[22] + kernel_img_mul_131[23] + 
                kernel_img_mul_131[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1055:1048] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1055:1048] <= kernel_img_sum_131[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1055:1048] <= 'd0;
end

wire  [39:0]  kernel_img_mul_132[0:24];
assign kernel_img_mul_132[0] = buffer_data_4[1047:1040] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_132[1] = buffer_data_4[1055:1048] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_132[2] = buffer_data_4[1063:1056] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_132[3] = buffer_data_4[1071:1064] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_132[4] = buffer_data_4[1079:1072] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_132[5] = buffer_data_3[1047:1040] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_132[6] = buffer_data_3[1055:1048] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_132[7] = buffer_data_3[1063:1056] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_132[8] = buffer_data_3[1071:1064] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_132[9] = buffer_data_3[1079:1072] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_132[10] = buffer_data_2[1047:1040] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_132[11] = buffer_data_2[1055:1048] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_132[12] = buffer_data_2[1063:1056] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_132[13] = buffer_data_2[1071:1064] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_132[14] = buffer_data_2[1079:1072] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_132[15] = buffer_data_1[1047:1040] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_132[16] = buffer_data_1[1055:1048] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_132[17] = buffer_data_1[1063:1056] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_132[18] = buffer_data_1[1071:1064] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_132[19] = buffer_data_1[1079:1072] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_132[20] = buffer_data_0[1047:1040] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_132[21] = buffer_data_0[1055:1048] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_132[22] = buffer_data_0[1063:1056] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_132[23] = buffer_data_0[1071:1064] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_132[24] = buffer_data_0[1079:1072] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_132 = kernel_img_mul_132[0] + kernel_img_mul_132[1] + kernel_img_mul_132[2] + 
                kernel_img_mul_132[3] + kernel_img_mul_132[4] + kernel_img_mul_132[5] + 
                kernel_img_mul_132[6] + kernel_img_mul_132[7] + kernel_img_mul_132[8] + 
                kernel_img_mul_132[9] + kernel_img_mul_132[10] + kernel_img_mul_132[11] + 
                kernel_img_mul_132[12] + kernel_img_mul_132[13] + kernel_img_mul_132[14] + 
                kernel_img_mul_132[15] + kernel_img_mul_132[16] + kernel_img_mul_132[17] + 
                kernel_img_mul_132[18] + kernel_img_mul_132[19] + kernel_img_mul_132[20] + 
                kernel_img_mul_132[21] + kernel_img_mul_132[22] + kernel_img_mul_132[23] + 
                kernel_img_mul_132[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1063:1056] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1063:1056] <= kernel_img_sum_132[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1063:1056] <= 'd0;
end

wire  [39:0]  kernel_img_mul_133[0:24];
assign kernel_img_mul_133[0] = buffer_data_4[1055:1048] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_133[1] = buffer_data_4[1063:1056] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_133[2] = buffer_data_4[1071:1064] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_133[3] = buffer_data_4[1079:1072] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_133[4] = buffer_data_4[1087:1080] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_133[5] = buffer_data_3[1055:1048] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_133[6] = buffer_data_3[1063:1056] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_133[7] = buffer_data_3[1071:1064] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_133[8] = buffer_data_3[1079:1072] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_133[9] = buffer_data_3[1087:1080] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_133[10] = buffer_data_2[1055:1048] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_133[11] = buffer_data_2[1063:1056] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_133[12] = buffer_data_2[1071:1064] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_133[13] = buffer_data_2[1079:1072] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_133[14] = buffer_data_2[1087:1080] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_133[15] = buffer_data_1[1055:1048] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_133[16] = buffer_data_1[1063:1056] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_133[17] = buffer_data_1[1071:1064] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_133[18] = buffer_data_1[1079:1072] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_133[19] = buffer_data_1[1087:1080] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_133[20] = buffer_data_0[1055:1048] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_133[21] = buffer_data_0[1063:1056] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_133[22] = buffer_data_0[1071:1064] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_133[23] = buffer_data_0[1079:1072] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_133[24] = buffer_data_0[1087:1080] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_133 = kernel_img_mul_133[0] + kernel_img_mul_133[1] + kernel_img_mul_133[2] + 
                kernel_img_mul_133[3] + kernel_img_mul_133[4] + kernel_img_mul_133[5] + 
                kernel_img_mul_133[6] + kernel_img_mul_133[7] + kernel_img_mul_133[8] + 
                kernel_img_mul_133[9] + kernel_img_mul_133[10] + kernel_img_mul_133[11] + 
                kernel_img_mul_133[12] + kernel_img_mul_133[13] + kernel_img_mul_133[14] + 
                kernel_img_mul_133[15] + kernel_img_mul_133[16] + kernel_img_mul_133[17] + 
                kernel_img_mul_133[18] + kernel_img_mul_133[19] + kernel_img_mul_133[20] + 
                kernel_img_mul_133[21] + kernel_img_mul_133[22] + kernel_img_mul_133[23] + 
                kernel_img_mul_133[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1071:1064] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1071:1064] <= kernel_img_sum_133[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1071:1064] <= 'd0;
end

wire  [39:0]  kernel_img_mul_134[0:24];
assign kernel_img_mul_134[0] = buffer_data_4[1063:1056] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_134[1] = buffer_data_4[1071:1064] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_134[2] = buffer_data_4[1079:1072] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_134[3] = buffer_data_4[1087:1080] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_134[4] = buffer_data_4[1095:1088] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_134[5] = buffer_data_3[1063:1056] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_134[6] = buffer_data_3[1071:1064] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_134[7] = buffer_data_3[1079:1072] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_134[8] = buffer_data_3[1087:1080] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_134[9] = buffer_data_3[1095:1088] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_134[10] = buffer_data_2[1063:1056] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_134[11] = buffer_data_2[1071:1064] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_134[12] = buffer_data_2[1079:1072] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_134[13] = buffer_data_2[1087:1080] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_134[14] = buffer_data_2[1095:1088] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_134[15] = buffer_data_1[1063:1056] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_134[16] = buffer_data_1[1071:1064] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_134[17] = buffer_data_1[1079:1072] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_134[18] = buffer_data_1[1087:1080] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_134[19] = buffer_data_1[1095:1088] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_134[20] = buffer_data_0[1063:1056] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_134[21] = buffer_data_0[1071:1064] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_134[22] = buffer_data_0[1079:1072] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_134[23] = buffer_data_0[1087:1080] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_134[24] = buffer_data_0[1095:1088] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_134 = kernel_img_mul_134[0] + kernel_img_mul_134[1] + kernel_img_mul_134[2] + 
                kernel_img_mul_134[3] + kernel_img_mul_134[4] + kernel_img_mul_134[5] + 
                kernel_img_mul_134[6] + kernel_img_mul_134[7] + kernel_img_mul_134[8] + 
                kernel_img_mul_134[9] + kernel_img_mul_134[10] + kernel_img_mul_134[11] + 
                kernel_img_mul_134[12] + kernel_img_mul_134[13] + kernel_img_mul_134[14] + 
                kernel_img_mul_134[15] + kernel_img_mul_134[16] + kernel_img_mul_134[17] + 
                kernel_img_mul_134[18] + kernel_img_mul_134[19] + kernel_img_mul_134[20] + 
                kernel_img_mul_134[21] + kernel_img_mul_134[22] + kernel_img_mul_134[23] + 
                kernel_img_mul_134[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1079:1072] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1079:1072] <= kernel_img_sum_134[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1079:1072] <= 'd0;
end

wire  [39:0]  kernel_img_mul_135[0:24];
assign kernel_img_mul_135[0] = buffer_data_4[1071:1064] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_135[1] = buffer_data_4[1079:1072] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_135[2] = buffer_data_4[1087:1080] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_135[3] = buffer_data_4[1095:1088] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_135[4] = buffer_data_4[1103:1096] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_135[5] = buffer_data_3[1071:1064] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_135[6] = buffer_data_3[1079:1072] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_135[7] = buffer_data_3[1087:1080] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_135[8] = buffer_data_3[1095:1088] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_135[9] = buffer_data_3[1103:1096] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_135[10] = buffer_data_2[1071:1064] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_135[11] = buffer_data_2[1079:1072] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_135[12] = buffer_data_2[1087:1080] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_135[13] = buffer_data_2[1095:1088] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_135[14] = buffer_data_2[1103:1096] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_135[15] = buffer_data_1[1071:1064] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_135[16] = buffer_data_1[1079:1072] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_135[17] = buffer_data_1[1087:1080] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_135[18] = buffer_data_1[1095:1088] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_135[19] = buffer_data_1[1103:1096] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_135[20] = buffer_data_0[1071:1064] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_135[21] = buffer_data_0[1079:1072] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_135[22] = buffer_data_0[1087:1080] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_135[23] = buffer_data_0[1095:1088] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_135[24] = buffer_data_0[1103:1096] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_135 = kernel_img_mul_135[0] + kernel_img_mul_135[1] + kernel_img_mul_135[2] + 
                kernel_img_mul_135[3] + kernel_img_mul_135[4] + kernel_img_mul_135[5] + 
                kernel_img_mul_135[6] + kernel_img_mul_135[7] + kernel_img_mul_135[8] + 
                kernel_img_mul_135[9] + kernel_img_mul_135[10] + kernel_img_mul_135[11] + 
                kernel_img_mul_135[12] + kernel_img_mul_135[13] + kernel_img_mul_135[14] + 
                kernel_img_mul_135[15] + kernel_img_mul_135[16] + kernel_img_mul_135[17] + 
                kernel_img_mul_135[18] + kernel_img_mul_135[19] + kernel_img_mul_135[20] + 
                kernel_img_mul_135[21] + kernel_img_mul_135[22] + kernel_img_mul_135[23] + 
                kernel_img_mul_135[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1087:1080] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1087:1080] <= kernel_img_sum_135[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1087:1080] <= 'd0;
end

wire  [39:0]  kernel_img_mul_136[0:24];
assign kernel_img_mul_136[0] = buffer_data_4[1079:1072] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_136[1] = buffer_data_4[1087:1080] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_136[2] = buffer_data_4[1095:1088] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_136[3] = buffer_data_4[1103:1096] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_136[4] = buffer_data_4[1111:1104] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_136[5] = buffer_data_3[1079:1072] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_136[6] = buffer_data_3[1087:1080] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_136[7] = buffer_data_3[1095:1088] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_136[8] = buffer_data_3[1103:1096] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_136[9] = buffer_data_3[1111:1104] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_136[10] = buffer_data_2[1079:1072] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_136[11] = buffer_data_2[1087:1080] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_136[12] = buffer_data_2[1095:1088] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_136[13] = buffer_data_2[1103:1096] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_136[14] = buffer_data_2[1111:1104] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_136[15] = buffer_data_1[1079:1072] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_136[16] = buffer_data_1[1087:1080] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_136[17] = buffer_data_1[1095:1088] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_136[18] = buffer_data_1[1103:1096] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_136[19] = buffer_data_1[1111:1104] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_136[20] = buffer_data_0[1079:1072] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_136[21] = buffer_data_0[1087:1080] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_136[22] = buffer_data_0[1095:1088] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_136[23] = buffer_data_0[1103:1096] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_136[24] = buffer_data_0[1111:1104] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_136 = kernel_img_mul_136[0] + kernel_img_mul_136[1] + kernel_img_mul_136[2] + 
                kernel_img_mul_136[3] + kernel_img_mul_136[4] + kernel_img_mul_136[5] + 
                kernel_img_mul_136[6] + kernel_img_mul_136[7] + kernel_img_mul_136[8] + 
                kernel_img_mul_136[9] + kernel_img_mul_136[10] + kernel_img_mul_136[11] + 
                kernel_img_mul_136[12] + kernel_img_mul_136[13] + kernel_img_mul_136[14] + 
                kernel_img_mul_136[15] + kernel_img_mul_136[16] + kernel_img_mul_136[17] + 
                kernel_img_mul_136[18] + kernel_img_mul_136[19] + kernel_img_mul_136[20] + 
                kernel_img_mul_136[21] + kernel_img_mul_136[22] + kernel_img_mul_136[23] + 
                kernel_img_mul_136[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1095:1088] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1095:1088] <= kernel_img_sum_136[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1095:1088] <= 'd0;
end

wire  [39:0]  kernel_img_mul_137[0:24];
assign kernel_img_mul_137[0] = buffer_data_4[1087:1080] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_137[1] = buffer_data_4[1095:1088] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_137[2] = buffer_data_4[1103:1096] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_137[3] = buffer_data_4[1111:1104] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_137[4] = buffer_data_4[1119:1112] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_137[5] = buffer_data_3[1087:1080] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_137[6] = buffer_data_3[1095:1088] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_137[7] = buffer_data_3[1103:1096] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_137[8] = buffer_data_3[1111:1104] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_137[9] = buffer_data_3[1119:1112] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_137[10] = buffer_data_2[1087:1080] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_137[11] = buffer_data_2[1095:1088] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_137[12] = buffer_data_2[1103:1096] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_137[13] = buffer_data_2[1111:1104] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_137[14] = buffer_data_2[1119:1112] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_137[15] = buffer_data_1[1087:1080] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_137[16] = buffer_data_1[1095:1088] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_137[17] = buffer_data_1[1103:1096] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_137[18] = buffer_data_1[1111:1104] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_137[19] = buffer_data_1[1119:1112] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_137[20] = buffer_data_0[1087:1080] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_137[21] = buffer_data_0[1095:1088] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_137[22] = buffer_data_0[1103:1096] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_137[23] = buffer_data_0[1111:1104] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_137[24] = buffer_data_0[1119:1112] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_137 = kernel_img_mul_137[0] + kernel_img_mul_137[1] + kernel_img_mul_137[2] + 
                kernel_img_mul_137[3] + kernel_img_mul_137[4] + kernel_img_mul_137[5] + 
                kernel_img_mul_137[6] + kernel_img_mul_137[7] + kernel_img_mul_137[8] + 
                kernel_img_mul_137[9] + kernel_img_mul_137[10] + kernel_img_mul_137[11] + 
                kernel_img_mul_137[12] + kernel_img_mul_137[13] + kernel_img_mul_137[14] + 
                kernel_img_mul_137[15] + kernel_img_mul_137[16] + kernel_img_mul_137[17] + 
                kernel_img_mul_137[18] + kernel_img_mul_137[19] + kernel_img_mul_137[20] + 
                kernel_img_mul_137[21] + kernel_img_mul_137[22] + kernel_img_mul_137[23] + 
                kernel_img_mul_137[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1103:1096] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1103:1096] <= kernel_img_sum_137[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1103:1096] <= 'd0;
end

wire  [39:0]  kernel_img_mul_138[0:24];
assign kernel_img_mul_138[0] = buffer_data_4[1095:1088] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_138[1] = buffer_data_4[1103:1096] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_138[2] = buffer_data_4[1111:1104] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_138[3] = buffer_data_4[1119:1112] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_138[4] = buffer_data_4[1127:1120] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_138[5] = buffer_data_3[1095:1088] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_138[6] = buffer_data_3[1103:1096] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_138[7] = buffer_data_3[1111:1104] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_138[8] = buffer_data_3[1119:1112] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_138[9] = buffer_data_3[1127:1120] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_138[10] = buffer_data_2[1095:1088] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_138[11] = buffer_data_2[1103:1096] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_138[12] = buffer_data_2[1111:1104] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_138[13] = buffer_data_2[1119:1112] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_138[14] = buffer_data_2[1127:1120] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_138[15] = buffer_data_1[1095:1088] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_138[16] = buffer_data_1[1103:1096] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_138[17] = buffer_data_1[1111:1104] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_138[18] = buffer_data_1[1119:1112] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_138[19] = buffer_data_1[1127:1120] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_138[20] = buffer_data_0[1095:1088] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_138[21] = buffer_data_0[1103:1096] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_138[22] = buffer_data_0[1111:1104] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_138[23] = buffer_data_0[1119:1112] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_138[24] = buffer_data_0[1127:1120] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_138 = kernel_img_mul_138[0] + kernel_img_mul_138[1] + kernel_img_mul_138[2] + 
                kernel_img_mul_138[3] + kernel_img_mul_138[4] + kernel_img_mul_138[5] + 
                kernel_img_mul_138[6] + kernel_img_mul_138[7] + kernel_img_mul_138[8] + 
                kernel_img_mul_138[9] + kernel_img_mul_138[10] + kernel_img_mul_138[11] + 
                kernel_img_mul_138[12] + kernel_img_mul_138[13] + kernel_img_mul_138[14] + 
                kernel_img_mul_138[15] + kernel_img_mul_138[16] + kernel_img_mul_138[17] + 
                kernel_img_mul_138[18] + kernel_img_mul_138[19] + kernel_img_mul_138[20] + 
                kernel_img_mul_138[21] + kernel_img_mul_138[22] + kernel_img_mul_138[23] + 
                kernel_img_mul_138[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1111:1104] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1111:1104] <= kernel_img_sum_138[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1111:1104] <= 'd0;
end

wire  [39:0]  kernel_img_mul_139[0:24];
assign kernel_img_mul_139[0] = buffer_data_4[1103:1096] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_139[1] = buffer_data_4[1111:1104] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_139[2] = buffer_data_4[1119:1112] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_139[3] = buffer_data_4[1127:1120] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_139[4] = buffer_data_4[1135:1128] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_139[5] = buffer_data_3[1103:1096] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_139[6] = buffer_data_3[1111:1104] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_139[7] = buffer_data_3[1119:1112] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_139[8] = buffer_data_3[1127:1120] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_139[9] = buffer_data_3[1135:1128] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_139[10] = buffer_data_2[1103:1096] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_139[11] = buffer_data_2[1111:1104] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_139[12] = buffer_data_2[1119:1112] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_139[13] = buffer_data_2[1127:1120] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_139[14] = buffer_data_2[1135:1128] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_139[15] = buffer_data_1[1103:1096] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_139[16] = buffer_data_1[1111:1104] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_139[17] = buffer_data_1[1119:1112] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_139[18] = buffer_data_1[1127:1120] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_139[19] = buffer_data_1[1135:1128] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_139[20] = buffer_data_0[1103:1096] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_139[21] = buffer_data_0[1111:1104] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_139[22] = buffer_data_0[1119:1112] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_139[23] = buffer_data_0[1127:1120] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_139[24] = buffer_data_0[1135:1128] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_139 = kernel_img_mul_139[0] + kernel_img_mul_139[1] + kernel_img_mul_139[2] + 
                kernel_img_mul_139[3] + kernel_img_mul_139[4] + kernel_img_mul_139[5] + 
                kernel_img_mul_139[6] + kernel_img_mul_139[7] + kernel_img_mul_139[8] + 
                kernel_img_mul_139[9] + kernel_img_mul_139[10] + kernel_img_mul_139[11] + 
                kernel_img_mul_139[12] + kernel_img_mul_139[13] + kernel_img_mul_139[14] + 
                kernel_img_mul_139[15] + kernel_img_mul_139[16] + kernel_img_mul_139[17] + 
                kernel_img_mul_139[18] + kernel_img_mul_139[19] + kernel_img_mul_139[20] + 
                kernel_img_mul_139[21] + kernel_img_mul_139[22] + kernel_img_mul_139[23] + 
                kernel_img_mul_139[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1119:1112] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1119:1112] <= kernel_img_sum_139[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1119:1112] <= 'd0;
end

wire  [39:0]  kernel_img_mul_140[0:24];
assign kernel_img_mul_140[0] = buffer_data_4[1111:1104] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_140[1] = buffer_data_4[1119:1112] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_140[2] = buffer_data_4[1127:1120] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_140[3] = buffer_data_4[1135:1128] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_140[4] = buffer_data_4[1143:1136] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_140[5] = buffer_data_3[1111:1104] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_140[6] = buffer_data_3[1119:1112] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_140[7] = buffer_data_3[1127:1120] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_140[8] = buffer_data_3[1135:1128] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_140[9] = buffer_data_3[1143:1136] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_140[10] = buffer_data_2[1111:1104] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_140[11] = buffer_data_2[1119:1112] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_140[12] = buffer_data_2[1127:1120] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_140[13] = buffer_data_2[1135:1128] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_140[14] = buffer_data_2[1143:1136] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_140[15] = buffer_data_1[1111:1104] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_140[16] = buffer_data_1[1119:1112] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_140[17] = buffer_data_1[1127:1120] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_140[18] = buffer_data_1[1135:1128] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_140[19] = buffer_data_1[1143:1136] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_140[20] = buffer_data_0[1111:1104] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_140[21] = buffer_data_0[1119:1112] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_140[22] = buffer_data_0[1127:1120] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_140[23] = buffer_data_0[1135:1128] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_140[24] = buffer_data_0[1143:1136] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_140 = kernel_img_mul_140[0] + kernel_img_mul_140[1] + kernel_img_mul_140[2] + 
                kernel_img_mul_140[3] + kernel_img_mul_140[4] + kernel_img_mul_140[5] + 
                kernel_img_mul_140[6] + kernel_img_mul_140[7] + kernel_img_mul_140[8] + 
                kernel_img_mul_140[9] + kernel_img_mul_140[10] + kernel_img_mul_140[11] + 
                kernel_img_mul_140[12] + kernel_img_mul_140[13] + kernel_img_mul_140[14] + 
                kernel_img_mul_140[15] + kernel_img_mul_140[16] + kernel_img_mul_140[17] + 
                kernel_img_mul_140[18] + kernel_img_mul_140[19] + kernel_img_mul_140[20] + 
                kernel_img_mul_140[21] + kernel_img_mul_140[22] + kernel_img_mul_140[23] + 
                kernel_img_mul_140[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1127:1120] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1127:1120] <= kernel_img_sum_140[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1127:1120] <= 'd0;
end

wire  [39:0]  kernel_img_mul_141[0:24];
assign kernel_img_mul_141[0] = buffer_data_4[1119:1112] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_141[1] = buffer_data_4[1127:1120] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_141[2] = buffer_data_4[1135:1128] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_141[3] = buffer_data_4[1143:1136] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_141[4] = buffer_data_4[1151:1144] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_141[5] = buffer_data_3[1119:1112] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_141[6] = buffer_data_3[1127:1120] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_141[7] = buffer_data_3[1135:1128] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_141[8] = buffer_data_3[1143:1136] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_141[9] = buffer_data_3[1151:1144] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_141[10] = buffer_data_2[1119:1112] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_141[11] = buffer_data_2[1127:1120] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_141[12] = buffer_data_2[1135:1128] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_141[13] = buffer_data_2[1143:1136] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_141[14] = buffer_data_2[1151:1144] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_141[15] = buffer_data_1[1119:1112] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_141[16] = buffer_data_1[1127:1120] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_141[17] = buffer_data_1[1135:1128] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_141[18] = buffer_data_1[1143:1136] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_141[19] = buffer_data_1[1151:1144] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_141[20] = buffer_data_0[1119:1112] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_141[21] = buffer_data_0[1127:1120] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_141[22] = buffer_data_0[1135:1128] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_141[23] = buffer_data_0[1143:1136] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_141[24] = buffer_data_0[1151:1144] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_141 = kernel_img_mul_141[0] + kernel_img_mul_141[1] + kernel_img_mul_141[2] + 
                kernel_img_mul_141[3] + kernel_img_mul_141[4] + kernel_img_mul_141[5] + 
                kernel_img_mul_141[6] + kernel_img_mul_141[7] + kernel_img_mul_141[8] + 
                kernel_img_mul_141[9] + kernel_img_mul_141[10] + kernel_img_mul_141[11] + 
                kernel_img_mul_141[12] + kernel_img_mul_141[13] + kernel_img_mul_141[14] + 
                kernel_img_mul_141[15] + kernel_img_mul_141[16] + kernel_img_mul_141[17] + 
                kernel_img_mul_141[18] + kernel_img_mul_141[19] + kernel_img_mul_141[20] + 
                kernel_img_mul_141[21] + kernel_img_mul_141[22] + kernel_img_mul_141[23] + 
                kernel_img_mul_141[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1135:1128] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1135:1128] <= kernel_img_sum_141[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1135:1128] <= 'd0;
end

wire  [39:0]  kernel_img_mul_142[0:24];
assign kernel_img_mul_142[0] = buffer_data_4[1127:1120] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_142[1] = buffer_data_4[1135:1128] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_142[2] = buffer_data_4[1143:1136] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_142[3] = buffer_data_4[1151:1144] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_142[4] = buffer_data_4[1159:1152] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_142[5] = buffer_data_3[1127:1120] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_142[6] = buffer_data_3[1135:1128] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_142[7] = buffer_data_3[1143:1136] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_142[8] = buffer_data_3[1151:1144] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_142[9] = buffer_data_3[1159:1152] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_142[10] = buffer_data_2[1127:1120] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_142[11] = buffer_data_2[1135:1128] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_142[12] = buffer_data_2[1143:1136] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_142[13] = buffer_data_2[1151:1144] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_142[14] = buffer_data_2[1159:1152] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_142[15] = buffer_data_1[1127:1120] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_142[16] = buffer_data_1[1135:1128] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_142[17] = buffer_data_1[1143:1136] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_142[18] = buffer_data_1[1151:1144] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_142[19] = buffer_data_1[1159:1152] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_142[20] = buffer_data_0[1127:1120] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_142[21] = buffer_data_0[1135:1128] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_142[22] = buffer_data_0[1143:1136] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_142[23] = buffer_data_0[1151:1144] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_142[24] = buffer_data_0[1159:1152] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_142 = kernel_img_mul_142[0] + kernel_img_mul_142[1] + kernel_img_mul_142[2] + 
                kernel_img_mul_142[3] + kernel_img_mul_142[4] + kernel_img_mul_142[5] + 
                kernel_img_mul_142[6] + kernel_img_mul_142[7] + kernel_img_mul_142[8] + 
                kernel_img_mul_142[9] + kernel_img_mul_142[10] + kernel_img_mul_142[11] + 
                kernel_img_mul_142[12] + kernel_img_mul_142[13] + kernel_img_mul_142[14] + 
                kernel_img_mul_142[15] + kernel_img_mul_142[16] + kernel_img_mul_142[17] + 
                kernel_img_mul_142[18] + kernel_img_mul_142[19] + kernel_img_mul_142[20] + 
                kernel_img_mul_142[21] + kernel_img_mul_142[22] + kernel_img_mul_142[23] + 
                kernel_img_mul_142[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1143:1136] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1143:1136] <= kernel_img_sum_142[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1143:1136] <= 'd0;
end

wire  [39:0]  kernel_img_mul_143[0:24];
assign kernel_img_mul_143[0] = buffer_data_4[1135:1128] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_143[1] = buffer_data_4[1143:1136] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_143[2] = buffer_data_4[1151:1144] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_143[3] = buffer_data_4[1159:1152] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_143[4] = buffer_data_4[1167:1160] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_143[5] = buffer_data_3[1135:1128] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_143[6] = buffer_data_3[1143:1136] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_143[7] = buffer_data_3[1151:1144] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_143[8] = buffer_data_3[1159:1152] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_143[9] = buffer_data_3[1167:1160] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_143[10] = buffer_data_2[1135:1128] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_143[11] = buffer_data_2[1143:1136] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_143[12] = buffer_data_2[1151:1144] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_143[13] = buffer_data_2[1159:1152] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_143[14] = buffer_data_2[1167:1160] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_143[15] = buffer_data_1[1135:1128] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_143[16] = buffer_data_1[1143:1136] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_143[17] = buffer_data_1[1151:1144] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_143[18] = buffer_data_1[1159:1152] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_143[19] = buffer_data_1[1167:1160] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_143[20] = buffer_data_0[1135:1128] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_143[21] = buffer_data_0[1143:1136] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_143[22] = buffer_data_0[1151:1144] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_143[23] = buffer_data_0[1159:1152] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_143[24] = buffer_data_0[1167:1160] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_143 = kernel_img_mul_143[0] + kernel_img_mul_143[1] + kernel_img_mul_143[2] + 
                kernel_img_mul_143[3] + kernel_img_mul_143[4] + kernel_img_mul_143[5] + 
                kernel_img_mul_143[6] + kernel_img_mul_143[7] + kernel_img_mul_143[8] + 
                kernel_img_mul_143[9] + kernel_img_mul_143[10] + kernel_img_mul_143[11] + 
                kernel_img_mul_143[12] + kernel_img_mul_143[13] + kernel_img_mul_143[14] + 
                kernel_img_mul_143[15] + kernel_img_mul_143[16] + kernel_img_mul_143[17] + 
                kernel_img_mul_143[18] + kernel_img_mul_143[19] + kernel_img_mul_143[20] + 
                kernel_img_mul_143[21] + kernel_img_mul_143[22] + kernel_img_mul_143[23] + 
                kernel_img_mul_143[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1151:1144] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1151:1144] <= kernel_img_sum_143[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1151:1144] <= 'd0;
end

wire  [39:0]  kernel_img_mul_144[0:24];
assign kernel_img_mul_144[0] = buffer_data_4[1143:1136] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_144[1] = buffer_data_4[1151:1144] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_144[2] = buffer_data_4[1159:1152] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_144[3] = buffer_data_4[1167:1160] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_144[4] = buffer_data_4[1175:1168] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_144[5] = buffer_data_3[1143:1136] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_144[6] = buffer_data_3[1151:1144] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_144[7] = buffer_data_3[1159:1152] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_144[8] = buffer_data_3[1167:1160] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_144[9] = buffer_data_3[1175:1168] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_144[10] = buffer_data_2[1143:1136] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_144[11] = buffer_data_2[1151:1144] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_144[12] = buffer_data_2[1159:1152] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_144[13] = buffer_data_2[1167:1160] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_144[14] = buffer_data_2[1175:1168] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_144[15] = buffer_data_1[1143:1136] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_144[16] = buffer_data_1[1151:1144] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_144[17] = buffer_data_1[1159:1152] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_144[18] = buffer_data_1[1167:1160] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_144[19] = buffer_data_1[1175:1168] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_144[20] = buffer_data_0[1143:1136] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_144[21] = buffer_data_0[1151:1144] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_144[22] = buffer_data_0[1159:1152] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_144[23] = buffer_data_0[1167:1160] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_144[24] = buffer_data_0[1175:1168] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_144 = kernel_img_mul_144[0] + kernel_img_mul_144[1] + kernel_img_mul_144[2] + 
                kernel_img_mul_144[3] + kernel_img_mul_144[4] + kernel_img_mul_144[5] + 
                kernel_img_mul_144[6] + kernel_img_mul_144[7] + kernel_img_mul_144[8] + 
                kernel_img_mul_144[9] + kernel_img_mul_144[10] + kernel_img_mul_144[11] + 
                kernel_img_mul_144[12] + kernel_img_mul_144[13] + kernel_img_mul_144[14] + 
                kernel_img_mul_144[15] + kernel_img_mul_144[16] + kernel_img_mul_144[17] + 
                kernel_img_mul_144[18] + kernel_img_mul_144[19] + kernel_img_mul_144[20] + 
                kernel_img_mul_144[21] + kernel_img_mul_144[22] + kernel_img_mul_144[23] + 
                kernel_img_mul_144[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1159:1152] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1159:1152] <= kernel_img_sum_144[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1159:1152] <= 'd0;
end

wire  [39:0]  kernel_img_mul_145[0:24];
assign kernel_img_mul_145[0] = buffer_data_4[1151:1144] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_145[1] = buffer_data_4[1159:1152] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_145[2] = buffer_data_4[1167:1160] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_145[3] = buffer_data_4[1175:1168] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_145[4] = buffer_data_4[1183:1176] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_145[5] = buffer_data_3[1151:1144] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_145[6] = buffer_data_3[1159:1152] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_145[7] = buffer_data_3[1167:1160] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_145[8] = buffer_data_3[1175:1168] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_145[9] = buffer_data_3[1183:1176] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_145[10] = buffer_data_2[1151:1144] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_145[11] = buffer_data_2[1159:1152] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_145[12] = buffer_data_2[1167:1160] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_145[13] = buffer_data_2[1175:1168] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_145[14] = buffer_data_2[1183:1176] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_145[15] = buffer_data_1[1151:1144] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_145[16] = buffer_data_1[1159:1152] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_145[17] = buffer_data_1[1167:1160] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_145[18] = buffer_data_1[1175:1168] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_145[19] = buffer_data_1[1183:1176] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_145[20] = buffer_data_0[1151:1144] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_145[21] = buffer_data_0[1159:1152] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_145[22] = buffer_data_0[1167:1160] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_145[23] = buffer_data_0[1175:1168] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_145[24] = buffer_data_0[1183:1176] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_145 = kernel_img_mul_145[0] + kernel_img_mul_145[1] + kernel_img_mul_145[2] + 
                kernel_img_mul_145[3] + kernel_img_mul_145[4] + kernel_img_mul_145[5] + 
                kernel_img_mul_145[6] + kernel_img_mul_145[7] + kernel_img_mul_145[8] + 
                kernel_img_mul_145[9] + kernel_img_mul_145[10] + kernel_img_mul_145[11] + 
                kernel_img_mul_145[12] + kernel_img_mul_145[13] + kernel_img_mul_145[14] + 
                kernel_img_mul_145[15] + kernel_img_mul_145[16] + kernel_img_mul_145[17] + 
                kernel_img_mul_145[18] + kernel_img_mul_145[19] + kernel_img_mul_145[20] + 
                kernel_img_mul_145[21] + kernel_img_mul_145[22] + kernel_img_mul_145[23] + 
                kernel_img_mul_145[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1167:1160] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1167:1160] <= kernel_img_sum_145[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1167:1160] <= 'd0;
end

wire  [39:0]  kernel_img_mul_146[0:24];
assign kernel_img_mul_146[0] = buffer_data_4[1159:1152] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_146[1] = buffer_data_4[1167:1160] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_146[2] = buffer_data_4[1175:1168] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_146[3] = buffer_data_4[1183:1176] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_146[4] = buffer_data_4[1191:1184] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_146[5] = buffer_data_3[1159:1152] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_146[6] = buffer_data_3[1167:1160] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_146[7] = buffer_data_3[1175:1168] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_146[8] = buffer_data_3[1183:1176] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_146[9] = buffer_data_3[1191:1184] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_146[10] = buffer_data_2[1159:1152] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_146[11] = buffer_data_2[1167:1160] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_146[12] = buffer_data_2[1175:1168] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_146[13] = buffer_data_2[1183:1176] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_146[14] = buffer_data_2[1191:1184] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_146[15] = buffer_data_1[1159:1152] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_146[16] = buffer_data_1[1167:1160] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_146[17] = buffer_data_1[1175:1168] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_146[18] = buffer_data_1[1183:1176] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_146[19] = buffer_data_1[1191:1184] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_146[20] = buffer_data_0[1159:1152] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_146[21] = buffer_data_0[1167:1160] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_146[22] = buffer_data_0[1175:1168] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_146[23] = buffer_data_0[1183:1176] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_146[24] = buffer_data_0[1191:1184] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_146 = kernel_img_mul_146[0] + kernel_img_mul_146[1] + kernel_img_mul_146[2] + 
                kernel_img_mul_146[3] + kernel_img_mul_146[4] + kernel_img_mul_146[5] + 
                kernel_img_mul_146[6] + kernel_img_mul_146[7] + kernel_img_mul_146[8] + 
                kernel_img_mul_146[9] + kernel_img_mul_146[10] + kernel_img_mul_146[11] + 
                kernel_img_mul_146[12] + kernel_img_mul_146[13] + kernel_img_mul_146[14] + 
                kernel_img_mul_146[15] + kernel_img_mul_146[16] + kernel_img_mul_146[17] + 
                kernel_img_mul_146[18] + kernel_img_mul_146[19] + kernel_img_mul_146[20] + 
                kernel_img_mul_146[21] + kernel_img_mul_146[22] + kernel_img_mul_146[23] + 
                kernel_img_mul_146[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1175:1168] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1175:1168] <= kernel_img_sum_146[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1175:1168] <= 'd0;
end

wire  [39:0]  kernel_img_mul_147[0:24];
assign kernel_img_mul_147[0] = buffer_data_4[1167:1160] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_147[1] = buffer_data_4[1175:1168] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_147[2] = buffer_data_4[1183:1176] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_147[3] = buffer_data_4[1191:1184] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_147[4] = buffer_data_4[1199:1192] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_147[5] = buffer_data_3[1167:1160] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_147[6] = buffer_data_3[1175:1168] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_147[7] = buffer_data_3[1183:1176] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_147[8] = buffer_data_3[1191:1184] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_147[9] = buffer_data_3[1199:1192] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_147[10] = buffer_data_2[1167:1160] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_147[11] = buffer_data_2[1175:1168] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_147[12] = buffer_data_2[1183:1176] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_147[13] = buffer_data_2[1191:1184] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_147[14] = buffer_data_2[1199:1192] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_147[15] = buffer_data_1[1167:1160] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_147[16] = buffer_data_1[1175:1168] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_147[17] = buffer_data_1[1183:1176] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_147[18] = buffer_data_1[1191:1184] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_147[19] = buffer_data_1[1199:1192] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_147[20] = buffer_data_0[1167:1160] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_147[21] = buffer_data_0[1175:1168] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_147[22] = buffer_data_0[1183:1176] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_147[23] = buffer_data_0[1191:1184] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_147[24] = buffer_data_0[1199:1192] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_147 = kernel_img_mul_147[0] + kernel_img_mul_147[1] + kernel_img_mul_147[2] + 
                kernel_img_mul_147[3] + kernel_img_mul_147[4] + kernel_img_mul_147[5] + 
                kernel_img_mul_147[6] + kernel_img_mul_147[7] + kernel_img_mul_147[8] + 
                kernel_img_mul_147[9] + kernel_img_mul_147[10] + kernel_img_mul_147[11] + 
                kernel_img_mul_147[12] + kernel_img_mul_147[13] + kernel_img_mul_147[14] + 
                kernel_img_mul_147[15] + kernel_img_mul_147[16] + kernel_img_mul_147[17] + 
                kernel_img_mul_147[18] + kernel_img_mul_147[19] + kernel_img_mul_147[20] + 
                kernel_img_mul_147[21] + kernel_img_mul_147[22] + kernel_img_mul_147[23] + 
                kernel_img_mul_147[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1183:1176] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1183:1176] <= kernel_img_sum_147[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1183:1176] <= 'd0;
end

wire  [39:0]  kernel_img_mul_148[0:24];
assign kernel_img_mul_148[0] = buffer_data_4[1175:1168] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_148[1] = buffer_data_4[1183:1176] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_148[2] = buffer_data_4[1191:1184] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_148[3] = buffer_data_4[1199:1192] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_148[4] = buffer_data_4[1207:1200] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_148[5] = buffer_data_3[1175:1168] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_148[6] = buffer_data_3[1183:1176] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_148[7] = buffer_data_3[1191:1184] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_148[8] = buffer_data_3[1199:1192] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_148[9] = buffer_data_3[1207:1200] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_148[10] = buffer_data_2[1175:1168] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_148[11] = buffer_data_2[1183:1176] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_148[12] = buffer_data_2[1191:1184] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_148[13] = buffer_data_2[1199:1192] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_148[14] = buffer_data_2[1207:1200] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_148[15] = buffer_data_1[1175:1168] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_148[16] = buffer_data_1[1183:1176] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_148[17] = buffer_data_1[1191:1184] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_148[18] = buffer_data_1[1199:1192] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_148[19] = buffer_data_1[1207:1200] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_148[20] = buffer_data_0[1175:1168] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_148[21] = buffer_data_0[1183:1176] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_148[22] = buffer_data_0[1191:1184] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_148[23] = buffer_data_0[1199:1192] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_148[24] = buffer_data_0[1207:1200] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_148 = kernel_img_mul_148[0] + kernel_img_mul_148[1] + kernel_img_mul_148[2] + 
                kernel_img_mul_148[3] + kernel_img_mul_148[4] + kernel_img_mul_148[5] + 
                kernel_img_mul_148[6] + kernel_img_mul_148[7] + kernel_img_mul_148[8] + 
                kernel_img_mul_148[9] + kernel_img_mul_148[10] + kernel_img_mul_148[11] + 
                kernel_img_mul_148[12] + kernel_img_mul_148[13] + kernel_img_mul_148[14] + 
                kernel_img_mul_148[15] + kernel_img_mul_148[16] + kernel_img_mul_148[17] + 
                kernel_img_mul_148[18] + kernel_img_mul_148[19] + kernel_img_mul_148[20] + 
                kernel_img_mul_148[21] + kernel_img_mul_148[22] + kernel_img_mul_148[23] + 
                kernel_img_mul_148[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1191:1184] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1191:1184] <= kernel_img_sum_148[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1191:1184] <= 'd0;
end

wire  [39:0]  kernel_img_mul_149[0:24];
assign kernel_img_mul_149[0] = buffer_data_4[1183:1176] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_149[1] = buffer_data_4[1191:1184] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_149[2] = buffer_data_4[1199:1192] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_149[3] = buffer_data_4[1207:1200] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_149[4] = buffer_data_4[1215:1208] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_149[5] = buffer_data_3[1183:1176] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_149[6] = buffer_data_3[1191:1184] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_149[7] = buffer_data_3[1199:1192] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_149[8] = buffer_data_3[1207:1200] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_149[9] = buffer_data_3[1215:1208] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_149[10] = buffer_data_2[1183:1176] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_149[11] = buffer_data_2[1191:1184] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_149[12] = buffer_data_2[1199:1192] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_149[13] = buffer_data_2[1207:1200] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_149[14] = buffer_data_2[1215:1208] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_149[15] = buffer_data_1[1183:1176] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_149[16] = buffer_data_1[1191:1184] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_149[17] = buffer_data_1[1199:1192] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_149[18] = buffer_data_1[1207:1200] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_149[19] = buffer_data_1[1215:1208] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_149[20] = buffer_data_0[1183:1176] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_149[21] = buffer_data_0[1191:1184] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_149[22] = buffer_data_0[1199:1192] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_149[23] = buffer_data_0[1207:1200] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_149[24] = buffer_data_0[1215:1208] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_149 = kernel_img_mul_149[0] + kernel_img_mul_149[1] + kernel_img_mul_149[2] + 
                kernel_img_mul_149[3] + kernel_img_mul_149[4] + kernel_img_mul_149[5] + 
                kernel_img_mul_149[6] + kernel_img_mul_149[7] + kernel_img_mul_149[8] + 
                kernel_img_mul_149[9] + kernel_img_mul_149[10] + kernel_img_mul_149[11] + 
                kernel_img_mul_149[12] + kernel_img_mul_149[13] + kernel_img_mul_149[14] + 
                kernel_img_mul_149[15] + kernel_img_mul_149[16] + kernel_img_mul_149[17] + 
                kernel_img_mul_149[18] + kernel_img_mul_149[19] + kernel_img_mul_149[20] + 
                kernel_img_mul_149[21] + kernel_img_mul_149[22] + kernel_img_mul_149[23] + 
                kernel_img_mul_149[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1199:1192] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1199:1192] <= kernel_img_sum_149[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1199:1192] <= 'd0;
end

wire  [39:0]  kernel_img_mul_150[0:24];
assign kernel_img_mul_150[0] = buffer_data_4[1191:1184] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_150[1] = buffer_data_4[1199:1192] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_150[2] = buffer_data_4[1207:1200] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_150[3] = buffer_data_4[1215:1208] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_150[4] = buffer_data_4[1223:1216] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_150[5] = buffer_data_3[1191:1184] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_150[6] = buffer_data_3[1199:1192] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_150[7] = buffer_data_3[1207:1200] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_150[8] = buffer_data_3[1215:1208] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_150[9] = buffer_data_3[1223:1216] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_150[10] = buffer_data_2[1191:1184] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_150[11] = buffer_data_2[1199:1192] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_150[12] = buffer_data_2[1207:1200] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_150[13] = buffer_data_2[1215:1208] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_150[14] = buffer_data_2[1223:1216] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_150[15] = buffer_data_1[1191:1184] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_150[16] = buffer_data_1[1199:1192] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_150[17] = buffer_data_1[1207:1200] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_150[18] = buffer_data_1[1215:1208] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_150[19] = buffer_data_1[1223:1216] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_150[20] = buffer_data_0[1191:1184] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_150[21] = buffer_data_0[1199:1192] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_150[22] = buffer_data_0[1207:1200] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_150[23] = buffer_data_0[1215:1208] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_150[24] = buffer_data_0[1223:1216] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_150 = kernel_img_mul_150[0] + kernel_img_mul_150[1] + kernel_img_mul_150[2] + 
                kernel_img_mul_150[3] + kernel_img_mul_150[4] + kernel_img_mul_150[5] + 
                kernel_img_mul_150[6] + kernel_img_mul_150[7] + kernel_img_mul_150[8] + 
                kernel_img_mul_150[9] + kernel_img_mul_150[10] + kernel_img_mul_150[11] + 
                kernel_img_mul_150[12] + kernel_img_mul_150[13] + kernel_img_mul_150[14] + 
                kernel_img_mul_150[15] + kernel_img_mul_150[16] + kernel_img_mul_150[17] + 
                kernel_img_mul_150[18] + kernel_img_mul_150[19] + kernel_img_mul_150[20] + 
                kernel_img_mul_150[21] + kernel_img_mul_150[22] + kernel_img_mul_150[23] + 
                kernel_img_mul_150[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1207:1200] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1207:1200] <= kernel_img_sum_150[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1207:1200] <= 'd0;
end

wire  [39:0]  kernel_img_mul_151[0:24];
assign kernel_img_mul_151[0] = buffer_data_4[1199:1192] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_151[1] = buffer_data_4[1207:1200] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_151[2] = buffer_data_4[1215:1208] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_151[3] = buffer_data_4[1223:1216] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_151[4] = buffer_data_4[1231:1224] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_151[5] = buffer_data_3[1199:1192] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_151[6] = buffer_data_3[1207:1200] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_151[7] = buffer_data_3[1215:1208] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_151[8] = buffer_data_3[1223:1216] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_151[9] = buffer_data_3[1231:1224] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_151[10] = buffer_data_2[1199:1192] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_151[11] = buffer_data_2[1207:1200] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_151[12] = buffer_data_2[1215:1208] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_151[13] = buffer_data_2[1223:1216] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_151[14] = buffer_data_2[1231:1224] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_151[15] = buffer_data_1[1199:1192] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_151[16] = buffer_data_1[1207:1200] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_151[17] = buffer_data_1[1215:1208] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_151[18] = buffer_data_1[1223:1216] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_151[19] = buffer_data_1[1231:1224] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_151[20] = buffer_data_0[1199:1192] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_151[21] = buffer_data_0[1207:1200] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_151[22] = buffer_data_0[1215:1208] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_151[23] = buffer_data_0[1223:1216] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_151[24] = buffer_data_0[1231:1224] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_151 = kernel_img_mul_151[0] + kernel_img_mul_151[1] + kernel_img_mul_151[2] + 
                kernel_img_mul_151[3] + kernel_img_mul_151[4] + kernel_img_mul_151[5] + 
                kernel_img_mul_151[6] + kernel_img_mul_151[7] + kernel_img_mul_151[8] + 
                kernel_img_mul_151[9] + kernel_img_mul_151[10] + kernel_img_mul_151[11] + 
                kernel_img_mul_151[12] + kernel_img_mul_151[13] + kernel_img_mul_151[14] + 
                kernel_img_mul_151[15] + kernel_img_mul_151[16] + kernel_img_mul_151[17] + 
                kernel_img_mul_151[18] + kernel_img_mul_151[19] + kernel_img_mul_151[20] + 
                kernel_img_mul_151[21] + kernel_img_mul_151[22] + kernel_img_mul_151[23] + 
                kernel_img_mul_151[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1215:1208] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1215:1208] <= kernel_img_sum_151[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1215:1208] <= 'd0;
end

wire  [39:0]  kernel_img_mul_152[0:24];
assign kernel_img_mul_152[0] = buffer_data_4[1207:1200] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_152[1] = buffer_data_4[1215:1208] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_152[2] = buffer_data_4[1223:1216] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_152[3] = buffer_data_4[1231:1224] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_152[4] = buffer_data_4[1239:1232] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_152[5] = buffer_data_3[1207:1200] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_152[6] = buffer_data_3[1215:1208] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_152[7] = buffer_data_3[1223:1216] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_152[8] = buffer_data_3[1231:1224] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_152[9] = buffer_data_3[1239:1232] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_152[10] = buffer_data_2[1207:1200] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_152[11] = buffer_data_2[1215:1208] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_152[12] = buffer_data_2[1223:1216] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_152[13] = buffer_data_2[1231:1224] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_152[14] = buffer_data_2[1239:1232] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_152[15] = buffer_data_1[1207:1200] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_152[16] = buffer_data_1[1215:1208] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_152[17] = buffer_data_1[1223:1216] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_152[18] = buffer_data_1[1231:1224] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_152[19] = buffer_data_1[1239:1232] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_152[20] = buffer_data_0[1207:1200] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_152[21] = buffer_data_0[1215:1208] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_152[22] = buffer_data_0[1223:1216] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_152[23] = buffer_data_0[1231:1224] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_152[24] = buffer_data_0[1239:1232] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_152 = kernel_img_mul_152[0] + kernel_img_mul_152[1] + kernel_img_mul_152[2] + 
                kernel_img_mul_152[3] + kernel_img_mul_152[4] + kernel_img_mul_152[5] + 
                kernel_img_mul_152[6] + kernel_img_mul_152[7] + kernel_img_mul_152[8] + 
                kernel_img_mul_152[9] + kernel_img_mul_152[10] + kernel_img_mul_152[11] + 
                kernel_img_mul_152[12] + kernel_img_mul_152[13] + kernel_img_mul_152[14] + 
                kernel_img_mul_152[15] + kernel_img_mul_152[16] + kernel_img_mul_152[17] + 
                kernel_img_mul_152[18] + kernel_img_mul_152[19] + kernel_img_mul_152[20] + 
                kernel_img_mul_152[21] + kernel_img_mul_152[22] + kernel_img_mul_152[23] + 
                kernel_img_mul_152[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1223:1216] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1223:1216] <= kernel_img_sum_152[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1223:1216] <= 'd0;
end

wire  [39:0]  kernel_img_mul_153[0:24];
assign kernel_img_mul_153[0] = buffer_data_4[1215:1208] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_153[1] = buffer_data_4[1223:1216] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_153[2] = buffer_data_4[1231:1224] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_153[3] = buffer_data_4[1239:1232] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_153[4] = buffer_data_4[1247:1240] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_153[5] = buffer_data_3[1215:1208] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_153[6] = buffer_data_3[1223:1216] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_153[7] = buffer_data_3[1231:1224] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_153[8] = buffer_data_3[1239:1232] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_153[9] = buffer_data_3[1247:1240] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_153[10] = buffer_data_2[1215:1208] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_153[11] = buffer_data_2[1223:1216] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_153[12] = buffer_data_2[1231:1224] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_153[13] = buffer_data_2[1239:1232] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_153[14] = buffer_data_2[1247:1240] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_153[15] = buffer_data_1[1215:1208] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_153[16] = buffer_data_1[1223:1216] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_153[17] = buffer_data_1[1231:1224] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_153[18] = buffer_data_1[1239:1232] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_153[19] = buffer_data_1[1247:1240] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_153[20] = buffer_data_0[1215:1208] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_153[21] = buffer_data_0[1223:1216] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_153[22] = buffer_data_0[1231:1224] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_153[23] = buffer_data_0[1239:1232] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_153[24] = buffer_data_0[1247:1240] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_153 = kernel_img_mul_153[0] + kernel_img_mul_153[1] + kernel_img_mul_153[2] + 
                kernel_img_mul_153[3] + kernel_img_mul_153[4] + kernel_img_mul_153[5] + 
                kernel_img_mul_153[6] + kernel_img_mul_153[7] + kernel_img_mul_153[8] + 
                kernel_img_mul_153[9] + kernel_img_mul_153[10] + kernel_img_mul_153[11] + 
                kernel_img_mul_153[12] + kernel_img_mul_153[13] + kernel_img_mul_153[14] + 
                kernel_img_mul_153[15] + kernel_img_mul_153[16] + kernel_img_mul_153[17] + 
                kernel_img_mul_153[18] + kernel_img_mul_153[19] + kernel_img_mul_153[20] + 
                kernel_img_mul_153[21] + kernel_img_mul_153[22] + kernel_img_mul_153[23] + 
                kernel_img_mul_153[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1231:1224] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1231:1224] <= kernel_img_sum_153[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1231:1224] <= 'd0;
end

wire  [39:0]  kernel_img_mul_154[0:24];
assign kernel_img_mul_154[0] = buffer_data_4[1223:1216] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_154[1] = buffer_data_4[1231:1224] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_154[2] = buffer_data_4[1239:1232] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_154[3] = buffer_data_4[1247:1240] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_154[4] = buffer_data_4[1255:1248] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_154[5] = buffer_data_3[1223:1216] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_154[6] = buffer_data_3[1231:1224] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_154[7] = buffer_data_3[1239:1232] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_154[8] = buffer_data_3[1247:1240] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_154[9] = buffer_data_3[1255:1248] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_154[10] = buffer_data_2[1223:1216] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_154[11] = buffer_data_2[1231:1224] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_154[12] = buffer_data_2[1239:1232] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_154[13] = buffer_data_2[1247:1240] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_154[14] = buffer_data_2[1255:1248] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_154[15] = buffer_data_1[1223:1216] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_154[16] = buffer_data_1[1231:1224] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_154[17] = buffer_data_1[1239:1232] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_154[18] = buffer_data_1[1247:1240] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_154[19] = buffer_data_1[1255:1248] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_154[20] = buffer_data_0[1223:1216] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_154[21] = buffer_data_0[1231:1224] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_154[22] = buffer_data_0[1239:1232] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_154[23] = buffer_data_0[1247:1240] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_154[24] = buffer_data_0[1255:1248] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_154 = kernel_img_mul_154[0] + kernel_img_mul_154[1] + kernel_img_mul_154[2] + 
                kernel_img_mul_154[3] + kernel_img_mul_154[4] + kernel_img_mul_154[5] + 
                kernel_img_mul_154[6] + kernel_img_mul_154[7] + kernel_img_mul_154[8] + 
                kernel_img_mul_154[9] + kernel_img_mul_154[10] + kernel_img_mul_154[11] + 
                kernel_img_mul_154[12] + kernel_img_mul_154[13] + kernel_img_mul_154[14] + 
                kernel_img_mul_154[15] + kernel_img_mul_154[16] + kernel_img_mul_154[17] + 
                kernel_img_mul_154[18] + kernel_img_mul_154[19] + kernel_img_mul_154[20] + 
                kernel_img_mul_154[21] + kernel_img_mul_154[22] + kernel_img_mul_154[23] + 
                kernel_img_mul_154[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1239:1232] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1239:1232] <= kernel_img_sum_154[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1239:1232] <= 'd0;
end

wire  [39:0]  kernel_img_mul_155[0:24];
assign kernel_img_mul_155[0] = buffer_data_4[1231:1224] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_155[1] = buffer_data_4[1239:1232] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_155[2] = buffer_data_4[1247:1240] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_155[3] = buffer_data_4[1255:1248] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_155[4] = buffer_data_4[1263:1256] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_155[5] = buffer_data_3[1231:1224] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_155[6] = buffer_data_3[1239:1232] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_155[7] = buffer_data_3[1247:1240] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_155[8] = buffer_data_3[1255:1248] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_155[9] = buffer_data_3[1263:1256] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_155[10] = buffer_data_2[1231:1224] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_155[11] = buffer_data_2[1239:1232] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_155[12] = buffer_data_2[1247:1240] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_155[13] = buffer_data_2[1255:1248] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_155[14] = buffer_data_2[1263:1256] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_155[15] = buffer_data_1[1231:1224] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_155[16] = buffer_data_1[1239:1232] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_155[17] = buffer_data_1[1247:1240] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_155[18] = buffer_data_1[1255:1248] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_155[19] = buffer_data_1[1263:1256] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_155[20] = buffer_data_0[1231:1224] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_155[21] = buffer_data_0[1239:1232] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_155[22] = buffer_data_0[1247:1240] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_155[23] = buffer_data_0[1255:1248] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_155[24] = buffer_data_0[1263:1256] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_155 = kernel_img_mul_155[0] + kernel_img_mul_155[1] + kernel_img_mul_155[2] + 
                kernel_img_mul_155[3] + kernel_img_mul_155[4] + kernel_img_mul_155[5] + 
                kernel_img_mul_155[6] + kernel_img_mul_155[7] + kernel_img_mul_155[8] + 
                kernel_img_mul_155[9] + kernel_img_mul_155[10] + kernel_img_mul_155[11] + 
                kernel_img_mul_155[12] + kernel_img_mul_155[13] + kernel_img_mul_155[14] + 
                kernel_img_mul_155[15] + kernel_img_mul_155[16] + kernel_img_mul_155[17] + 
                kernel_img_mul_155[18] + kernel_img_mul_155[19] + kernel_img_mul_155[20] + 
                kernel_img_mul_155[21] + kernel_img_mul_155[22] + kernel_img_mul_155[23] + 
                kernel_img_mul_155[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1247:1240] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1247:1240] <= kernel_img_sum_155[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1247:1240] <= 'd0;
end

wire  [39:0]  kernel_img_mul_156[0:24];
assign kernel_img_mul_156[0] = buffer_data_4[1239:1232] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_156[1] = buffer_data_4[1247:1240] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_156[2] = buffer_data_4[1255:1248] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_156[3] = buffer_data_4[1263:1256] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_156[4] = buffer_data_4[1271:1264] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_156[5] = buffer_data_3[1239:1232] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_156[6] = buffer_data_3[1247:1240] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_156[7] = buffer_data_3[1255:1248] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_156[8] = buffer_data_3[1263:1256] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_156[9] = buffer_data_3[1271:1264] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_156[10] = buffer_data_2[1239:1232] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_156[11] = buffer_data_2[1247:1240] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_156[12] = buffer_data_2[1255:1248] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_156[13] = buffer_data_2[1263:1256] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_156[14] = buffer_data_2[1271:1264] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_156[15] = buffer_data_1[1239:1232] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_156[16] = buffer_data_1[1247:1240] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_156[17] = buffer_data_1[1255:1248] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_156[18] = buffer_data_1[1263:1256] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_156[19] = buffer_data_1[1271:1264] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_156[20] = buffer_data_0[1239:1232] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_156[21] = buffer_data_0[1247:1240] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_156[22] = buffer_data_0[1255:1248] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_156[23] = buffer_data_0[1263:1256] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_156[24] = buffer_data_0[1271:1264] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_156 = kernel_img_mul_156[0] + kernel_img_mul_156[1] + kernel_img_mul_156[2] + 
                kernel_img_mul_156[3] + kernel_img_mul_156[4] + kernel_img_mul_156[5] + 
                kernel_img_mul_156[6] + kernel_img_mul_156[7] + kernel_img_mul_156[8] + 
                kernel_img_mul_156[9] + kernel_img_mul_156[10] + kernel_img_mul_156[11] + 
                kernel_img_mul_156[12] + kernel_img_mul_156[13] + kernel_img_mul_156[14] + 
                kernel_img_mul_156[15] + kernel_img_mul_156[16] + kernel_img_mul_156[17] + 
                kernel_img_mul_156[18] + kernel_img_mul_156[19] + kernel_img_mul_156[20] + 
                kernel_img_mul_156[21] + kernel_img_mul_156[22] + kernel_img_mul_156[23] + 
                kernel_img_mul_156[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1255:1248] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1255:1248] <= kernel_img_sum_156[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1255:1248] <= 'd0;
end

wire  [39:0]  kernel_img_mul_157[0:24];
assign kernel_img_mul_157[0] = buffer_data_4[1247:1240] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_157[1] = buffer_data_4[1255:1248] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_157[2] = buffer_data_4[1263:1256] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_157[3] = buffer_data_4[1271:1264] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_157[4] = buffer_data_4[1279:1272] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_157[5] = buffer_data_3[1247:1240] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_157[6] = buffer_data_3[1255:1248] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_157[7] = buffer_data_3[1263:1256] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_157[8] = buffer_data_3[1271:1264] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_157[9] = buffer_data_3[1279:1272] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_157[10] = buffer_data_2[1247:1240] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_157[11] = buffer_data_2[1255:1248] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_157[12] = buffer_data_2[1263:1256] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_157[13] = buffer_data_2[1271:1264] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_157[14] = buffer_data_2[1279:1272] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_157[15] = buffer_data_1[1247:1240] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_157[16] = buffer_data_1[1255:1248] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_157[17] = buffer_data_1[1263:1256] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_157[18] = buffer_data_1[1271:1264] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_157[19] = buffer_data_1[1279:1272] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_157[20] = buffer_data_0[1247:1240] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_157[21] = buffer_data_0[1255:1248] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_157[22] = buffer_data_0[1263:1256] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_157[23] = buffer_data_0[1271:1264] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_157[24] = buffer_data_0[1279:1272] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_157 = kernel_img_mul_157[0] + kernel_img_mul_157[1] + kernel_img_mul_157[2] + 
                kernel_img_mul_157[3] + kernel_img_mul_157[4] + kernel_img_mul_157[5] + 
                kernel_img_mul_157[6] + kernel_img_mul_157[7] + kernel_img_mul_157[8] + 
                kernel_img_mul_157[9] + kernel_img_mul_157[10] + kernel_img_mul_157[11] + 
                kernel_img_mul_157[12] + kernel_img_mul_157[13] + kernel_img_mul_157[14] + 
                kernel_img_mul_157[15] + kernel_img_mul_157[16] + kernel_img_mul_157[17] + 
                kernel_img_mul_157[18] + kernel_img_mul_157[19] + kernel_img_mul_157[20] + 
                kernel_img_mul_157[21] + kernel_img_mul_157[22] + kernel_img_mul_157[23] + 
                kernel_img_mul_157[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1263:1256] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1263:1256] <= kernel_img_sum_157[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1263:1256] <= 'd0;
end

wire  [39:0]  kernel_img_mul_158[0:24];
assign kernel_img_mul_158[0] = buffer_data_4[1255:1248] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_158[1] = buffer_data_4[1263:1256] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_158[2] = buffer_data_4[1271:1264] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_158[3] = buffer_data_4[1279:1272] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_158[4] = buffer_data_4[1287:1280] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_158[5] = buffer_data_3[1255:1248] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_158[6] = buffer_data_3[1263:1256] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_158[7] = buffer_data_3[1271:1264] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_158[8] = buffer_data_3[1279:1272] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_158[9] = buffer_data_3[1287:1280] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_158[10] = buffer_data_2[1255:1248] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_158[11] = buffer_data_2[1263:1256] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_158[12] = buffer_data_2[1271:1264] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_158[13] = buffer_data_2[1279:1272] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_158[14] = buffer_data_2[1287:1280] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_158[15] = buffer_data_1[1255:1248] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_158[16] = buffer_data_1[1263:1256] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_158[17] = buffer_data_1[1271:1264] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_158[18] = buffer_data_1[1279:1272] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_158[19] = buffer_data_1[1287:1280] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_158[20] = buffer_data_0[1255:1248] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_158[21] = buffer_data_0[1263:1256] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_158[22] = buffer_data_0[1271:1264] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_158[23] = buffer_data_0[1279:1272] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_158[24] = buffer_data_0[1287:1280] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_158 = kernel_img_mul_158[0] + kernel_img_mul_158[1] + kernel_img_mul_158[2] + 
                kernel_img_mul_158[3] + kernel_img_mul_158[4] + kernel_img_mul_158[5] + 
                kernel_img_mul_158[6] + kernel_img_mul_158[7] + kernel_img_mul_158[8] + 
                kernel_img_mul_158[9] + kernel_img_mul_158[10] + kernel_img_mul_158[11] + 
                kernel_img_mul_158[12] + kernel_img_mul_158[13] + kernel_img_mul_158[14] + 
                kernel_img_mul_158[15] + kernel_img_mul_158[16] + kernel_img_mul_158[17] + 
                kernel_img_mul_158[18] + kernel_img_mul_158[19] + kernel_img_mul_158[20] + 
                kernel_img_mul_158[21] + kernel_img_mul_158[22] + kernel_img_mul_158[23] + 
                kernel_img_mul_158[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1271:1264] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1271:1264] <= kernel_img_sum_158[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1271:1264] <= 'd0;
end

wire  [39:0]  kernel_img_mul_159[0:24];
assign kernel_img_mul_159[0] = buffer_data_4[1263:1256] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_159[1] = buffer_data_4[1271:1264] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_159[2] = buffer_data_4[1279:1272] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_159[3] = buffer_data_4[1287:1280] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_159[4] = buffer_data_4[1295:1288] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_159[5] = buffer_data_3[1263:1256] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_159[6] = buffer_data_3[1271:1264] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_159[7] = buffer_data_3[1279:1272] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_159[8] = buffer_data_3[1287:1280] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_159[9] = buffer_data_3[1295:1288] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_159[10] = buffer_data_2[1263:1256] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_159[11] = buffer_data_2[1271:1264] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_159[12] = buffer_data_2[1279:1272] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_159[13] = buffer_data_2[1287:1280] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_159[14] = buffer_data_2[1295:1288] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_159[15] = buffer_data_1[1263:1256] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_159[16] = buffer_data_1[1271:1264] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_159[17] = buffer_data_1[1279:1272] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_159[18] = buffer_data_1[1287:1280] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_159[19] = buffer_data_1[1295:1288] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_159[20] = buffer_data_0[1263:1256] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_159[21] = buffer_data_0[1271:1264] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_159[22] = buffer_data_0[1279:1272] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_159[23] = buffer_data_0[1287:1280] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_159[24] = buffer_data_0[1295:1288] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_159 = kernel_img_mul_159[0] + kernel_img_mul_159[1] + kernel_img_mul_159[2] + 
                kernel_img_mul_159[3] + kernel_img_mul_159[4] + kernel_img_mul_159[5] + 
                kernel_img_mul_159[6] + kernel_img_mul_159[7] + kernel_img_mul_159[8] + 
                kernel_img_mul_159[9] + kernel_img_mul_159[10] + kernel_img_mul_159[11] + 
                kernel_img_mul_159[12] + kernel_img_mul_159[13] + kernel_img_mul_159[14] + 
                kernel_img_mul_159[15] + kernel_img_mul_159[16] + kernel_img_mul_159[17] + 
                kernel_img_mul_159[18] + kernel_img_mul_159[19] + kernel_img_mul_159[20] + 
                kernel_img_mul_159[21] + kernel_img_mul_159[22] + kernel_img_mul_159[23] + 
                kernel_img_mul_159[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1279:1272] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1279:1272] <= kernel_img_sum_159[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1279:1272] <= 'd0;
end

wire  [39:0]  kernel_img_mul_160[0:24];
assign kernel_img_mul_160[0] = buffer_data_4[1271:1264] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_160[1] = buffer_data_4[1279:1272] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_160[2] = buffer_data_4[1287:1280] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_160[3] = buffer_data_4[1295:1288] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_160[4] = buffer_data_4[1303:1296] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_160[5] = buffer_data_3[1271:1264] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_160[6] = buffer_data_3[1279:1272] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_160[7] = buffer_data_3[1287:1280] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_160[8] = buffer_data_3[1295:1288] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_160[9] = buffer_data_3[1303:1296] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_160[10] = buffer_data_2[1271:1264] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_160[11] = buffer_data_2[1279:1272] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_160[12] = buffer_data_2[1287:1280] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_160[13] = buffer_data_2[1295:1288] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_160[14] = buffer_data_2[1303:1296] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_160[15] = buffer_data_1[1271:1264] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_160[16] = buffer_data_1[1279:1272] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_160[17] = buffer_data_1[1287:1280] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_160[18] = buffer_data_1[1295:1288] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_160[19] = buffer_data_1[1303:1296] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_160[20] = buffer_data_0[1271:1264] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_160[21] = buffer_data_0[1279:1272] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_160[22] = buffer_data_0[1287:1280] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_160[23] = buffer_data_0[1295:1288] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_160[24] = buffer_data_0[1303:1296] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_160 = kernel_img_mul_160[0] + kernel_img_mul_160[1] + kernel_img_mul_160[2] + 
                kernel_img_mul_160[3] + kernel_img_mul_160[4] + kernel_img_mul_160[5] + 
                kernel_img_mul_160[6] + kernel_img_mul_160[7] + kernel_img_mul_160[8] + 
                kernel_img_mul_160[9] + kernel_img_mul_160[10] + kernel_img_mul_160[11] + 
                kernel_img_mul_160[12] + kernel_img_mul_160[13] + kernel_img_mul_160[14] + 
                kernel_img_mul_160[15] + kernel_img_mul_160[16] + kernel_img_mul_160[17] + 
                kernel_img_mul_160[18] + kernel_img_mul_160[19] + kernel_img_mul_160[20] + 
                kernel_img_mul_160[21] + kernel_img_mul_160[22] + kernel_img_mul_160[23] + 
                kernel_img_mul_160[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1287:1280] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1287:1280] <= kernel_img_sum_160[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1287:1280] <= 'd0;
end

wire  [39:0]  kernel_img_mul_161[0:24];
assign kernel_img_mul_161[0] = buffer_data_4[1279:1272] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_161[1] = buffer_data_4[1287:1280] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_161[2] = buffer_data_4[1295:1288] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_161[3] = buffer_data_4[1303:1296] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_161[4] = buffer_data_4[1311:1304] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_161[5] = buffer_data_3[1279:1272] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_161[6] = buffer_data_3[1287:1280] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_161[7] = buffer_data_3[1295:1288] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_161[8] = buffer_data_3[1303:1296] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_161[9] = buffer_data_3[1311:1304] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_161[10] = buffer_data_2[1279:1272] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_161[11] = buffer_data_2[1287:1280] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_161[12] = buffer_data_2[1295:1288] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_161[13] = buffer_data_2[1303:1296] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_161[14] = buffer_data_2[1311:1304] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_161[15] = buffer_data_1[1279:1272] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_161[16] = buffer_data_1[1287:1280] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_161[17] = buffer_data_1[1295:1288] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_161[18] = buffer_data_1[1303:1296] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_161[19] = buffer_data_1[1311:1304] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_161[20] = buffer_data_0[1279:1272] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_161[21] = buffer_data_0[1287:1280] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_161[22] = buffer_data_0[1295:1288] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_161[23] = buffer_data_0[1303:1296] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_161[24] = buffer_data_0[1311:1304] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_161 = kernel_img_mul_161[0] + kernel_img_mul_161[1] + kernel_img_mul_161[2] + 
                kernel_img_mul_161[3] + kernel_img_mul_161[4] + kernel_img_mul_161[5] + 
                kernel_img_mul_161[6] + kernel_img_mul_161[7] + kernel_img_mul_161[8] + 
                kernel_img_mul_161[9] + kernel_img_mul_161[10] + kernel_img_mul_161[11] + 
                kernel_img_mul_161[12] + kernel_img_mul_161[13] + kernel_img_mul_161[14] + 
                kernel_img_mul_161[15] + kernel_img_mul_161[16] + kernel_img_mul_161[17] + 
                kernel_img_mul_161[18] + kernel_img_mul_161[19] + kernel_img_mul_161[20] + 
                kernel_img_mul_161[21] + kernel_img_mul_161[22] + kernel_img_mul_161[23] + 
                kernel_img_mul_161[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1295:1288] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1295:1288] <= kernel_img_sum_161[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1295:1288] <= 'd0;
end

wire  [39:0]  kernel_img_mul_162[0:24];
assign kernel_img_mul_162[0] = buffer_data_4[1287:1280] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_162[1] = buffer_data_4[1295:1288] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_162[2] = buffer_data_4[1303:1296] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_162[3] = buffer_data_4[1311:1304] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_162[4] = buffer_data_4[1319:1312] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_162[5] = buffer_data_3[1287:1280] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_162[6] = buffer_data_3[1295:1288] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_162[7] = buffer_data_3[1303:1296] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_162[8] = buffer_data_3[1311:1304] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_162[9] = buffer_data_3[1319:1312] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_162[10] = buffer_data_2[1287:1280] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_162[11] = buffer_data_2[1295:1288] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_162[12] = buffer_data_2[1303:1296] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_162[13] = buffer_data_2[1311:1304] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_162[14] = buffer_data_2[1319:1312] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_162[15] = buffer_data_1[1287:1280] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_162[16] = buffer_data_1[1295:1288] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_162[17] = buffer_data_1[1303:1296] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_162[18] = buffer_data_1[1311:1304] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_162[19] = buffer_data_1[1319:1312] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_162[20] = buffer_data_0[1287:1280] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_162[21] = buffer_data_0[1295:1288] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_162[22] = buffer_data_0[1303:1296] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_162[23] = buffer_data_0[1311:1304] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_162[24] = buffer_data_0[1319:1312] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_162 = kernel_img_mul_162[0] + kernel_img_mul_162[1] + kernel_img_mul_162[2] + 
                kernel_img_mul_162[3] + kernel_img_mul_162[4] + kernel_img_mul_162[5] + 
                kernel_img_mul_162[6] + kernel_img_mul_162[7] + kernel_img_mul_162[8] + 
                kernel_img_mul_162[9] + kernel_img_mul_162[10] + kernel_img_mul_162[11] + 
                kernel_img_mul_162[12] + kernel_img_mul_162[13] + kernel_img_mul_162[14] + 
                kernel_img_mul_162[15] + kernel_img_mul_162[16] + kernel_img_mul_162[17] + 
                kernel_img_mul_162[18] + kernel_img_mul_162[19] + kernel_img_mul_162[20] + 
                kernel_img_mul_162[21] + kernel_img_mul_162[22] + kernel_img_mul_162[23] + 
                kernel_img_mul_162[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1303:1296] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1303:1296] <= kernel_img_sum_162[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1303:1296] <= 'd0;
end

wire  [39:0]  kernel_img_mul_163[0:24];
assign kernel_img_mul_163[0] = buffer_data_4[1295:1288] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_163[1] = buffer_data_4[1303:1296] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_163[2] = buffer_data_4[1311:1304] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_163[3] = buffer_data_4[1319:1312] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_163[4] = buffer_data_4[1327:1320] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_163[5] = buffer_data_3[1295:1288] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_163[6] = buffer_data_3[1303:1296] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_163[7] = buffer_data_3[1311:1304] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_163[8] = buffer_data_3[1319:1312] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_163[9] = buffer_data_3[1327:1320] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_163[10] = buffer_data_2[1295:1288] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_163[11] = buffer_data_2[1303:1296] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_163[12] = buffer_data_2[1311:1304] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_163[13] = buffer_data_2[1319:1312] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_163[14] = buffer_data_2[1327:1320] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_163[15] = buffer_data_1[1295:1288] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_163[16] = buffer_data_1[1303:1296] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_163[17] = buffer_data_1[1311:1304] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_163[18] = buffer_data_1[1319:1312] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_163[19] = buffer_data_1[1327:1320] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_163[20] = buffer_data_0[1295:1288] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_163[21] = buffer_data_0[1303:1296] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_163[22] = buffer_data_0[1311:1304] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_163[23] = buffer_data_0[1319:1312] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_163[24] = buffer_data_0[1327:1320] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_163 = kernel_img_mul_163[0] + kernel_img_mul_163[1] + kernel_img_mul_163[2] + 
                kernel_img_mul_163[3] + kernel_img_mul_163[4] + kernel_img_mul_163[5] + 
                kernel_img_mul_163[6] + kernel_img_mul_163[7] + kernel_img_mul_163[8] + 
                kernel_img_mul_163[9] + kernel_img_mul_163[10] + kernel_img_mul_163[11] + 
                kernel_img_mul_163[12] + kernel_img_mul_163[13] + kernel_img_mul_163[14] + 
                kernel_img_mul_163[15] + kernel_img_mul_163[16] + kernel_img_mul_163[17] + 
                kernel_img_mul_163[18] + kernel_img_mul_163[19] + kernel_img_mul_163[20] + 
                kernel_img_mul_163[21] + kernel_img_mul_163[22] + kernel_img_mul_163[23] + 
                kernel_img_mul_163[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1311:1304] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1311:1304] <= kernel_img_sum_163[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1311:1304] <= 'd0;
end

wire  [39:0]  kernel_img_mul_164[0:24];
assign kernel_img_mul_164[0] = buffer_data_4[1303:1296] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_164[1] = buffer_data_4[1311:1304] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_164[2] = buffer_data_4[1319:1312] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_164[3] = buffer_data_4[1327:1320] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_164[4] = buffer_data_4[1335:1328] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_164[5] = buffer_data_3[1303:1296] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_164[6] = buffer_data_3[1311:1304] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_164[7] = buffer_data_3[1319:1312] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_164[8] = buffer_data_3[1327:1320] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_164[9] = buffer_data_3[1335:1328] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_164[10] = buffer_data_2[1303:1296] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_164[11] = buffer_data_2[1311:1304] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_164[12] = buffer_data_2[1319:1312] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_164[13] = buffer_data_2[1327:1320] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_164[14] = buffer_data_2[1335:1328] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_164[15] = buffer_data_1[1303:1296] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_164[16] = buffer_data_1[1311:1304] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_164[17] = buffer_data_1[1319:1312] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_164[18] = buffer_data_1[1327:1320] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_164[19] = buffer_data_1[1335:1328] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_164[20] = buffer_data_0[1303:1296] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_164[21] = buffer_data_0[1311:1304] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_164[22] = buffer_data_0[1319:1312] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_164[23] = buffer_data_0[1327:1320] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_164[24] = buffer_data_0[1335:1328] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_164 = kernel_img_mul_164[0] + kernel_img_mul_164[1] + kernel_img_mul_164[2] + 
                kernel_img_mul_164[3] + kernel_img_mul_164[4] + kernel_img_mul_164[5] + 
                kernel_img_mul_164[6] + kernel_img_mul_164[7] + kernel_img_mul_164[8] + 
                kernel_img_mul_164[9] + kernel_img_mul_164[10] + kernel_img_mul_164[11] + 
                kernel_img_mul_164[12] + kernel_img_mul_164[13] + kernel_img_mul_164[14] + 
                kernel_img_mul_164[15] + kernel_img_mul_164[16] + kernel_img_mul_164[17] + 
                kernel_img_mul_164[18] + kernel_img_mul_164[19] + kernel_img_mul_164[20] + 
                kernel_img_mul_164[21] + kernel_img_mul_164[22] + kernel_img_mul_164[23] + 
                kernel_img_mul_164[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1319:1312] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1319:1312] <= kernel_img_sum_164[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1319:1312] <= 'd0;
end

wire  [39:0]  kernel_img_mul_165[0:24];
assign kernel_img_mul_165[0] = buffer_data_4[1311:1304] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_165[1] = buffer_data_4[1319:1312] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_165[2] = buffer_data_4[1327:1320] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_165[3] = buffer_data_4[1335:1328] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_165[4] = buffer_data_4[1343:1336] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_165[5] = buffer_data_3[1311:1304] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_165[6] = buffer_data_3[1319:1312] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_165[7] = buffer_data_3[1327:1320] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_165[8] = buffer_data_3[1335:1328] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_165[9] = buffer_data_3[1343:1336] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_165[10] = buffer_data_2[1311:1304] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_165[11] = buffer_data_2[1319:1312] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_165[12] = buffer_data_2[1327:1320] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_165[13] = buffer_data_2[1335:1328] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_165[14] = buffer_data_2[1343:1336] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_165[15] = buffer_data_1[1311:1304] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_165[16] = buffer_data_1[1319:1312] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_165[17] = buffer_data_1[1327:1320] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_165[18] = buffer_data_1[1335:1328] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_165[19] = buffer_data_1[1343:1336] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_165[20] = buffer_data_0[1311:1304] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_165[21] = buffer_data_0[1319:1312] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_165[22] = buffer_data_0[1327:1320] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_165[23] = buffer_data_0[1335:1328] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_165[24] = buffer_data_0[1343:1336] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_165 = kernel_img_mul_165[0] + kernel_img_mul_165[1] + kernel_img_mul_165[2] + 
                kernel_img_mul_165[3] + kernel_img_mul_165[4] + kernel_img_mul_165[5] + 
                kernel_img_mul_165[6] + kernel_img_mul_165[7] + kernel_img_mul_165[8] + 
                kernel_img_mul_165[9] + kernel_img_mul_165[10] + kernel_img_mul_165[11] + 
                kernel_img_mul_165[12] + kernel_img_mul_165[13] + kernel_img_mul_165[14] + 
                kernel_img_mul_165[15] + kernel_img_mul_165[16] + kernel_img_mul_165[17] + 
                kernel_img_mul_165[18] + kernel_img_mul_165[19] + kernel_img_mul_165[20] + 
                kernel_img_mul_165[21] + kernel_img_mul_165[22] + kernel_img_mul_165[23] + 
                kernel_img_mul_165[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1327:1320] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1327:1320] <= kernel_img_sum_165[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1327:1320] <= 'd0;
end

wire  [39:0]  kernel_img_mul_166[0:24];
assign kernel_img_mul_166[0] = buffer_data_4[1319:1312] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_166[1] = buffer_data_4[1327:1320] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_166[2] = buffer_data_4[1335:1328] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_166[3] = buffer_data_4[1343:1336] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_166[4] = buffer_data_4[1351:1344] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_166[5] = buffer_data_3[1319:1312] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_166[6] = buffer_data_3[1327:1320] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_166[7] = buffer_data_3[1335:1328] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_166[8] = buffer_data_3[1343:1336] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_166[9] = buffer_data_3[1351:1344] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_166[10] = buffer_data_2[1319:1312] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_166[11] = buffer_data_2[1327:1320] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_166[12] = buffer_data_2[1335:1328] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_166[13] = buffer_data_2[1343:1336] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_166[14] = buffer_data_2[1351:1344] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_166[15] = buffer_data_1[1319:1312] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_166[16] = buffer_data_1[1327:1320] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_166[17] = buffer_data_1[1335:1328] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_166[18] = buffer_data_1[1343:1336] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_166[19] = buffer_data_1[1351:1344] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_166[20] = buffer_data_0[1319:1312] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_166[21] = buffer_data_0[1327:1320] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_166[22] = buffer_data_0[1335:1328] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_166[23] = buffer_data_0[1343:1336] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_166[24] = buffer_data_0[1351:1344] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_166 = kernel_img_mul_166[0] + kernel_img_mul_166[1] + kernel_img_mul_166[2] + 
                kernel_img_mul_166[3] + kernel_img_mul_166[4] + kernel_img_mul_166[5] + 
                kernel_img_mul_166[6] + kernel_img_mul_166[7] + kernel_img_mul_166[8] + 
                kernel_img_mul_166[9] + kernel_img_mul_166[10] + kernel_img_mul_166[11] + 
                kernel_img_mul_166[12] + kernel_img_mul_166[13] + kernel_img_mul_166[14] + 
                kernel_img_mul_166[15] + kernel_img_mul_166[16] + kernel_img_mul_166[17] + 
                kernel_img_mul_166[18] + kernel_img_mul_166[19] + kernel_img_mul_166[20] + 
                kernel_img_mul_166[21] + kernel_img_mul_166[22] + kernel_img_mul_166[23] + 
                kernel_img_mul_166[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1335:1328] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1335:1328] <= kernel_img_sum_166[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1335:1328] <= 'd0;
end

wire  [39:0]  kernel_img_mul_167[0:24];
assign kernel_img_mul_167[0] = buffer_data_4[1327:1320] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_167[1] = buffer_data_4[1335:1328] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_167[2] = buffer_data_4[1343:1336] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_167[3] = buffer_data_4[1351:1344] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_167[4] = buffer_data_4[1359:1352] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_167[5] = buffer_data_3[1327:1320] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_167[6] = buffer_data_3[1335:1328] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_167[7] = buffer_data_3[1343:1336] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_167[8] = buffer_data_3[1351:1344] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_167[9] = buffer_data_3[1359:1352] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_167[10] = buffer_data_2[1327:1320] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_167[11] = buffer_data_2[1335:1328] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_167[12] = buffer_data_2[1343:1336] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_167[13] = buffer_data_2[1351:1344] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_167[14] = buffer_data_2[1359:1352] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_167[15] = buffer_data_1[1327:1320] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_167[16] = buffer_data_1[1335:1328] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_167[17] = buffer_data_1[1343:1336] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_167[18] = buffer_data_1[1351:1344] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_167[19] = buffer_data_1[1359:1352] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_167[20] = buffer_data_0[1327:1320] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_167[21] = buffer_data_0[1335:1328] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_167[22] = buffer_data_0[1343:1336] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_167[23] = buffer_data_0[1351:1344] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_167[24] = buffer_data_0[1359:1352] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_167 = kernel_img_mul_167[0] + kernel_img_mul_167[1] + kernel_img_mul_167[2] + 
                kernel_img_mul_167[3] + kernel_img_mul_167[4] + kernel_img_mul_167[5] + 
                kernel_img_mul_167[6] + kernel_img_mul_167[7] + kernel_img_mul_167[8] + 
                kernel_img_mul_167[9] + kernel_img_mul_167[10] + kernel_img_mul_167[11] + 
                kernel_img_mul_167[12] + kernel_img_mul_167[13] + kernel_img_mul_167[14] + 
                kernel_img_mul_167[15] + kernel_img_mul_167[16] + kernel_img_mul_167[17] + 
                kernel_img_mul_167[18] + kernel_img_mul_167[19] + kernel_img_mul_167[20] + 
                kernel_img_mul_167[21] + kernel_img_mul_167[22] + kernel_img_mul_167[23] + 
                kernel_img_mul_167[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1343:1336] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1343:1336] <= kernel_img_sum_167[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1343:1336] <= 'd0;
end

wire  [39:0]  kernel_img_mul_168[0:24];
assign kernel_img_mul_168[0] = buffer_data_4[1335:1328] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_168[1] = buffer_data_4[1343:1336] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_168[2] = buffer_data_4[1351:1344] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_168[3] = buffer_data_4[1359:1352] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_168[4] = buffer_data_4[1367:1360] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_168[5] = buffer_data_3[1335:1328] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_168[6] = buffer_data_3[1343:1336] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_168[7] = buffer_data_3[1351:1344] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_168[8] = buffer_data_3[1359:1352] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_168[9] = buffer_data_3[1367:1360] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_168[10] = buffer_data_2[1335:1328] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_168[11] = buffer_data_2[1343:1336] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_168[12] = buffer_data_2[1351:1344] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_168[13] = buffer_data_2[1359:1352] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_168[14] = buffer_data_2[1367:1360] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_168[15] = buffer_data_1[1335:1328] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_168[16] = buffer_data_1[1343:1336] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_168[17] = buffer_data_1[1351:1344] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_168[18] = buffer_data_1[1359:1352] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_168[19] = buffer_data_1[1367:1360] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_168[20] = buffer_data_0[1335:1328] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_168[21] = buffer_data_0[1343:1336] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_168[22] = buffer_data_0[1351:1344] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_168[23] = buffer_data_0[1359:1352] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_168[24] = buffer_data_0[1367:1360] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_168 = kernel_img_mul_168[0] + kernel_img_mul_168[1] + kernel_img_mul_168[2] + 
                kernel_img_mul_168[3] + kernel_img_mul_168[4] + kernel_img_mul_168[5] + 
                kernel_img_mul_168[6] + kernel_img_mul_168[7] + kernel_img_mul_168[8] + 
                kernel_img_mul_168[9] + kernel_img_mul_168[10] + kernel_img_mul_168[11] + 
                kernel_img_mul_168[12] + kernel_img_mul_168[13] + kernel_img_mul_168[14] + 
                kernel_img_mul_168[15] + kernel_img_mul_168[16] + kernel_img_mul_168[17] + 
                kernel_img_mul_168[18] + kernel_img_mul_168[19] + kernel_img_mul_168[20] + 
                kernel_img_mul_168[21] + kernel_img_mul_168[22] + kernel_img_mul_168[23] + 
                kernel_img_mul_168[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1351:1344] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1351:1344] <= kernel_img_sum_168[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1351:1344] <= 'd0;
end

wire  [39:0]  kernel_img_mul_169[0:24];
assign kernel_img_mul_169[0] = buffer_data_4[1343:1336] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_169[1] = buffer_data_4[1351:1344] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_169[2] = buffer_data_4[1359:1352] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_169[3] = buffer_data_4[1367:1360] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_169[4] = buffer_data_4[1375:1368] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_169[5] = buffer_data_3[1343:1336] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_169[6] = buffer_data_3[1351:1344] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_169[7] = buffer_data_3[1359:1352] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_169[8] = buffer_data_3[1367:1360] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_169[9] = buffer_data_3[1375:1368] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_169[10] = buffer_data_2[1343:1336] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_169[11] = buffer_data_2[1351:1344] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_169[12] = buffer_data_2[1359:1352] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_169[13] = buffer_data_2[1367:1360] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_169[14] = buffer_data_2[1375:1368] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_169[15] = buffer_data_1[1343:1336] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_169[16] = buffer_data_1[1351:1344] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_169[17] = buffer_data_1[1359:1352] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_169[18] = buffer_data_1[1367:1360] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_169[19] = buffer_data_1[1375:1368] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_169[20] = buffer_data_0[1343:1336] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_169[21] = buffer_data_0[1351:1344] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_169[22] = buffer_data_0[1359:1352] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_169[23] = buffer_data_0[1367:1360] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_169[24] = buffer_data_0[1375:1368] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_169 = kernel_img_mul_169[0] + kernel_img_mul_169[1] + kernel_img_mul_169[2] + 
                kernel_img_mul_169[3] + kernel_img_mul_169[4] + kernel_img_mul_169[5] + 
                kernel_img_mul_169[6] + kernel_img_mul_169[7] + kernel_img_mul_169[8] + 
                kernel_img_mul_169[9] + kernel_img_mul_169[10] + kernel_img_mul_169[11] + 
                kernel_img_mul_169[12] + kernel_img_mul_169[13] + kernel_img_mul_169[14] + 
                kernel_img_mul_169[15] + kernel_img_mul_169[16] + kernel_img_mul_169[17] + 
                kernel_img_mul_169[18] + kernel_img_mul_169[19] + kernel_img_mul_169[20] + 
                kernel_img_mul_169[21] + kernel_img_mul_169[22] + kernel_img_mul_169[23] + 
                kernel_img_mul_169[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1359:1352] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1359:1352] <= kernel_img_sum_169[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1359:1352] <= 'd0;
end

wire  [39:0]  kernel_img_mul_170[0:24];
assign kernel_img_mul_170[0] = buffer_data_4[1351:1344] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_170[1] = buffer_data_4[1359:1352] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_170[2] = buffer_data_4[1367:1360] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_170[3] = buffer_data_4[1375:1368] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_170[4] = buffer_data_4[1383:1376] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_170[5] = buffer_data_3[1351:1344] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_170[6] = buffer_data_3[1359:1352] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_170[7] = buffer_data_3[1367:1360] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_170[8] = buffer_data_3[1375:1368] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_170[9] = buffer_data_3[1383:1376] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_170[10] = buffer_data_2[1351:1344] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_170[11] = buffer_data_2[1359:1352] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_170[12] = buffer_data_2[1367:1360] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_170[13] = buffer_data_2[1375:1368] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_170[14] = buffer_data_2[1383:1376] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_170[15] = buffer_data_1[1351:1344] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_170[16] = buffer_data_1[1359:1352] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_170[17] = buffer_data_1[1367:1360] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_170[18] = buffer_data_1[1375:1368] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_170[19] = buffer_data_1[1383:1376] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_170[20] = buffer_data_0[1351:1344] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_170[21] = buffer_data_0[1359:1352] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_170[22] = buffer_data_0[1367:1360] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_170[23] = buffer_data_0[1375:1368] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_170[24] = buffer_data_0[1383:1376] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_170 = kernel_img_mul_170[0] + kernel_img_mul_170[1] + kernel_img_mul_170[2] + 
                kernel_img_mul_170[3] + kernel_img_mul_170[4] + kernel_img_mul_170[5] + 
                kernel_img_mul_170[6] + kernel_img_mul_170[7] + kernel_img_mul_170[8] + 
                kernel_img_mul_170[9] + kernel_img_mul_170[10] + kernel_img_mul_170[11] + 
                kernel_img_mul_170[12] + kernel_img_mul_170[13] + kernel_img_mul_170[14] + 
                kernel_img_mul_170[15] + kernel_img_mul_170[16] + kernel_img_mul_170[17] + 
                kernel_img_mul_170[18] + kernel_img_mul_170[19] + kernel_img_mul_170[20] + 
                kernel_img_mul_170[21] + kernel_img_mul_170[22] + kernel_img_mul_170[23] + 
                kernel_img_mul_170[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1367:1360] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1367:1360] <= kernel_img_sum_170[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1367:1360] <= 'd0;
end

wire  [39:0]  kernel_img_mul_171[0:24];
assign kernel_img_mul_171[0] = buffer_data_4[1359:1352] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_171[1] = buffer_data_4[1367:1360] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_171[2] = buffer_data_4[1375:1368] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_171[3] = buffer_data_4[1383:1376] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_171[4] = buffer_data_4[1391:1384] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_171[5] = buffer_data_3[1359:1352] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_171[6] = buffer_data_3[1367:1360] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_171[7] = buffer_data_3[1375:1368] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_171[8] = buffer_data_3[1383:1376] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_171[9] = buffer_data_3[1391:1384] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_171[10] = buffer_data_2[1359:1352] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_171[11] = buffer_data_2[1367:1360] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_171[12] = buffer_data_2[1375:1368] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_171[13] = buffer_data_2[1383:1376] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_171[14] = buffer_data_2[1391:1384] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_171[15] = buffer_data_1[1359:1352] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_171[16] = buffer_data_1[1367:1360] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_171[17] = buffer_data_1[1375:1368] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_171[18] = buffer_data_1[1383:1376] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_171[19] = buffer_data_1[1391:1384] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_171[20] = buffer_data_0[1359:1352] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_171[21] = buffer_data_0[1367:1360] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_171[22] = buffer_data_0[1375:1368] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_171[23] = buffer_data_0[1383:1376] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_171[24] = buffer_data_0[1391:1384] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_171 = kernel_img_mul_171[0] + kernel_img_mul_171[1] + kernel_img_mul_171[2] + 
                kernel_img_mul_171[3] + kernel_img_mul_171[4] + kernel_img_mul_171[5] + 
                kernel_img_mul_171[6] + kernel_img_mul_171[7] + kernel_img_mul_171[8] + 
                kernel_img_mul_171[9] + kernel_img_mul_171[10] + kernel_img_mul_171[11] + 
                kernel_img_mul_171[12] + kernel_img_mul_171[13] + kernel_img_mul_171[14] + 
                kernel_img_mul_171[15] + kernel_img_mul_171[16] + kernel_img_mul_171[17] + 
                kernel_img_mul_171[18] + kernel_img_mul_171[19] + kernel_img_mul_171[20] + 
                kernel_img_mul_171[21] + kernel_img_mul_171[22] + kernel_img_mul_171[23] + 
                kernel_img_mul_171[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1375:1368] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1375:1368] <= kernel_img_sum_171[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1375:1368] <= 'd0;
end

wire  [39:0]  kernel_img_mul_172[0:24];
assign kernel_img_mul_172[0] = buffer_data_4[1367:1360] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_172[1] = buffer_data_4[1375:1368] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_172[2] = buffer_data_4[1383:1376] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_172[3] = buffer_data_4[1391:1384] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_172[4] = buffer_data_4[1399:1392] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_172[5] = buffer_data_3[1367:1360] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_172[6] = buffer_data_3[1375:1368] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_172[7] = buffer_data_3[1383:1376] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_172[8] = buffer_data_3[1391:1384] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_172[9] = buffer_data_3[1399:1392] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_172[10] = buffer_data_2[1367:1360] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_172[11] = buffer_data_2[1375:1368] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_172[12] = buffer_data_2[1383:1376] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_172[13] = buffer_data_2[1391:1384] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_172[14] = buffer_data_2[1399:1392] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_172[15] = buffer_data_1[1367:1360] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_172[16] = buffer_data_1[1375:1368] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_172[17] = buffer_data_1[1383:1376] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_172[18] = buffer_data_1[1391:1384] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_172[19] = buffer_data_1[1399:1392] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_172[20] = buffer_data_0[1367:1360] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_172[21] = buffer_data_0[1375:1368] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_172[22] = buffer_data_0[1383:1376] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_172[23] = buffer_data_0[1391:1384] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_172[24] = buffer_data_0[1399:1392] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_172 = kernel_img_mul_172[0] + kernel_img_mul_172[1] + kernel_img_mul_172[2] + 
                kernel_img_mul_172[3] + kernel_img_mul_172[4] + kernel_img_mul_172[5] + 
                kernel_img_mul_172[6] + kernel_img_mul_172[7] + kernel_img_mul_172[8] + 
                kernel_img_mul_172[9] + kernel_img_mul_172[10] + kernel_img_mul_172[11] + 
                kernel_img_mul_172[12] + kernel_img_mul_172[13] + kernel_img_mul_172[14] + 
                kernel_img_mul_172[15] + kernel_img_mul_172[16] + kernel_img_mul_172[17] + 
                kernel_img_mul_172[18] + kernel_img_mul_172[19] + kernel_img_mul_172[20] + 
                kernel_img_mul_172[21] + kernel_img_mul_172[22] + kernel_img_mul_172[23] + 
                kernel_img_mul_172[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1383:1376] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1383:1376] <= kernel_img_sum_172[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1383:1376] <= 'd0;
end

wire  [39:0]  kernel_img_mul_173[0:24];
assign kernel_img_mul_173[0] = buffer_data_4[1375:1368] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_173[1] = buffer_data_4[1383:1376] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_173[2] = buffer_data_4[1391:1384] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_173[3] = buffer_data_4[1399:1392] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_173[4] = buffer_data_4[1407:1400] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_173[5] = buffer_data_3[1375:1368] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_173[6] = buffer_data_3[1383:1376] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_173[7] = buffer_data_3[1391:1384] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_173[8] = buffer_data_3[1399:1392] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_173[9] = buffer_data_3[1407:1400] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_173[10] = buffer_data_2[1375:1368] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_173[11] = buffer_data_2[1383:1376] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_173[12] = buffer_data_2[1391:1384] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_173[13] = buffer_data_2[1399:1392] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_173[14] = buffer_data_2[1407:1400] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_173[15] = buffer_data_1[1375:1368] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_173[16] = buffer_data_1[1383:1376] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_173[17] = buffer_data_1[1391:1384] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_173[18] = buffer_data_1[1399:1392] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_173[19] = buffer_data_1[1407:1400] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_173[20] = buffer_data_0[1375:1368] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_173[21] = buffer_data_0[1383:1376] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_173[22] = buffer_data_0[1391:1384] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_173[23] = buffer_data_0[1399:1392] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_173[24] = buffer_data_0[1407:1400] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_173 = kernel_img_mul_173[0] + kernel_img_mul_173[1] + kernel_img_mul_173[2] + 
                kernel_img_mul_173[3] + kernel_img_mul_173[4] + kernel_img_mul_173[5] + 
                kernel_img_mul_173[6] + kernel_img_mul_173[7] + kernel_img_mul_173[8] + 
                kernel_img_mul_173[9] + kernel_img_mul_173[10] + kernel_img_mul_173[11] + 
                kernel_img_mul_173[12] + kernel_img_mul_173[13] + kernel_img_mul_173[14] + 
                kernel_img_mul_173[15] + kernel_img_mul_173[16] + kernel_img_mul_173[17] + 
                kernel_img_mul_173[18] + kernel_img_mul_173[19] + kernel_img_mul_173[20] + 
                kernel_img_mul_173[21] + kernel_img_mul_173[22] + kernel_img_mul_173[23] + 
                kernel_img_mul_173[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1391:1384] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1391:1384] <= kernel_img_sum_173[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1391:1384] <= 'd0;
end

wire  [39:0]  kernel_img_mul_174[0:24];
assign kernel_img_mul_174[0] = buffer_data_4[1383:1376] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_174[1] = buffer_data_4[1391:1384] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_174[2] = buffer_data_4[1399:1392] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_174[3] = buffer_data_4[1407:1400] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_174[4] = buffer_data_4[1415:1408] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_174[5] = buffer_data_3[1383:1376] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_174[6] = buffer_data_3[1391:1384] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_174[7] = buffer_data_3[1399:1392] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_174[8] = buffer_data_3[1407:1400] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_174[9] = buffer_data_3[1415:1408] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_174[10] = buffer_data_2[1383:1376] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_174[11] = buffer_data_2[1391:1384] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_174[12] = buffer_data_2[1399:1392] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_174[13] = buffer_data_2[1407:1400] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_174[14] = buffer_data_2[1415:1408] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_174[15] = buffer_data_1[1383:1376] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_174[16] = buffer_data_1[1391:1384] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_174[17] = buffer_data_1[1399:1392] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_174[18] = buffer_data_1[1407:1400] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_174[19] = buffer_data_1[1415:1408] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_174[20] = buffer_data_0[1383:1376] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_174[21] = buffer_data_0[1391:1384] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_174[22] = buffer_data_0[1399:1392] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_174[23] = buffer_data_0[1407:1400] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_174[24] = buffer_data_0[1415:1408] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_174 = kernel_img_mul_174[0] + kernel_img_mul_174[1] + kernel_img_mul_174[2] + 
                kernel_img_mul_174[3] + kernel_img_mul_174[4] + kernel_img_mul_174[5] + 
                kernel_img_mul_174[6] + kernel_img_mul_174[7] + kernel_img_mul_174[8] + 
                kernel_img_mul_174[9] + kernel_img_mul_174[10] + kernel_img_mul_174[11] + 
                kernel_img_mul_174[12] + kernel_img_mul_174[13] + kernel_img_mul_174[14] + 
                kernel_img_mul_174[15] + kernel_img_mul_174[16] + kernel_img_mul_174[17] + 
                kernel_img_mul_174[18] + kernel_img_mul_174[19] + kernel_img_mul_174[20] + 
                kernel_img_mul_174[21] + kernel_img_mul_174[22] + kernel_img_mul_174[23] + 
                kernel_img_mul_174[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1399:1392] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1399:1392] <= kernel_img_sum_174[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1399:1392] <= 'd0;
end

wire  [39:0]  kernel_img_mul_175[0:24];
assign kernel_img_mul_175[0] = buffer_data_4[1391:1384] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_175[1] = buffer_data_4[1399:1392] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_175[2] = buffer_data_4[1407:1400] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_175[3] = buffer_data_4[1415:1408] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_175[4] = buffer_data_4[1423:1416] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_175[5] = buffer_data_3[1391:1384] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_175[6] = buffer_data_3[1399:1392] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_175[7] = buffer_data_3[1407:1400] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_175[8] = buffer_data_3[1415:1408] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_175[9] = buffer_data_3[1423:1416] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_175[10] = buffer_data_2[1391:1384] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_175[11] = buffer_data_2[1399:1392] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_175[12] = buffer_data_2[1407:1400] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_175[13] = buffer_data_2[1415:1408] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_175[14] = buffer_data_2[1423:1416] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_175[15] = buffer_data_1[1391:1384] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_175[16] = buffer_data_1[1399:1392] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_175[17] = buffer_data_1[1407:1400] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_175[18] = buffer_data_1[1415:1408] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_175[19] = buffer_data_1[1423:1416] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_175[20] = buffer_data_0[1391:1384] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_175[21] = buffer_data_0[1399:1392] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_175[22] = buffer_data_0[1407:1400] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_175[23] = buffer_data_0[1415:1408] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_175[24] = buffer_data_0[1423:1416] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_175 = kernel_img_mul_175[0] + kernel_img_mul_175[1] + kernel_img_mul_175[2] + 
                kernel_img_mul_175[3] + kernel_img_mul_175[4] + kernel_img_mul_175[5] + 
                kernel_img_mul_175[6] + kernel_img_mul_175[7] + kernel_img_mul_175[8] + 
                kernel_img_mul_175[9] + kernel_img_mul_175[10] + kernel_img_mul_175[11] + 
                kernel_img_mul_175[12] + kernel_img_mul_175[13] + kernel_img_mul_175[14] + 
                kernel_img_mul_175[15] + kernel_img_mul_175[16] + kernel_img_mul_175[17] + 
                kernel_img_mul_175[18] + kernel_img_mul_175[19] + kernel_img_mul_175[20] + 
                kernel_img_mul_175[21] + kernel_img_mul_175[22] + kernel_img_mul_175[23] + 
                kernel_img_mul_175[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1407:1400] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1407:1400] <= kernel_img_sum_175[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1407:1400] <= 'd0;
end

wire  [39:0]  kernel_img_mul_176[0:24];
assign kernel_img_mul_176[0] = buffer_data_4[1399:1392] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_176[1] = buffer_data_4[1407:1400] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_176[2] = buffer_data_4[1415:1408] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_176[3] = buffer_data_4[1423:1416] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_176[4] = buffer_data_4[1431:1424] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_176[5] = buffer_data_3[1399:1392] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_176[6] = buffer_data_3[1407:1400] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_176[7] = buffer_data_3[1415:1408] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_176[8] = buffer_data_3[1423:1416] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_176[9] = buffer_data_3[1431:1424] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_176[10] = buffer_data_2[1399:1392] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_176[11] = buffer_data_2[1407:1400] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_176[12] = buffer_data_2[1415:1408] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_176[13] = buffer_data_2[1423:1416] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_176[14] = buffer_data_2[1431:1424] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_176[15] = buffer_data_1[1399:1392] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_176[16] = buffer_data_1[1407:1400] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_176[17] = buffer_data_1[1415:1408] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_176[18] = buffer_data_1[1423:1416] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_176[19] = buffer_data_1[1431:1424] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_176[20] = buffer_data_0[1399:1392] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_176[21] = buffer_data_0[1407:1400] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_176[22] = buffer_data_0[1415:1408] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_176[23] = buffer_data_0[1423:1416] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_176[24] = buffer_data_0[1431:1424] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_176 = kernel_img_mul_176[0] + kernel_img_mul_176[1] + kernel_img_mul_176[2] + 
                kernel_img_mul_176[3] + kernel_img_mul_176[4] + kernel_img_mul_176[5] + 
                kernel_img_mul_176[6] + kernel_img_mul_176[7] + kernel_img_mul_176[8] + 
                kernel_img_mul_176[9] + kernel_img_mul_176[10] + kernel_img_mul_176[11] + 
                kernel_img_mul_176[12] + kernel_img_mul_176[13] + kernel_img_mul_176[14] + 
                kernel_img_mul_176[15] + kernel_img_mul_176[16] + kernel_img_mul_176[17] + 
                kernel_img_mul_176[18] + kernel_img_mul_176[19] + kernel_img_mul_176[20] + 
                kernel_img_mul_176[21] + kernel_img_mul_176[22] + kernel_img_mul_176[23] + 
                kernel_img_mul_176[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1415:1408] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1415:1408] <= kernel_img_sum_176[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1415:1408] <= 'd0;
end

wire  [39:0]  kernel_img_mul_177[0:24];
assign kernel_img_mul_177[0] = buffer_data_4[1407:1400] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_177[1] = buffer_data_4[1415:1408] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_177[2] = buffer_data_4[1423:1416] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_177[3] = buffer_data_4[1431:1424] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_177[4] = buffer_data_4[1439:1432] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_177[5] = buffer_data_3[1407:1400] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_177[6] = buffer_data_3[1415:1408] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_177[7] = buffer_data_3[1423:1416] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_177[8] = buffer_data_3[1431:1424] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_177[9] = buffer_data_3[1439:1432] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_177[10] = buffer_data_2[1407:1400] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_177[11] = buffer_data_2[1415:1408] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_177[12] = buffer_data_2[1423:1416] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_177[13] = buffer_data_2[1431:1424] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_177[14] = buffer_data_2[1439:1432] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_177[15] = buffer_data_1[1407:1400] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_177[16] = buffer_data_1[1415:1408] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_177[17] = buffer_data_1[1423:1416] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_177[18] = buffer_data_1[1431:1424] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_177[19] = buffer_data_1[1439:1432] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_177[20] = buffer_data_0[1407:1400] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_177[21] = buffer_data_0[1415:1408] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_177[22] = buffer_data_0[1423:1416] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_177[23] = buffer_data_0[1431:1424] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_177[24] = buffer_data_0[1439:1432] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_177 = kernel_img_mul_177[0] + kernel_img_mul_177[1] + kernel_img_mul_177[2] + 
                kernel_img_mul_177[3] + kernel_img_mul_177[4] + kernel_img_mul_177[5] + 
                kernel_img_mul_177[6] + kernel_img_mul_177[7] + kernel_img_mul_177[8] + 
                kernel_img_mul_177[9] + kernel_img_mul_177[10] + kernel_img_mul_177[11] + 
                kernel_img_mul_177[12] + kernel_img_mul_177[13] + kernel_img_mul_177[14] + 
                kernel_img_mul_177[15] + kernel_img_mul_177[16] + kernel_img_mul_177[17] + 
                kernel_img_mul_177[18] + kernel_img_mul_177[19] + kernel_img_mul_177[20] + 
                kernel_img_mul_177[21] + kernel_img_mul_177[22] + kernel_img_mul_177[23] + 
                kernel_img_mul_177[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1423:1416] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1423:1416] <= kernel_img_sum_177[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1423:1416] <= 'd0;
end

wire  [39:0]  kernel_img_mul_178[0:24];
assign kernel_img_mul_178[0] = buffer_data_4[1415:1408] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_178[1] = buffer_data_4[1423:1416] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_178[2] = buffer_data_4[1431:1424] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_178[3] = buffer_data_4[1439:1432] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_178[4] = buffer_data_4[1447:1440] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_178[5] = buffer_data_3[1415:1408] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_178[6] = buffer_data_3[1423:1416] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_178[7] = buffer_data_3[1431:1424] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_178[8] = buffer_data_3[1439:1432] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_178[9] = buffer_data_3[1447:1440] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_178[10] = buffer_data_2[1415:1408] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_178[11] = buffer_data_2[1423:1416] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_178[12] = buffer_data_2[1431:1424] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_178[13] = buffer_data_2[1439:1432] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_178[14] = buffer_data_2[1447:1440] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_178[15] = buffer_data_1[1415:1408] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_178[16] = buffer_data_1[1423:1416] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_178[17] = buffer_data_1[1431:1424] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_178[18] = buffer_data_1[1439:1432] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_178[19] = buffer_data_1[1447:1440] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_178[20] = buffer_data_0[1415:1408] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_178[21] = buffer_data_0[1423:1416] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_178[22] = buffer_data_0[1431:1424] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_178[23] = buffer_data_0[1439:1432] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_178[24] = buffer_data_0[1447:1440] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_178 = kernel_img_mul_178[0] + kernel_img_mul_178[1] + kernel_img_mul_178[2] + 
                kernel_img_mul_178[3] + kernel_img_mul_178[4] + kernel_img_mul_178[5] + 
                kernel_img_mul_178[6] + kernel_img_mul_178[7] + kernel_img_mul_178[8] + 
                kernel_img_mul_178[9] + kernel_img_mul_178[10] + kernel_img_mul_178[11] + 
                kernel_img_mul_178[12] + kernel_img_mul_178[13] + kernel_img_mul_178[14] + 
                kernel_img_mul_178[15] + kernel_img_mul_178[16] + kernel_img_mul_178[17] + 
                kernel_img_mul_178[18] + kernel_img_mul_178[19] + kernel_img_mul_178[20] + 
                kernel_img_mul_178[21] + kernel_img_mul_178[22] + kernel_img_mul_178[23] + 
                kernel_img_mul_178[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1431:1424] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1431:1424] <= kernel_img_sum_178[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1431:1424] <= 'd0;
end

wire  [39:0]  kernel_img_mul_179[0:24];
assign kernel_img_mul_179[0] = buffer_data_4[1423:1416] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_179[1] = buffer_data_4[1431:1424] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_179[2] = buffer_data_4[1439:1432] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_179[3] = buffer_data_4[1447:1440] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_179[4] = buffer_data_4[1455:1448] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_179[5] = buffer_data_3[1423:1416] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_179[6] = buffer_data_3[1431:1424] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_179[7] = buffer_data_3[1439:1432] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_179[8] = buffer_data_3[1447:1440] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_179[9] = buffer_data_3[1455:1448] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_179[10] = buffer_data_2[1423:1416] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_179[11] = buffer_data_2[1431:1424] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_179[12] = buffer_data_2[1439:1432] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_179[13] = buffer_data_2[1447:1440] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_179[14] = buffer_data_2[1455:1448] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_179[15] = buffer_data_1[1423:1416] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_179[16] = buffer_data_1[1431:1424] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_179[17] = buffer_data_1[1439:1432] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_179[18] = buffer_data_1[1447:1440] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_179[19] = buffer_data_1[1455:1448] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_179[20] = buffer_data_0[1423:1416] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_179[21] = buffer_data_0[1431:1424] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_179[22] = buffer_data_0[1439:1432] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_179[23] = buffer_data_0[1447:1440] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_179[24] = buffer_data_0[1455:1448] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_179 = kernel_img_mul_179[0] + kernel_img_mul_179[1] + kernel_img_mul_179[2] + 
                kernel_img_mul_179[3] + kernel_img_mul_179[4] + kernel_img_mul_179[5] + 
                kernel_img_mul_179[6] + kernel_img_mul_179[7] + kernel_img_mul_179[8] + 
                kernel_img_mul_179[9] + kernel_img_mul_179[10] + kernel_img_mul_179[11] + 
                kernel_img_mul_179[12] + kernel_img_mul_179[13] + kernel_img_mul_179[14] + 
                kernel_img_mul_179[15] + kernel_img_mul_179[16] + kernel_img_mul_179[17] + 
                kernel_img_mul_179[18] + kernel_img_mul_179[19] + kernel_img_mul_179[20] + 
                kernel_img_mul_179[21] + kernel_img_mul_179[22] + kernel_img_mul_179[23] + 
                kernel_img_mul_179[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1439:1432] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1439:1432] <= kernel_img_sum_179[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1439:1432] <= 'd0;
end

wire  [39:0]  kernel_img_mul_180[0:24];
assign kernel_img_mul_180[0] = buffer_data_4[1431:1424] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_180[1] = buffer_data_4[1439:1432] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_180[2] = buffer_data_4[1447:1440] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_180[3] = buffer_data_4[1455:1448] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_180[4] = buffer_data_4[1463:1456] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_180[5] = buffer_data_3[1431:1424] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_180[6] = buffer_data_3[1439:1432] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_180[7] = buffer_data_3[1447:1440] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_180[8] = buffer_data_3[1455:1448] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_180[9] = buffer_data_3[1463:1456] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_180[10] = buffer_data_2[1431:1424] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_180[11] = buffer_data_2[1439:1432] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_180[12] = buffer_data_2[1447:1440] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_180[13] = buffer_data_2[1455:1448] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_180[14] = buffer_data_2[1463:1456] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_180[15] = buffer_data_1[1431:1424] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_180[16] = buffer_data_1[1439:1432] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_180[17] = buffer_data_1[1447:1440] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_180[18] = buffer_data_1[1455:1448] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_180[19] = buffer_data_1[1463:1456] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_180[20] = buffer_data_0[1431:1424] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_180[21] = buffer_data_0[1439:1432] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_180[22] = buffer_data_0[1447:1440] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_180[23] = buffer_data_0[1455:1448] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_180[24] = buffer_data_0[1463:1456] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_180 = kernel_img_mul_180[0] + kernel_img_mul_180[1] + kernel_img_mul_180[2] + 
                kernel_img_mul_180[3] + kernel_img_mul_180[4] + kernel_img_mul_180[5] + 
                kernel_img_mul_180[6] + kernel_img_mul_180[7] + kernel_img_mul_180[8] + 
                kernel_img_mul_180[9] + kernel_img_mul_180[10] + kernel_img_mul_180[11] + 
                kernel_img_mul_180[12] + kernel_img_mul_180[13] + kernel_img_mul_180[14] + 
                kernel_img_mul_180[15] + kernel_img_mul_180[16] + kernel_img_mul_180[17] + 
                kernel_img_mul_180[18] + kernel_img_mul_180[19] + kernel_img_mul_180[20] + 
                kernel_img_mul_180[21] + kernel_img_mul_180[22] + kernel_img_mul_180[23] + 
                kernel_img_mul_180[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1447:1440] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1447:1440] <= kernel_img_sum_180[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1447:1440] <= 'd0;
end

wire  [39:0]  kernel_img_mul_181[0:24];
assign kernel_img_mul_181[0] = buffer_data_4[1439:1432] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_181[1] = buffer_data_4[1447:1440] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_181[2] = buffer_data_4[1455:1448] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_181[3] = buffer_data_4[1463:1456] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_181[4] = buffer_data_4[1471:1464] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_181[5] = buffer_data_3[1439:1432] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_181[6] = buffer_data_3[1447:1440] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_181[7] = buffer_data_3[1455:1448] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_181[8] = buffer_data_3[1463:1456] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_181[9] = buffer_data_3[1471:1464] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_181[10] = buffer_data_2[1439:1432] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_181[11] = buffer_data_2[1447:1440] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_181[12] = buffer_data_2[1455:1448] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_181[13] = buffer_data_2[1463:1456] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_181[14] = buffer_data_2[1471:1464] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_181[15] = buffer_data_1[1439:1432] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_181[16] = buffer_data_1[1447:1440] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_181[17] = buffer_data_1[1455:1448] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_181[18] = buffer_data_1[1463:1456] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_181[19] = buffer_data_1[1471:1464] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_181[20] = buffer_data_0[1439:1432] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_181[21] = buffer_data_0[1447:1440] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_181[22] = buffer_data_0[1455:1448] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_181[23] = buffer_data_0[1463:1456] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_181[24] = buffer_data_0[1471:1464] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_181 = kernel_img_mul_181[0] + kernel_img_mul_181[1] + kernel_img_mul_181[2] + 
                kernel_img_mul_181[3] + kernel_img_mul_181[4] + kernel_img_mul_181[5] + 
                kernel_img_mul_181[6] + kernel_img_mul_181[7] + kernel_img_mul_181[8] + 
                kernel_img_mul_181[9] + kernel_img_mul_181[10] + kernel_img_mul_181[11] + 
                kernel_img_mul_181[12] + kernel_img_mul_181[13] + kernel_img_mul_181[14] + 
                kernel_img_mul_181[15] + kernel_img_mul_181[16] + kernel_img_mul_181[17] + 
                kernel_img_mul_181[18] + kernel_img_mul_181[19] + kernel_img_mul_181[20] + 
                kernel_img_mul_181[21] + kernel_img_mul_181[22] + kernel_img_mul_181[23] + 
                kernel_img_mul_181[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1455:1448] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1455:1448] <= kernel_img_sum_181[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1455:1448] <= 'd0;
end

wire  [39:0]  kernel_img_mul_182[0:24];
assign kernel_img_mul_182[0] = buffer_data_4[1447:1440] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_182[1] = buffer_data_4[1455:1448] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_182[2] = buffer_data_4[1463:1456] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_182[3] = buffer_data_4[1471:1464] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_182[4] = buffer_data_4[1479:1472] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_182[5] = buffer_data_3[1447:1440] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_182[6] = buffer_data_3[1455:1448] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_182[7] = buffer_data_3[1463:1456] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_182[8] = buffer_data_3[1471:1464] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_182[9] = buffer_data_3[1479:1472] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_182[10] = buffer_data_2[1447:1440] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_182[11] = buffer_data_2[1455:1448] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_182[12] = buffer_data_2[1463:1456] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_182[13] = buffer_data_2[1471:1464] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_182[14] = buffer_data_2[1479:1472] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_182[15] = buffer_data_1[1447:1440] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_182[16] = buffer_data_1[1455:1448] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_182[17] = buffer_data_1[1463:1456] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_182[18] = buffer_data_1[1471:1464] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_182[19] = buffer_data_1[1479:1472] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_182[20] = buffer_data_0[1447:1440] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_182[21] = buffer_data_0[1455:1448] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_182[22] = buffer_data_0[1463:1456] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_182[23] = buffer_data_0[1471:1464] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_182[24] = buffer_data_0[1479:1472] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_182 = kernel_img_mul_182[0] + kernel_img_mul_182[1] + kernel_img_mul_182[2] + 
                kernel_img_mul_182[3] + kernel_img_mul_182[4] + kernel_img_mul_182[5] + 
                kernel_img_mul_182[6] + kernel_img_mul_182[7] + kernel_img_mul_182[8] + 
                kernel_img_mul_182[9] + kernel_img_mul_182[10] + kernel_img_mul_182[11] + 
                kernel_img_mul_182[12] + kernel_img_mul_182[13] + kernel_img_mul_182[14] + 
                kernel_img_mul_182[15] + kernel_img_mul_182[16] + kernel_img_mul_182[17] + 
                kernel_img_mul_182[18] + kernel_img_mul_182[19] + kernel_img_mul_182[20] + 
                kernel_img_mul_182[21] + kernel_img_mul_182[22] + kernel_img_mul_182[23] + 
                kernel_img_mul_182[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1463:1456] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1463:1456] <= kernel_img_sum_182[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1463:1456] <= 'd0;
end

wire  [39:0]  kernel_img_mul_183[0:24];
assign kernel_img_mul_183[0] = buffer_data_4[1455:1448] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_183[1] = buffer_data_4[1463:1456] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_183[2] = buffer_data_4[1471:1464] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_183[3] = buffer_data_4[1479:1472] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_183[4] = buffer_data_4[1487:1480] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_183[5] = buffer_data_3[1455:1448] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_183[6] = buffer_data_3[1463:1456] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_183[7] = buffer_data_3[1471:1464] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_183[8] = buffer_data_3[1479:1472] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_183[9] = buffer_data_3[1487:1480] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_183[10] = buffer_data_2[1455:1448] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_183[11] = buffer_data_2[1463:1456] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_183[12] = buffer_data_2[1471:1464] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_183[13] = buffer_data_2[1479:1472] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_183[14] = buffer_data_2[1487:1480] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_183[15] = buffer_data_1[1455:1448] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_183[16] = buffer_data_1[1463:1456] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_183[17] = buffer_data_1[1471:1464] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_183[18] = buffer_data_1[1479:1472] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_183[19] = buffer_data_1[1487:1480] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_183[20] = buffer_data_0[1455:1448] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_183[21] = buffer_data_0[1463:1456] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_183[22] = buffer_data_0[1471:1464] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_183[23] = buffer_data_0[1479:1472] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_183[24] = buffer_data_0[1487:1480] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_183 = kernel_img_mul_183[0] + kernel_img_mul_183[1] + kernel_img_mul_183[2] + 
                kernel_img_mul_183[3] + kernel_img_mul_183[4] + kernel_img_mul_183[5] + 
                kernel_img_mul_183[6] + kernel_img_mul_183[7] + kernel_img_mul_183[8] + 
                kernel_img_mul_183[9] + kernel_img_mul_183[10] + kernel_img_mul_183[11] + 
                kernel_img_mul_183[12] + kernel_img_mul_183[13] + kernel_img_mul_183[14] + 
                kernel_img_mul_183[15] + kernel_img_mul_183[16] + kernel_img_mul_183[17] + 
                kernel_img_mul_183[18] + kernel_img_mul_183[19] + kernel_img_mul_183[20] + 
                kernel_img_mul_183[21] + kernel_img_mul_183[22] + kernel_img_mul_183[23] + 
                kernel_img_mul_183[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1471:1464] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1471:1464] <= kernel_img_sum_183[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1471:1464] <= 'd0;
end

wire  [39:0]  kernel_img_mul_184[0:24];
assign kernel_img_mul_184[0] = buffer_data_4[1463:1456] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_184[1] = buffer_data_4[1471:1464] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_184[2] = buffer_data_4[1479:1472] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_184[3] = buffer_data_4[1487:1480] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_184[4] = buffer_data_4[1495:1488] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_184[5] = buffer_data_3[1463:1456] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_184[6] = buffer_data_3[1471:1464] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_184[7] = buffer_data_3[1479:1472] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_184[8] = buffer_data_3[1487:1480] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_184[9] = buffer_data_3[1495:1488] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_184[10] = buffer_data_2[1463:1456] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_184[11] = buffer_data_2[1471:1464] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_184[12] = buffer_data_2[1479:1472] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_184[13] = buffer_data_2[1487:1480] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_184[14] = buffer_data_2[1495:1488] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_184[15] = buffer_data_1[1463:1456] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_184[16] = buffer_data_1[1471:1464] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_184[17] = buffer_data_1[1479:1472] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_184[18] = buffer_data_1[1487:1480] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_184[19] = buffer_data_1[1495:1488] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_184[20] = buffer_data_0[1463:1456] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_184[21] = buffer_data_0[1471:1464] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_184[22] = buffer_data_0[1479:1472] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_184[23] = buffer_data_0[1487:1480] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_184[24] = buffer_data_0[1495:1488] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_184 = kernel_img_mul_184[0] + kernel_img_mul_184[1] + kernel_img_mul_184[2] + 
                kernel_img_mul_184[3] + kernel_img_mul_184[4] + kernel_img_mul_184[5] + 
                kernel_img_mul_184[6] + kernel_img_mul_184[7] + kernel_img_mul_184[8] + 
                kernel_img_mul_184[9] + kernel_img_mul_184[10] + kernel_img_mul_184[11] + 
                kernel_img_mul_184[12] + kernel_img_mul_184[13] + kernel_img_mul_184[14] + 
                kernel_img_mul_184[15] + kernel_img_mul_184[16] + kernel_img_mul_184[17] + 
                kernel_img_mul_184[18] + kernel_img_mul_184[19] + kernel_img_mul_184[20] + 
                kernel_img_mul_184[21] + kernel_img_mul_184[22] + kernel_img_mul_184[23] + 
                kernel_img_mul_184[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1479:1472] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1479:1472] <= kernel_img_sum_184[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1479:1472] <= 'd0;
end

wire  [39:0]  kernel_img_mul_185[0:24];
assign kernel_img_mul_185[0] = buffer_data_4[1471:1464] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_185[1] = buffer_data_4[1479:1472] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_185[2] = buffer_data_4[1487:1480] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_185[3] = buffer_data_4[1495:1488] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_185[4] = buffer_data_4[1503:1496] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_185[5] = buffer_data_3[1471:1464] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_185[6] = buffer_data_3[1479:1472] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_185[7] = buffer_data_3[1487:1480] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_185[8] = buffer_data_3[1495:1488] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_185[9] = buffer_data_3[1503:1496] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_185[10] = buffer_data_2[1471:1464] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_185[11] = buffer_data_2[1479:1472] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_185[12] = buffer_data_2[1487:1480] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_185[13] = buffer_data_2[1495:1488] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_185[14] = buffer_data_2[1503:1496] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_185[15] = buffer_data_1[1471:1464] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_185[16] = buffer_data_1[1479:1472] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_185[17] = buffer_data_1[1487:1480] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_185[18] = buffer_data_1[1495:1488] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_185[19] = buffer_data_1[1503:1496] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_185[20] = buffer_data_0[1471:1464] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_185[21] = buffer_data_0[1479:1472] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_185[22] = buffer_data_0[1487:1480] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_185[23] = buffer_data_0[1495:1488] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_185[24] = buffer_data_0[1503:1496] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_185 = kernel_img_mul_185[0] + kernel_img_mul_185[1] + kernel_img_mul_185[2] + 
                kernel_img_mul_185[3] + kernel_img_mul_185[4] + kernel_img_mul_185[5] + 
                kernel_img_mul_185[6] + kernel_img_mul_185[7] + kernel_img_mul_185[8] + 
                kernel_img_mul_185[9] + kernel_img_mul_185[10] + kernel_img_mul_185[11] + 
                kernel_img_mul_185[12] + kernel_img_mul_185[13] + kernel_img_mul_185[14] + 
                kernel_img_mul_185[15] + kernel_img_mul_185[16] + kernel_img_mul_185[17] + 
                kernel_img_mul_185[18] + kernel_img_mul_185[19] + kernel_img_mul_185[20] + 
                kernel_img_mul_185[21] + kernel_img_mul_185[22] + kernel_img_mul_185[23] + 
                kernel_img_mul_185[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1487:1480] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1487:1480] <= kernel_img_sum_185[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1487:1480] <= 'd0;
end

wire  [39:0]  kernel_img_mul_186[0:24];
assign kernel_img_mul_186[0] = buffer_data_4[1479:1472] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_186[1] = buffer_data_4[1487:1480] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_186[2] = buffer_data_4[1495:1488] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_186[3] = buffer_data_4[1503:1496] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_186[4] = buffer_data_4[1511:1504] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_186[5] = buffer_data_3[1479:1472] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_186[6] = buffer_data_3[1487:1480] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_186[7] = buffer_data_3[1495:1488] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_186[8] = buffer_data_3[1503:1496] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_186[9] = buffer_data_3[1511:1504] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_186[10] = buffer_data_2[1479:1472] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_186[11] = buffer_data_2[1487:1480] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_186[12] = buffer_data_2[1495:1488] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_186[13] = buffer_data_2[1503:1496] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_186[14] = buffer_data_2[1511:1504] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_186[15] = buffer_data_1[1479:1472] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_186[16] = buffer_data_1[1487:1480] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_186[17] = buffer_data_1[1495:1488] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_186[18] = buffer_data_1[1503:1496] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_186[19] = buffer_data_1[1511:1504] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_186[20] = buffer_data_0[1479:1472] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_186[21] = buffer_data_0[1487:1480] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_186[22] = buffer_data_0[1495:1488] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_186[23] = buffer_data_0[1503:1496] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_186[24] = buffer_data_0[1511:1504] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_186 = kernel_img_mul_186[0] + kernel_img_mul_186[1] + kernel_img_mul_186[2] + 
                kernel_img_mul_186[3] + kernel_img_mul_186[4] + kernel_img_mul_186[5] + 
                kernel_img_mul_186[6] + kernel_img_mul_186[7] + kernel_img_mul_186[8] + 
                kernel_img_mul_186[9] + kernel_img_mul_186[10] + kernel_img_mul_186[11] + 
                kernel_img_mul_186[12] + kernel_img_mul_186[13] + kernel_img_mul_186[14] + 
                kernel_img_mul_186[15] + kernel_img_mul_186[16] + kernel_img_mul_186[17] + 
                kernel_img_mul_186[18] + kernel_img_mul_186[19] + kernel_img_mul_186[20] + 
                kernel_img_mul_186[21] + kernel_img_mul_186[22] + kernel_img_mul_186[23] + 
                kernel_img_mul_186[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1495:1488] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1495:1488] <= kernel_img_sum_186[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1495:1488] <= 'd0;
end

wire  [39:0]  kernel_img_mul_187[0:24];
assign kernel_img_mul_187[0] = buffer_data_4[1487:1480] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_187[1] = buffer_data_4[1495:1488] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_187[2] = buffer_data_4[1503:1496] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_187[3] = buffer_data_4[1511:1504] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_187[4] = buffer_data_4[1519:1512] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_187[5] = buffer_data_3[1487:1480] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_187[6] = buffer_data_3[1495:1488] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_187[7] = buffer_data_3[1503:1496] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_187[8] = buffer_data_3[1511:1504] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_187[9] = buffer_data_3[1519:1512] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_187[10] = buffer_data_2[1487:1480] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_187[11] = buffer_data_2[1495:1488] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_187[12] = buffer_data_2[1503:1496] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_187[13] = buffer_data_2[1511:1504] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_187[14] = buffer_data_2[1519:1512] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_187[15] = buffer_data_1[1487:1480] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_187[16] = buffer_data_1[1495:1488] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_187[17] = buffer_data_1[1503:1496] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_187[18] = buffer_data_1[1511:1504] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_187[19] = buffer_data_1[1519:1512] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_187[20] = buffer_data_0[1487:1480] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_187[21] = buffer_data_0[1495:1488] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_187[22] = buffer_data_0[1503:1496] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_187[23] = buffer_data_0[1511:1504] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_187[24] = buffer_data_0[1519:1512] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_187 = kernel_img_mul_187[0] + kernel_img_mul_187[1] + kernel_img_mul_187[2] + 
                kernel_img_mul_187[3] + kernel_img_mul_187[4] + kernel_img_mul_187[5] + 
                kernel_img_mul_187[6] + kernel_img_mul_187[7] + kernel_img_mul_187[8] + 
                kernel_img_mul_187[9] + kernel_img_mul_187[10] + kernel_img_mul_187[11] + 
                kernel_img_mul_187[12] + kernel_img_mul_187[13] + kernel_img_mul_187[14] + 
                kernel_img_mul_187[15] + kernel_img_mul_187[16] + kernel_img_mul_187[17] + 
                kernel_img_mul_187[18] + kernel_img_mul_187[19] + kernel_img_mul_187[20] + 
                kernel_img_mul_187[21] + kernel_img_mul_187[22] + kernel_img_mul_187[23] + 
                kernel_img_mul_187[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1503:1496] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1503:1496] <= kernel_img_sum_187[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1503:1496] <= 'd0;
end

wire  [39:0]  kernel_img_mul_188[0:24];
assign kernel_img_mul_188[0] = buffer_data_4[1495:1488] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_188[1] = buffer_data_4[1503:1496] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_188[2] = buffer_data_4[1511:1504] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_188[3] = buffer_data_4[1519:1512] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_188[4] = buffer_data_4[1527:1520] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_188[5] = buffer_data_3[1495:1488] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_188[6] = buffer_data_3[1503:1496] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_188[7] = buffer_data_3[1511:1504] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_188[8] = buffer_data_3[1519:1512] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_188[9] = buffer_data_3[1527:1520] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_188[10] = buffer_data_2[1495:1488] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_188[11] = buffer_data_2[1503:1496] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_188[12] = buffer_data_2[1511:1504] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_188[13] = buffer_data_2[1519:1512] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_188[14] = buffer_data_2[1527:1520] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_188[15] = buffer_data_1[1495:1488] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_188[16] = buffer_data_1[1503:1496] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_188[17] = buffer_data_1[1511:1504] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_188[18] = buffer_data_1[1519:1512] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_188[19] = buffer_data_1[1527:1520] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_188[20] = buffer_data_0[1495:1488] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_188[21] = buffer_data_0[1503:1496] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_188[22] = buffer_data_0[1511:1504] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_188[23] = buffer_data_0[1519:1512] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_188[24] = buffer_data_0[1527:1520] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_188 = kernel_img_mul_188[0] + kernel_img_mul_188[1] + kernel_img_mul_188[2] + 
                kernel_img_mul_188[3] + kernel_img_mul_188[4] + kernel_img_mul_188[5] + 
                kernel_img_mul_188[6] + kernel_img_mul_188[7] + kernel_img_mul_188[8] + 
                kernel_img_mul_188[9] + kernel_img_mul_188[10] + kernel_img_mul_188[11] + 
                kernel_img_mul_188[12] + kernel_img_mul_188[13] + kernel_img_mul_188[14] + 
                kernel_img_mul_188[15] + kernel_img_mul_188[16] + kernel_img_mul_188[17] + 
                kernel_img_mul_188[18] + kernel_img_mul_188[19] + kernel_img_mul_188[20] + 
                kernel_img_mul_188[21] + kernel_img_mul_188[22] + kernel_img_mul_188[23] + 
                kernel_img_mul_188[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1511:1504] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1511:1504] <= kernel_img_sum_188[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1511:1504] <= 'd0;
end

wire  [39:0]  kernel_img_mul_189[0:24];
assign kernel_img_mul_189[0] = buffer_data_4[1503:1496] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_189[1] = buffer_data_4[1511:1504] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_189[2] = buffer_data_4[1519:1512] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_189[3] = buffer_data_4[1527:1520] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_189[4] = buffer_data_4[1535:1528] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_189[5] = buffer_data_3[1503:1496] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_189[6] = buffer_data_3[1511:1504] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_189[7] = buffer_data_3[1519:1512] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_189[8] = buffer_data_3[1527:1520] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_189[9] = buffer_data_3[1535:1528] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_189[10] = buffer_data_2[1503:1496] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_189[11] = buffer_data_2[1511:1504] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_189[12] = buffer_data_2[1519:1512] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_189[13] = buffer_data_2[1527:1520] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_189[14] = buffer_data_2[1535:1528] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_189[15] = buffer_data_1[1503:1496] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_189[16] = buffer_data_1[1511:1504] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_189[17] = buffer_data_1[1519:1512] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_189[18] = buffer_data_1[1527:1520] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_189[19] = buffer_data_1[1535:1528] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_189[20] = buffer_data_0[1503:1496] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_189[21] = buffer_data_0[1511:1504] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_189[22] = buffer_data_0[1519:1512] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_189[23] = buffer_data_0[1527:1520] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_189[24] = buffer_data_0[1535:1528] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_189 = kernel_img_mul_189[0] + kernel_img_mul_189[1] + kernel_img_mul_189[2] + 
                kernel_img_mul_189[3] + kernel_img_mul_189[4] + kernel_img_mul_189[5] + 
                kernel_img_mul_189[6] + kernel_img_mul_189[7] + kernel_img_mul_189[8] + 
                kernel_img_mul_189[9] + kernel_img_mul_189[10] + kernel_img_mul_189[11] + 
                kernel_img_mul_189[12] + kernel_img_mul_189[13] + kernel_img_mul_189[14] + 
                kernel_img_mul_189[15] + kernel_img_mul_189[16] + kernel_img_mul_189[17] + 
                kernel_img_mul_189[18] + kernel_img_mul_189[19] + kernel_img_mul_189[20] + 
                kernel_img_mul_189[21] + kernel_img_mul_189[22] + kernel_img_mul_189[23] + 
                kernel_img_mul_189[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1519:1512] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1519:1512] <= kernel_img_sum_189[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1519:1512] <= 'd0;
end

wire  [39:0]  kernel_img_mul_190[0:24];
assign kernel_img_mul_190[0] = buffer_data_4[1511:1504] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_190[1] = buffer_data_4[1519:1512] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_190[2] = buffer_data_4[1527:1520] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_190[3] = buffer_data_4[1535:1528] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_190[4] = buffer_data_4[1543:1536] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_190[5] = buffer_data_3[1511:1504] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_190[6] = buffer_data_3[1519:1512] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_190[7] = buffer_data_3[1527:1520] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_190[8] = buffer_data_3[1535:1528] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_190[9] = buffer_data_3[1543:1536] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_190[10] = buffer_data_2[1511:1504] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_190[11] = buffer_data_2[1519:1512] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_190[12] = buffer_data_2[1527:1520] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_190[13] = buffer_data_2[1535:1528] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_190[14] = buffer_data_2[1543:1536] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_190[15] = buffer_data_1[1511:1504] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_190[16] = buffer_data_1[1519:1512] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_190[17] = buffer_data_1[1527:1520] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_190[18] = buffer_data_1[1535:1528] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_190[19] = buffer_data_1[1543:1536] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_190[20] = buffer_data_0[1511:1504] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_190[21] = buffer_data_0[1519:1512] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_190[22] = buffer_data_0[1527:1520] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_190[23] = buffer_data_0[1535:1528] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_190[24] = buffer_data_0[1543:1536] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_190 = kernel_img_mul_190[0] + kernel_img_mul_190[1] + kernel_img_mul_190[2] + 
                kernel_img_mul_190[3] + kernel_img_mul_190[4] + kernel_img_mul_190[5] + 
                kernel_img_mul_190[6] + kernel_img_mul_190[7] + kernel_img_mul_190[8] + 
                kernel_img_mul_190[9] + kernel_img_mul_190[10] + kernel_img_mul_190[11] + 
                kernel_img_mul_190[12] + kernel_img_mul_190[13] + kernel_img_mul_190[14] + 
                kernel_img_mul_190[15] + kernel_img_mul_190[16] + kernel_img_mul_190[17] + 
                kernel_img_mul_190[18] + kernel_img_mul_190[19] + kernel_img_mul_190[20] + 
                kernel_img_mul_190[21] + kernel_img_mul_190[22] + kernel_img_mul_190[23] + 
                kernel_img_mul_190[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1527:1520] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1527:1520] <= kernel_img_sum_190[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1527:1520] <= 'd0;
end

wire  [39:0]  kernel_img_mul_191[0:24];
assign kernel_img_mul_191[0] = buffer_data_4[1519:1512] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_191[1] = buffer_data_4[1527:1520] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_191[2] = buffer_data_4[1535:1528] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_191[3] = buffer_data_4[1543:1536] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_191[4] = buffer_data_4[1551:1544] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_191[5] = buffer_data_3[1519:1512] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_191[6] = buffer_data_3[1527:1520] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_191[7] = buffer_data_3[1535:1528] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_191[8] = buffer_data_3[1543:1536] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_191[9] = buffer_data_3[1551:1544] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_191[10] = buffer_data_2[1519:1512] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_191[11] = buffer_data_2[1527:1520] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_191[12] = buffer_data_2[1535:1528] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_191[13] = buffer_data_2[1543:1536] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_191[14] = buffer_data_2[1551:1544] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_191[15] = buffer_data_1[1519:1512] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_191[16] = buffer_data_1[1527:1520] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_191[17] = buffer_data_1[1535:1528] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_191[18] = buffer_data_1[1543:1536] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_191[19] = buffer_data_1[1551:1544] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_191[20] = buffer_data_0[1519:1512] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_191[21] = buffer_data_0[1527:1520] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_191[22] = buffer_data_0[1535:1528] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_191[23] = buffer_data_0[1543:1536] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_191[24] = buffer_data_0[1551:1544] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_191 = kernel_img_mul_191[0] + kernel_img_mul_191[1] + kernel_img_mul_191[2] + 
                kernel_img_mul_191[3] + kernel_img_mul_191[4] + kernel_img_mul_191[5] + 
                kernel_img_mul_191[6] + kernel_img_mul_191[7] + kernel_img_mul_191[8] + 
                kernel_img_mul_191[9] + kernel_img_mul_191[10] + kernel_img_mul_191[11] + 
                kernel_img_mul_191[12] + kernel_img_mul_191[13] + kernel_img_mul_191[14] + 
                kernel_img_mul_191[15] + kernel_img_mul_191[16] + kernel_img_mul_191[17] + 
                kernel_img_mul_191[18] + kernel_img_mul_191[19] + kernel_img_mul_191[20] + 
                kernel_img_mul_191[21] + kernel_img_mul_191[22] + kernel_img_mul_191[23] + 
                kernel_img_mul_191[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1535:1528] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1535:1528] <= kernel_img_sum_191[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1535:1528] <= 'd0;
end

wire  [39:0]  kernel_img_mul_192[0:24];
assign kernel_img_mul_192[0] = buffer_data_4[1527:1520] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_192[1] = buffer_data_4[1535:1528] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_192[2] = buffer_data_4[1543:1536] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_192[3] = buffer_data_4[1551:1544] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_192[4] = buffer_data_4[1559:1552] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_192[5] = buffer_data_3[1527:1520] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_192[6] = buffer_data_3[1535:1528] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_192[7] = buffer_data_3[1543:1536] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_192[8] = buffer_data_3[1551:1544] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_192[9] = buffer_data_3[1559:1552] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_192[10] = buffer_data_2[1527:1520] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_192[11] = buffer_data_2[1535:1528] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_192[12] = buffer_data_2[1543:1536] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_192[13] = buffer_data_2[1551:1544] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_192[14] = buffer_data_2[1559:1552] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_192[15] = buffer_data_1[1527:1520] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_192[16] = buffer_data_1[1535:1528] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_192[17] = buffer_data_1[1543:1536] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_192[18] = buffer_data_1[1551:1544] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_192[19] = buffer_data_1[1559:1552] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_192[20] = buffer_data_0[1527:1520] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_192[21] = buffer_data_0[1535:1528] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_192[22] = buffer_data_0[1543:1536] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_192[23] = buffer_data_0[1551:1544] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_192[24] = buffer_data_0[1559:1552] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_192 = kernel_img_mul_192[0] + kernel_img_mul_192[1] + kernel_img_mul_192[2] + 
                kernel_img_mul_192[3] + kernel_img_mul_192[4] + kernel_img_mul_192[5] + 
                kernel_img_mul_192[6] + kernel_img_mul_192[7] + kernel_img_mul_192[8] + 
                kernel_img_mul_192[9] + kernel_img_mul_192[10] + kernel_img_mul_192[11] + 
                kernel_img_mul_192[12] + kernel_img_mul_192[13] + kernel_img_mul_192[14] + 
                kernel_img_mul_192[15] + kernel_img_mul_192[16] + kernel_img_mul_192[17] + 
                kernel_img_mul_192[18] + kernel_img_mul_192[19] + kernel_img_mul_192[20] + 
                kernel_img_mul_192[21] + kernel_img_mul_192[22] + kernel_img_mul_192[23] + 
                kernel_img_mul_192[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1543:1536] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1543:1536] <= kernel_img_sum_192[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1543:1536] <= 'd0;
end

wire  [39:0]  kernel_img_mul_193[0:24];
assign kernel_img_mul_193[0] = buffer_data_4[1535:1528] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_193[1] = buffer_data_4[1543:1536] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_193[2] = buffer_data_4[1551:1544] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_193[3] = buffer_data_4[1559:1552] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_193[4] = buffer_data_4[1567:1560] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_193[5] = buffer_data_3[1535:1528] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_193[6] = buffer_data_3[1543:1536] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_193[7] = buffer_data_3[1551:1544] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_193[8] = buffer_data_3[1559:1552] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_193[9] = buffer_data_3[1567:1560] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_193[10] = buffer_data_2[1535:1528] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_193[11] = buffer_data_2[1543:1536] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_193[12] = buffer_data_2[1551:1544] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_193[13] = buffer_data_2[1559:1552] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_193[14] = buffer_data_2[1567:1560] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_193[15] = buffer_data_1[1535:1528] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_193[16] = buffer_data_1[1543:1536] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_193[17] = buffer_data_1[1551:1544] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_193[18] = buffer_data_1[1559:1552] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_193[19] = buffer_data_1[1567:1560] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_193[20] = buffer_data_0[1535:1528] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_193[21] = buffer_data_0[1543:1536] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_193[22] = buffer_data_0[1551:1544] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_193[23] = buffer_data_0[1559:1552] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_193[24] = buffer_data_0[1567:1560] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_193 = kernel_img_mul_193[0] + kernel_img_mul_193[1] + kernel_img_mul_193[2] + 
                kernel_img_mul_193[3] + kernel_img_mul_193[4] + kernel_img_mul_193[5] + 
                kernel_img_mul_193[6] + kernel_img_mul_193[7] + kernel_img_mul_193[8] + 
                kernel_img_mul_193[9] + kernel_img_mul_193[10] + kernel_img_mul_193[11] + 
                kernel_img_mul_193[12] + kernel_img_mul_193[13] + kernel_img_mul_193[14] + 
                kernel_img_mul_193[15] + kernel_img_mul_193[16] + kernel_img_mul_193[17] + 
                kernel_img_mul_193[18] + kernel_img_mul_193[19] + kernel_img_mul_193[20] + 
                kernel_img_mul_193[21] + kernel_img_mul_193[22] + kernel_img_mul_193[23] + 
                kernel_img_mul_193[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1551:1544] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1551:1544] <= kernel_img_sum_193[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1551:1544] <= 'd0;
end

wire  [39:0]  kernel_img_mul_194[0:24];
assign kernel_img_mul_194[0] = buffer_data_4[1543:1536] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_194[1] = buffer_data_4[1551:1544] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_194[2] = buffer_data_4[1559:1552] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_194[3] = buffer_data_4[1567:1560] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_194[4] = buffer_data_4[1575:1568] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_194[5] = buffer_data_3[1543:1536] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_194[6] = buffer_data_3[1551:1544] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_194[7] = buffer_data_3[1559:1552] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_194[8] = buffer_data_3[1567:1560] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_194[9] = buffer_data_3[1575:1568] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_194[10] = buffer_data_2[1543:1536] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_194[11] = buffer_data_2[1551:1544] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_194[12] = buffer_data_2[1559:1552] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_194[13] = buffer_data_2[1567:1560] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_194[14] = buffer_data_2[1575:1568] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_194[15] = buffer_data_1[1543:1536] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_194[16] = buffer_data_1[1551:1544] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_194[17] = buffer_data_1[1559:1552] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_194[18] = buffer_data_1[1567:1560] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_194[19] = buffer_data_1[1575:1568] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_194[20] = buffer_data_0[1543:1536] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_194[21] = buffer_data_0[1551:1544] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_194[22] = buffer_data_0[1559:1552] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_194[23] = buffer_data_0[1567:1560] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_194[24] = buffer_data_0[1575:1568] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_194 = kernel_img_mul_194[0] + kernel_img_mul_194[1] + kernel_img_mul_194[2] + 
                kernel_img_mul_194[3] + kernel_img_mul_194[4] + kernel_img_mul_194[5] + 
                kernel_img_mul_194[6] + kernel_img_mul_194[7] + kernel_img_mul_194[8] + 
                kernel_img_mul_194[9] + kernel_img_mul_194[10] + kernel_img_mul_194[11] + 
                kernel_img_mul_194[12] + kernel_img_mul_194[13] + kernel_img_mul_194[14] + 
                kernel_img_mul_194[15] + kernel_img_mul_194[16] + kernel_img_mul_194[17] + 
                kernel_img_mul_194[18] + kernel_img_mul_194[19] + kernel_img_mul_194[20] + 
                kernel_img_mul_194[21] + kernel_img_mul_194[22] + kernel_img_mul_194[23] + 
                kernel_img_mul_194[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1559:1552] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1559:1552] <= kernel_img_sum_194[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1559:1552] <= 'd0;
end

wire  [39:0]  kernel_img_mul_195[0:24];
assign kernel_img_mul_195[0] = buffer_data_4[1551:1544] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_195[1] = buffer_data_4[1559:1552] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_195[2] = buffer_data_4[1567:1560] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_195[3] = buffer_data_4[1575:1568] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_195[4] = buffer_data_4[1583:1576] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_195[5] = buffer_data_3[1551:1544] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_195[6] = buffer_data_3[1559:1552] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_195[7] = buffer_data_3[1567:1560] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_195[8] = buffer_data_3[1575:1568] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_195[9] = buffer_data_3[1583:1576] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_195[10] = buffer_data_2[1551:1544] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_195[11] = buffer_data_2[1559:1552] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_195[12] = buffer_data_2[1567:1560] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_195[13] = buffer_data_2[1575:1568] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_195[14] = buffer_data_2[1583:1576] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_195[15] = buffer_data_1[1551:1544] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_195[16] = buffer_data_1[1559:1552] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_195[17] = buffer_data_1[1567:1560] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_195[18] = buffer_data_1[1575:1568] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_195[19] = buffer_data_1[1583:1576] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_195[20] = buffer_data_0[1551:1544] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_195[21] = buffer_data_0[1559:1552] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_195[22] = buffer_data_0[1567:1560] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_195[23] = buffer_data_0[1575:1568] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_195[24] = buffer_data_0[1583:1576] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_195 = kernel_img_mul_195[0] + kernel_img_mul_195[1] + kernel_img_mul_195[2] + 
                kernel_img_mul_195[3] + kernel_img_mul_195[4] + kernel_img_mul_195[5] + 
                kernel_img_mul_195[6] + kernel_img_mul_195[7] + kernel_img_mul_195[8] + 
                kernel_img_mul_195[9] + kernel_img_mul_195[10] + kernel_img_mul_195[11] + 
                kernel_img_mul_195[12] + kernel_img_mul_195[13] + kernel_img_mul_195[14] + 
                kernel_img_mul_195[15] + kernel_img_mul_195[16] + kernel_img_mul_195[17] + 
                kernel_img_mul_195[18] + kernel_img_mul_195[19] + kernel_img_mul_195[20] + 
                kernel_img_mul_195[21] + kernel_img_mul_195[22] + kernel_img_mul_195[23] + 
                kernel_img_mul_195[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1567:1560] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1567:1560] <= kernel_img_sum_195[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1567:1560] <= 'd0;
end

wire  [39:0]  kernel_img_mul_196[0:24];
assign kernel_img_mul_196[0] = buffer_data_4[1559:1552] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_196[1] = buffer_data_4[1567:1560] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_196[2] = buffer_data_4[1575:1568] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_196[3] = buffer_data_4[1583:1576] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_196[4] = buffer_data_4[1591:1584] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_196[5] = buffer_data_3[1559:1552] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_196[6] = buffer_data_3[1567:1560] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_196[7] = buffer_data_3[1575:1568] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_196[8] = buffer_data_3[1583:1576] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_196[9] = buffer_data_3[1591:1584] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_196[10] = buffer_data_2[1559:1552] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_196[11] = buffer_data_2[1567:1560] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_196[12] = buffer_data_2[1575:1568] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_196[13] = buffer_data_2[1583:1576] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_196[14] = buffer_data_2[1591:1584] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_196[15] = buffer_data_1[1559:1552] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_196[16] = buffer_data_1[1567:1560] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_196[17] = buffer_data_1[1575:1568] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_196[18] = buffer_data_1[1583:1576] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_196[19] = buffer_data_1[1591:1584] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_196[20] = buffer_data_0[1559:1552] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_196[21] = buffer_data_0[1567:1560] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_196[22] = buffer_data_0[1575:1568] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_196[23] = buffer_data_0[1583:1576] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_196[24] = buffer_data_0[1591:1584] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_196 = kernel_img_mul_196[0] + kernel_img_mul_196[1] + kernel_img_mul_196[2] + 
                kernel_img_mul_196[3] + kernel_img_mul_196[4] + kernel_img_mul_196[5] + 
                kernel_img_mul_196[6] + kernel_img_mul_196[7] + kernel_img_mul_196[8] + 
                kernel_img_mul_196[9] + kernel_img_mul_196[10] + kernel_img_mul_196[11] + 
                kernel_img_mul_196[12] + kernel_img_mul_196[13] + kernel_img_mul_196[14] + 
                kernel_img_mul_196[15] + kernel_img_mul_196[16] + kernel_img_mul_196[17] + 
                kernel_img_mul_196[18] + kernel_img_mul_196[19] + kernel_img_mul_196[20] + 
                kernel_img_mul_196[21] + kernel_img_mul_196[22] + kernel_img_mul_196[23] + 
                kernel_img_mul_196[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1575:1568] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1575:1568] <= kernel_img_sum_196[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1575:1568] <= 'd0;
end

wire  [39:0]  kernel_img_mul_197[0:24];
assign kernel_img_mul_197[0] = buffer_data_4[1567:1560] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_197[1] = buffer_data_4[1575:1568] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_197[2] = buffer_data_4[1583:1576] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_197[3] = buffer_data_4[1591:1584] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_197[4] = buffer_data_4[1599:1592] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_197[5] = buffer_data_3[1567:1560] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_197[6] = buffer_data_3[1575:1568] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_197[7] = buffer_data_3[1583:1576] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_197[8] = buffer_data_3[1591:1584] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_197[9] = buffer_data_3[1599:1592] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_197[10] = buffer_data_2[1567:1560] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_197[11] = buffer_data_2[1575:1568] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_197[12] = buffer_data_2[1583:1576] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_197[13] = buffer_data_2[1591:1584] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_197[14] = buffer_data_2[1599:1592] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_197[15] = buffer_data_1[1567:1560] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_197[16] = buffer_data_1[1575:1568] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_197[17] = buffer_data_1[1583:1576] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_197[18] = buffer_data_1[1591:1584] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_197[19] = buffer_data_1[1599:1592] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_197[20] = buffer_data_0[1567:1560] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_197[21] = buffer_data_0[1575:1568] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_197[22] = buffer_data_0[1583:1576] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_197[23] = buffer_data_0[1591:1584] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_197[24] = buffer_data_0[1599:1592] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_197 = kernel_img_mul_197[0] + kernel_img_mul_197[1] + kernel_img_mul_197[2] + 
                kernel_img_mul_197[3] + kernel_img_mul_197[4] + kernel_img_mul_197[5] + 
                kernel_img_mul_197[6] + kernel_img_mul_197[7] + kernel_img_mul_197[8] + 
                kernel_img_mul_197[9] + kernel_img_mul_197[10] + kernel_img_mul_197[11] + 
                kernel_img_mul_197[12] + kernel_img_mul_197[13] + kernel_img_mul_197[14] + 
                kernel_img_mul_197[15] + kernel_img_mul_197[16] + kernel_img_mul_197[17] + 
                kernel_img_mul_197[18] + kernel_img_mul_197[19] + kernel_img_mul_197[20] + 
                kernel_img_mul_197[21] + kernel_img_mul_197[22] + kernel_img_mul_197[23] + 
                kernel_img_mul_197[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1583:1576] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1583:1576] <= kernel_img_sum_197[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1583:1576] <= 'd0;
end

wire  [39:0]  kernel_img_mul_198[0:24];
assign kernel_img_mul_198[0] = buffer_data_4[1575:1568] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_198[1] = buffer_data_4[1583:1576] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_198[2] = buffer_data_4[1591:1584] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_198[3] = buffer_data_4[1599:1592] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_198[4] = buffer_data_4[1607:1600] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_198[5] = buffer_data_3[1575:1568] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_198[6] = buffer_data_3[1583:1576] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_198[7] = buffer_data_3[1591:1584] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_198[8] = buffer_data_3[1599:1592] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_198[9] = buffer_data_3[1607:1600] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_198[10] = buffer_data_2[1575:1568] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_198[11] = buffer_data_2[1583:1576] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_198[12] = buffer_data_2[1591:1584] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_198[13] = buffer_data_2[1599:1592] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_198[14] = buffer_data_2[1607:1600] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_198[15] = buffer_data_1[1575:1568] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_198[16] = buffer_data_1[1583:1576] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_198[17] = buffer_data_1[1591:1584] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_198[18] = buffer_data_1[1599:1592] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_198[19] = buffer_data_1[1607:1600] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_198[20] = buffer_data_0[1575:1568] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_198[21] = buffer_data_0[1583:1576] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_198[22] = buffer_data_0[1591:1584] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_198[23] = buffer_data_0[1599:1592] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_198[24] = buffer_data_0[1607:1600] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_198 = kernel_img_mul_198[0] + kernel_img_mul_198[1] + kernel_img_mul_198[2] + 
                kernel_img_mul_198[3] + kernel_img_mul_198[4] + kernel_img_mul_198[5] + 
                kernel_img_mul_198[6] + kernel_img_mul_198[7] + kernel_img_mul_198[8] + 
                kernel_img_mul_198[9] + kernel_img_mul_198[10] + kernel_img_mul_198[11] + 
                kernel_img_mul_198[12] + kernel_img_mul_198[13] + kernel_img_mul_198[14] + 
                kernel_img_mul_198[15] + kernel_img_mul_198[16] + kernel_img_mul_198[17] + 
                kernel_img_mul_198[18] + kernel_img_mul_198[19] + kernel_img_mul_198[20] + 
                kernel_img_mul_198[21] + kernel_img_mul_198[22] + kernel_img_mul_198[23] + 
                kernel_img_mul_198[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1591:1584] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1591:1584] <= kernel_img_sum_198[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1591:1584] <= 'd0;
end

wire  [39:0]  kernel_img_mul_199[0:24];
assign kernel_img_mul_199[0] = buffer_data_4[1583:1576] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_199[1] = buffer_data_4[1591:1584] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_199[2] = buffer_data_4[1599:1592] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_199[3] = buffer_data_4[1607:1600] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_199[4] = buffer_data_4[1615:1608] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_199[5] = buffer_data_3[1583:1576] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_199[6] = buffer_data_3[1591:1584] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_199[7] = buffer_data_3[1599:1592] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_199[8] = buffer_data_3[1607:1600] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_199[9] = buffer_data_3[1615:1608] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_199[10] = buffer_data_2[1583:1576] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_199[11] = buffer_data_2[1591:1584] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_199[12] = buffer_data_2[1599:1592] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_199[13] = buffer_data_2[1607:1600] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_199[14] = buffer_data_2[1615:1608] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_199[15] = buffer_data_1[1583:1576] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_199[16] = buffer_data_1[1591:1584] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_199[17] = buffer_data_1[1599:1592] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_199[18] = buffer_data_1[1607:1600] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_199[19] = buffer_data_1[1615:1608] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_199[20] = buffer_data_0[1583:1576] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_199[21] = buffer_data_0[1591:1584] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_199[22] = buffer_data_0[1599:1592] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_199[23] = buffer_data_0[1607:1600] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_199[24] = buffer_data_0[1615:1608] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_199 = kernel_img_mul_199[0] + kernel_img_mul_199[1] + kernel_img_mul_199[2] + 
                kernel_img_mul_199[3] + kernel_img_mul_199[4] + kernel_img_mul_199[5] + 
                kernel_img_mul_199[6] + kernel_img_mul_199[7] + kernel_img_mul_199[8] + 
                kernel_img_mul_199[9] + kernel_img_mul_199[10] + kernel_img_mul_199[11] + 
                kernel_img_mul_199[12] + kernel_img_mul_199[13] + kernel_img_mul_199[14] + 
                kernel_img_mul_199[15] + kernel_img_mul_199[16] + kernel_img_mul_199[17] + 
                kernel_img_mul_199[18] + kernel_img_mul_199[19] + kernel_img_mul_199[20] + 
                kernel_img_mul_199[21] + kernel_img_mul_199[22] + kernel_img_mul_199[23] + 
                kernel_img_mul_199[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1599:1592] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1599:1592] <= kernel_img_sum_199[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1599:1592] <= 'd0;
end

wire  [39:0]  kernel_img_mul_200[0:24];
assign kernel_img_mul_200[0] = buffer_data_4[1591:1584] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_200[1] = buffer_data_4[1599:1592] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_200[2] = buffer_data_4[1607:1600] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_200[3] = buffer_data_4[1615:1608] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_200[4] = buffer_data_4[1623:1616] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_200[5] = buffer_data_3[1591:1584] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_200[6] = buffer_data_3[1599:1592] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_200[7] = buffer_data_3[1607:1600] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_200[8] = buffer_data_3[1615:1608] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_200[9] = buffer_data_3[1623:1616] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_200[10] = buffer_data_2[1591:1584] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_200[11] = buffer_data_2[1599:1592] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_200[12] = buffer_data_2[1607:1600] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_200[13] = buffer_data_2[1615:1608] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_200[14] = buffer_data_2[1623:1616] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_200[15] = buffer_data_1[1591:1584] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_200[16] = buffer_data_1[1599:1592] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_200[17] = buffer_data_1[1607:1600] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_200[18] = buffer_data_1[1615:1608] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_200[19] = buffer_data_1[1623:1616] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_200[20] = buffer_data_0[1591:1584] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_200[21] = buffer_data_0[1599:1592] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_200[22] = buffer_data_0[1607:1600] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_200[23] = buffer_data_0[1615:1608] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_200[24] = buffer_data_0[1623:1616] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_200 = kernel_img_mul_200[0] + kernel_img_mul_200[1] + kernel_img_mul_200[2] + 
                kernel_img_mul_200[3] + kernel_img_mul_200[4] + kernel_img_mul_200[5] + 
                kernel_img_mul_200[6] + kernel_img_mul_200[7] + kernel_img_mul_200[8] + 
                kernel_img_mul_200[9] + kernel_img_mul_200[10] + kernel_img_mul_200[11] + 
                kernel_img_mul_200[12] + kernel_img_mul_200[13] + kernel_img_mul_200[14] + 
                kernel_img_mul_200[15] + kernel_img_mul_200[16] + kernel_img_mul_200[17] + 
                kernel_img_mul_200[18] + kernel_img_mul_200[19] + kernel_img_mul_200[20] + 
                kernel_img_mul_200[21] + kernel_img_mul_200[22] + kernel_img_mul_200[23] + 
                kernel_img_mul_200[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1607:1600] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1607:1600] <= kernel_img_sum_200[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1607:1600] <= 'd0;
end

wire  [39:0]  kernel_img_mul_201[0:24];
assign kernel_img_mul_201[0] = buffer_data_4[1599:1592] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_201[1] = buffer_data_4[1607:1600] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_201[2] = buffer_data_4[1615:1608] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_201[3] = buffer_data_4[1623:1616] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_201[4] = buffer_data_4[1631:1624] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_201[5] = buffer_data_3[1599:1592] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_201[6] = buffer_data_3[1607:1600] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_201[7] = buffer_data_3[1615:1608] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_201[8] = buffer_data_3[1623:1616] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_201[9] = buffer_data_3[1631:1624] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_201[10] = buffer_data_2[1599:1592] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_201[11] = buffer_data_2[1607:1600] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_201[12] = buffer_data_2[1615:1608] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_201[13] = buffer_data_2[1623:1616] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_201[14] = buffer_data_2[1631:1624] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_201[15] = buffer_data_1[1599:1592] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_201[16] = buffer_data_1[1607:1600] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_201[17] = buffer_data_1[1615:1608] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_201[18] = buffer_data_1[1623:1616] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_201[19] = buffer_data_1[1631:1624] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_201[20] = buffer_data_0[1599:1592] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_201[21] = buffer_data_0[1607:1600] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_201[22] = buffer_data_0[1615:1608] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_201[23] = buffer_data_0[1623:1616] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_201[24] = buffer_data_0[1631:1624] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_201 = kernel_img_mul_201[0] + kernel_img_mul_201[1] + kernel_img_mul_201[2] + 
                kernel_img_mul_201[3] + kernel_img_mul_201[4] + kernel_img_mul_201[5] + 
                kernel_img_mul_201[6] + kernel_img_mul_201[7] + kernel_img_mul_201[8] + 
                kernel_img_mul_201[9] + kernel_img_mul_201[10] + kernel_img_mul_201[11] + 
                kernel_img_mul_201[12] + kernel_img_mul_201[13] + kernel_img_mul_201[14] + 
                kernel_img_mul_201[15] + kernel_img_mul_201[16] + kernel_img_mul_201[17] + 
                kernel_img_mul_201[18] + kernel_img_mul_201[19] + kernel_img_mul_201[20] + 
                kernel_img_mul_201[21] + kernel_img_mul_201[22] + kernel_img_mul_201[23] + 
                kernel_img_mul_201[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1615:1608] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1615:1608] <= kernel_img_sum_201[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1615:1608] <= 'd0;
end

wire  [39:0]  kernel_img_mul_202[0:24];
assign kernel_img_mul_202[0] = buffer_data_4[1607:1600] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_202[1] = buffer_data_4[1615:1608] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_202[2] = buffer_data_4[1623:1616] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_202[3] = buffer_data_4[1631:1624] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_202[4] = buffer_data_4[1639:1632] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_202[5] = buffer_data_3[1607:1600] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_202[6] = buffer_data_3[1615:1608] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_202[7] = buffer_data_3[1623:1616] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_202[8] = buffer_data_3[1631:1624] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_202[9] = buffer_data_3[1639:1632] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_202[10] = buffer_data_2[1607:1600] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_202[11] = buffer_data_2[1615:1608] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_202[12] = buffer_data_2[1623:1616] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_202[13] = buffer_data_2[1631:1624] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_202[14] = buffer_data_2[1639:1632] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_202[15] = buffer_data_1[1607:1600] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_202[16] = buffer_data_1[1615:1608] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_202[17] = buffer_data_1[1623:1616] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_202[18] = buffer_data_1[1631:1624] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_202[19] = buffer_data_1[1639:1632] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_202[20] = buffer_data_0[1607:1600] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_202[21] = buffer_data_0[1615:1608] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_202[22] = buffer_data_0[1623:1616] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_202[23] = buffer_data_0[1631:1624] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_202[24] = buffer_data_0[1639:1632] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_202 = kernel_img_mul_202[0] + kernel_img_mul_202[1] + kernel_img_mul_202[2] + 
                kernel_img_mul_202[3] + kernel_img_mul_202[4] + kernel_img_mul_202[5] + 
                kernel_img_mul_202[6] + kernel_img_mul_202[7] + kernel_img_mul_202[8] + 
                kernel_img_mul_202[9] + kernel_img_mul_202[10] + kernel_img_mul_202[11] + 
                kernel_img_mul_202[12] + kernel_img_mul_202[13] + kernel_img_mul_202[14] + 
                kernel_img_mul_202[15] + kernel_img_mul_202[16] + kernel_img_mul_202[17] + 
                kernel_img_mul_202[18] + kernel_img_mul_202[19] + kernel_img_mul_202[20] + 
                kernel_img_mul_202[21] + kernel_img_mul_202[22] + kernel_img_mul_202[23] + 
                kernel_img_mul_202[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1623:1616] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1623:1616] <= kernel_img_sum_202[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1623:1616] <= 'd0;
end

wire  [39:0]  kernel_img_mul_203[0:24];
assign kernel_img_mul_203[0] = buffer_data_4[1615:1608] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_203[1] = buffer_data_4[1623:1616] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_203[2] = buffer_data_4[1631:1624] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_203[3] = buffer_data_4[1639:1632] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_203[4] = buffer_data_4[1647:1640] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_203[5] = buffer_data_3[1615:1608] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_203[6] = buffer_data_3[1623:1616] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_203[7] = buffer_data_3[1631:1624] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_203[8] = buffer_data_3[1639:1632] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_203[9] = buffer_data_3[1647:1640] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_203[10] = buffer_data_2[1615:1608] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_203[11] = buffer_data_2[1623:1616] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_203[12] = buffer_data_2[1631:1624] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_203[13] = buffer_data_2[1639:1632] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_203[14] = buffer_data_2[1647:1640] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_203[15] = buffer_data_1[1615:1608] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_203[16] = buffer_data_1[1623:1616] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_203[17] = buffer_data_1[1631:1624] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_203[18] = buffer_data_1[1639:1632] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_203[19] = buffer_data_1[1647:1640] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_203[20] = buffer_data_0[1615:1608] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_203[21] = buffer_data_0[1623:1616] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_203[22] = buffer_data_0[1631:1624] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_203[23] = buffer_data_0[1639:1632] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_203[24] = buffer_data_0[1647:1640] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_203 = kernel_img_mul_203[0] + kernel_img_mul_203[1] + kernel_img_mul_203[2] + 
                kernel_img_mul_203[3] + kernel_img_mul_203[4] + kernel_img_mul_203[5] + 
                kernel_img_mul_203[6] + kernel_img_mul_203[7] + kernel_img_mul_203[8] + 
                kernel_img_mul_203[9] + kernel_img_mul_203[10] + kernel_img_mul_203[11] + 
                kernel_img_mul_203[12] + kernel_img_mul_203[13] + kernel_img_mul_203[14] + 
                kernel_img_mul_203[15] + kernel_img_mul_203[16] + kernel_img_mul_203[17] + 
                kernel_img_mul_203[18] + kernel_img_mul_203[19] + kernel_img_mul_203[20] + 
                kernel_img_mul_203[21] + kernel_img_mul_203[22] + kernel_img_mul_203[23] + 
                kernel_img_mul_203[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1631:1624] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1631:1624] <= kernel_img_sum_203[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1631:1624] <= 'd0;
end

wire  [39:0]  kernel_img_mul_204[0:24];
assign kernel_img_mul_204[0] = buffer_data_4[1623:1616] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_204[1] = buffer_data_4[1631:1624] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_204[2] = buffer_data_4[1639:1632] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_204[3] = buffer_data_4[1647:1640] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_204[4] = buffer_data_4[1655:1648] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_204[5] = buffer_data_3[1623:1616] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_204[6] = buffer_data_3[1631:1624] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_204[7] = buffer_data_3[1639:1632] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_204[8] = buffer_data_3[1647:1640] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_204[9] = buffer_data_3[1655:1648] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_204[10] = buffer_data_2[1623:1616] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_204[11] = buffer_data_2[1631:1624] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_204[12] = buffer_data_2[1639:1632] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_204[13] = buffer_data_2[1647:1640] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_204[14] = buffer_data_2[1655:1648] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_204[15] = buffer_data_1[1623:1616] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_204[16] = buffer_data_1[1631:1624] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_204[17] = buffer_data_1[1639:1632] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_204[18] = buffer_data_1[1647:1640] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_204[19] = buffer_data_1[1655:1648] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_204[20] = buffer_data_0[1623:1616] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_204[21] = buffer_data_0[1631:1624] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_204[22] = buffer_data_0[1639:1632] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_204[23] = buffer_data_0[1647:1640] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_204[24] = buffer_data_0[1655:1648] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_204 = kernel_img_mul_204[0] + kernel_img_mul_204[1] + kernel_img_mul_204[2] + 
                kernel_img_mul_204[3] + kernel_img_mul_204[4] + kernel_img_mul_204[5] + 
                kernel_img_mul_204[6] + kernel_img_mul_204[7] + kernel_img_mul_204[8] + 
                kernel_img_mul_204[9] + kernel_img_mul_204[10] + kernel_img_mul_204[11] + 
                kernel_img_mul_204[12] + kernel_img_mul_204[13] + kernel_img_mul_204[14] + 
                kernel_img_mul_204[15] + kernel_img_mul_204[16] + kernel_img_mul_204[17] + 
                kernel_img_mul_204[18] + kernel_img_mul_204[19] + kernel_img_mul_204[20] + 
                kernel_img_mul_204[21] + kernel_img_mul_204[22] + kernel_img_mul_204[23] + 
                kernel_img_mul_204[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1639:1632] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1639:1632] <= kernel_img_sum_204[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1639:1632] <= 'd0;
end

wire  [39:0]  kernel_img_mul_205[0:24];
assign kernel_img_mul_205[0] = buffer_data_4[1631:1624] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_205[1] = buffer_data_4[1639:1632] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_205[2] = buffer_data_4[1647:1640] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_205[3] = buffer_data_4[1655:1648] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_205[4] = buffer_data_4[1663:1656] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_205[5] = buffer_data_3[1631:1624] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_205[6] = buffer_data_3[1639:1632] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_205[7] = buffer_data_3[1647:1640] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_205[8] = buffer_data_3[1655:1648] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_205[9] = buffer_data_3[1663:1656] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_205[10] = buffer_data_2[1631:1624] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_205[11] = buffer_data_2[1639:1632] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_205[12] = buffer_data_2[1647:1640] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_205[13] = buffer_data_2[1655:1648] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_205[14] = buffer_data_2[1663:1656] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_205[15] = buffer_data_1[1631:1624] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_205[16] = buffer_data_1[1639:1632] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_205[17] = buffer_data_1[1647:1640] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_205[18] = buffer_data_1[1655:1648] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_205[19] = buffer_data_1[1663:1656] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_205[20] = buffer_data_0[1631:1624] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_205[21] = buffer_data_0[1639:1632] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_205[22] = buffer_data_0[1647:1640] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_205[23] = buffer_data_0[1655:1648] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_205[24] = buffer_data_0[1663:1656] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_205 = kernel_img_mul_205[0] + kernel_img_mul_205[1] + kernel_img_mul_205[2] + 
                kernel_img_mul_205[3] + kernel_img_mul_205[4] + kernel_img_mul_205[5] + 
                kernel_img_mul_205[6] + kernel_img_mul_205[7] + kernel_img_mul_205[8] + 
                kernel_img_mul_205[9] + kernel_img_mul_205[10] + kernel_img_mul_205[11] + 
                kernel_img_mul_205[12] + kernel_img_mul_205[13] + kernel_img_mul_205[14] + 
                kernel_img_mul_205[15] + kernel_img_mul_205[16] + kernel_img_mul_205[17] + 
                kernel_img_mul_205[18] + kernel_img_mul_205[19] + kernel_img_mul_205[20] + 
                kernel_img_mul_205[21] + kernel_img_mul_205[22] + kernel_img_mul_205[23] + 
                kernel_img_mul_205[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1647:1640] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1647:1640] <= kernel_img_sum_205[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1647:1640] <= 'd0;
end

wire  [39:0]  kernel_img_mul_206[0:24];
assign kernel_img_mul_206[0] = buffer_data_4[1639:1632] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_206[1] = buffer_data_4[1647:1640] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_206[2] = buffer_data_4[1655:1648] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_206[3] = buffer_data_4[1663:1656] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_206[4] = buffer_data_4[1671:1664] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_206[5] = buffer_data_3[1639:1632] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_206[6] = buffer_data_3[1647:1640] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_206[7] = buffer_data_3[1655:1648] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_206[8] = buffer_data_3[1663:1656] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_206[9] = buffer_data_3[1671:1664] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_206[10] = buffer_data_2[1639:1632] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_206[11] = buffer_data_2[1647:1640] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_206[12] = buffer_data_2[1655:1648] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_206[13] = buffer_data_2[1663:1656] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_206[14] = buffer_data_2[1671:1664] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_206[15] = buffer_data_1[1639:1632] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_206[16] = buffer_data_1[1647:1640] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_206[17] = buffer_data_1[1655:1648] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_206[18] = buffer_data_1[1663:1656] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_206[19] = buffer_data_1[1671:1664] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_206[20] = buffer_data_0[1639:1632] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_206[21] = buffer_data_0[1647:1640] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_206[22] = buffer_data_0[1655:1648] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_206[23] = buffer_data_0[1663:1656] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_206[24] = buffer_data_0[1671:1664] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_206 = kernel_img_mul_206[0] + kernel_img_mul_206[1] + kernel_img_mul_206[2] + 
                kernel_img_mul_206[3] + kernel_img_mul_206[4] + kernel_img_mul_206[5] + 
                kernel_img_mul_206[6] + kernel_img_mul_206[7] + kernel_img_mul_206[8] + 
                kernel_img_mul_206[9] + kernel_img_mul_206[10] + kernel_img_mul_206[11] + 
                kernel_img_mul_206[12] + kernel_img_mul_206[13] + kernel_img_mul_206[14] + 
                kernel_img_mul_206[15] + kernel_img_mul_206[16] + kernel_img_mul_206[17] + 
                kernel_img_mul_206[18] + kernel_img_mul_206[19] + kernel_img_mul_206[20] + 
                kernel_img_mul_206[21] + kernel_img_mul_206[22] + kernel_img_mul_206[23] + 
                kernel_img_mul_206[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1655:1648] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1655:1648] <= kernel_img_sum_206[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1655:1648] <= 'd0;
end

wire  [39:0]  kernel_img_mul_207[0:24];
assign kernel_img_mul_207[0] = buffer_data_4[1647:1640] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_207[1] = buffer_data_4[1655:1648] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_207[2] = buffer_data_4[1663:1656] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_207[3] = buffer_data_4[1671:1664] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_207[4] = buffer_data_4[1679:1672] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_207[5] = buffer_data_3[1647:1640] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_207[6] = buffer_data_3[1655:1648] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_207[7] = buffer_data_3[1663:1656] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_207[8] = buffer_data_3[1671:1664] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_207[9] = buffer_data_3[1679:1672] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_207[10] = buffer_data_2[1647:1640] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_207[11] = buffer_data_2[1655:1648] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_207[12] = buffer_data_2[1663:1656] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_207[13] = buffer_data_2[1671:1664] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_207[14] = buffer_data_2[1679:1672] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_207[15] = buffer_data_1[1647:1640] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_207[16] = buffer_data_1[1655:1648] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_207[17] = buffer_data_1[1663:1656] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_207[18] = buffer_data_1[1671:1664] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_207[19] = buffer_data_1[1679:1672] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_207[20] = buffer_data_0[1647:1640] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_207[21] = buffer_data_0[1655:1648] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_207[22] = buffer_data_0[1663:1656] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_207[23] = buffer_data_0[1671:1664] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_207[24] = buffer_data_0[1679:1672] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_207 = kernel_img_mul_207[0] + kernel_img_mul_207[1] + kernel_img_mul_207[2] + 
                kernel_img_mul_207[3] + kernel_img_mul_207[4] + kernel_img_mul_207[5] + 
                kernel_img_mul_207[6] + kernel_img_mul_207[7] + kernel_img_mul_207[8] + 
                kernel_img_mul_207[9] + kernel_img_mul_207[10] + kernel_img_mul_207[11] + 
                kernel_img_mul_207[12] + kernel_img_mul_207[13] + kernel_img_mul_207[14] + 
                kernel_img_mul_207[15] + kernel_img_mul_207[16] + kernel_img_mul_207[17] + 
                kernel_img_mul_207[18] + kernel_img_mul_207[19] + kernel_img_mul_207[20] + 
                kernel_img_mul_207[21] + kernel_img_mul_207[22] + kernel_img_mul_207[23] + 
                kernel_img_mul_207[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1663:1656] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1663:1656] <= kernel_img_sum_207[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1663:1656] <= 'd0;
end

wire  [39:0]  kernel_img_mul_208[0:24];
assign kernel_img_mul_208[0] = buffer_data_4[1655:1648] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_208[1] = buffer_data_4[1663:1656] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_208[2] = buffer_data_4[1671:1664] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_208[3] = buffer_data_4[1679:1672] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_208[4] = buffer_data_4[1687:1680] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_208[5] = buffer_data_3[1655:1648] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_208[6] = buffer_data_3[1663:1656] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_208[7] = buffer_data_3[1671:1664] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_208[8] = buffer_data_3[1679:1672] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_208[9] = buffer_data_3[1687:1680] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_208[10] = buffer_data_2[1655:1648] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_208[11] = buffer_data_2[1663:1656] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_208[12] = buffer_data_2[1671:1664] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_208[13] = buffer_data_2[1679:1672] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_208[14] = buffer_data_2[1687:1680] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_208[15] = buffer_data_1[1655:1648] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_208[16] = buffer_data_1[1663:1656] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_208[17] = buffer_data_1[1671:1664] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_208[18] = buffer_data_1[1679:1672] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_208[19] = buffer_data_1[1687:1680] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_208[20] = buffer_data_0[1655:1648] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_208[21] = buffer_data_0[1663:1656] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_208[22] = buffer_data_0[1671:1664] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_208[23] = buffer_data_0[1679:1672] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_208[24] = buffer_data_0[1687:1680] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_208 = kernel_img_mul_208[0] + kernel_img_mul_208[1] + kernel_img_mul_208[2] + 
                kernel_img_mul_208[3] + kernel_img_mul_208[4] + kernel_img_mul_208[5] + 
                kernel_img_mul_208[6] + kernel_img_mul_208[7] + kernel_img_mul_208[8] + 
                kernel_img_mul_208[9] + kernel_img_mul_208[10] + kernel_img_mul_208[11] + 
                kernel_img_mul_208[12] + kernel_img_mul_208[13] + kernel_img_mul_208[14] + 
                kernel_img_mul_208[15] + kernel_img_mul_208[16] + kernel_img_mul_208[17] + 
                kernel_img_mul_208[18] + kernel_img_mul_208[19] + kernel_img_mul_208[20] + 
                kernel_img_mul_208[21] + kernel_img_mul_208[22] + kernel_img_mul_208[23] + 
                kernel_img_mul_208[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1671:1664] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1671:1664] <= kernel_img_sum_208[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1671:1664] <= 'd0;
end

wire  [39:0]  kernel_img_mul_209[0:24];
assign kernel_img_mul_209[0] = buffer_data_4[1663:1656] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_209[1] = buffer_data_4[1671:1664] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_209[2] = buffer_data_4[1679:1672] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_209[3] = buffer_data_4[1687:1680] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_209[4] = buffer_data_4[1695:1688] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_209[5] = buffer_data_3[1663:1656] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_209[6] = buffer_data_3[1671:1664] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_209[7] = buffer_data_3[1679:1672] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_209[8] = buffer_data_3[1687:1680] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_209[9] = buffer_data_3[1695:1688] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_209[10] = buffer_data_2[1663:1656] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_209[11] = buffer_data_2[1671:1664] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_209[12] = buffer_data_2[1679:1672] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_209[13] = buffer_data_2[1687:1680] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_209[14] = buffer_data_2[1695:1688] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_209[15] = buffer_data_1[1663:1656] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_209[16] = buffer_data_1[1671:1664] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_209[17] = buffer_data_1[1679:1672] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_209[18] = buffer_data_1[1687:1680] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_209[19] = buffer_data_1[1695:1688] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_209[20] = buffer_data_0[1663:1656] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_209[21] = buffer_data_0[1671:1664] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_209[22] = buffer_data_0[1679:1672] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_209[23] = buffer_data_0[1687:1680] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_209[24] = buffer_data_0[1695:1688] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_209 = kernel_img_mul_209[0] + kernel_img_mul_209[1] + kernel_img_mul_209[2] + 
                kernel_img_mul_209[3] + kernel_img_mul_209[4] + kernel_img_mul_209[5] + 
                kernel_img_mul_209[6] + kernel_img_mul_209[7] + kernel_img_mul_209[8] + 
                kernel_img_mul_209[9] + kernel_img_mul_209[10] + kernel_img_mul_209[11] + 
                kernel_img_mul_209[12] + kernel_img_mul_209[13] + kernel_img_mul_209[14] + 
                kernel_img_mul_209[15] + kernel_img_mul_209[16] + kernel_img_mul_209[17] + 
                kernel_img_mul_209[18] + kernel_img_mul_209[19] + kernel_img_mul_209[20] + 
                kernel_img_mul_209[21] + kernel_img_mul_209[22] + kernel_img_mul_209[23] + 
                kernel_img_mul_209[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1679:1672] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1679:1672] <= kernel_img_sum_209[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1679:1672] <= 'd0;
end

wire  [39:0]  kernel_img_mul_210[0:24];
assign kernel_img_mul_210[0] = buffer_data_4[1671:1664] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_210[1] = buffer_data_4[1679:1672] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_210[2] = buffer_data_4[1687:1680] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_210[3] = buffer_data_4[1695:1688] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_210[4] = buffer_data_4[1703:1696] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_210[5] = buffer_data_3[1671:1664] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_210[6] = buffer_data_3[1679:1672] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_210[7] = buffer_data_3[1687:1680] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_210[8] = buffer_data_3[1695:1688] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_210[9] = buffer_data_3[1703:1696] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_210[10] = buffer_data_2[1671:1664] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_210[11] = buffer_data_2[1679:1672] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_210[12] = buffer_data_2[1687:1680] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_210[13] = buffer_data_2[1695:1688] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_210[14] = buffer_data_2[1703:1696] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_210[15] = buffer_data_1[1671:1664] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_210[16] = buffer_data_1[1679:1672] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_210[17] = buffer_data_1[1687:1680] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_210[18] = buffer_data_1[1695:1688] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_210[19] = buffer_data_1[1703:1696] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_210[20] = buffer_data_0[1671:1664] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_210[21] = buffer_data_0[1679:1672] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_210[22] = buffer_data_0[1687:1680] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_210[23] = buffer_data_0[1695:1688] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_210[24] = buffer_data_0[1703:1696] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_210 = kernel_img_mul_210[0] + kernel_img_mul_210[1] + kernel_img_mul_210[2] + 
                kernel_img_mul_210[3] + kernel_img_mul_210[4] + kernel_img_mul_210[5] + 
                kernel_img_mul_210[6] + kernel_img_mul_210[7] + kernel_img_mul_210[8] + 
                kernel_img_mul_210[9] + kernel_img_mul_210[10] + kernel_img_mul_210[11] + 
                kernel_img_mul_210[12] + kernel_img_mul_210[13] + kernel_img_mul_210[14] + 
                kernel_img_mul_210[15] + kernel_img_mul_210[16] + kernel_img_mul_210[17] + 
                kernel_img_mul_210[18] + kernel_img_mul_210[19] + kernel_img_mul_210[20] + 
                kernel_img_mul_210[21] + kernel_img_mul_210[22] + kernel_img_mul_210[23] + 
                kernel_img_mul_210[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1687:1680] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1687:1680] <= kernel_img_sum_210[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1687:1680] <= 'd0;
end

wire  [39:0]  kernel_img_mul_211[0:24];
assign kernel_img_mul_211[0] = buffer_data_4[1679:1672] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_211[1] = buffer_data_4[1687:1680] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_211[2] = buffer_data_4[1695:1688] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_211[3] = buffer_data_4[1703:1696] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_211[4] = buffer_data_4[1711:1704] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_211[5] = buffer_data_3[1679:1672] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_211[6] = buffer_data_3[1687:1680] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_211[7] = buffer_data_3[1695:1688] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_211[8] = buffer_data_3[1703:1696] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_211[9] = buffer_data_3[1711:1704] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_211[10] = buffer_data_2[1679:1672] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_211[11] = buffer_data_2[1687:1680] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_211[12] = buffer_data_2[1695:1688] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_211[13] = buffer_data_2[1703:1696] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_211[14] = buffer_data_2[1711:1704] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_211[15] = buffer_data_1[1679:1672] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_211[16] = buffer_data_1[1687:1680] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_211[17] = buffer_data_1[1695:1688] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_211[18] = buffer_data_1[1703:1696] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_211[19] = buffer_data_1[1711:1704] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_211[20] = buffer_data_0[1679:1672] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_211[21] = buffer_data_0[1687:1680] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_211[22] = buffer_data_0[1695:1688] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_211[23] = buffer_data_0[1703:1696] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_211[24] = buffer_data_0[1711:1704] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_211 = kernel_img_mul_211[0] + kernel_img_mul_211[1] + kernel_img_mul_211[2] + 
                kernel_img_mul_211[3] + kernel_img_mul_211[4] + kernel_img_mul_211[5] + 
                kernel_img_mul_211[6] + kernel_img_mul_211[7] + kernel_img_mul_211[8] + 
                kernel_img_mul_211[9] + kernel_img_mul_211[10] + kernel_img_mul_211[11] + 
                kernel_img_mul_211[12] + kernel_img_mul_211[13] + kernel_img_mul_211[14] + 
                kernel_img_mul_211[15] + kernel_img_mul_211[16] + kernel_img_mul_211[17] + 
                kernel_img_mul_211[18] + kernel_img_mul_211[19] + kernel_img_mul_211[20] + 
                kernel_img_mul_211[21] + kernel_img_mul_211[22] + kernel_img_mul_211[23] + 
                kernel_img_mul_211[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1695:1688] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1695:1688] <= kernel_img_sum_211[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1695:1688] <= 'd0;
end

wire  [39:0]  kernel_img_mul_212[0:24];
assign kernel_img_mul_212[0] = buffer_data_4[1687:1680] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_212[1] = buffer_data_4[1695:1688] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_212[2] = buffer_data_4[1703:1696] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_212[3] = buffer_data_4[1711:1704] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_212[4] = buffer_data_4[1719:1712] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_212[5] = buffer_data_3[1687:1680] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_212[6] = buffer_data_3[1695:1688] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_212[7] = buffer_data_3[1703:1696] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_212[8] = buffer_data_3[1711:1704] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_212[9] = buffer_data_3[1719:1712] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_212[10] = buffer_data_2[1687:1680] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_212[11] = buffer_data_2[1695:1688] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_212[12] = buffer_data_2[1703:1696] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_212[13] = buffer_data_2[1711:1704] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_212[14] = buffer_data_2[1719:1712] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_212[15] = buffer_data_1[1687:1680] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_212[16] = buffer_data_1[1695:1688] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_212[17] = buffer_data_1[1703:1696] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_212[18] = buffer_data_1[1711:1704] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_212[19] = buffer_data_1[1719:1712] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_212[20] = buffer_data_0[1687:1680] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_212[21] = buffer_data_0[1695:1688] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_212[22] = buffer_data_0[1703:1696] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_212[23] = buffer_data_0[1711:1704] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_212[24] = buffer_data_0[1719:1712] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_212 = kernel_img_mul_212[0] + kernel_img_mul_212[1] + kernel_img_mul_212[2] + 
                kernel_img_mul_212[3] + kernel_img_mul_212[4] + kernel_img_mul_212[5] + 
                kernel_img_mul_212[6] + kernel_img_mul_212[7] + kernel_img_mul_212[8] + 
                kernel_img_mul_212[9] + kernel_img_mul_212[10] + kernel_img_mul_212[11] + 
                kernel_img_mul_212[12] + kernel_img_mul_212[13] + kernel_img_mul_212[14] + 
                kernel_img_mul_212[15] + kernel_img_mul_212[16] + kernel_img_mul_212[17] + 
                kernel_img_mul_212[18] + kernel_img_mul_212[19] + kernel_img_mul_212[20] + 
                kernel_img_mul_212[21] + kernel_img_mul_212[22] + kernel_img_mul_212[23] + 
                kernel_img_mul_212[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1703:1696] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1703:1696] <= kernel_img_sum_212[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1703:1696] <= 'd0;
end

wire  [39:0]  kernel_img_mul_213[0:24];
assign kernel_img_mul_213[0] = buffer_data_4[1695:1688] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_213[1] = buffer_data_4[1703:1696] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_213[2] = buffer_data_4[1711:1704] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_213[3] = buffer_data_4[1719:1712] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_213[4] = buffer_data_4[1727:1720] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_213[5] = buffer_data_3[1695:1688] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_213[6] = buffer_data_3[1703:1696] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_213[7] = buffer_data_3[1711:1704] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_213[8] = buffer_data_3[1719:1712] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_213[9] = buffer_data_3[1727:1720] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_213[10] = buffer_data_2[1695:1688] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_213[11] = buffer_data_2[1703:1696] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_213[12] = buffer_data_2[1711:1704] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_213[13] = buffer_data_2[1719:1712] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_213[14] = buffer_data_2[1727:1720] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_213[15] = buffer_data_1[1695:1688] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_213[16] = buffer_data_1[1703:1696] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_213[17] = buffer_data_1[1711:1704] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_213[18] = buffer_data_1[1719:1712] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_213[19] = buffer_data_1[1727:1720] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_213[20] = buffer_data_0[1695:1688] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_213[21] = buffer_data_0[1703:1696] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_213[22] = buffer_data_0[1711:1704] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_213[23] = buffer_data_0[1719:1712] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_213[24] = buffer_data_0[1727:1720] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_213 = kernel_img_mul_213[0] + kernel_img_mul_213[1] + kernel_img_mul_213[2] + 
                kernel_img_mul_213[3] + kernel_img_mul_213[4] + kernel_img_mul_213[5] + 
                kernel_img_mul_213[6] + kernel_img_mul_213[7] + kernel_img_mul_213[8] + 
                kernel_img_mul_213[9] + kernel_img_mul_213[10] + kernel_img_mul_213[11] + 
                kernel_img_mul_213[12] + kernel_img_mul_213[13] + kernel_img_mul_213[14] + 
                kernel_img_mul_213[15] + kernel_img_mul_213[16] + kernel_img_mul_213[17] + 
                kernel_img_mul_213[18] + kernel_img_mul_213[19] + kernel_img_mul_213[20] + 
                kernel_img_mul_213[21] + kernel_img_mul_213[22] + kernel_img_mul_213[23] + 
                kernel_img_mul_213[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1711:1704] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1711:1704] <= kernel_img_sum_213[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1711:1704] <= 'd0;
end

wire  [39:0]  kernel_img_mul_214[0:24];
assign kernel_img_mul_214[0] = buffer_data_4[1703:1696] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_214[1] = buffer_data_4[1711:1704] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_214[2] = buffer_data_4[1719:1712] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_214[3] = buffer_data_4[1727:1720] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_214[4] = buffer_data_4[1735:1728] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_214[5] = buffer_data_3[1703:1696] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_214[6] = buffer_data_3[1711:1704] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_214[7] = buffer_data_3[1719:1712] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_214[8] = buffer_data_3[1727:1720] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_214[9] = buffer_data_3[1735:1728] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_214[10] = buffer_data_2[1703:1696] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_214[11] = buffer_data_2[1711:1704] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_214[12] = buffer_data_2[1719:1712] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_214[13] = buffer_data_2[1727:1720] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_214[14] = buffer_data_2[1735:1728] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_214[15] = buffer_data_1[1703:1696] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_214[16] = buffer_data_1[1711:1704] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_214[17] = buffer_data_1[1719:1712] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_214[18] = buffer_data_1[1727:1720] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_214[19] = buffer_data_1[1735:1728] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_214[20] = buffer_data_0[1703:1696] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_214[21] = buffer_data_0[1711:1704] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_214[22] = buffer_data_0[1719:1712] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_214[23] = buffer_data_0[1727:1720] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_214[24] = buffer_data_0[1735:1728] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_214 = kernel_img_mul_214[0] + kernel_img_mul_214[1] + kernel_img_mul_214[2] + 
                kernel_img_mul_214[3] + kernel_img_mul_214[4] + kernel_img_mul_214[5] + 
                kernel_img_mul_214[6] + kernel_img_mul_214[7] + kernel_img_mul_214[8] + 
                kernel_img_mul_214[9] + kernel_img_mul_214[10] + kernel_img_mul_214[11] + 
                kernel_img_mul_214[12] + kernel_img_mul_214[13] + kernel_img_mul_214[14] + 
                kernel_img_mul_214[15] + kernel_img_mul_214[16] + kernel_img_mul_214[17] + 
                kernel_img_mul_214[18] + kernel_img_mul_214[19] + kernel_img_mul_214[20] + 
                kernel_img_mul_214[21] + kernel_img_mul_214[22] + kernel_img_mul_214[23] + 
                kernel_img_mul_214[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1719:1712] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1719:1712] <= kernel_img_sum_214[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1719:1712] <= 'd0;
end

wire  [39:0]  kernel_img_mul_215[0:24];
assign kernel_img_mul_215[0] = buffer_data_4[1711:1704] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_215[1] = buffer_data_4[1719:1712] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_215[2] = buffer_data_4[1727:1720] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_215[3] = buffer_data_4[1735:1728] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_215[4] = buffer_data_4[1743:1736] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_215[5] = buffer_data_3[1711:1704] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_215[6] = buffer_data_3[1719:1712] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_215[7] = buffer_data_3[1727:1720] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_215[8] = buffer_data_3[1735:1728] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_215[9] = buffer_data_3[1743:1736] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_215[10] = buffer_data_2[1711:1704] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_215[11] = buffer_data_2[1719:1712] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_215[12] = buffer_data_2[1727:1720] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_215[13] = buffer_data_2[1735:1728] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_215[14] = buffer_data_2[1743:1736] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_215[15] = buffer_data_1[1711:1704] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_215[16] = buffer_data_1[1719:1712] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_215[17] = buffer_data_1[1727:1720] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_215[18] = buffer_data_1[1735:1728] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_215[19] = buffer_data_1[1743:1736] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_215[20] = buffer_data_0[1711:1704] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_215[21] = buffer_data_0[1719:1712] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_215[22] = buffer_data_0[1727:1720] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_215[23] = buffer_data_0[1735:1728] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_215[24] = buffer_data_0[1743:1736] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_215 = kernel_img_mul_215[0] + kernel_img_mul_215[1] + kernel_img_mul_215[2] + 
                kernel_img_mul_215[3] + kernel_img_mul_215[4] + kernel_img_mul_215[5] + 
                kernel_img_mul_215[6] + kernel_img_mul_215[7] + kernel_img_mul_215[8] + 
                kernel_img_mul_215[9] + kernel_img_mul_215[10] + kernel_img_mul_215[11] + 
                kernel_img_mul_215[12] + kernel_img_mul_215[13] + kernel_img_mul_215[14] + 
                kernel_img_mul_215[15] + kernel_img_mul_215[16] + kernel_img_mul_215[17] + 
                kernel_img_mul_215[18] + kernel_img_mul_215[19] + kernel_img_mul_215[20] + 
                kernel_img_mul_215[21] + kernel_img_mul_215[22] + kernel_img_mul_215[23] + 
                kernel_img_mul_215[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1727:1720] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1727:1720] <= kernel_img_sum_215[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1727:1720] <= 'd0;
end

wire  [39:0]  kernel_img_mul_216[0:24];
assign kernel_img_mul_216[0] = buffer_data_4[1719:1712] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_216[1] = buffer_data_4[1727:1720] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_216[2] = buffer_data_4[1735:1728] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_216[3] = buffer_data_4[1743:1736] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_216[4] = buffer_data_4[1751:1744] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_216[5] = buffer_data_3[1719:1712] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_216[6] = buffer_data_3[1727:1720] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_216[7] = buffer_data_3[1735:1728] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_216[8] = buffer_data_3[1743:1736] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_216[9] = buffer_data_3[1751:1744] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_216[10] = buffer_data_2[1719:1712] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_216[11] = buffer_data_2[1727:1720] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_216[12] = buffer_data_2[1735:1728] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_216[13] = buffer_data_2[1743:1736] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_216[14] = buffer_data_2[1751:1744] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_216[15] = buffer_data_1[1719:1712] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_216[16] = buffer_data_1[1727:1720] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_216[17] = buffer_data_1[1735:1728] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_216[18] = buffer_data_1[1743:1736] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_216[19] = buffer_data_1[1751:1744] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_216[20] = buffer_data_0[1719:1712] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_216[21] = buffer_data_0[1727:1720] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_216[22] = buffer_data_0[1735:1728] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_216[23] = buffer_data_0[1743:1736] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_216[24] = buffer_data_0[1751:1744] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_216 = kernel_img_mul_216[0] + kernel_img_mul_216[1] + kernel_img_mul_216[2] + 
                kernel_img_mul_216[3] + kernel_img_mul_216[4] + kernel_img_mul_216[5] + 
                kernel_img_mul_216[6] + kernel_img_mul_216[7] + kernel_img_mul_216[8] + 
                kernel_img_mul_216[9] + kernel_img_mul_216[10] + kernel_img_mul_216[11] + 
                kernel_img_mul_216[12] + kernel_img_mul_216[13] + kernel_img_mul_216[14] + 
                kernel_img_mul_216[15] + kernel_img_mul_216[16] + kernel_img_mul_216[17] + 
                kernel_img_mul_216[18] + kernel_img_mul_216[19] + kernel_img_mul_216[20] + 
                kernel_img_mul_216[21] + kernel_img_mul_216[22] + kernel_img_mul_216[23] + 
                kernel_img_mul_216[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1735:1728] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1735:1728] <= kernel_img_sum_216[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1735:1728] <= 'd0;
end

wire  [39:0]  kernel_img_mul_217[0:24];
assign kernel_img_mul_217[0] = buffer_data_4[1727:1720] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_217[1] = buffer_data_4[1735:1728] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_217[2] = buffer_data_4[1743:1736] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_217[3] = buffer_data_4[1751:1744] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_217[4] = buffer_data_4[1759:1752] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_217[5] = buffer_data_3[1727:1720] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_217[6] = buffer_data_3[1735:1728] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_217[7] = buffer_data_3[1743:1736] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_217[8] = buffer_data_3[1751:1744] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_217[9] = buffer_data_3[1759:1752] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_217[10] = buffer_data_2[1727:1720] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_217[11] = buffer_data_2[1735:1728] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_217[12] = buffer_data_2[1743:1736] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_217[13] = buffer_data_2[1751:1744] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_217[14] = buffer_data_2[1759:1752] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_217[15] = buffer_data_1[1727:1720] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_217[16] = buffer_data_1[1735:1728] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_217[17] = buffer_data_1[1743:1736] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_217[18] = buffer_data_1[1751:1744] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_217[19] = buffer_data_1[1759:1752] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_217[20] = buffer_data_0[1727:1720] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_217[21] = buffer_data_0[1735:1728] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_217[22] = buffer_data_0[1743:1736] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_217[23] = buffer_data_0[1751:1744] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_217[24] = buffer_data_0[1759:1752] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_217 = kernel_img_mul_217[0] + kernel_img_mul_217[1] + kernel_img_mul_217[2] + 
                kernel_img_mul_217[3] + kernel_img_mul_217[4] + kernel_img_mul_217[5] + 
                kernel_img_mul_217[6] + kernel_img_mul_217[7] + kernel_img_mul_217[8] + 
                kernel_img_mul_217[9] + kernel_img_mul_217[10] + kernel_img_mul_217[11] + 
                kernel_img_mul_217[12] + kernel_img_mul_217[13] + kernel_img_mul_217[14] + 
                kernel_img_mul_217[15] + kernel_img_mul_217[16] + kernel_img_mul_217[17] + 
                kernel_img_mul_217[18] + kernel_img_mul_217[19] + kernel_img_mul_217[20] + 
                kernel_img_mul_217[21] + kernel_img_mul_217[22] + kernel_img_mul_217[23] + 
                kernel_img_mul_217[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1743:1736] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1743:1736] <= kernel_img_sum_217[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1743:1736] <= 'd0;
end

wire  [39:0]  kernel_img_mul_218[0:24];
assign kernel_img_mul_218[0] = buffer_data_4[1735:1728] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_218[1] = buffer_data_4[1743:1736] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_218[2] = buffer_data_4[1751:1744] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_218[3] = buffer_data_4[1759:1752] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_218[4] = buffer_data_4[1767:1760] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_218[5] = buffer_data_3[1735:1728] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_218[6] = buffer_data_3[1743:1736] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_218[7] = buffer_data_3[1751:1744] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_218[8] = buffer_data_3[1759:1752] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_218[9] = buffer_data_3[1767:1760] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_218[10] = buffer_data_2[1735:1728] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_218[11] = buffer_data_2[1743:1736] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_218[12] = buffer_data_2[1751:1744] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_218[13] = buffer_data_2[1759:1752] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_218[14] = buffer_data_2[1767:1760] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_218[15] = buffer_data_1[1735:1728] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_218[16] = buffer_data_1[1743:1736] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_218[17] = buffer_data_1[1751:1744] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_218[18] = buffer_data_1[1759:1752] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_218[19] = buffer_data_1[1767:1760] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_218[20] = buffer_data_0[1735:1728] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_218[21] = buffer_data_0[1743:1736] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_218[22] = buffer_data_0[1751:1744] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_218[23] = buffer_data_0[1759:1752] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_218[24] = buffer_data_0[1767:1760] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_218 = kernel_img_mul_218[0] + kernel_img_mul_218[1] + kernel_img_mul_218[2] + 
                kernel_img_mul_218[3] + kernel_img_mul_218[4] + kernel_img_mul_218[5] + 
                kernel_img_mul_218[6] + kernel_img_mul_218[7] + kernel_img_mul_218[8] + 
                kernel_img_mul_218[9] + kernel_img_mul_218[10] + kernel_img_mul_218[11] + 
                kernel_img_mul_218[12] + kernel_img_mul_218[13] + kernel_img_mul_218[14] + 
                kernel_img_mul_218[15] + kernel_img_mul_218[16] + kernel_img_mul_218[17] + 
                kernel_img_mul_218[18] + kernel_img_mul_218[19] + kernel_img_mul_218[20] + 
                kernel_img_mul_218[21] + kernel_img_mul_218[22] + kernel_img_mul_218[23] + 
                kernel_img_mul_218[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1751:1744] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1751:1744] <= kernel_img_sum_218[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1751:1744] <= 'd0;
end

wire  [39:0]  kernel_img_mul_219[0:24];
assign kernel_img_mul_219[0] = buffer_data_4[1743:1736] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_219[1] = buffer_data_4[1751:1744] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_219[2] = buffer_data_4[1759:1752] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_219[3] = buffer_data_4[1767:1760] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_219[4] = buffer_data_4[1775:1768] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_219[5] = buffer_data_3[1743:1736] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_219[6] = buffer_data_3[1751:1744] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_219[7] = buffer_data_3[1759:1752] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_219[8] = buffer_data_3[1767:1760] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_219[9] = buffer_data_3[1775:1768] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_219[10] = buffer_data_2[1743:1736] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_219[11] = buffer_data_2[1751:1744] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_219[12] = buffer_data_2[1759:1752] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_219[13] = buffer_data_2[1767:1760] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_219[14] = buffer_data_2[1775:1768] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_219[15] = buffer_data_1[1743:1736] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_219[16] = buffer_data_1[1751:1744] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_219[17] = buffer_data_1[1759:1752] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_219[18] = buffer_data_1[1767:1760] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_219[19] = buffer_data_1[1775:1768] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_219[20] = buffer_data_0[1743:1736] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_219[21] = buffer_data_0[1751:1744] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_219[22] = buffer_data_0[1759:1752] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_219[23] = buffer_data_0[1767:1760] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_219[24] = buffer_data_0[1775:1768] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_219 = kernel_img_mul_219[0] + kernel_img_mul_219[1] + kernel_img_mul_219[2] + 
                kernel_img_mul_219[3] + kernel_img_mul_219[4] + kernel_img_mul_219[5] + 
                kernel_img_mul_219[6] + kernel_img_mul_219[7] + kernel_img_mul_219[8] + 
                kernel_img_mul_219[9] + kernel_img_mul_219[10] + kernel_img_mul_219[11] + 
                kernel_img_mul_219[12] + kernel_img_mul_219[13] + kernel_img_mul_219[14] + 
                kernel_img_mul_219[15] + kernel_img_mul_219[16] + kernel_img_mul_219[17] + 
                kernel_img_mul_219[18] + kernel_img_mul_219[19] + kernel_img_mul_219[20] + 
                kernel_img_mul_219[21] + kernel_img_mul_219[22] + kernel_img_mul_219[23] + 
                kernel_img_mul_219[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1759:1752] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1759:1752] <= kernel_img_sum_219[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1759:1752] <= 'd0;
end

wire  [39:0]  kernel_img_mul_220[0:24];
assign kernel_img_mul_220[0] = buffer_data_4[1751:1744] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_220[1] = buffer_data_4[1759:1752] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_220[2] = buffer_data_4[1767:1760] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_220[3] = buffer_data_4[1775:1768] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_220[4] = buffer_data_4[1783:1776] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_220[5] = buffer_data_3[1751:1744] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_220[6] = buffer_data_3[1759:1752] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_220[7] = buffer_data_3[1767:1760] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_220[8] = buffer_data_3[1775:1768] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_220[9] = buffer_data_3[1783:1776] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_220[10] = buffer_data_2[1751:1744] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_220[11] = buffer_data_2[1759:1752] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_220[12] = buffer_data_2[1767:1760] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_220[13] = buffer_data_2[1775:1768] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_220[14] = buffer_data_2[1783:1776] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_220[15] = buffer_data_1[1751:1744] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_220[16] = buffer_data_1[1759:1752] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_220[17] = buffer_data_1[1767:1760] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_220[18] = buffer_data_1[1775:1768] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_220[19] = buffer_data_1[1783:1776] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_220[20] = buffer_data_0[1751:1744] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_220[21] = buffer_data_0[1759:1752] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_220[22] = buffer_data_0[1767:1760] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_220[23] = buffer_data_0[1775:1768] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_220[24] = buffer_data_0[1783:1776] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_220 = kernel_img_mul_220[0] + kernel_img_mul_220[1] + kernel_img_mul_220[2] + 
                kernel_img_mul_220[3] + kernel_img_mul_220[4] + kernel_img_mul_220[5] + 
                kernel_img_mul_220[6] + kernel_img_mul_220[7] + kernel_img_mul_220[8] + 
                kernel_img_mul_220[9] + kernel_img_mul_220[10] + kernel_img_mul_220[11] + 
                kernel_img_mul_220[12] + kernel_img_mul_220[13] + kernel_img_mul_220[14] + 
                kernel_img_mul_220[15] + kernel_img_mul_220[16] + kernel_img_mul_220[17] + 
                kernel_img_mul_220[18] + kernel_img_mul_220[19] + kernel_img_mul_220[20] + 
                kernel_img_mul_220[21] + kernel_img_mul_220[22] + kernel_img_mul_220[23] + 
                kernel_img_mul_220[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1767:1760] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1767:1760] <= kernel_img_sum_220[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1767:1760] <= 'd0;
end

wire  [39:0]  kernel_img_mul_221[0:24];
assign kernel_img_mul_221[0] = buffer_data_4[1759:1752] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_221[1] = buffer_data_4[1767:1760] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_221[2] = buffer_data_4[1775:1768] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_221[3] = buffer_data_4[1783:1776] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_221[4] = buffer_data_4[1791:1784] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_221[5] = buffer_data_3[1759:1752] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_221[6] = buffer_data_3[1767:1760] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_221[7] = buffer_data_3[1775:1768] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_221[8] = buffer_data_3[1783:1776] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_221[9] = buffer_data_3[1791:1784] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_221[10] = buffer_data_2[1759:1752] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_221[11] = buffer_data_2[1767:1760] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_221[12] = buffer_data_2[1775:1768] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_221[13] = buffer_data_2[1783:1776] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_221[14] = buffer_data_2[1791:1784] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_221[15] = buffer_data_1[1759:1752] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_221[16] = buffer_data_1[1767:1760] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_221[17] = buffer_data_1[1775:1768] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_221[18] = buffer_data_1[1783:1776] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_221[19] = buffer_data_1[1791:1784] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_221[20] = buffer_data_0[1759:1752] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_221[21] = buffer_data_0[1767:1760] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_221[22] = buffer_data_0[1775:1768] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_221[23] = buffer_data_0[1783:1776] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_221[24] = buffer_data_0[1791:1784] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_221 = kernel_img_mul_221[0] + kernel_img_mul_221[1] + kernel_img_mul_221[2] + 
                kernel_img_mul_221[3] + kernel_img_mul_221[4] + kernel_img_mul_221[5] + 
                kernel_img_mul_221[6] + kernel_img_mul_221[7] + kernel_img_mul_221[8] + 
                kernel_img_mul_221[9] + kernel_img_mul_221[10] + kernel_img_mul_221[11] + 
                kernel_img_mul_221[12] + kernel_img_mul_221[13] + kernel_img_mul_221[14] + 
                kernel_img_mul_221[15] + kernel_img_mul_221[16] + kernel_img_mul_221[17] + 
                kernel_img_mul_221[18] + kernel_img_mul_221[19] + kernel_img_mul_221[20] + 
                kernel_img_mul_221[21] + kernel_img_mul_221[22] + kernel_img_mul_221[23] + 
                kernel_img_mul_221[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1775:1768] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1775:1768] <= kernel_img_sum_221[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1775:1768] <= 'd0;
end

wire  [39:0]  kernel_img_mul_222[0:24];
assign kernel_img_mul_222[0] = buffer_data_4[1767:1760] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_222[1] = buffer_data_4[1775:1768] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_222[2] = buffer_data_4[1783:1776] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_222[3] = buffer_data_4[1791:1784] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_222[4] = buffer_data_4[1799:1792] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_222[5] = buffer_data_3[1767:1760] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_222[6] = buffer_data_3[1775:1768] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_222[7] = buffer_data_3[1783:1776] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_222[8] = buffer_data_3[1791:1784] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_222[9] = buffer_data_3[1799:1792] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_222[10] = buffer_data_2[1767:1760] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_222[11] = buffer_data_2[1775:1768] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_222[12] = buffer_data_2[1783:1776] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_222[13] = buffer_data_2[1791:1784] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_222[14] = buffer_data_2[1799:1792] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_222[15] = buffer_data_1[1767:1760] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_222[16] = buffer_data_1[1775:1768] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_222[17] = buffer_data_1[1783:1776] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_222[18] = buffer_data_1[1791:1784] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_222[19] = buffer_data_1[1799:1792] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_222[20] = buffer_data_0[1767:1760] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_222[21] = buffer_data_0[1775:1768] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_222[22] = buffer_data_0[1783:1776] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_222[23] = buffer_data_0[1791:1784] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_222[24] = buffer_data_0[1799:1792] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_222 = kernel_img_mul_222[0] + kernel_img_mul_222[1] + kernel_img_mul_222[2] + 
                kernel_img_mul_222[3] + kernel_img_mul_222[4] + kernel_img_mul_222[5] + 
                kernel_img_mul_222[6] + kernel_img_mul_222[7] + kernel_img_mul_222[8] + 
                kernel_img_mul_222[9] + kernel_img_mul_222[10] + kernel_img_mul_222[11] + 
                kernel_img_mul_222[12] + kernel_img_mul_222[13] + kernel_img_mul_222[14] + 
                kernel_img_mul_222[15] + kernel_img_mul_222[16] + kernel_img_mul_222[17] + 
                kernel_img_mul_222[18] + kernel_img_mul_222[19] + kernel_img_mul_222[20] + 
                kernel_img_mul_222[21] + kernel_img_mul_222[22] + kernel_img_mul_222[23] + 
                kernel_img_mul_222[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1783:1776] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1783:1776] <= kernel_img_sum_222[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1783:1776] <= 'd0;
end

wire  [39:0]  kernel_img_mul_223[0:24];
assign kernel_img_mul_223[0] = buffer_data_4[1775:1768] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_223[1] = buffer_data_4[1783:1776] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_223[2] = buffer_data_4[1791:1784] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_223[3] = buffer_data_4[1799:1792] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_223[4] = buffer_data_4[1807:1800] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_223[5] = buffer_data_3[1775:1768] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_223[6] = buffer_data_3[1783:1776] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_223[7] = buffer_data_3[1791:1784] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_223[8] = buffer_data_3[1799:1792] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_223[9] = buffer_data_3[1807:1800] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_223[10] = buffer_data_2[1775:1768] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_223[11] = buffer_data_2[1783:1776] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_223[12] = buffer_data_2[1791:1784] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_223[13] = buffer_data_2[1799:1792] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_223[14] = buffer_data_2[1807:1800] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_223[15] = buffer_data_1[1775:1768] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_223[16] = buffer_data_1[1783:1776] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_223[17] = buffer_data_1[1791:1784] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_223[18] = buffer_data_1[1799:1792] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_223[19] = buffer_data_1[1807:1800] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_223[20] = buffer_data_0[1775:1768] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_223[21] = buffer_data_0[1783:1776] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_223[22] = buffer_data_0[1791:1784] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_223[23] = buffer_data_0[1799:1792] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_223[24] = buffer_data_0[1807:1800] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_223 = kernel_img_mul_223[0] + kernel_img_mul_223[1] + kernel_img_mul_223[2] + 
                kernel_img_mul_223[3] + kernel_img_mul_223[4] + kernel_img_mul_223[5] + 
                kernel_img_mul_223[6] + kernel_img_mul_223[7] + kernel_img_mul_223[8] + 
                kernel_img_mul_223[9] + kernel_img_mul_223[10] + kernel_img_mul_223[11] + 
                kernel_img_mul_223[12] + kernel_img_mul_223[13] + kernel_img_mul_223[14] + 
                kernel_img_mul_223[15] + kernel_img_mul_223[16] + kernel_img_mul_223[17] + 
                kernel_img_mul_223[18] + kernel_img_mul_223[19] + kernel_img_mul_223[20] + 
                kernel_img_mul_223[21] + kernel_img_mul_223[22] + kernel_img_mul_223[23] + 
                kernel_img_mul_223[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1791:1784] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1791:1784] <= kernel_img_sum_223[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1791:1784] <= 'd0;
end

wire  [39:0]  kernel_img_mul_224[0:24];
assign kernel_img_mul_224[0] = buffer_data_4[1783:1776] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_224[1] = buffer_data_4[1791:1784] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_224[2] = buffer_data_4[1799:1792] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_224[3] = buffer_data_4[1807:1800] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_224[4] = buffer_data_4[1815:1808] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_224[5] = buffer_data_3[1783:1776] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_224[6] = buffer_data_3[1791:1784] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_224[7] = buffer_data_3[1799:1792] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_224[8] = buffer_data_3[1807:1800] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_224[9] = buffer_data_3[1815:1808] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_224[10] = buffer_data_2[1783:1776] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_224[11] = buffer_data_2[1791:1784] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_224[12] = buffer_data_2[1799:1792] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_224[13] = buffer_data_2[1807:1800] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_224[14] = buffer_data_2[1815:1808] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_224[15] = buffer_data_1[1783:1776] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_224[16] = buffer_data_1[1791:1784] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_224[17] = buffer_data_1[1799:1792] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_224[18] = buffer_data_1[1807:1800] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_224[19] = buffer_data_1[1815:1808] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_224[20] = buffer_data_0[1783:1776] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_224[21] = buffer_data_0[1791:1784] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_224[22] = buffer_data_0[1799:1792] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_224[23] = buffer_data_0[1807:1800] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_224[24] = buffer_data_0[1815:1808] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_224 = kernel_img_mul_224[0] + kernel_img_mul_224[1] + kernel_img_mul_224[2] + 
                kernel_img_mul_224[3] + kernel_img_mul_224[4] + kernel_img_mul_224[5] + 
                kernel_img_mul_224[6] + kernel_img_mul_224[7] + kernel_img_mul_224[8] + 
                kernel_img_mul_224[9] + kernel_img_mul_224[10] + kernel_img_mul_224[11] + 
                kernel_img_mul_224[12] + kernel_img_mul_224[13] + kernel_img_mul_224[14] + 
                kernel_img_mul_224[15] + kernel_img_mul_224[16] + kernel_img_mul_224[17] + 
                kernel_img_mul_224[18] + kernel_img_mul_224[19] + kernel_img_mul_224[20] + 
                kernel_img_mul_224[21] + kernel_img_mul_224[22] + kernel_img_mul_224[23] + 
                kernel_img_mul_224[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1799:1792] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1799:1792] <= kernel_img_sum_224[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1799:1792] <= 'd0;
end

wire  [39:0]  kernel_img_mul_225[0:24];
assign kernel_img_mul_225[0] = buffer_data_4[1791:1784] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_225[1] = buffer_data_4[1799:1792] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_225[2] = buffer_data_4[1807:1800] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_225[3] = buffer_data_4[1815:1808] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_225[4] = buffer_data_4[1823:1816] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_225[5] = buffer_data_3[1791:1784] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_225[6] = buffer_data_3[1799:1792] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_225[7] = buffer_data_3[1807:1800] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_225[8] = buffer_data_3[1815:1808] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_225[9] = buffer_data_3[1823:1816] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_225[10] = buffer_data_2[1791:1784] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_225[11] = buffer_data_2[1799:1792] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_225[12] = buffer_data_2[1807:1800] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_225[13] = buffer_data_2[1815:1808] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_225[14] = buffer_data_2[1823:1816] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_225[15] = buffer_data_1[1791:1784] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_225[16] = buffer_data_1[1799:1792] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_225[17] = buffer_data_1[1807:1800] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_225[18] = buffer_data_1[1815:1808] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_225[19] = buffer_data_1[1823:1816] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_225[20] = buffer_data_0[1791:1784] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_225[21] = buffer_data_0[1799:1792] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_225[22] = buffer_data_0[1807:1800] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_225[23] = buffer_data_0[1815:1808] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_225[24] = buffer_data_0[1823:1816] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_225 = kernel_img_mul_225[0] + kernel_img_mul_225[1] + kernel_img_mul_225[2] + 
                kernel_img_mul_225[3] + kernel_img_mul_225[4] + kernel_img_mul_225[5] + 
                kernel_img_mul_225[6] + kernel_img_mul_225[7] + kernel_img_mul_225[8] + 
                kernel_img_mul_225[9] + kernel_img_mul_225[10] + kernel_img_mul_225[11] + 
                kernel_img_mul_225[12] + kernel_img_mul_225[13] + kernel_img_mul_225[14] + 
                kernel_img_mul_225[15] + kernel_img_mul_225[16] + kernel_img_mul_225[17] + 
                kernel_img_mul_225[18] + kernel_img_mul_225[19] + kernel_img_mul_225[20] + 
                kernel_img_mul_225[21] + kernel_img_mul_225[22] + kernel_img_mul_225[23] + 
                kernel_img_mul_225[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1807:1800] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1807:1800] <= kernel_img_sum_225[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1807:1800] <= 'd0;
end

wire  [39:0]  kernel_img_mul_226[0:24];
assign kernel_img_mul_226[0] = buffer_data_4[1799:1792] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_226[1] = buffer_data_4[1807:1800] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_226[2] = buffer_data_4[1815:1808] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_226[3] = buffer_data_4[1823:1816] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_226[4] = buffer_data_4[1831:1824] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_226[5] = buffer_data_3[1799:1792] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_226[6] = buffer_data_3[1807:1800] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_226[7] = buffer_data_3[1815:1808] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_226[8] = buffer_data_3[1823:1816] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_226[9] = buffer_data_3[1831:1824] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_226[10] = buffer_data_2[1799:1792] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_226[11] = buffer_data_2[1807:1800] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_226[12] = buffer_data_2[1815:1808] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_226[13] = buffer_data_2[1823:1816] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_226[14] = buffer_data_2[1831:1824] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_226[15] = buffer_data_1[1799:1792] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_226[16] = buffer_data_1[1807:1800] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_226[17] = buffer_data_1[1815:1808] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_226[18] = buffer_data_1[1823:1816] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_226[19] = buffer_data_1[1831:1824] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_226[20] = buffer_data_0[1799:1792] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_226[21] = buffer_data_0[1807:1800] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_226[22] = buffer_data_0[1815:1808] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_226[23] = buffer_data_0[1823:1816] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_226[24] = buffer_data_0[1831:1824] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_226 = kernel_img_mul_226[0] + kernel_img_mul_226[1] + kernel_img_mul_226[2] + 
                kernel_img_mul_226[3] + kernel_img_mul_226[4] + kernel_img_mul_226[5] + 
                kernel_img_mul_226[6] + kernel_img_mul_226[7] + kernel_img_mul_226[8] + 
                kernel_img_mul_226[9] + kernel_img_mul_226[10] + kernel_img_mul_226[11] + 
                kernel_img_mul_226[12] + kernel_img_mul_226[13] + kernel_img_mul_226[14] + 
                kernel_img_mul_226[15] + kernel_img_mul_226[16] + kernel_img_mul_226[17] + 
                kernel_img_mul_226[18] + kernel_img_mul_226[19] + kernel_img_mul_226[20] + 
                kernel_img_mul_226[21] + kernel_img_mul_226[22] + kernel_img_mul_226[23] + 
                kernel_img_mul_226[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1815:1808] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1815:1808] <= kernel_img_sum_226[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1815:1808] <= 'd0;
end

wire  [39:0]  kernel_img_mul_227[0:24];
assign kernel_img_mul_227[0] = buffer_data_4[1807:1800] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_227[1] = buffer_data_4[1815:1808] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_227[2] = buffer_data_4[1823:1816] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_227[3] = buffer_data_4[1831:1824] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_227[4] = buffer_data_4[1839:1832] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_227[5] = buffer_data_3[1807:1800] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_227[6] = buffer_data_3[1815:1808] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_227[7] = buffer_data_3[1823:1816] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_227[8] = buffer_data_3[1831:1824] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_227[9] = buffer_data_3[1839:1832] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_227[10] = buffer_data_2[1807:1800] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_227[11] = buffer_data_2[1815:1808] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_227[12] = buffer_data_2[1823:1816] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_227[13] = buffer_data_2[1831:1824] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_227[14] = buffer_data_2[1839:1832] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_227[15] = buffer_data_1[1807:1800] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_227[16] = buffer_data_1[1815:1808] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_227[17] = buffer_data_1[1823:1816] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_227[18] = buffer_data_1[1831:1824] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_227[19] = buffer_data_1[1839:1832] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_227[20] = buffer_data_0[1807:1800] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_227[21] = buffer_data_0[1815:1808] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_227[22] = buffer_data_0[1823:1816] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_227[23] = buffer_data_0[1831:1824] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_227[24] = buffer_data_0[1839:1832] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_227 = kernel_img_mul_227[0] + kernel_img_mul_227[1] + kernel_img_mul_227[2] + 
                kernel_img_mul_227[3] + kernel_img_mul_227[4] + kernel_img_mul_227[5] + 
                kernel_img_mul_227[6] + kernel_img_mul_227[7] + kernel_img_mul_227[8] + 
                kernel_img_mul_227[9] + kernel_img_mul_227[10] + kernel_img_mul_227[11] + 
                kernel_img_mul_227[12] + kernel_img_mul_227[13] + kernel_img_mul_227[14] + 
                kernel_img_mul_227[15] + kernel_img_mul_227[16] + kernel_img_mul_227[17] + 
                kernel_img_mul_227[18] + kernel_img_mul_227[19] + kernel_img_mul_227[20] + 
                kernel_img_mul_227[21] + kernel_img_mul_227[22] + kernel_img_mul_227[23] + 
                kernel_img_mul_227[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1823:1816] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1823:1816] <= kernel_img_sum_227[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1823:1816] <= 'd0;
end

wire  [39:0]  kernel_img_mul_228[0:24];
assign kernel_img_mul_228[0] = buffer_data_4[1815:1808] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_228[1] = buffer_data_4[1823:1816] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_228[2] = buffer_data_4[1831:1824] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_228[3] = buffer_data_4[1839:1832] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_228[4] = buffer_data_4[1847:1840] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_228[5] = buffer_data_3[1815:1808] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_228[6] = buffer_data_3[1823:1816] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_228[7] = buffer_data_3[1831:1824] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_228[8] = buffer_data_3[1839:1832] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_228[9] = buffer_data_3[1847:1840] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_228[10] = buffer_data_2[1815:1808] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_228[11] = buffer_data_2[1823:1816] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_228[12] = buffer_data_2[1831:1824] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_228[13] = buffer_data_2[1839:1832] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_228[14] = buffer_data_2[1847:1840] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_228[15] = buffer_data_1[1815:1808] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_228[16] = buffer_data_1[1823:1816] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_228[17] = buffer_data_1[1831:1824] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_228[18] = buffer_data_1[1839:1832] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_228[19] = buffer_data_1[1847:1840] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_228[20] = buffer_data_0[1815:1808] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_228[21] = buffer_data_0[1823:1816] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_228[22] = buffer_data_0[1831:1824] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_228[23] = buffer_data_0[1839:1832] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_228[24] = buffer_data_0[1847:1840] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_228 = kernel_img_mul_228[0] + kernel_img_mul_228[1] + kernel_img_mul_228[2] + 
                kernel_img_mul_228[3] + kernel_img_mul_228[4] + kernel_img_mul_228[5] + 
                kernel_img_mul_228[6] + kernel_img_mul_228[7] + kernel_img_mul_228[8] + 
                kernel_img_mul_228[9] + kernel_img_mul_228[10] + kernel_img_mul_228[11] + 
                kernel_img_mul_228[12] + kernel_img_mul_228[13] + kernel_img_mul_228[14] + 
                kernel_img_mul_228[15] + kernel_img_mul_228[16] + kernel_img_mul_228[17] + 
                kernel_img_mul_228[18] + kernel_img_mul_228[19] + kernel_img_mul_228[20] + 
                kernel_img_mul_228[21] + kernel_img_mul_228[22] + kernel_img_mul_228[23] + 
                kernel_img_mul_228[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1831:1824] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1831:1824] <= kernel_img_sum_228[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1831:1824] <= 'd0;
end

wire  [39:0]  kernel_img_mul_229[0:24];
assign kernel_img_mul_229[0] = buffer_data_4[1823:1816] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_229[1] = buffer_data_4[1831:1824] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_229[2] = buffer_data_4[1839:1832] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_229[3] = buffer_data_4[1847:1840] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_229[4] = buffer_data_4[1855:1848] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_229[5] = buffer_data_3[1823:1816] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_229[6] = buffer_data_3[1831:1824] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_229[7] = buffer_data_3[1839:1832] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_229[8] = buffer_data_3[1847:1840] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_229[9] = buffer_data_3[1855:1848] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_229[10] = buffer_data_2[1823:1816] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_229[11] = buffer_data_2[1831:1824] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_229[12] = buffer_data_2[1839:1832] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_229[13] = buffer_data_2[1847:1840] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_229[14] = buffer_data_2[1855:1848] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_229[15] = buffer_data_1[1823:1816] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_229[16] = buffer_data_1[1831:1824] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_229[17] = buffer_data_1[1839:1832] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_229[18] = buffer_data_1[1847:1840] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_229[19] = buffer_data_1[1855:1848] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_229[20] = buffer_data_0[1823:1816] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_229[21] = buffer_data_0[1831:1824] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_229[22] = buffer_data_0[1839:1832] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_229[23] = buffer_data_0[1847:1840] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_229[24] = buffer_data_0[1855:1848] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_229 = kernel_img_mul_229[0] + kernel_img_mul_229[1] + kernel_img_mul_229[2] + 
                kernel_img_mul_229[3] + kernel_img_mul_229[4] + kernel_img_mul_229[5] + 
                kernel_img_mul_229[6] + kernel_img_mul_229[7] + kernel_img_mul_229[8] + 
                kernel_img_mul_229[9] + kernel_img_mul_229[10] + kernel_img_mul_229[11] + 
                kernel_img_mul_229[12] + kernel_img_mul_229[13] + kernel_img_mul_229[14] + 
                kernel_img_mul_229[15] + kernel_img_mul_229[16] + kernel_img_mul_229[17] + 
                kernel_img_mul_229[18] + kernel_img_mul_229[19] + kernel_img_mul_229[20] + 
                kernel_img_mul_229[21] + kernel_img_mul_229[22] + kernel_img_mul_229[23] + 
                kernel_img_mul_229[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1839:1832] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1839:1832] <= kernel_img_sum_229[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1839:1832] <= 'd0;
end

wire  [39:0]  kernel_img_mul_230[0:24];
assign kernel_img_mul_230[0] = buffer_data_4[1831:1824] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_230[1] = buffer_data_4[1839:1832] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_230[2] = buffer_data_4[1847:1840] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_230[3] = buffer_data_4[1855:1848] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_230[4] = buffer_data_4[1863:1856] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_230[5] = buffer_data_3[1831:1824] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_230[6] = buffer_data_3[1839:1832] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_230[7] = buffer_data_3[1847:1840] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_230[8] = buffer_data_3[1855:1848] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_230[9] = buffer_data_3[1863:1856] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_230[10] = buffer_data_2[1831:1824] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_230[11] = buffer_data_2[1839:1832] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_230[12] = buffer_data_2[1847:1840] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_230[13] = buffer_data_2[1855:1848] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_230[14] = buffer_data_2[1863:1856] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_230[15] = buffer_data_1[1831:1824] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_230[16] = buffer_data_1[1839:1832] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_230[17] = buffer_data_1[1847:1840] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_230[18] = buffer_data_1[1855:1848] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_230[19] = buffer_data_1[1863:1856] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_230[20] = buffer_data_0[1831:1824] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_230[21] = buffer_data_0[1839:1832] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_230[22] = buffer_data_0[1847:1840] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_230[23] = buffer_data_0[1855:1848] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_230[24] = buffer_data_0[1863:1856] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_230 = kernel_img_mul_230[0] + kernel_img_mul_230[1] + kernel_img_mul_230[2] + 
                kernel_img_mul_230[3] + kernel_img_mul_230[4] + kernel_img_mul_230[5] + 
                kernel_img_mul_230[6] + kernel_img_mul_230[7] + kernel_img_mul_230[8] + 
                kernel_img_mul_230[9] + kernel_img_mul_230[10] + kernel_img_mul_230[11] + 
                kernel_img_mul_230[12] + kernel_img_mul_230[13] + kernel_img_mul_230[14] + 
                kernel_img_mul_230[15] + kernel_img_mul_230[16] + kernel_img_mul_230[17] + 
                kernel_img_mul_230[18] + kernel_img_mul_230[19] + kernel_img_mul_230[20] + 
                kernel_img_mul_230[21] + kernel_img_mul_230[22] + kernel_img_mul_230[23] + 
                kernel_img_mul_230[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1847:1840] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1847:1840] <= kernel_img_sum_230[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1847:1840] <= 'd0;
end

wire  [39:0]  kernel_img_mul_231[0:24];
assign kernel_img_mul_231[0] = buffer_data_4[1839:1832] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_231[1] = buffer_data_4[1847:1840] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_231[2] = buffer_data_4[1855:1848] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_231[3] = buffer_data_4[1863:1856] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_231[4] = buffer_data_4[1871:1864] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_231[5] = buffer_data_3[1839:1832] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_231[6] = buffer_data_3[1847:1840] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_231[7] = buffer_data_3[1855:1848] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_231[8] = buffer_data_3[1863:1856] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_231[9] = buffer_data_3[1871:1864] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_231[10] = buffer_data_2[1839:1832] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_231[11] = buffer_data_2[1847:1840] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_231[12] = buffer_data_2[1855:1848] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_231[13] = buffer_data_2[1863:1856] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_231[14] = buffer_data_2[1871:1864] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_231[15] = buffer_data_1[1839:1832] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_231[16] = buffer_data_1[1847:1840] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_231[17] = buffer_data_1[1855:1848] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_231[18] = buffer_data_1[1863:1856] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_231[19] = buffer_data_1[1871:1864] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_231[20] = buffer_data_0[1839:1832] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_231[21] = buffer_data_0[1847:1840] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_231[22] = buffer_data_0[1855:1848] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_231[23] = buffer_data_0[1863:1856] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_231[24] = buffer_data_0[1871:1864] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_231 = kernel_img_mul_231[0] + kernel_img_mul_231[1] + kernel_img_mul_231[2] + 
                kernel_img_mul_231[3] + kernel_img_mul_231[4] + kernel_img_mul_231[5] + 
                kernel_img_mul_231[6] + kernel_img_mul_231[7] + kernel_img_mul_231[8] + 
                kernel_img_mul_231[9] + kernel_img_mul_231[10] + kernel_img_mul_231[11] + 
                kernel_img_mul_231[12] + kernel_img_mul_231[13] + kernel_img_mul_231[14] + 
                kernel_img_mul_231[15] + kernel_img_mul_231[16] + kernel_img_mul_231[17] + 
                kernel_img_mul_231[18] + kernel_img_mul_231[19] + kernel_img_mul_231[20] + 
                kernel_img_mul_231[21] + kernel_img_mul_231[22] + kernel_img_mul_231[23] + 
                kernel_img_mul_231[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1855:1848] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1855:1848] <= kernel_img_sum_231[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1855:1848] <= 'd0;
end

wire  [39:0]  kernel_img_mul_232[0:24];
assign kernel_img_mul_232[0] = buffer_data_4[1847:1840] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_232[1] = buffer_data_4[1855:1848] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_232[2] = buffer_data_4[1863:1856] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_232[3] = buffer_data_4[1871:1864] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_232[4] = buffer_data_4[1879:1872] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_232[5] = buffer_data_3[1847:1840] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_232[6] = buffer_data_3[1855:1848] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_232[7] = buffer_data_3[1863:1856] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_232[8] = buffer_data_3[1871:1864] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_232[9] = buffer_data_3[1879:1872] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_232[10] = buffer_data_2[1847:1840] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_232[11] = buffer_data_2[1855:1848] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_232[12] = buffer_data_2[1863:1856] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_232[13] = buffer_data_2[1871:1864] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_232[14] = buffer_data_2[1879:1872] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_232[15] = buffer_data_1[1847:1840] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_232[16] = buffer_data_1[1855:1848] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_232[17] = buffer_data_1[1863:1856] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_232[18] = buffer_data_1[1871:1864] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_232[19] = buffer_data_1[1879:1872] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_232[20] = buffer_data_0[1847:1840] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_232[21] = buffer_data_0[1855:1848] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_232[22] = buffer_data_0[1863:1856] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_232[23] = buffer_data_0[1871:1864] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_232[24] = buffer_data_0[1879:1872] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_232 = kernel_img_mul_232[0] + kernel_img_mul_232[1] + kernel_img_mul_232[2] + 
                kernel_img_mul_232[3] + kernel_img_mul_232[4] + kernel_img_mul_232[5] + 
                kernel_img_mul_232[6] + kernel_img_mul_232[7] + kernel_img_mul_232[8] + 
                kernel_img_mul_232[9] + kernel_img_mul_232[10] + kernel_img_mul_232[11] + 
                kernel_img_mul_232[12] + kernel_img_mul_232[13] + kernel_img_mul_232[14] + 
                kernel_img_mul_232[15] + kernel_img_mul_232[16] + kernel_img_mul_232[17] + 
                kernel_img_mul_232[18] + kernel_img_mul_232[19] + kernel_img_mul_232[20] + 
                kernel_img_mul_232[21] + kernel_img_mul_232[22] + kernel_img_mul_232[23] + 
                kernel_img_mul_232[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1863:1856] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1863:1856] <= kernel_img_sum_232[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1863:1856] <= 'd0;
end

wire  [39:0]  kernel_img_mul_233[0:24];
assign kernel_img_mul_233[0] = buffer_data_4[1855:1848] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_233[1] = buffer_data_4[1863:1856] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_233[2] = buffer_data_4[1871:1864] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_233[3] = buffer_data_4[1879:1872] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_233[4] = buffer_data_4[1887:1880] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_233[5] = buffer_data_3[1855:1848] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_233[6] = buffer_data_3[1863:1856] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_233[7] = buffer_data_3[1871:1864] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_233[8] = buffer_data_3[1879:1872] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_233[9] = buffer_data_3[1887:1880] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_233[10] = buffer_data_2[1855:1848] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_233[11] = buffer_data_2[1863:1856] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_233[12] = buffer_data_2[1871:1864] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_233[13] = buffer_data_2[1879:1872] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_233[14] = buffer_data_2[1887:1880] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_233[15] = buffer_data_1[1855:1848] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_233[16] = buffer_data_1[1863:1856] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_233[17] = buffer_data_1[1871:1864] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_233[18] = buffer_data_1[1879:1872] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_233[19] = buffer_data_1[1887:1880] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_233[20] = buffer_data_0[1855:1848] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_233[21] = buffer_data_0[1863:1856] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_233[22] = buffer_data_0[1871:1864] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_233[23] = buffer_data_0[1879:1872] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_233[24] = buffer_data_0[1887:1880] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_233 = kernel_img_mul_233[0] + kernel_img_mul_233[1] + kernel_img_mul_233[2] + 
                kernel_img_mul_233[3] + kernel_img_mul_233[4] + kernel_img_mul_233[5] + 
                kernel_img_mul_233[6] + kernel_img_mul_233[7] + kernel_img_mul_233[8] + 
                kernel_img_mul_233[9] + kernel_img_mul_233[10] + kernel_img_mul_233[11] + 
                kernel_img_mul_233[12] + kernel_img_mul_233[13] + kernel_img_mul_233[14] + 
                kernel_img_mul_233[15] + kernel_img_mul_233[16] + kernel_img_mul_233[17] + 
                kernel_img_mul_233[18] + kernel_img_mul_233[19] + kernel_img_mul_233[20] + 
                kernel_img_mul_233[21] + kernel_img_mul_233[22] + kernel_img_mul_233[23] + 
                kernel_img_mul_233[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1871:1864] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1871:1864] <= kernel_img_sum_233[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1871:1864] <= 'd0;
end

wire  [39:0]  kernel_img_mul_234[0:24];
assign kernel_img_mul_234[0] = buffer_data_4[1863:1856] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_234[1] = buffer_data_4[1871:1864] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_234[2] = buffer_data_4[1879:1872] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_234[3] = buffer_data_4[1887:1880] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_234[4] = buffer_data_4[1895:1888] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_234[5] = buffer_data_3[1863:1856] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_234[6] = buffer_data_3[1871:1864] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_234[7] = buffer_data_3[1879:1872] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_234[8] = buffer_data_3[1887:1880] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_234[9] = buffer_data_3[1895:1888] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_234[10] = buffer_data_2[1863:1856] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_234[11] = buffer_data_2[1871:1864] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_234[12] = buffer_data_2[1879:1872] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_234[13] = buffer_data_2[1887:1880] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_234[14] = buffer_data_2[1895:1888] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_234[15] = buffer_data_1[1863:1856] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_234[16] = buffer_data_1[1871:1864] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_234[17] = buffer_data_1[1879:1872] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_234[18] = buffer_data_1[1887:1880] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_234[19] = buffer_data_1[1895:1888] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_234[20] = buffer_data_0[1863:1856] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_234[21] = buffer_data_0[1871:1864] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_234[22] = buffer_data_0[1879:1872] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_234[23] = buffer_data_0[1887:1880] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_234[24] = buffer_data_0[1895:1888] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_234 = kernel_img_mul_234[0] + kernel_img_mul_234[1] + kernel_img_mul_234[2] + 
                kernel_img_mul_234[3] + kernel_img_mul_234[4] + kernel_img_mul_234[5] + 
                kernel_img_mul_234[6] + kernel_img_mul_234[7] + kernel_img_mul_234[8] + 
                kernel_img_mul_234[9] + kernel_img_mul_234[10] + kernel_img_mul_234[11] + 
                kernel_img_mul_234[12] + kernel_img_mul_234[13] + kernel_img_mul_234[14] + 
                kernel_img_mul_234[15] + kernel_img_mul_234[16] + kernel_img_mul_234[17] + 
                kernel_img_mul_234[18] + kernel_img_mul_234[19] + kernel_img_mul_234[20] + 
                kernel_img_mul_234[21] + kernel_img_mul_234[22] + kernel_img_mul_234[23] + 
                kernel_img_mul_234[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1879:1872] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1879:1872] <= kernel_img_sum_234[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1879:1872] <= 'd0;
end

wire  [39:0]  kernel_img_mul_235[0:24];
assign kernel_img_mul_235[0] = buffer_data_4[1871:1864] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_235[1] = buffer_data_4[1879:1872] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_235[2] = buffer_data_4[1887:1880] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_235[3] = buffer_data_4[1895:1888] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_235[4] = buffer_data_4[1903:1896] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_235[5] = buffer_data_3[1871:1864] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_235[6] = buffer_data_3[1879:1872] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_235[7] = buffer_data_3[1887:1880] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_235[8] = buffer_data_3[1895:1888] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_235[9] = buffer_data_3[1903:1896] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_235[10] = buffer_data_2[1871:1864] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_235[11] = buffer_data_2[1879:1872] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_235[12] = buffer_data_2[1887:1880] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_235[13] = buffer_data_2[1895:1888] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_235[14] = buffer_data_2[1903:1896] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_235[15] = buffer_data_1[1871:1864] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_235[16] = buffer_data_1[1879:1872] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_235[17] = buffer_data_1[1887:1880] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_235[18] = buffer_data_1[1895:1888] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_235[19] = buffer_data_1[1903:1896] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_235[20] = buffer_data_0[1871:1864] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_235[21] = buffer_data_0[1879:1872] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_235[22] = buffer_data_0[1887:1880] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_235[23] = buffer_data_0[1895:1888] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_235[24] = buffer_data_0[1903:1896] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_235 = kernel_img_mul_235[0] + kernel_img_mul_235[1] + kernel_img_mul_235[2] + 
                kernel_img_mul_235[3] + kernel_img_mul_235[4] + kernel_img_mul_235[5] + 
                kernel_img_mul_235[6] + kernel_img_mul_235[7] + kernel_img_mul_235[8] + 
                kernel_img_mul_235[9] + kernel_img_mul_235[10] + kernel_img_mul_235[11] + 
                kernel_img_mul_235[12] + kernel_img_mul_235[13] + kernel_img_mul_235[14] + 
                kernel_img_mul_235[15] + kernel_img_mul_235[16] + kernel_img_mul_235[17] + 
                kernel_img_mul_235[18] + kernel_img_mul_235[19] + kernel_img_mul_235[20] + 
                kernel_img_mul_235[21] + kernel_img_mul_235[22] + kernel_img_mul_235[23] + 
                kernel_img_mul_235[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1887:1880] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1887:1880] <= kernel_img_sum_235[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1887:1880] <= 'd0;
end

wire  [39:0]  kernel_img_mul_236[0:24];
assign kernel_img_mul_236[0] = buffer_data_4[1879:1872] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_236[1] = buffer_data_4[1887:1880] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_236[2] = buffer_data_4[1895:1888] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_236[3] = buffer_data_4[1903:1896] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_236[4] = buffer_data_4[1911:1904] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_236[5] = buffer_data_3[1879:1872] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_236[6] = buffer_data_3[1887:1880] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_236[7] = buffer_data_3[1895:1888] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_236[8] = buffer_data_3[1903:1896] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_236[9] = buffer_data_3[1911:1904] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_236[10] = buffer_data_2[1879:1872] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_236[11] = buffer_data_2[1887:1880] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_236[12] = buffer_data_2[1895:1888] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_236[13] = buffer_data_2[1903:1896] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_236[14] = buffer_data_2[1911:1904] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_236[15] = buffer_data_1[1879:1872] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_236[16] = buffer_data_1[1887:1880] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_236[17] = buffer_data_1[1895:1888] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_236[18] = buffer_data_1[1903:1896] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_236[19] = buffer_data_1[1911:1904] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_236[20] = buffer_data_0[1879:1872] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_236[21] = buffer_data_0[1887:1880] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_236[22] = buffer_data_0[1895:1888] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_236[23] = buffer_data_0[1903:1896] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_236[24] = buffer_data_0[1911:1904] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_236 = kernel_img_mul_236[0] + kernel_img_mul_236[1] + kernel_img_mul_236[2] + 
                kernel_img_mul_236[3] + kernel_img_mul_236[4] + kernel_img_mul_236[5] + 
                kernel_img_mul_236[6] + kernel_img_mul_236[7] + kernel_img_mul_236[8] + 
                kernel_img_mul_236[9] + kernel_img_mul_236[10] + kernel_img_mul_236[11] + 
                kernel_img_mul_236[12] + kernel_img_mul_236[13] + kernel_img_mul_236[14] + 
                kernel_img_mul_236[15] + kernel_img_mul_236[16] + kernel_img_mul_236[17] + 
                kernel_img_mul_236[18] + kernel_img_mul_236[19] + kernel_img_mul_236[20] + 
                kernel_img_mul_236[21] + kernel_img_mul_236[22] + kernel_img_mul_236[23] + 
                kernel_img_mul_236[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1895:1888] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1895:1888] <= kernel_img_sum_236[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1895:1888] <= 'd0;
end

wire  [39:0]  kernel_img_mul_237[0:24];
assign kernel_img_mul_237[0] = buffer_data_4[1887:1880] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_237[1] = buffer_data_4[1895:1888] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_237[2] = buffer_data_4[1903:1896] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_237[3] = buffer_data_4[1911:1904] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_237[4] = buffer_data_4[1919:1912] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_237[5] = buffer_data_3[1887:1880] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_237[6] = buffer_data_3[1895:1888] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_237[7] = buffer_data_3[1903:1896] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_237[8] = buffer_data_3[1911:1904] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_237[9] = buffer_data_3[1919:1912] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_237[10] = buffer_data_2[1887:1880] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_237[11] = buffer_data_2[1895:1888] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_237[12] = buffer_data_2[1903:1896] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_237[13] = buffer_data_2[1911:1904] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_237[14] = buffer_data_2[1919:1912] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_237[15] = buffer_data_1[1887:1880] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_237[16] = buffer_data_1[1895:1888] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_237[17] = buffer_data_1[1903:1896] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_237[18] = buffer_data_1[1911:1904] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_237[19] = buffer_data_1[1919:1912] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_237[20] = buffer_data_0[1887:1880] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_237[21] = buffer_data_0[1895:1888] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_237[22] = buffer_data_0[1903:1896] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_237[23] = buffer_data_0[1911:1904] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_237[24] = buffer_data_0[1919:1912] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_237 = kernel_img_mul_237[0] + kernel_img_mul_237[1] + kernel_img_mul_237[2] + 
                kernel_img_mul_237[3] + kernel_img_mul_237[4] + kernel_img_mul_237[5] + 
                kernel_img_mul_237[6] + kernel_img_mul_237[7] + kernel_img_mul_237[8] + 
                kernel_img_mul_237[9] + kernel_img_mul_237[10] + kernel_img_mul_237[11] + 
                kernel_img_mul_237[12] + kernel_img_mul_237[13] + kernel_img_mul_237[14] + 
                kernel_img_mul_237[15] + kernel_img_mul_237[16] + kernel_img_mul_237[17] + 
                kernel_img_mul_237[18] + kernel_img_mul_237[19] + kernel_img_mul_237[20] + 
                kernel_img_mul_237[21] + kernel_img_mul_237[22] + kernel_img_mul_237[23] + 
                kernel_img_mul_237[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1903:1896] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1903:1896] <= kernel_img_sum_237[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1903:1896] <= 'd0;
end

wire  [39:0]  kernel_img_mul_238[0:24];
assign kernel_img_mul_238[0] = buffer_data_4[1895:1888] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_238[1] = buffer_data_4[1903:1896] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_238[2] = buffer_data_4[1911:1904] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_238[3] = buffer_data_4[1919:1912] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_238[4] = buffer_data_4[1927:1920] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_238[5] = buffer_data_3[1895:1888] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_238[6] = buffer_data_3[1903:1896] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_238[7] = buffer_data_3[1911:1904] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_238[8] = buffer_data_3[1919:1912] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_238[9] = buffer_data_3[1927:1920] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_238[10] = buffer_data_2[1895:1888] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_238[11] = buffer_data_2[1903:1896] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_238[12] = buffer_data_2[1911:1904] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_238[13] = buffer_data_2[1919:1912] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_238[14] = buffer_data_2[1927:1920] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_238[15] = buffer_data_1[1895:1888] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_238[16] = buffer_data_1[1903:1896] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_238[17] = buffer_data_1[1911:1904] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_238[18] = buffer_data_1[1919:1912] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_238[19] = buffer_data_1[1927:1920] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_238[20] = buffer_data_0[1895:1888] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_238[21] = buffer_data_0[1903:1896] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_238[22] = buffer_data_0[1911:1904] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_238[23] = buffer_data_0[1919:1912] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_238[24] = buffer_data_0[1927:1920] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_238 = kernel_img_mul_238[0] + kernel_img_mul_238[1] + kernel_img_mul_238[2] + 
                kernel_img_mul_238[3] + kernel_img_mul_238[4] + kernel_img_mul_238[5] + 
                kernel_img_mul_238[6] + kernel_img_mul_238[7] + kernel_img_mul_238[8] + 
                kernel_img_mul_238[9] + kernel_img_mul_238[10] + kernel_img_mul_238[11] + 
                kernel_img_mul_238[12] + kernel_img_mul_238[13] + kernel_img_mul_238[14] + 
                kernel_img_mul_238[15] + kernel_img_mul_238[16] + kernel_img_mul_238[17] + 
                kernel_img_mul_238[18] + kernel_img_mul_238[19] + kernel_img_mul_238[20] + 
                kernel_img_mul_238[21] + kernel_img_mul_238[22] + kernel_img_mul_238[23] + 
                kernel_img_mul_238[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1911:1904] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1911:1904] <= kernel_img_sum_238[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1911:1904] <= 'd0;
end

wire  [39:0]  kernel_img_mul_239[0:24];
assign kernel_img_mul_239[0] = buffer_data_4[1903:1896] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_239[1] = buffer_data_4[1911:1904] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_239[2] = buffer_data_4[1919:1912] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_239[3] = buffer_data_4[1927:1920] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_239[4] = buffer_data_4[1935:1928] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_239[5] = buffer_data_3[1903:1896] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_239[6] = buffer_data_3[1911:1904] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_239[7] = buffer_data_3[1919:1912] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_239[8] = buffer_data_3[1927:1920] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_239[9] = buffer_data_3[1935:1928] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_239[10] = buffer_data_2[1903:1896] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_239[11] = buffer_data_2[1911:1904] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_239[12] = buffer_data_2[1919:1912] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_239[13] = buffer_data_2[1927:1920] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_239[14] = buffer_data_2[1935:1928] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_239[15] = buffer_data_1[1903:1896] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_239[16] = buffer_data_1[1911:1904] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_239[17] = buffer_data_1[1919:1912] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_239[18] = buffer_data_1[1927:1920] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_239[19] = buffer_data_1[1935:1928] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_239[20] = buffer_data_0[1903:1896] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_239[21] = buffer_data_0[1911:1904] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_239[22] = buffer_data_0[1919:1912] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_239[23] = buffer_data_0[1927:1920] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_239[24] = buffer_data_0[1935:1928] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_239 = kernel_img_mul_239[0] + kernel_img_mul_239[1] + kernel_img_mul_239[2] + 
                kernel_img_mul_239[3] + kernel_img_mul_239[4] + kernel_img_mul_239[5] + 
                kernel_img_mul_239[6] + kernel_img_mul_239[7] + kernel_img_mul_239[8] + 
                kernel_img_mul_239[9] + kernel_img_mul_239[10] + kernel_img_mul_239[11] + 
                kernel_img_mul_239[12] + kernel_img_mul_239[13] + kernel_img_mul_239[14] + 
                kernel_img_mul_239[15] + kernel_img_mul_239[16] + kernel_img_mul_239[17] + 
                kernel_img_mul_239[18] + kernel_img_mul_239[19] + kernel_img_mul_239[20] + 
                kernel_img_mul_239[21] + kernel_img_mul_239[22] + kernel_img_mul_239[23] + 
                kernel_img_mul_239[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1919:1912] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1919:1912] <= kernel_img_sum_239[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1919:1912] <= 'd0;
end

wire  [39:0]  kernel_img_mul_240[0:24];
assign kernel_img_mul_240[0] = buffer_data_4[1911:1904] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_240[1] = buffer_data_4[1919:1912] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_240[2] = buffer_data_4[1927:1920] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_240[3] = buffer_data_4[1935:1928] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_240[4] = buffer_data_4[1943:1936] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_240[5] = buffer_data_3[1911:1904] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_240[6] = buffer_data_3[1919:1912] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_240[7] = buffer_data_3[1927:1920] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_240[8] = buffer_data_3[1935:1928] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_240[9] = buffer_data_3[1943:1936] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_240[10] = buffer_data_2[1911:1904] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_240[11] = buffer_data_2[1919:1912] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_240[12] = buffer_data_2[1927:1920] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_240[13] = buffer_data_2[1935:1928] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_240[14] = buffer_data_2[1943:1936] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_240[15] = buffer_data_1[1911:1904] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_240[16] = buffer_data_1[1919:1912] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_240[17] = buffer_data_1[1927:1920] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_240[18] = buffer_data_1[1935:1928] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_240[19] = buffer_data_1[1943:1936] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_240[20] = buffer_data_0[1911:1904] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_240[21] = buffer_data_0[1919:1912] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_240[22] = buffer_data_0[1927:1920] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_240[23] = buffer_data_0[1935:1928] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_240[24] = buffer_data_0[1943:1936] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_240 = kernel_img_mul_240[0] + kernel_img_mul_240[1] + kernel_img_mul_240[2] + 
                kernel_img_mul_240[3] + kernel_img_mul_240[4] + kernel_img_mul_240[5] + 
                kernel_img_mul_240[6] + kernel_img_mul_240[7] + kernel_img_mul_240[8] + 
                kernel_img_mul_240[9] + kernel_img_mul_240[10] + kernel_img_mul_240[11] + 
                kernel_img_mul_240[12] + kernel_img_mul_240[13] + kernel_img_mul_240[14] + 
                kernel_img_mul_240[15] + kernel_img_mul_240[16] + kernel_img_mul_240[17] + 
                kernel_img_mul_240[18] + kernel_img_mul_240[19] + kernel_img_mul_240[20] + 
                kernel_img_mul_240[21] + kernel_img_mul_240[22] + kernel_img_mul_240[23] + 
                kernel_img_mul_240[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1927:1920] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1927:1920] <= kernel_img_sum_240[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1927:1920] <= 'd0;
end

wire  [39:0]  kernel_img_mul_241[0:24];
assign kernel_img_mul_241[0] = buffer_data_4[1919:1912] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_241[1] = buffer_data_4[1927:1920] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_241[2] = buffer_data_4[1935:1928] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_241[3] = buffer_data_4[1943:1936] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_241[4] = buffer_data_4[1951:1944] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_241[5] = buffer_data_3[1919:1912] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_241[6] = buffer_data_3[1927:1920] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_241[7] = buffer_data_3[1935:1928] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_241[8] = buffer_data_3[1943:1936] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_241[9] = buffer_data_3[1951:1944] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_241[10] = buffer_data_2[1919:1912] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_241[11] = buffer_data_2[1927:1920] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_241[12] = buffer_data_2[1935:1928] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_241[13] = buffer_data_2[1943:1936] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_241[14] = buffer_data_2[1951:1944] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_241[15] = buffer_data_1[1919:1912] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_241[16] = buffer_data_1[1927:1920] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_241[17] = buffer_data_1[1935:1928] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_241[18] = buffer_data_1[1943:1936] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_241[19] = buffer_data_1[1951:1944] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_241[20] = buffer_data_0[1919:1912] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_241[21] = buffer_data_0[1927:1920] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_241[22] = buffer_data_0[1935:1928] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_241[23] = buffer_data_0[1943:1936] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_241[24] = buffer_data_0[1951:1944] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_241 = kernel_img_mul_241[0] + kernel_img_mul_241[1] + kernel_img_mul_241[2] + 
                kernel_img_mul_241[3] + kernel_img_mul_241[4] + kernel_img_mul_241[5] + 
                kernel_img_mul_241[6] + kernel_img_mul_241[7] + kernel_img_mul_241[8] + 
                kernel_img_mul_241[9] + kernel_img_mul_241[10] + kernel_img_mul_241[11] + 
                kernel_img_mul_241[12] + kernel_img_mul_241[13] + kernel_img_mul_241[14] + 
                kernel_img_mul_241[15] + kernel_img_mul_241[16] + kernel_img_mul_241[17] + 
                kernel_img_mul_241[18] + kernel_img_mul_241[19] + kernel_img_mul_241[20] + 
                kernel_img_mul_241[21] + kernel_img_mul_241[22] + kernel_img_mul_241[23] + 
                kernel_img_mul_241[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1935:1928] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1935:1928] <= kernel_img_sum_241[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1935:1928] <= 'd0;
end

wire  [39:0]  kernel_img_mul_242[0:24];
assign kernel_img_mul_242[0] = buffer_data_4[1927:1920] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_242[1] = buffer_data_4[1935:1928] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_242[2] = buffer_data_4[1943:1936] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_242[3] = buffer_data_4[1951:1944] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_242[4] = buffer_data_4[1959:1952] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_242[5] = buffer_data_3[1927:1920] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_242[6] = buffer_data_3[1935:1928] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_242[7] = buffer_data_3[1943:1936] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_242[8] = buffer_data_3[1951:1944] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_242[9] = buffer_data_3[1959:1952] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_242[10] = buffer_data_2[1927:1920] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_242[11] = buffer_data_2[1935:1928] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_242[12] = buffer_data_2[1943:1936] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_242[13] = buffer_data_2[1951:1944] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_242[14] = buffer_data_2[1959:1952] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_242[15] = buffer_data_1[1927:1920] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_242[16] = buffer_data_1[1935:1928] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_242[17] = buffer_data_1[1943:1936] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_242[18] = buffer_data_1[1951:1944] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_242[19] = buffer_data_1[1959:1952] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_242[20] = buffer_data_0[1927:1920] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_242[21] = buffer_data_0[1935:1928] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_242[22] = buffer_data_0[1943:1936] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_242[23] = buffer_data_0[1951:1944] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_242[24] = buffer_data_0[1959:1952] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_242 = kernel_img_mul_242[0] + kernel_img_mul_242[1] + kernel_img_mul_242[2] + 
                kernel_img_mul_242[3] + kernel_img_mul_242[4] + kernel_img_mul_242[5] + 
                kernel_img_mul_242[6] + kernel_img_mul_242[7] + kernel_img_mul_242[8] + 
                kernel_img_mul_242[9] + kernel_img_mul_242[10] + kernel_img_mul_242[11] + 
                kernel_img_mul_242[12] + kernel_img_mul_242[13] + kernel_img_mul_242[14] + 
                kernel_img_mul_242[15] + kernel_img_mul_242[16] + kernel_img_mul_242[17] + 
                kernel_img_mul_242[18] + kernel_img_mul_242[19] + kernel_img_mul_242[20] + 
                kernel_img_mul_242[21] + kernel_img_mul_242[22] + kernel_img_mul_242[23] + 
                kernel_img_mul_242[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1943:1936] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1943:1936] <= kernel_img_sum_242[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1943:1936] <= 'd0;
end

wire  [39:0]  kernel_img_mul_243[0:24];
assign kernel_img_mul_243[0] = buffer_data_4[1935:1928] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_243[1] = buffer_data_4[1943:1936] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_243[2] = buffer_data_4[1951:1944] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_243[3] = buffer_data_4[1959:1952] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_243[4] = buffer_data_4[1967:1960] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_243[5] = buffer_data_3[1935:1928] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_243[6] = buffer_data_3[1943:1936] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_243[7] = buffer_data_3[1951:1944] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_243[8] = buffer_data_3[1959:1952] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_243[9] = buffer_data_3[1967:1960] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_243[10] = buffer_data_2[1935:1928] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_243[11] = buffer_data_2[1943:1936] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_243[12] = buffer_data_2[1951:1944] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_243[13] = buffer_data_2[1959:1952] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_243[14] = buffer_data_2[1967:1960] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_243[15] = buffer_data_1[1935:1928] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_243[16] = buffer_data_1[1943:1936] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_243[17] = buffer_data_1[1951:1944] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_243[18] = buffer_data_1[1959:1952] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_243[19] = buffer_data_1[1967:1960] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_243[20] = buffer_data_0[1935:1928] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_243[21] = buffer_data_0[1943:1936] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_243[22] = buffer_data_0[1951:1944] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_243[23] = buffer_data_0[1959:1952] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_243[24] = buffer_data_0[1967:1960] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_243 = kernel_img_mul_243[0] + kernel_img_mul_243[1] + kernel_img_mul_243[2] + 
                kernel_img_mul_243[3] + kernel_img_mul_243[4] + kernel_img_mul_243[5] + 
                kernel_img_mul_243[6] + kernel_img_mul_243[7] + kernel_img_mul_243[8] + 
                kernel_img_mul_243[9] + kernel_img_mul_243[10] + kernel_img_mul_243[11] + 
                kernel_img_mul_243[12] + kernel_img_mul_243[13] + kernel_img_mul_243[14] + 
                kernel_img_mul_243[15] + kernel_img_mul_243[16] + kernel_img_mul_243[17] + 
                kernel_img_mul_243[18] + kernel_img_mul_243[19] + kernel_img_mul_243[20] + 
                kernel_img_mul_243[21] + kernel_img_mul_243[22] + kernel_img_mul_243[23] + 
                kernel_img_mul_243[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1951:1944] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1951:1944] <= kernel_img_sum_243[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1951:1944] <= 'd0;
end

wire  [39:0]  kernel_img_mul_244[0:24];
assign kernel_img_mul_244[0] = buffer_data_4[1943:1936] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_244[1] = buffer_data_4[1951:1944] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_244[2] = buffer_data_4[1959:1952] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_244[3] = buffer_data_4[1967:1960] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_244[4] = buffer_data_4[1975:1968] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_244[5] = buffer_data_3[1943:1936] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_244[6] = buffer_data_3[1951:1944] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_244[7] = buffer_data_3[1959:1952] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_244[8] = buffer_data_3[1967:1960] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_244[9] = buffer_data_3[1975:1968] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_244[10] = buffer_data_2[1943:1936] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_244[11] = buffer_data_2[1951:1944] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_244[12] = buffer_data_2[1959:1952] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_244[13] = buffer_data_2[1967:1960] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_244[14] = buffer_data_2[1975:1968] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_244[15] = buffer_data_1[1943:1936] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_244[16] = buffer_data_1[1951:1944] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_244[17] = buffer_data_1[1959:1952] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_244[18] = buffer_data_1[1967:1960] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_244[19] = buffer_data_1[1975:1968] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_244[20] = buffer_data_0[1943:1936] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_244[21] = buffer_data_0[1951:1944] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_244[22] = buffer_data_0[1959:1952] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_244[23] = buffer_data_0[1967:1960] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_244[24] = buffer_data_0[1975:1968] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_244 = kernel_img_mul_244[0] + kernel_img_mul_244[1] + kernel_img_mul_244[2] + 
                kernel_img_mul_244[3] + kernel_img_mul_244[4] + kernel_img_mul_244[5] + 
                kernel_img_mul_244[6] + kernel_img_mul_244[7] + kernel_img_mul_244[8] + 
                kernel_img_mul_244[9] + kernel_img_mul_244[10] + kernel_img_mul_244[11] + 
                kernel_img_mul_244[12] + kernel_img_mul_244[13] + kernel_img_mul_244[14] + 
                kernel_img_mul_244[15] + kernel_img_mul_244[16] + kernel_img_mul_244[17] + 
                kernel_img_mul_244[18] + kernel_img_mul_244[19] + kernel_img_mul_244[20] + 
                kernel_img_mul_244[21] + kernel_img_mul_244[22] + kernel_img_mul_244[23] + 
                kernel_img_mul_244[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1959:1952] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1959:1952] <= kernel_img_sum_244[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1959:1952] <= 'd0;
end

wire  [39:0]  kernel_img_mul_245[0:24];
assign kernel_img_mul_245[0] = buffer_data_4[1951:1944] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_245[1] = buffer_data_4[1959:1952] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_245[2] = buffer_data_4[1967:1960] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_245[3] = buffer_data_4[1975:1968] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_245[4] = buffer_data_4[1983:1976] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_245[5] = buffer_data_3[1951:1944] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_245[6] = buffer_data_3[1959:1952] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_245[7] = buffer_data_3[1967:1960] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_245[8] = buffer_data_3[1975:1968] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_245[9] = buffer_data_3[1983:1976] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_245[10] = buffer_data_2[1951:1944] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_245[11] = buffer_data_2[1959:1952] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_245[12] = buffer_data_2[1967:1960] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_245[13] = buffer_data_2[1975:1968] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_245[14] = buffer_data_2[1983:1976] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_245[15] = buffer_data_1[1951:1944] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_245[16] = buffer_data_1[1959:1952] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_245[17] = buffer_data_1[1967:1960] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_245[18] = buffer_data_1[1975:1968] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_245[19] = buffer_data_1[1983:1976] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_245[20] = buffer_data_0[1951:1944] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_245[21] = buffer_data_0[1959:1952] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_245[22] = buffer_data_0[1967:1960] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_245[23] = buffer_data_0[1975:1968] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_245[24] = buffer_data_0[1983:1976] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_245 = kernel_img_mul_245[0] + kernel_img_mul_245[1] + kernel_img_mul_245[2] + 
                kernel_img_mul_245[3] + kernel_img_mul_245[4] + kernel_img_mul_245[5] + 
                kernel_img_mul_245[6] + kernel_img_mul_245[7] + kernel_img_mul_245[8] + 
                kernel_img_mul_245[9] + kernel_img_mul_245[10] + kernel_img_mul_245[11] + 
                kernel_img_mul_245[12] + kernel_img_mul_245[13] + kernel_img_mul_245[14] + 
                kernel_img_mul_245[15] + kernel_img_mul_245[16] + kernel_img_mul_245[17] + 
                kernel_img_mul_245[18] + kernel_img_mul_245[19] + kernel_img_mul_245[20] + 
                kernel_img_mul_245[21] + kernel_img_mul_245[22] + kernel_img_mul_245[23] + 
                kernel_img_mul_245[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1967:1960] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1967:1960] <= kernel_img_sum_245[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1967:1960] <= 'd0;
end

wire  [39:0]  kernel_img_mul_246[0:24];
assign kernel_img_mul_246[0] = buffer_data_4[1959:1952] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_246[1] = buffer_data_4[1967:1960] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_246[2] = buffer_data_4[1975:1968] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_246[3] = buffer_data_4[1983:1976] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_246[4] = buffer_data_4[1991:1984] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_246[5] = buffer_data_3[1959:1952] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_246[6] = buffer_data_3[1967:1960] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_246[7] = buffer_data_3[1975:1968] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_246[8] = buffer_data_3[1983:1976] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_246[9] = buffer_data_3[1991:1984] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_246[10] = buffer_data_2[1959:1952] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_246[11] = buffer_data_2[1967:1960] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_246[12] = buffer_data_2[1975:1968] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_246[13] = buffer_data_2[1983:1976] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_246[14] = buffer_data_2[1991:1984] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_246[15] = buffer_data_1[1959:1952] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_246[16] = buffer_data_1[1967:1960] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_246[17] = buffer_data_1[1975:1968] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_246[18] = buffer_data_1[1983:1976] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_246[19] = buffer_data_1[1991:1984] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_246[20] = buffer_data_0[1959:1952] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_246[21] = buffer_data_0[1967:1960] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_246[22] = buffer_data_0[1975:1968] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_246[23] = buffer_data_0[1983:1976] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_246[24] = buffer_data_0[1991:1984] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_246 = kernel_img_mul_246[0] + kernel_img_mul_246[1] + kernel_img_mul_246[2] + 
                kernel_img_mul_246[3] + kernel_img_mul_246[4] + kernel_img_mul_246[5] + 
                kernel_img_mul_246[6] + kernel_img_mul_246[7] + kernel_img_mul_246[8] + 
                kernel_img_mul_246[9] + kernel_img_mul_246[10] + kernel_img_mul_246[11] + 
                kernel_img_mul_246[12] + kernel_img_mul_246[13] + kernel_img_mul_246[14] + 
                kernel_img_mul_246[15] + kernel_img_mul_246[16] + kernel_img_mul_246[17] + 
                kernel_img_mul_246[18] + kernel_img_mul_246[19] + kernel_img_mul_246[20] + 
                kernel_img_mul_246[21] + kernel_img_mul_246[22] + kernel_img_mul_246[23] + 
                kernel_img_mul_246[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1975:1968] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1975:1968] <= kernel_img_sum_246[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1975:1968] <= 'd0;
end

wire  [39:0]  kernel_img_mul_247[0:24];
assign kernel_img_mul_247[0] = buffer_data_4[1967:1960] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_247[1] = buffer_data_4[1975:1968] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_247[2] = buffer_data_4[1983:1976] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_247[3] = buffer_data_4[1991:1984] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_247[4] = buffer_data_4[1999:1992] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_247[5] = buffer_data_3[1967:1960] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_247[6] = buffer_data_3[1975:1968] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_247[7] = buffer_data_3[1983:1976] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_247[8] = buffer_data_3[1991:1984] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_247[9] = buffer_data_3[1999:1992] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_247[10] = buffer_data_2[1967:1960] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_247[11] = buffer_data_2[1975:1968] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_247[12] = buffer_data_2[1983:1976] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_247[13] = buffer_data_2[1991:1984] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_247[14] = buffer_data_2[1999:1992] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_247[15] = buffer_data_1[1967:1960] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_247[16] = buffer_data_1[1975:1968] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_247[17] = buffer_data_1[1983:1976] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_247[18] = buffer_data_1[1991:1984] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_247[19] = buffer_data_1[1999:1992] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_247[20] = buffer_data_0[1967:1960] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_247[21] = buffer_data_0[1975:1968] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_247[22] = buffer_data_0[1983:1976] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_247[23] = buffer_data_0[1991:1984] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_247[24] = buffer_data_0[1999:1992] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_247 = kernel_img_mul_247[0] + kernel_img_mul_247[1] + kernel_img_mul_247[2] + 
                kernel_img_mul_247[3] + kernel_img_mul_247[4] + kernel_img_mul_247[5] + 
                kernel_img_mul_247[6] + kernel_img_mul_247[7] + kernel_img_mul_247[8] + 
                kernel_img_mul_247[9] + kernel_img_mul_247[10] + kernel_img_mul_247[11] + 
                kernel_img_mul_247[12] + kernel_img_mul_247[13] + kernel_img_mul_247[14] + 
                kernel_img_mul_247[15] + kernel_img_mul_247[16] + kernel_img_mul_247[17] + 
                kernel_img_mul_247[18] + kernel_img_mul_247[19] + kernel_img_mul_247[20] + 
                kernel_img_mul_247[21] + kernel_img_mul_247[22] + kernel_img_mul_247[23] + 
                kernel_img_mul_247[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1983:1976] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1983:1976] <= kernel_img_sum_247[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1983:1976] <= 'd0;
end

wire  [39:0]  kernel_img_mul_248[0:24];
assign kernel_img_mul_248[0] = buffer_data_4[1975:1968] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_248[1] = buffer_data_4[1983:1976] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_248[2] = buffer_data_4[1991:1984] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_248[3] = buffer_data_4[1999:1992] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_248[4] = buffer_data_4[2007:2000] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_248[5] = buffer_data_3[1975:1968] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_248[6] = buffer_data_3[1983:1976] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_248[7] = buffer_data_3[1991:1984] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_248[8] = buffer_data_3[1999:1992] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_248[9] = buffer_data_3[2007:2000] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_248[10] = buffer_data_2[1975:1968] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_248[11] = buffer_data_2[1983:1976] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_248[12] = buffer_data_2[1991:1984] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_248[13] = buffer_data_2[1999:1992] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_248[14] = buffer_data_2[2007:2000] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_248[15] = buffer_data_1[1975:1968] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_248[16] = buffer_data_1[1983:1976] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_248[17] = buffer_data_1[1991:1984] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_248[18] = buffer_data_1[1999:1992] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_248[19] = buffer_data_1[2007:2000] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_248[20] = buffer_data_0[1975:1968] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_248[21] = buffer_data_0[1983:1976] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_248[22] = buffer_data_0[1991:1984] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_248[23] = buffer_data_0[1999:1992] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_248[24] = buffer_data_0[2007:2000] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_248 = kernel_img_mul_248[0] + kernel_img_mul_248[1] + kernel_img_mul_248[2] + 
                kernel_img_mul_248[3] + kernel_img_mul_248[4] + kernel_img_mul_248[5] + 
                kernel_img_mul_248[6] + kernel_img_mul_248[7] + kernel_img_mul_248[8] + 
                kernel_img_mul_248[9] + kernel_img_mul_248[10] + kernel_img_mul_248[11] + 
                kernel_img_mul_248[12] + kernel_img_mul_248[13] + kernel_img_mul_248[14] + 
                kernel_img_mul_248[15] + kernel_img_mul_248[16] + kernel_img_mul_248[17] + 
                kernel_img_mul_248[18] + kernel_img_mul_248[19] + kernel_img_mul_248[20] + 
                kernel_img_mul_248[21] + kernel_img_mul_248[22] + kernel_img_mul_248[23] + 
                kernel_img_mul_248[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1991:1984] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1991:1984] <= kernel_img_sum_248[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1991:1984] <= 'd0;
end

wire  [39:0]  kernel_img_mul_249[0:24];
assign kernel_img_mul_249[0] = buffer_data_4[1983:1976] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_249[1] = buffer_data_4[1991:1984] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_249[2] = buffer_data_4[1999:1992] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_249[3] = buffer_data_4[2007:2000] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_249[4] = buffer_data_4[2015:2008] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_249[5] = buffer_data_3[1983:1976] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_249[6] = buffer_data_3[1991:1984] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_249[7] = buffer_data_3[1999:1992] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_249[8] = buffer_data_3[2007:2000] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_249[9] = buffer_data_3[2015:2008] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_249[10] = buffer_data_2[1983:1976] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_249[11] = buffer_data_2[1991:1984] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_249[12] = buffer_data_2[1999:1992] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_249[13] = buffer_data_2[2007:2000] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_249[14] = buffer_data_2[2015:2008] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_249[15] = buffer_data_1[1983:1976] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_249[16] = buffer_data_1[1991:1984] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_249[17] = buffer_data_1[1999:1992] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_249[18] = buffer_data_1[2007:2000] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_249[19] = buffer_data_1[2015:2008] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_249[20] = buffer_data_0[1983:1976] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_249[21] = buffer_data_0[1991:1984] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_249[22] = buffer_data_0[1999:1992] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_249[23] = buffer_data_0[2007:2000] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_249[24] = buffer_data_0[2015:2008] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_249 = kernel_img_mul_249[0] + kernel_img_mul_249[1] + kernel_img_mul_249[2] + 
                kernel_img_mul_249[3] + kernel_img_mul_249[4] + kernel_img_mul_249[5] + 
                kernel_img_mul_249[6] + kernel_img_mul_249[7] + kernel_img_mul_249[8] + 
                kernel_img_mul_249[9] + kernel_img_mul_249[10] + kernel_img_mul_249[11] + 
                kernel_img_mul_249[12] + kernel_img_mul_249[13] + kernel_img_mul_249[14] + 
                kernel_img_mul_249[15] + kernel_img_mul_249[16] + kernel_img_mul_249[17] + 
                kernel_img_mul_249[18] + kernel_img_mul_249[19] + kernel_img_mul_249[20] + 
                kernel_img_mul_249[21] + kernel_img_mul_249[22] + kernel_img_mul_249[23] + 
                kernel_img_mul_249[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[1999:1992] <= 'd0;
  else if (current_state==ST_START)
    blur_din[1999:1992] <= kernel_img_sum_249[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1999:1992] <= 'd0;
end

wire  [39:0]  kernel_img_mul_250[0:24];
assign kernel_img_mul_250[0] = buffer_data_4[1991:1984] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_250[1] = buffer_data_4[1999:1992] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_250[2] = buffer_data_4[2007:2000] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_250[3] = buffer_data_4[2015:2008] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_250[4] = buffer_data_4[2023:2016] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_250[5] = buffer_data_3[1991:1984] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_250[6] = buffer_data_3[1999:1992] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_250[7] = buffer_data_3[2007:2000] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_250[8] = buffer_data_3[2015:2008] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_250[9] = buffer_data_3[2023:2016] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_250[10] = buffer_data_2[1991:1984] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_250[11] = buffer_data_2[1999:1992] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_250[12] = buffer_data_2[2007:2000] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_250[13] = buffer_data_2[2015:2008] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_250[14] = buffer_data_2[2023:2016] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_250[15] = buffer_data_1[1991:1984] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_250[16] = buffer_data_1[1999:1992] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_250[17] = buffer_data_1[2007:2000] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_250[18] = buffer_data_1[2015:2008] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_250[19] = buffer_data_1[2023:2016] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_250[20] = buffer_data_0[1991:1984] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_250[21] = buffer_data_0[1999:1992] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_250[22] = buffer_data_0[2007:2000] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_250[23] = buffer_data_0[2015:2008] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_250[24] = buffer_data_0[2023:2016] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_250 = kernel_img_mul_250[0] + kernel_img_mul_250[1] + kernel_img_mul_250[2] + 
                kernel_img_mul_250[3] + kernel_img_mul_250[4] + kernel_img_mul_250[5] + 
                kernel_img_mul_250[6] + kernel_img_mul_250[7] + kernel_img_mul_250[8] + 
                kernel_img_mul_250[9] + kernel_img_mul_250[10] + kernel_img_mul_250[11] + 
                kernel_img_mul_250[12] + kernel_img_mul_250[13] + kernel_img_mul_250[14] + 
                kernel_img_mul_250[15] + kernel_img_mul_250[16] + kernel_img_mul_250[17] + 
                kernel_img_mul_250[18] + kernel_img_mul_250[19] + kernel_img_mul_250[20] + 
                kernel_img_mul_250[21] + kernel_img_mul_250[22] + kernel_img_mul_250[23] + 
                kernel_img_mul_250[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2007:2000] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2007:2000] <= kernel_img_sum_250[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2007:2000] <= 'd0;
end

wire  [39:0]  kernel_img_mul_251[0:24];
assign kernel_img_mul_251[0] = buffer_data_4[1999:1992] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_251[1] = buffer_data_4[2007:2000] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_251[2] = buffer_data_4[2015:2008] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_251[3] = buffer_data_4[2023:2016] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_251[4] = buffer_data_4[2031:2024] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_251[5] = buffer_data_3[1999:1992] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_251[6] = buffer_data_3[2007:2000] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_251[7] = buffer_data_3[2015:2008] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_251[8] = buffer_data_3[2023:2016] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_251[9] = buffer_data_3[2031:2024] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_251[10] = buffer_data_2[1999:1992] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_251[11] = buffer_data_2[2007:2000] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_251[12] = buffer_data_2[2015:2008] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_251[13] = buffer_data_2[2023:2016] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_251[14] = buffer_data_2[2031:2024] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_251[15] = buffer_data_1[1999:1992] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_251[16] = buffer_data_1[2007:2000] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_251[17] = buffer_data_1[2015:2008] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_251[18] = buffer_data_1[2023:2016] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_251[19] = buffer_data_1[2031:2024] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_251[20] = buffer_data_0[1999:1992] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_251[21] = buffer_data_0[2007:2000] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_251[22] = buffer_data_0[2015:2008] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_251[23] = buffer_data_0[2023:2016] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_251[24] = buffer_data_0[2031:2024] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_251 = kernel_img_mul_251[0] + kernel_img_mul_251[1] + kernel_img_mul_251[2] + 
                kernel_img_mul_251[3] + kernel_img_mul_251[4] + kernel_img_mul_251[5] + 
                kernel_img_mul_251[6] + kernel_img_mul_251[7] + kernel_img_mul_251[8] + 
                kernel_img_mul_251[9] + kernel_img_mul_251[10] + kernel_img_mul_251[11] + 
                kernel_img_mul_251[12] + kernel_img_mul_251[13] + kernel_img_mul_251[14] + 
                kernel_img_mul_251[15] + kernel_img_mul_251[16] + kernel_img_mul_251[17] + 
                kernel_img_mul_251[18] + kernel_img_mul_251[19] + kernel_img_mul_251[20] + 
                kernel_img_mul_251[21] + kernel_img_mul_251[22] + kernel_img_mul_251[23] + 
                kernel_img_mul_251[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2015:2008] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2015:2008] <= kernel_img_sum_251[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2015:2008] <= 'd0;
end

wire  [39:0]  kernel_img_mul_252[0:24];
assign kernel_img_mul_252[0] = buffer_data_4[2007:2000] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_252[1] = buffer_data_4[2015:2008] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_252[2] = buffer_data_4[2023:2016] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_252[3] = buffer_data_4[2031:2024] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_252[4] = buffer_data_4[2039:2032] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_252[5] = buffer_data_3[2007:2000] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_252[6] = buffer_data_3[2015:2008] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_252[7] = buffer_data_3[2023:2016] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_252[8] = buffer_data_3[2031:2024] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_252[9] = buffer_data_3[2039:2032] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_252[10] = buffer_data_2[2007:2000] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_252[11] = buffer_data_2[2015:2008] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_252[12] = buffer_data_2[2023:2016] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_252[13] = buffer_data_2[2031:2024] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_252[14] = buffer_data_2[2039:2032] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_252[15] = buffer_data_1[2007:2000] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_252[16] = buffer_data_1[2015:2008] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_252[17] = buffer_data_1[2023:2016] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_252[18] = buffer_data_1[2031:2024] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_252[19] = buffer_data_1[2039:2032] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_252[20] = buffer_data_0[2007:2000] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_252[21] = buffer_data_0[2015:2008] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_252[22] = buffer_data_0[2023:2016] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_252[23] = buffer_data_0[2031:2024] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_252[24] = buffer_data_0[2039:2032] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_252 = kernel_img_mul_252[0] + kernel_img_mul_252[1] + kernel_img_mul_252[2] + 
                kernel_img_mul_252[3] + kernel_img_mul_252[4] + kernel_img_mul_252[5] + 
                kernel_img_mul_252[6] + kernel_img_mul_252[7] + kernel_img_mul_252[8] + 
                kernel_img_mul_252[9] + kernel_img_mul_252[10] + kernel_img_mul_252[11] + 
                kernel_img_mul_252[12] + kernel_img_mul_252[13] + kernel_img_mul_252[14] + 
                kernel_img_mul_252[15] + kernel_img_mul_252[16] + kernel_img_mul_252[17] + 
                kernel_img_mul_252[18] + kernel_img_mul_252[19] + kernel_img_mul_252[20] + 
                kernel_img_mul_252[21] + kernel_img_mul_252[22] + kernel_img_mul_252[23] + 
                kernel_img_mul_252[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2023:2016] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2023:2016] <= kernel_img_sum_252[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2023:2016] <= 'd0;
end

wire  [39:0]  kernel_img_mul_253[0:24];
assign kernel_img_mul_253[0] = buffer_data_4[2015:2008] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_253[1] = buffer_data_4[2023:2016] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_253[2] = buffer_data_4[2031:2024] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_253[3] = buffer_data_4[2039:2032] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_253[4] = buffer_data_4[2047:2040] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_253[5] = buffer_data_3[2015:2008] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_253[6] = buffer_data_3[2023:2016] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_253[7] = buffer_data_3[2031:2024] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_253[8] = buffer_data_3[2039:2032] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_253[9] = buffer_data_3[2047:2040] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_253[10] = buffer_data_2[2015:2008] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_253[11] = buffer_data_2[2023:2016] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_253[12] = buffer_data_2[2031:2024] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_253[13] = buffer_data_2[2039:2032] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_253[14] = buffer_data_2[2047:2040] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_253[15] = buffer_data_1[2015:2008] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_253[16] = buffer_data_1[2023:2016] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_253[17] = buffer_data_1[2031:2024] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_253[18] = buffer_data_1[2039:2032] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_253[19] = buffer_data_1[2047:2040] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_253[20] = buffer_data_0[2015:2008] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_253[21] = buffer_data_0[2023:2016] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_253[22] = buffer_data_0[2031:2024] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_253[23] = buffer_data_0[2039:2032] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_253[24] = buffer_data_0[2047:2040] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_253 = kernel_img_mul_253[0] + kernel_img_mul_253[1] + kernel_img_mul_253[2] + 
                kernel_img_mul_253[3] + kernel_img_mul_253[4] + kernel_img_mul_253[5] + 
                kernel_img_mul_253[6] + kernel_img_mul_253[7] + kernel_img_mul_253[8] + 
                kernel_img_mul_253[9] + kernel_img_mul_253[10] + kernel_img_mul_253[11] + 
                kernel_img_mul_253[12] + kernel_img_mul_253[13] + kernel_img_mul_253[14] + 
                kernel_img_mul_253[15] + kernel_img_mul_253[16] + kernel_img_mul_253[17] + 
                kernel_img_mul_253[18] + kernel_img_mul_253[19] + kernel_img_mul_253[20] + 
                kernel_img_mul_253[21] + kernel_img_mul_253[22] + kernel_img_mul_253[23] + 
                kernel_img_mul_253[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2031:2024] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2031:2024] <= kernel_img_sum_253[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2031:2024] <= 'd0;
end

wire  [39:0]  kernel_img_mul_254[0:24];
assign kernel_img_mul_254[0] = buffer_data_4[2023:2016] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_254[1] = buffer_data_4[2031:2024] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_254[2] = buffer_data_4[2039:2032] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_254[3] = buffer_data_4[2047:2040] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_254[4] = buffer_data_4[2055:2048] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_254[5] = buffer_data_3[2023:2016] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_254[6] = buffer_data_3[2031:2024] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_254[7] = buffer_data_3[2039:2032] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_254[8] = buffer_data_3[2047:2040] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_254[9] = buffer_data_3[2055:2048] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_254[10] = buffer_data_2[2023:2016] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_254[11] = buffer_data_2[2031:2024] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_254[12] = buffer_data_2[2039:2032] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_254[13] = buffer_data_2[2047:2040] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_254[14] = buffer_data_2[2055:2048] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_254[15] = buffer_data_1[2023:2016] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_254[16] = buffer_data_1[2031:2024] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_254[17] = buffer_data_1[2039:2032] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_254[18] = buffer_data_1[2047:2040] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_254[19] = buffer_data_1[2055:2048] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_254[20] = buffer_data_0[2023:2016] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_254[21] = buffer_data_0[2031:2024] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_254[22] = buffer_data_0[2039:2032] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_254[23] = buffer_data_0[2047:2040] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_254[24] = buffer_data_0[2055:2048] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_254 = kernel_img_mul_254[0] + kernel_img_mul_254[1] + kernel_img_mul_254[2] + 
                kernel_img_mul_254[3] + kernel_img_mul_254[4] + kernel_img_mul_254[5] + 
                kernel_img_mul_254[6] + kernel_img_mul_254[7] + kernel_img_mul_254[8] + 
                kernel_img_mul_254[9] + kernel_img_mul_254[10] + kernel_img_mul_254[11] + 
                kernel_img_mul_254[12] + kernel_img_mul_254[13] + kernel_img_mul_254[14] + 
                kernel_img_mul_254[15] + kernel_img_mul_254[16] + kernel_img_mul_254[17] + 
                kernel_img_mul_254[18] + kernel_img_mul_254[19] + kernel_img_mul_254[20] + 
                kernel_img_mul_254[21] + kernel_img_mul_254[22] + kernel_img_mul_254[23] + 
                kernel_img_mul_254[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2039:2032] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2039:2032] <= kernel_img_sum_254[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2039:2032] <= 'd0;
end

wire  [39:0]  kernel_img_mul_255[0:24];
assign kernel_img_mul_255[0] = buffer_data_4[2031:2024] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_255[1] = buffer_data_4[2039:2032] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_255[2] = buffer_data_4[2047:2040] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_255[3] = buffer_data_4[2055:2048] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_255[4] = buffer_data_4[2063:2056] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_255[5] = buffer_data_3[2031:2024] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_255[6] = buffer_data_3[2039:2032] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_255[7] = buffer_data_3[2047:2040] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_255[8] = buffer_data_3[2055:2048] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_255[9] = buffer_data_3[2063:2056] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_255[10] = buffer_data_2[2031:2024] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_255[11] = buffer_data_2[2039:2032] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_255[12] = buffer_data_2[2047:2040] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_255[13] = buffer_data_2[2055:2048] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_255[14] = buffer_data_2[2063:2056] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_255[15] = buffer_data_1[2031:2024] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_255[16] = buffer_data_1[2039:2032] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_255[17] = buffer_data_1[2047:2040] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_255[18] = buffer_data_1[2055:2048] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_255[19] = buffer_data_1[2063:2056] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_255[20] = buffer_data_0[2031:2024] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_255[21] = buffer_data_0[2039:2032] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_255[22] = buffer_data_0[2047:2040] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_255[23] = buffer_data_0[2055:2048] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_255[24] = buffer_data_0[2063:2056] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_255 = kernel_img_mul_255[0] + kernel_img_mul_255[1] + kernel_img_mul_255[2] + 
                kernel_img_mul_255[3] + kernel_img_mul_255[4] + kernel_img_mul_255[5] + 
                kernel_img_mul_255[6] + kernel_img_mul_255[7] + kernel_img_mul_255[8] + 
                kernel_img_mul_255[9] + kernel_img_mul_255[10] + kernel_img_mul_255[11] + 
                kernel_img_mul_255[12] + kernel_img_mul_255[13] + kernel_img_mul_255[14] + 
                kernel_img_mul_255[15] + kernel_img_mul_255[16] + kernel_img_mul_255[17] + 
                kernel_img_mul_255[18] + kernel_img_mul_255[19] + kernel_img_mul_255[20] + 
                kernel_img_mul_255[21] + kernel_img_mul_255[22] + kernel_img_mul_255[23] + 
                kernel_img_mul_255[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2047:2040] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2047:2040] <= kernel_img_sum_255[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2047:2040] <= 'd0;
end

wire  [39:0]  kernel_img_mul_256[0:24];
assign kernel_img_mul_256[0] = buffer_data_4[2039:2032] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_256[1] = buffer_data_4[2047:2040] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_256[2] = buffer_data_4[2055:2048] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_256[3] = buffer_data_4[2063:2056] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_256[4] = buffer_data_4[2071:2064] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_256[5] = buffer_data_3[2039:2032] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_256[6] = buffer_data_3[2047:2040] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_256[7] = buffer_data_3[2055:2048] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_256[8] = buffer_data_3[2063:2056] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_256[9] = buffer_data_3[2071:2064] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_256[10] = buffer_data_2[2039:2032] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_256[11] = buffer_data_2[2047:2040] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_256[12] = buffer_data_2[2055:2048] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_256[13] = buffer_data_2[2063:2056] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_256[14] = buffer_data_2[2071:2064] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_256[15] = buffer_data_1[2039:2032] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_256[16] = buffer_data_1[2047:2040] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_256[17] = buffer_data_1[2055:2048] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_256[18] = buffer_data_1[2063:2056] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_256[19] = buffer_data_1[2071:2064] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_256[20] = buffer_data_0[2039:2032] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_256[21] = buffer_data_0[2047:2040] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_256[22] = buffer_data_0[2055:2048] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_256[23] = buffer_data_0[2063:2056] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_256[24] = buffer_data_0[2071:2064] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_256 = kernel_img_mul_256[0] + kernel_img_mul_256[1] + kernel_img_mul_256[2] + 
                kernel_img_mul_256[3] + kernel_img_mul_256[4] + kernel_img_mul_256[5] + 
                kernel_img_mul_256[6] + kernel_img_mul_256[7] + kernel_img_mul_256[8] + 
                kernel_img_mul_256[9] + kernel_img_mul_256[10] + kernel_img_mul_256[11] + 
                kernel_img_mul_256[12] + kernel_img_mul_256[13] + kernel_img_mul_256[14] + 
                kernel_img_mul_256[15] + kernel_img_mul_256[16] + kernel_img_mul_256[17] + 
                kernel_img_mul_256[18] + kernel_img_mul_256[19] + kernel_img_mul_256[20] + 
                kernel_img_mul_256[21] + kernel_img_mul_256[22] + kernel_img_mul_256[23] + 
                kernel_img_mul_256[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2055:2048] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2055:2048] <= kernel_img_sum_256[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2055:2048] <= 'd0;
end

wire  [39:0]  kernel_img_mul_257[0:24];
assign kernel_img_mul_257[0] = buffer_data_4[2047:2040] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_257[1] = buffer_data_4[2055:2048] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_257[2] = buffer_data_4[2063:2056] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_257[3] = buffer_data_4[2071:2064] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_257[4] = buffer_data_4[2079:2072] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_257[5] = buffer_data_3[2047:2040] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_257[6] = buffer_data_3[2055:2048] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_257[7] = buffer_data_3[2063:2056] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_257[8] = buffer_data_3[2071:2064] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_257[9] = buffer_data_3[2079:2072] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_257[10] = buffer_data_2[2047:2040] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_257[11] = buffer_data_2[2055:2048] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_257[12] = buffer_data_2[2063:2056] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_257[13] = buffer_data_2[2071:2064] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_257[14] = buffer_data_2[2079:2072] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_257[15] = buffer_data_1[2047:2040] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_257[16] = buffer_data_1[2055:2048] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_257[17] = buffer_data_1[2063:2056] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_257[18] = buffer_data_1[2071:2064] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_257[19] = buffer_data_1[2079:2072] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_257[20] = buffer_data_0[2047:2040] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_257[21] = buffer_data_0[2055:2048] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_257[22] = buffer_data_0[2063:2056] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_257[23] = buffer_data_0[2071:2064] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_257[24] = buffer_data_0[2079:2072] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_257 = kernel_img_mul_257[0] + kernel_img_mul_257[1] + kernel_img_mul_257[2] + 
                kernel_img_mul_257[3] + kernel_img_mul_257[4] + kernel_img_mul_257[5] + 
                kernel_img_mul_257[6] + kernel_img_mul_257[7] + kernel_img_mul_257[8] + 
                kernel_img_mul_257[9] + kernel_img_mul_257[10] + kernel_img_mul_257[11] + 
                kernel_img_mul_257[12] + kernel_img_mul_257[13] + kernel_img_mul_257[14] + 
                kernel_img_mul_257[15] + kernel_img_mul_257[16] + kernel_img_mul_257[17] + 
                kernel_img_mul_257[18] + kernel_img_mul_257[19] + kernel_img_mul_257[20] + 
                kernel_img_mul_257[21] + kernel_img_mul_257[22] + kernel_img_mul_257[23] + 
                kernel_img_mul_257[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2063:2056] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2063:2056] <= kernel_img_sum_257[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2063:2056] <= 'd0;
end

wire  [39:0]  kernel_img_mul_258[0:24];
assign kernel_img_mul_258[0] = buffer_data_4[2055:2048] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_258[1] = buffer_data_4[2063:2056] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_258[2] = buffer_data_4[2071:2064] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_258[3] = buffer_data_4[2079:2072] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_258[4] = buffer_data_4[2087:2080] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_258[5] = buffer_data_3[2055:2048] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_258[6] = buffer_data_3[2063:2056] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_258[7] = buffer_data_3[2071:2064] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_258[8] = buffer_data_3[2079:2072] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_258[9] = buffer_data_3[2087:2080] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_258[10] = buffer_data_2[2055:2048] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_258[11] = buffer_data_2[2063:2056] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_258[12] = buffer_data_2[2071:2064] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_258[13] = buffer_data_2[2079:2072] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_258[14] = buffer_data_2[2087:2080] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_258[15] = buffer_data_1[2055:2048] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_258[16] = buffer_data_1[2063:2056] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_258[17] = buffer_data_1[2071:2064] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_258[18] = buffer_data_1[2079:2072] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_258[19] = buffer_data_1[2087:2080] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_258[20] = buffer_data_0[2055:2048] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_258[21] = buffer_data_0[2063:2056] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_258[22] = buffer_data_0[2071:2064] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_258[23] = buffer_data_0[2079:2072] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_258[24] = buffer_data_0[2087:2080] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_258 = kernel_img_mul_258[0] + kernel_img_mul_258[1] + kernel_img_mul_258[2] + 
                kernel_img_mul_258[3] + kernel_img_mul_258[4] + kernel_img_mul_258[5] + 
                kernel_img_mul_258[6] + kernel_img_mul_258[7] + kernel_img_mul_258[8] + 
                kernel_img_mul_258[9] + kernel_img_mul_258[10] + kernel_img_mul_258[11] + 
                kernel_img_mul_258[12] + kernel_img_mul_258[13] + kernel_img_mul_258[14] + 
                kernel_img_mul_258[15] + kernel_img_mul_258[16] + kernel_img_mul_258[17] + 
                kernel_img_mul_258[18] + kernel_img_mul_258[19] + kernel_img_mul_258[20] + 
                kernel_img_mul_258[21] + kernel_img_mul_258[22] + kernel_img_mul_258[23] + 
                kernel_img_mul_258[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2071:2064] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2071:2064] <= kernel_img_sum_258[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2071:2064] <= 'd0;
end

wire  [39:0]  kernel_img_mul_259[0:24];
assign kernel_img_mul_259[0] = buffer_data_4[2063:2056] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_259[1] = buffer_data_4[2071:2064] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_259[2] = buffer_data_4[2079:2072] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_259[3] = buffer_data_4[2087:2080] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_259[4] = buffer_data_4[2095:2088] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_259[5] = buffer_data_3[2063:2056] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_259[6] = buffer_data_3[2071:2064] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_259[7] = buffer_data_3[2079:2072] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_259[8] = buffer_data_3[2087:2080] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_259[9] = buffer_data_3[2095:2088] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_259[10] = buffer_data_2[2063:2056] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_259[11] = buffer_data_2[2071:2064] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_259[12] = buffer_data_2[2079:2072] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_259[13] = buffer_data_2[2087:2080] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_259[14] = buffer_data_2[2095:2088] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_259[15] = buffer_data_1[2063:2056] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_259[16] = buffer_data_1[2071:2064] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_259[17] = buffer_data_1[2079:2072] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_259[18] = buffer_data_1[2087:2080] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_259[19] = buffer_data_1[2095:2088] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_259[20] = buffer_data_0[2063:2056] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_259[21] = buffer_data_0[2071:2064] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_259[22] = buffer_data_0[2079:2072] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_259[23] = buffer_data_0[2087:2080] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_259[24] = buffer_data_0[2095:2088] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_259 = kernel_img_mul_259[0] + kernel_img_mul_259[1] + kernel_img_mul_259[2] + 
                kernel_img_mul_259[3] + kernel_img_mul_259[4] + kernel_img_mul_259[5] + 
                kernel_img_mul_259[6] + kernel_img_mul_259[7] + kernel_img_mul_259[8] + 
                kernel_img_mul_259[9] + kernel_img_mul_259[10] + kernel_img_mul_259[11] + 
                kernel_img_mul_259[12] + kernel_img_mul_259[13] + kernel_img_mul_259[14] + 
                kernel_img_mul_259[15] + kernel_img_mul_259[16] + kernel_img_mul_259[17] + 
                kernel_img_mul_259[18] + kernel_img_mul_259[19] + kernel_img_mul_259[20] + 
                kernel_img_mul_259[21] + kernel_img_mul_259[22] + kernel_img_mul_259[23] + 
                kernel_img_mul_259[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2079:2072] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2079:2072] <= kernel_img_sum_259[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2079:2072] <= 'd0;
end

wire  [39:0]  kernel_img_mul_260[0:24];
assign kernel_img_mul_260[0] = buffer_data_4[2071:2064] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_260[1] = buffer_data_4[2079:2072] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_260[2] = buffer_data_4[2087:2080] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_260[3] = buffer_data_4[2095:2088] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_260[4] = buffer_data_4[2103:2096] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_260[5] = buffer_data_3[2071:2064] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_260[6] = buffer_data_3[2079:2072] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_260[7] = buffer_data_3[2087:2080] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_260[8] = buffer_data_3[2095:2088] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_260[9] = buffer_data_3[2103:2096] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_260[10] = buffer_data_2[2071:2064] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_260[11] = buffer_data_2[2079:2072] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_260[12] = buffer_data_2[2087:2080] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_260[13] = buffer_data_2[2095:2088] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_260[14] = buffer_data_2[2103:2096] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_260[15] = buffer_data_1[2071:2064] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_260[16] = buffer_data_1[2079:2072] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_260[17] = buffer_data_1[2087:2080] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_260[18] = buffer_data_1[2095:2088] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_260[19] = buffer_data_1[2103:2096] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_260[20] = buffer_data_0[2071:2064] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_260[21] = buffer_data_0[2079:2072] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_260[22] = buffer_data_0[2087:2080] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_260[23] = buffer_data_0[2095:2088] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_260[24] = buffer_data_0[2103:2096] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_260 = kernel_img_mul_260[0] + kernel_img_mul_260[1] + kernel_img_mul_260[2] + 
                kernel_img_mul_260[3] + kernel_img_mul_260[4] + kernel_img_mul_260[5] + 
                kernel_img_mul_260[6] + kernel_img_mul_260[7] + kernel_img_mul_260[8] + 
                kernel_img_mul_260[9] + kernel_img_mul_260[10] + kernel_img_mul_260[11] + 
                kernel_img_mul_260[12] + kernel_img_mul_260[13] + kernel_img_mul_260[14] + 
                kernel_img_mul_260[15] + kernel_img_mul_260[16] + kernel_img_mul_260[17] + 
                kernel_img_mul_260[18] + kernel_img_mul_260[19] + kernel_img_mul_260[20] + 
                kernel_img_mul_260[21] + kernel_img_mul_260[22] + kernel_img_mul_260[23] + 
                kernel_img_mul_260[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2087:2080] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2087:2080] <= kernel_img_sum_260[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2087:2080] <= 'd0;
end

wire  [39:0]  kernel_img_mul_261[0:24];
assign kernel_img_mul_261[0] = buffer_data_4[2079:2072] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_261[1] = buffer_data_4[2087:2080] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_261[2] = buffer_data_4[2095:2088] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_261[3] = buffer_data_4[2103:2096] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_261[4] = buffer_data_4[2111:2104] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_261[5] = buffer_data_3[2079:2072] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_261[6] = buffer_data_3[2087:2080] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_261[7] = buffer_data_3[2095:2088] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_261[8] = buffer_data_3[2103:2096] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_261[9] = buffer_data_3[2111:2104] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_261[10] = buffer_data_2[2079:2072] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_261[11] = buffer_data_2[2087:2080] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_261[12] = buffer_data_2[2095:2088] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_261[13] = buffer_data_2[2103:2096] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_261[14] = buffer_data_2[2111:2104] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_261[15] = buffer_data_1[2079:2072] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_261[16] = buffer_data_1[2087:2080] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_261[17] = buffer_data_1[2095:2088] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_261[18] = buffer_data_1[2103:2096] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_261[19] = buffer_data_1[2111:2104] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_261[20] = buffer_data_0[2079:2072] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_261[21] = buffer_data_0[2087:2080] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_261[22] = buffer_data_0[2095:2088] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_261[23] = buffer_data_0[2103:2096] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_261[24] = buffer_data_0[2111:2104] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_261 = kernel_img_mul_261[0] + kernel_img_mul_261[1] + kernel_img_mul_261[2] + 
                kernel_img_mul_261[3] + kernel_img_mul_261[4] + kernel_img_mul_261[5] + 
                kernel_img_mul_261[6] + kernel_img_mul_261[7] + kernel_img_mul_261[8] + 
                kernel_img_mul_261[9] + kernel_img_mul_261[10] + kernel_img_mul_261[11] + 
                kernel_img_mul_261[12] + kernel_img_mul_261[13] + kernel_img_mul_261[14] + 
                kernel_img_mul_261[15] + kernel_img_mul_261[16] + kernel_img_mul_261[17] + 
                kernel_img_mul_261[18] + kernel_img_mul_261[19] + kernel_img_mul_261[20] + 
                kernel_img_mul_261[21] + kernel_img_mul_261[22] + kernel_img_mul_261[23] + 
                kernel_img_mul_261[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2095:2088] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2095:2088] <= kernel_img_sum_261[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2095:2088] <= 'd0;
end

wire  [39:0]  kernel_img_mul_262[0:24];
assign kernel_img_mul_262[0] = buffer_data_4[2087:2080] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_262[1] = buffer_data_4[2095:2088] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_262[2] = buffer_data_4[2103:2096] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_262[3] = buffer_data_4[2111:2104] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_262[4] = buffer_data_4[2119:2112] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_262[5] = buffer_data_3[2087:2080] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_262[6] = buffer_data_3[2095:2088] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_262[7] = buffer_data_3[2103:2096] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_262[8] = buffer_data_3[2111:2104] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_262[9] = buffer_data_3[2119:2112] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_262[10] = buffer_data_2[2087:2080] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_262[11] = buffer_data_2[2095:2088] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_262[12] = buffer_data_2[2103:2096] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_262[13] = buffer_data_2[2111:2104] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_262[14] = buffer_data_2[2119:2112] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_262[15] = buffer_data_1[2087:2080] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_262[16] = buffer_data_1[2095:2088] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_262[17] = buffer_data_1[2103:2096] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_262[18] = buffer_data_1[2111:2104] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_262[19] = buffer_data_1[2119:2112] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_262[20] = buffer_data_0[2087:2080] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_262[21] = buffer_data_0[2095:2088] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_262[22] = buffer_data_0[2103:2096] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_262[23] = buffer_data_0[2111:2104] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_262[24] = buffer_data_0[2119:2112] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_262 = kernel_img_mul_262[0] + kernel_img_mul_262[1] + kernel_img_mul_262[2] + 
                kernel_img_mul_262[3] + kernel_img_mul_262[4] + kernel_img_mul_262[5] + 
                kernel_img_mul_262[6] + kernel_img_mul_262[7] + kernel_img_mul_262[8] + 
                kernel_img_mul_262[9] + kernel_img_mul_262[10] + kernel_img_mul_262[11] + 
                kernel_img_mul_262[12] + kernel_img_mul_262[13] + kernel_img_mul_262[14] + 
                kernel_img_mul_262[15] + kernel_img_mul_262[16] + kernel_img_mul_262[17] + 
                kernel_img_mul_262[18] + kernel_img_mul_262[19] + kernel_img_mul_262[20] + 
                kernel_img_mul_262[21] + kernel_img_mul_262[22] + kernel_img_mul_262[23] + 
                kernel_img_mul_262[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2103:2096] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2103:2096] <= kernel_img_sum_262[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2103:2096] <= 'd0;
end

wire  [39:0]  kernel_img_mul_263[0:24];
assign kernel_img_mul_263[0] = buffer_data_4[2095:2088] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_263[1] = buffer_data_4[2103:2096] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_263[2] = buffer_data_4[2111:2104] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_263[3] = buffer_data_4[2119:2112] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_263[4] = buffer_data_4[2127:2120] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_263[5] = buffer_data_3[2095:2088] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_263[6] = buffer_data_3[2103:2096] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_263[7] = buffer_data_3[2111:2104] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_263[8] = buffer_data_3[2119:2112] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_263[9] = buffer_data_3[2127:2120] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_263[10] = buffer_data_2[2095:2088] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_263[11] = buffer_data_2[2103:2096] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_263[12] = buffer_data_2[2111:2104] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_263[13] = buffer_data_2[2119:2112] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_263[14] = buffer_data_2[2127:2120] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_263[15] = buffer_data_1[2095:2088] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_263[16] = buffer_data_1[2103:2096] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_263[17] = buffer_data_1[2111:2104] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_263[18] = buffer_data_1[2119:2112] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_263[19] = buffer_data_1[2127:2120] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_263[20] = buffer_data_0[2095:2088] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_263[21] = buffer_data_0[2103:2096] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_263[22] = buffer_data_0[2111:2104] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_263[23] = buffer_data_0[2119:2112] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_263[24] = buffer_data_0[2127:2120] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_263 = kernel_img_mul_263[0] + kernel_img_mul_263[1] + kernel_img_mul_263[2] + 
                kernel_img_mul_263[3] + kernel_img_mul_263[4] + kernel_img_mul_263[5] + 
                kernel_img_mul_263[6] + kernel_img_mul_263[7] + kernel_img_mul_263[8] + 
                kernel_img_mul_263[9] + kernel_img_mul_263[10] + kernel_img_mul_263[11] + 
                kernel_img_mul_263[12] + kernel_img_mul_263[13] + kernel_img_mul_263[14] + 
                kernel_img_mul_263[15] + kernel_img_mul_263[16] + kernel_img_mul_263[17] + 
                kernel_img_mul_263[18] + kernel_img_mul_263[19] + kernel_img_mul_263[20] + 
                kernel_img_mul_263[21] + kernel_img_mul_263[22] + kernel_img_mul_263[23] + 
                kernel_img_mul_263[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2111:2104] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2111:2104] <= kernel_img_sum_263[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2111:2104] <= 'd0;
end

wire  [39:0]  kernel_img_mul_264[0:24];
assign kernel_img_mul_264[0] = buffer_data_4[2103:2096] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_264[1] = buffer_data_4[2111:2104] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_264[2] = buffer_data_4[2119:2112] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_264[3] = buffer_data_4[2127:2120] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_264[4] = buffer_data_4[2135:2128] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_264[5] = buffer_data_3[2103:2096] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_264[6] = buffer_data_3[2111:2104] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_264[7] = buffer_data_3[2119:2112] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_264[8] = buffer_data_3[2127:2120] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_264[9] = buffer_data_3[2135:2128] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_264[10] = buffer_data_2[2103:2096] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_264[11] = buffer_data_2[2111:2104] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_264[12] = buffer_data_2[2119:2112] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_264[13] = buffer_data_2[2127:2120] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_264[14] = buffer_data_2[2135:2128] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_264[15] = buffer_data_1[2103:2096] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_264[16] = buffer_data_1[2111:2104] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_264[17] = buffer_data_1[2119:2112] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_264[18] = buffer_data_1[2127:2120] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_264[19] = buffer_data_1[2135:2128] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_264[20] = buffer_data_0[2103:2096] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_264[21] = buffer_data_0[2111:2104] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_264[22] = buffer_data_0[2119:2112] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_264[23] = buffer_data_0[2127:2120] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_264[24] = buffer_data_0[2135:2128] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_264 = kernel_img_mul_264[0] + kernel_img_mul_264[1] + kernel_img_mul_264[2] + 
                kernel_img_mul_264[3] + kernel_img_mul_264[4] + kernel_img_mul_264[5] + 
                kernel_img_mul_264[6] + kernel_img_mul_264[7] + kernel_img_mul_264[8] + 
                kernel_img_mul_264[9] + kernel_img_mul_264[10] + kernel_img_mul_264[11] + 
                kernel_img_mul_264[12] + kernel_img_mul_264[13] + kernel_img_mul_264[14] + 
                kernel_img_mul_264[15] + kernel_img_mul_264[16] + kernel_img_mul_264[17] + 
                kernel_img_mul_264[18] + kernel_img_mul_264[19] + kernel_img_mul_264[20] + 
                kernel_img_mul_264[21] + kernel_img_mul_264[22] + kernel_img_mul_264[23] + 
                kernel_img_mul_264[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2119:2112] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2119:2112] <= kernel_img_sum_264[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2119:2112] <= 'd0;
end

wire  [39:0]  kernel_img_mul_265[0:24];
assign kernel_img_mul_265[0] = buffer_data_4[2111:2104] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_265[1] = buffer_data_4[2119:2112] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_265[2] = buffer_data_4[2127:2120] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_265[3] = buffer_data_4[2135:2128] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_265[4] = buffer_data_4[2143:2136] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_265[5] = buffer_data_3[2111:2104] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_265[6] = buffer_data_3[2119:2112] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_265[7] = buffer_data_3[2127:2120] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_265[8] = buffer_data_3[2135:2128] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_265[9] = buffer_data_3[2143:2136] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_265[10] = buffer_data_2[2111:2104] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_265[11] = buffer_data_2[2119:2112] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_265[12] = buffer_data_2[2127:2120] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_265[13] = buffer_data_2[2135:2128] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_265[14] = buffer_data_2[2143:2136] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_265[15] = buffer_data_1[2111:2104] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_265[16] = buffer_data_1[2119:2112] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_265[17] = buffer_data_1[2127:2120] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_265[18] = buffer_data_1[2135:2128] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_265[19] = buffer_data_1[2143:2136] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_265[20] = buffer_data_0[2111:2104] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_265[21] = buffer_data_0[2119:2112] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_265[22] = buffer_data_0[2127:2120] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_265[23] = buffer_data_0[2135:2128] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_265[24] = buffer_data_0[2143:2136] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_265 = kernel_img_mul_265[0] + kernel_img_mul_265[1] + kernel_img_mul_265[2] + 
                kernel_img_mul_265[3] + kernel_img_mul_265[4] + kernel_img_mul_265[5] + 
                kernel_img_mul_265[6] + kernel_img_mul_265[7] + kernel_img_mul_265[8] + 
                kernel_img_mul_265[9] + kernel_img_mul_265[10] + kernel_img_mul_265[11] + 
                kernel_img_mul_265[12] + kernel_img_mul_265[13] + kernel_img_mul_265[14] + 
                kernel_img_mul_265[15] + kernel_img_mul_265[16] + kernel_img_mul_265[17] + 
                kernel_img_mul_265[18] + kernel_img_mul_265[19] + kernel_img_mul_265[20] + 
                kernel_img_mul_265[21] + kernel_img_mul_265[22] + kernel_img_mul_265[23] + 
                kernel_img_mul_265[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2127:2120] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2127:2120] <= kernel_img_sum_265[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2127:2120] <= 'd0;
end

wire  [39:0]  kernel_img_mul_266[0:24];
assign kernel_img_mul_266[0] = buffer_data_4[2119:2112] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_266[1] = buffer_data_4[2127:2120] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_266[2] = buffer_data_4[2135:2128] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_266[3] = buffer_data_4[2143:2136] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_266[4] = buffer_data_4[2151:2144] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_266[5] = buffer_data_3[2119:2112] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_266[6] = buffer_data_3[2127:2120] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_266[7] = buffer_data_3[2135:2128] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_266[8] = buffer_data_3[2143:2136] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_266[9] = buffer_data_3[2151:2144] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_266[10] = buffer_data_2[2119:2112] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_266[11] = buffer_data_2[2127:2120] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_266[12] = buffer_data_2[2135:2128] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_266[13] = buffer_data_2[2143:2136] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_266[14] = buffer_data_2[2151:2144] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_266[15] = buffer_data_1[2119:2112] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_266[16] = buffer_data_1[2127:2120] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_266[17] = buffer_data_1[2135:2128] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_266[18] = buffer_data_1[2143:2136] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_266[19] = buffer_data_1[2151:2144] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_266[20] = buffer_data_0[2119:2112] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_266[21] = buffer_data_0[2127:2120] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_266[22] = buffer_data_0[2135:2128] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_266[23] = buffer_data_0[2143:2136] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_266[24] = buffer_data_0[2151:2144] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_266 = kernel_img_mul_266[0] + kernel_img_mul_266[1] + kernel_img_mul_266[2] + 
                kernel_img_mul_266[3] + kernel_img_mul_266[4] + kernel_img_mul_266[5] + 
                kernel_img_mul_266[6] + kernel_img_mul_266[7] + kernel_img_mul_266[8] + 
                kernel_img_mul_266[9] + kernel_img_mul_266[10] + kernel_img_mul_266[11] + 
                kernel_img_mul_266[12] + kernel_img_mul_266[13] + kernel_img_mul_266[14] + 
                kernel_img_mul_266[15] + kernel_img_mul_266[16] + kernel_img_mul_266[17] + 
                kernel_img_mul_266[18] + kernel_img_mul_266[19] + kernel_img_mul_266[20] + 
                kernel_img_mul_266[21] + kernel_img_mul_266[22] + kernel_img_mul_266[23] + 
                kernel_img_mul_266[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2135:2128] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2135:2128] <= kernel_img_sum_266[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2135:2128] <= 'd0;
end

wire  [39:0]  kernel_img_mul_267[0:24];
assign kernel_img_mul_267[0] = buffer_data_4[2127:2120] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_267[1] = buffer_data_4[2135:2128] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_267[2] = buffer_data_4[2143:2136] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_267[3] = buffer_data_4[2151:2144] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_267[4] = buffer_data_4[2159:2152] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_267[5] = buffer_data_3[2127:2120] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_267[6] = buffer_data_3[2135:2128] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_267[7] = buffer_data_3[2143:2136] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_267[8] = buffer_data_3[2151:2144] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_267[9] = buffer_data_3[2159:2152] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_267[10] = buffer_data_2[2127:2120] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_267[11] = buffer_data_2[2135:2128] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_267[12] = buffer_data_2[2143:2136] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_267[13] = buffer_data_2[2151:2144] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_267[14] = buffer_data_2[2159:2152] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_267[15] = buffer_data_1[2127:2120] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_267[16] = buffer_data_1[2135:2128] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_267[17] = buffer_data_1[2143:2136] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_267[18] = buffer_data_1[2151:2144] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_267[19] = buffer_data_1[2159:2152] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_267[20] = buffer_data_0[2127:2120] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_267[21] = buffer_data_0[2135:2128] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_267[22] = buffer_data_0[2143:2136] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_267[23] = buffer_data_0[2151:2144] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_267[24] = buffer_data_0[2159:2152] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_267 = kernel_img_mul_267[0] + kernel_img_mul_267[1] + kernel_img_mul_267[2] + 
                kernel_img_mul_267[3] + kernel_img_mul_267[4] + kernel_img_mul_267[5] + 
                kernel_img_mul_267[6] + kernel_img_mul_267[7] + kernel_img_mul_267[8] + 
                kernel_img_mul_267[9] + kernel_img_mul_267[10] + kernel_img_mul_267[11] + 
                kernel_img_mul_267[12] + kernel_img_mul_267[13] + kernel_img_mul_267[14] + 
                kernel_img_mul_267[15] + kernel_img_mul_267[16] + kernel_img_mul_267[17] + 
                kernel_img_mul_267[18] + kernel_img_mul_267[19] + kernel_img_mul_267[20] + 
                kernel_img_mul_267[21] + kernel_img_mul_267[22] + kernel_img_mul_267[23] + 
                kernel_img_mul_267[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2143:2136] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2143:2136] <= kernel_img_sum_267[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2143:2136] <= 'd0;
end

wire  [39:0]  kernel_img_mul_268[0:24];
assign kernel_img_mul_268[0] = buffer_data_4[2135:2128] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_268[1] = buffer_data_4[2143:2136] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_268[2] = buffer_data_4[2151:2144] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_268[3] = buffer_data_4[2159:2152] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_268[4] = buffer_data_4[2167:2160] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_268[5] = buffer_data_3[2135:2128] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_268[6] = buffer_data_3[2143:2136] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_268[7] = buffer_data_3[2151:2144] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_268[8] = buffer_data_3[2159:2152] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_268[9] = buffer_data_3[2167:2160] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_268[10] = buffer_data_2[2135:2128] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_268[11] = buffer_data_2[2143:2136] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_268[12] = buffer_data_2[2151:2144] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_268[13] = buffer_data_2[2159:2152] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_268[14] = buffer_data_2[2167:2160] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_268[15] = buffer_data_1[2135:2128] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_268[16] = buffer_data_1[2143:2136] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_268[17] = buffer_data_1[2151:2144] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_268[18] = buffer_data_1[2159:2152] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_268[19] = buffer_data_1[2167:2160] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_268[20] = buffer_data_0[2135:2128] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_268[21] = buffer_data_0[2143:2136] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_268[22] = buffer_data_0[2151:2144] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_268[23] = buffer_data_0[2159:2152] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_268[24] = buffer_data_0[2167:2160] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_268 = kernel_img_mul_268[0] + kernel_img_mul_268[1] + kernel_img_mul_268[2] + 
                kernel_img_mul_268[3] + kernel_img_mul_268[4] + kernel_img_mul_268[5] + 
                kernel_img_mul_268[6] + kernel_img_mul_268[7] + kernel_img_mul_268[8] + 
                kernel_img_mul_268[9] + kernel_img_mul_268[10] + kernel_img_mul_268[11] + 
                kernel_img_mul_268[12] + kernel_img_mul_268[13] + kernel_img_mul_268[14] + 
                kernel_img_mul_268[15] + kernel_img_mul_268[16] + kernel_img_mul_268[17] + 
                kernel_img_mul_268[18] + kernel_img_mul_268[19] + kernel_img_mul_268[20] + 
                kernel_img_mul_268[21] + kernel_img_mul_268[22] + kernel_img_mul_268[23] + 
                kernel_img_mul_268[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2151:2144] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2151:2144] <= kernel_img_sum_268[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2151:2144] <= 'd0;
end

wire  [39:0]  kernel_img_mul_269[0:24];
assign kernel_img_mul_269[0] = buffer_data_4[2143:2136] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_269[1] = buffer_data_4[2151:2144] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_269[2] = buffer_data_4[2159:2152] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_269[3] = buffer_data_4[2167:2160] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_269[4] = buffer_data_4[2175:2168] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_269[5] = buffer_data_3[2143:2136] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_269[6] = buffer_data_3[2151:2144] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_269[7] = buffer_data_3[2159:2152] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_269[8] = buffer_data_3[2167:2160] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_269[9] = buffer_data_3[2175:2168] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_269[10] = buffer_data_2[2143:2136] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_269[11] = buffer_data_2[2151:2144] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_269[12] = buffer_data_2[2159:2152] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_269[13] = buffer_data_2[2167:2160] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_269[14] = buffer_data_2[2175:2168] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_269[15] = buffer_data_1[2143:2136] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_269[16] = buffer_data_1[2151:2144] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_269[17] = buffer_data_1[2159:2152] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_269[18] = buffer_data_1[2167:2160] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_269[19] = buffer_data_1[2175:2168] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_269[20] = buffer_data_0[2143:2136] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_269[21] = buffer_data_0[2151:2144] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_269[22] = buffer_data_0[2159:2152] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_269[23] = buffer_data_0[2167:2160] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_269[24] = buffer_data_0[2175:2168] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_269 = kernel_img_mul_269[0] + kernel_img_mul_269[1] + kernel_img_mul_269[2] + 
                kernel_img_mul_269[3] + kernel_img_mul_269[4] + kernel_img_mul_269[5] + 
                kernel_img_mul_269[6] + kernel_img_mul_269[7] + kernel_img_mul_269[8] + 
                kernel_img_mul_269[9] + kernel_img_mul_269[10] + kernel_img_mul_269[11] + 
                kernel_img_mul_269[12] + kernel_img_mul_269[13] + kernel_img_mul_269[14] + 
                kernel_img_mul_269[15] + kernel_img_mul_269[16] + kernel_img_mul_269[17] + 
                kernel_img_mul_269[18] + kernel_img_mul_269[19] + kernel_img_mul_269[20] + 
                kernel_img_mul_269[21] + kernel_img_mul_269[22] + kernel_img_mul_269[23] + 
                kernel_img_mul_269[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2159:2152] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2159:2152] <= kernel_img_sum_269[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2159:2152] <= 'd0;
end

wire  [39:0]  kernel_img_mul_270[0:24];
assign kernel_img_mul_270[0] = buffer_data_4[2151:2144] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_270[1] = buffer_data_4[2159:2152] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_270[2] = buffer_data_4[2167:2160] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_270[3] = buffer_data_4[2175:2168] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_270[4] = buffer_data_4[2183:2176] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_270[5] = buffer_data_3[2151:2144] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_270[6] = buffer_data_3[2159:2152] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_270[7] = buffer_data_3[2167:2160] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_270[8] = buffer_data_3[2175:2168] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_270[9] = buffer_data_3[2183:2176] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_270[10] = buffer_data_2[2151:2144] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_270[11] = buffer_data_2[2159:2152] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_270[12] = buffer_data_2[2167:2160] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_270[13] = buffer_data_2[2175:2168] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_270[14] = buffer_data_2[2183:2176] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_270[15] = buffer_data_1[2151:2144] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_270[16] = buffer_data_1[2159:2152] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_270[17] = buffer_data_1[2167:2160] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_270[18] = buffer_data_1[2175:2168] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_270[19] = buffer_data_1[2183:2176] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_270[20] = buffer_data_0[2151:2144] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_270[21] = buffer_data_0[2159:2152] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_270[22] = buffer_data_0[2167:2160] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_270[23] = buffer_data_0[2175:2168] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_270[24] = buffer_data_0[2183:2176] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_270 = kernel_img_mul_270[0] + kernel_img_mul_270[1] + kernel_img_mul_270[2] + 
                kernel_img_mul_270[3] + kernel_img_mul_270[4] + kernel_img_mul_270[5] + 
                kernel_img_mul_270[6] + kernel_img_mul_270[7] + kernel_img_mul_270[8] + 
                kernel_img_mul_270[9] + kernel_img_mul_270[10] + kernel_img_mul_270[11] + 
                kernel_img_mul_270[12] + kernel_img_mul_270[13] + kernel_img_mul_270[14] + 
                kernel_img_mul_270[15] + kernel_img_mul_270[16] + kernel_img_mul_270[17] + 
                kernel_img_mul_270[18] + kernel_img_mul_270[19] + kernel_img_mul_270[20] + 
                kernel_img_mul_270[21] + kernel_img_mul_270[22] + kernel_img_mul_270[23] + 
                kernel_img_mul_270[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2167:2160] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2167:2160] <= kernel_img_sum_270[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2167:2160] <= 'd0;
end

wire  [39:0]  kernel_img_mul_271[0:24];
assign kernel_img_mul_271[0] = buffer_data_4[2159:2152] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_271[1] = buffer_data_4[2167:2160] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_271[2] = buffer_data_4[2175:2168] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_271[3] = buffer_data_4[2183:2176] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_271[4] = buffer_data_4[2191:2184] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_271[5] = buffer_data_3[2159:2152] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_271[6] = buffer_data_3[2167:2160] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_271[7] = buffer_data_3[2175:2168] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_271[8] = buffer_data_3[2183:2176] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_271[9] = buffer_data_3[2191:2184] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_271[10] = buffer_data_2[2159:2152] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_271[11] = buffer_data_2[2167:2160] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_271[12] = buffer_data_2[2175:2168] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_271[13] = buffer_data_2[2183:2176] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_271[14] = buffer_data_2[2191:2184] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_271[15] = buffer_data_1[2159:2152] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_271[16] = buffer_data_1[2167:2160] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_271[17] = buffer_data_1[2175:2168] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_271[18] = buffer_data_1[2183:2176] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_271[19] = buffer_data_1[2191:2184] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_271[20] = buffer_data_0[2159:2152] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_271[21] = buffer_data_0[2167:2160] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_271[22] = buffer_data_0[2175:2168] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_271[23] = buffer_data_0[2183:2176] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_271[24] = buffer_data_0[2191:2184] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_271 = kernel_img_mul_271[0] + kernel_img_mul_271[1] + kernel_img_mul_271[2] + 
                kernel_img_mul_271[3] + kernel_img_mul_271[4] + kernel_img_mul_271[5] + 
                kernel_img_mul_271[6] + kernel_img_mul_271[7] + kernel_img_mul_271[8] + 
                kernel_img_mul_271[9] + kernel_img_mul_271[10] + kernel_img_mul_271[11] + 
                kernel_img_mul_271[12] + kernel_img_mul_271[13] + kernel_img_mul_271[14] + 
                kernel_img_mul_271[15] + kernel_img_mul_271[16] + kernel_img_mul_271[17] + 
                kernel_img_mul_271[18] + kernel_img_mul_271[19] + kernel_img_mul_271[20] + 
                kernel_img_mul_271[21] + kernel_img_mul_271[22] + kernel_img_mul_271[23] + 
                kernel_img_mul_271[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2175:2168] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2175:2168] <= kernel_img_sum_271[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2175:2168] <= 'd0;
end

wire  [39:0]  kernel_img_mul_272[0:24];
assign kernel_img_mul_272[0] = buffer_data_4[2167:2160] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_272[1] = buffer_data_4[2175:2168] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_272[2] = buffer_data_4[2183:2176] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_272[3] = buffer_data_4[2191:2184] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_272[4] = buffer_data_4[2199:2192] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_272[5] = buffer_data_3[2167:2160] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_272[6] = buffer_data_3[2175:2168] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_272[7] = buffer_data_3[2183:2176] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_272[8] = buffer_data_3[2191:2184] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_272[9] = buffer_data_3[2199:2192] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_272[10] = buffer_data_2[2167:2160] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_272[11] = buffer_data_2[2175:2168] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_272[12] = buffer_data_2[2183:2176] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_272[13] = buffer_data_2[2191:2184] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_272[14] = buffer_data_2[2199:2192] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_272[15] = buffer_data_1[2167:2160] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_272[16] = buffer_data_1[2175:2168] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_272[17] = buffer_data_1[2183:2176] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_272[18] = buffer_data_1[2191:2184] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_272[19] = buffer_data_1[2199:2192] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_272[20] = buffer_data_0[2167:2160] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_272[21] = buffer_data_0[2175:2168] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_272[22] = buffer_data_0[2183:2176] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_272[23] = buffer_data_0[2191:2184] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_272[24] = buffer_data_0[2199:2192] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_272 = kernel_img_mul_272[0] + kernel_img_mul_272[1] + kernel_img_mul_272[2] + 
                kernel_img_mul_272[3] + kernel_img_mul_272[4] + kernel_img_mul_272[5] + 
                kernel_img_mul_272[6] + kernel_img_mul_272[7] + kernel_img_mul_272[8] + 
                kernel_img_mul_272[9] + kernel_img_mul_272[10] + kernel_img_mul_272[11] + 
                kernel_img_mul_272[12] + kernel_img_mul_272[13] + kernel_img_mul_272[14] + 
                kernel_img_mul_272[15] + kernel_img_mul_272[16] + kernel_img_mul_272[17] + 
                kernel_img_mul_272[18] + kernel_img_mul_272[19] + kernel_img_mul_272[20] + 
                kernel_img_mul_272[21] + kernel_img_mul_272[22] + kernel_img_mul_272[23] + 
                kernel_img_mul_272[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2183:2176] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2183:2176] <= kernel_img_sum_272[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2183:2176] <= 'd0;
end

wire  [39:0]  kernel_img_mul_273[0:24];
assign kernel_img_mul_273[0] = buffer_data_4[2175:2168] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_273[1] = buffer_data_4[2183:2176] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_273[2] = buffer_data_4[2191:2184] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_273[3] = buffer_data_4[2199:2192] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_273[4] = buffer_data_4[2207:2200] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_273[5] = buffer_data_3[2175:2168] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_273[6] = buffer_data_3[2183:2176] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_273[7] = buffer_data_3[2191:2184] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_273[8] = buffer_data_3[2199:2192] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_273[9] = buffer_data_3[2207:2200] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_273[10] = buffer_data_2[2175:2168] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_273[11] = buffer_data_2[2183:2176] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_273[12] = buffer_data_2[2191:2184] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_273[13] = buffer_data_2[2199:2192] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_273[14] = buffer_data_2[2207:2200] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_273[15] = buffer_data_1[2175:2168] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_273[16] = buffer_data_1[2183:2176] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_273[17] = buffer_data_1[2191:2184] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_273[18] = buffer_data_1[2199:2192] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_273[19] = buffer_data_1[2207:2200] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_273[20] = buffer_data_0[2175:2168] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_273[21] = buffer_data_0[2183:2176] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_273[22] = buffer_data_0[2191:2184] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_273[23] = buffer_data_0[2199:2192] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_273[24] = buffer_data_0[2207:2200] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_273 = kernel_img_mul_273[0] + kernel_img_mul_273[1] + kernel_img_mul_273[2] + 
                kernel_img_mul_273[3] + kernel_img_mul_273[4] + kernel_img_mul_273[5] + 
                kernel_img_mul_273[6] + kernel_img_mul_273[7] + kernel_img_mul_273[8] + 
                kernel_img_mul_273[9] + kernel_img_mul_273[10] + kernel_img_mul_273[11] + 
                kernel_img_mul_273[12] + kernel_img_mul_273[13] + kernel_img_mul_273[14] + 
                kernel_img_mul_273[15] + kernel_img_mul_273[16] + kernel_img_mul_273[17] + 
                kernel_img_mul_273[18] + kernel_img_mul_273[19] + kernel_img_mul_273[20] + 
                kernel_img_mul_273[21] + kernel_img_mul_273[22] + kernel_img_mul_273[23] + 
                kernel_img_mul_273[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2191:2184] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2191:2184] <= kernel_img_sum_273[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2191:2184] <= 'd0;
end

wire  [39:0]  kernel_img_mul_274[0:24];
assign kernel_img_mul_274[0] = buffer_data_4[2183:2176] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_274[1] = buffer_data_4[2191:2184] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_274[2] = buffer_data_4[2199:2192] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_274[3] = buffer_data_4[2207:2200] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_274[4] = buffer_data_4[2215:2208] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_274[5] = buffer_data_3[2183:2176] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_274[6] = buffer_data_3[2191:2184] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_274[7] = buffer_data_3[2199:2192] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_274[8] = buffer_data_3[2207:2200] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_274[9] = buffer_data_3[2215:2208] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_274[10] = buffer_data_2[2183:2176] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_274[11] = buffer_data_2[2191:2184] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_274[12] = buffer_data_2[2199:2192] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_274[13] = buffer_data_2[2207:2200] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_274[14] = buffer_data_2[2215:2208] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_274[15] = buffer_data_1[2183:2176] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_274[16] = buffer_data_1[2191:2184] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_274[17] = buffer_data_1[2199:2192] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_274[18] = buffer_data_1[2207:2200] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_274[19] = buffer_data_1[2215:2208] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_274[20] = buffer_data_0[2183:2176] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_274[21] = buffer_data_0[2191:2184] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_274[22] = buffer_data_0[2199:2192] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_274[23] = buffer_data_0[2207:2200] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_274[24] = buffer_data_0[2215:2208] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_274 = kernel_img_mul_274[0] + kernel_img_mul_274[1] + kernel_img_mul_274[2] + 
                kernel_img_mul_274[3] + kernel_img_mul_274[4] + kernel_img_mul_274[5] + 
                kernel_img_mul_274[6] + kernel_img_mul_274[7] + kernel_img_mul_274[8] + 
                kernel_img_mul_274[9] + kernel_img_mul_274[10] + kernel_img_mul_274[11] + 
                kernel_img_mul_274[12] + kernel_img_mul_274[13] + kernel_img_mul_274[14] + 
                kernel_img_mul_274[15] + kernel_img_mul_274[16] + kernel_img_mul_274[17] + 
                kernel_img_mul_274[18] + kernel_img_mul_274[19] + kernel_img_mul_274[20] + 
                kernel_img_mul_274[21] + kernel_img_mul_274[22] + kernel_img_mul_274[23] + 
                kernel_img_mul_274[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2199:2192] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2199:2192] <= kernel_img_sum_274[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2199:2192] <= 'd0;
end

wire  [39:0]  kernel_img_mul_275[0:24];
assign kernel_img_mul_275[0] = buffer_data_4[2191:2184] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_275[1] = buffer_data_4[2199:2192] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_275[2] = buffer_data_4[2207:2200] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_275[3] = buffer_data_4[2215:2208] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_275[4] = buffer_data_4[2223:2216] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_275[5] = buffer_data_3[2191:2184] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_275[6] = buffer_data_3[2199:2192] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_275[7] = buffer_data_3[2207:2200] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_275[8] = buffer_data_3[2215:2208] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_275[9] = buffer_data_3[2223:2216] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_275[10] = buffer_data_2[2191:2184] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_275[11] = buffer_data_2[2199:2192] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_275[12] = buffer_data_2[2207:2200] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_275[13] = buffer_data_2[2215:2208] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_275[14] = buffer_data_2[2223:2216] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_275[15] = buffer_data_1[2191:2184] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_275[16] = buffer_data_1[2199:2192] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_275[17] = buffer_data_1[2207:2200] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_275[18] = buffer_data_1[2215:2208] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_275[19] = buffer_data_1[2223:2216] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_275[20] = buffer_data_0[2191:2184] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_275[21] = buffer_data_0[2199:2192] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_275[22] = buffer_data_0[2207:2200] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_275[23] = buffer_data_0[2215:2208] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_275[24] = buffer_data_0[2223:2216] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_275 = kernel_img_mul_275[0] + kernel_img_mul_275[1] + kernel_img_mul_275[2] + 
                kernel_img_mul_275[3] + kernel_img_mul_275[4] + kernel_img_mul_275[5] + 
                kernel_img_mul_275[6] + kernel_img_mul_275[7] + kernel_img_mul_275[8] + 
                kernel_img_mul_275[9] + kernel_img_mul_275[10] + kernel_img_mul_275[11] + 
                kernel_img_mul_275[12] + kernel_img_mul_275[13] + kernel_img_mul_275[14] + 
                kernel_img_mul_275[15] + kernel_img_mul_275[16] + kernel_img_mul_275[17] + 
                kernel_img_mul_275[18] + kernel_img_mul_275[19] + kernel_img_mul_275[20] + 
                kernel_img_mul_275[21] + kernel_img_mul_275[22] + kernel_img_mul_275[23] + 
                kernel_img_mul_275[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2207:2200] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2207:2200] <= kernel_img_sum_275[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2207:2200] <= 'd0;
end

wire  [39:0]  kernel_img_mul_276[0:24];
assign kernel_img_mul_276[0] = buffer_data_4[2199:2192] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_276[1] = buffer_data_4[2207:2200] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_276[2] = buffer_data_4[2215:2208] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_276[3] = buffer_data_4[2223:2216] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_276[4] = buffer_data_4[2231:2224] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_276[5] = buffer_data_3[2199:2192] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_276[6] = buffer_data_3[2207:2200] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_276[7] = buffer_data_3[2215:2208] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_276[8] = buffer_data_3[2223:2216] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_276[9] = buffer_data_3[2231:2224] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_276[10] = buffer_data_2[2199:2192] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_276[11] = buffer_data_2[2207:2200] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_276[12] = buffer_data_2[2215:2208] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_276[13] = buffer_data_2[2223:2216] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_276[14] = buffer_data_2[2231:2224] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_276[15] = buffer_data_1[2199:2192] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_276[16] = buffer_data_1[2207:2200] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_276[17] = buffer_data_1[2215:2208] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_276[18] = buffer_data_1[2223:2216] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_276[19] = buffer_data_1[2231:2224] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_276[20] = buffer_data_0[2199:2192] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_276[21] = buffer_data_0[2207:2200] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_276[22] = buffer_data_0[2215:2208] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_276[23] = buffer_data_0[2223:2216] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_276[24] = buffer_data_0[2231:2224] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_276 = kernel_img_mul_276[0] + kernel_img_mul_276[1] + kernel_img_mul_276[2] + 
                kernel_img_mul_276[3] + kernel_img_mul_276[4] + kernel_img_mul_276[5] + 
                kernel_img_mul_276[6] + kernel_img_mul_276[7] + kernel_img_mul_276[8] + 
                kernel_img_mul_276[9] + kernel_img_mul_276[10] + kernel_img_mul_276[11] + 
                kernel_img_mul_276[12] + kernel_img_mul_276[13] + kernel_img_mul_276[14] + 
                kernel_img_mul_276[15] + kernel_img_mul_276[16] + kernel_img_mul_276[17] + 
                kernel_img_mul_276[18] + kernel_img_mul_276[19] + kernel_img_mul_276[20] + 
                kernel_img_mul_276[21] + kernel_img_mul_276[22] + kernel_img_mul_276[23] + 
                kernel_img_mul_276[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2215:2208] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2215:2208] <= kernel_img_sum_276[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2215:2208] <= 'd0;
end

wire  [39:0]  kernel_img_mul_277[0:24];
assign kernel_img_mul_277[0] = buffer_data_4[2207:2200] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_277[1] = buffer_data_4[2215:2208] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_277[2] = buffer_data_4[2223:2216] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_277[3] = buffer_data_4[2231:2224] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_277[4] = buffer_data_4[2239:2232] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_277[5] = buffer_data_3[2207:2200] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_277[6] = buffer_data_3[2215:2208] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_277[7] = buffer_data_3[2223:2216] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_277[8] = buffer_data_3[2231:2224] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_277[9] = buffer_data_3[2239:2232] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_277[10] = buffer_data_2[2207:2200] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_277[11] = buffer_data_2[2215:2208] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_277[12] = buffer_data_2[2223:2216] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_277[13] = buffer_data_2[2231:2224] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_277[14] = buffer_data_2[2239:2232] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_277[15] = buffer_data_1[2207:2200] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_277[16] = buffer_data_1[2215:2208] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_277[17] = buffer_data_1[2223:2216] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_277[18] = buffer_data_1[2231:2224] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_277[19] = buffer_data_1[2239:2232] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_277[20] = buffer_data_0[2207:2200] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_277[21] = buffer_data_0[2215:2208] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_277[22] = buffer_data_0[2223:2216] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_277[23] = buffer_data_0[2231:2224] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_277[24] = buffer_data_0[2239:2232] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_277 = kernel_img_mul_277[0] + kernel_img_mul_277[1] + kernel_img_mul_277[2] + 
                kernel_img_mul_277[3] + kernel_img_mul_277[4] + kernel_img_mul_277[5] + 
                kernel_img_mul_277[6] + kernel_img_mul_277[7] + kernel_img_mul_277[8] + 
                kernel_img_mul_277[9] + kernel_img_mul_277[10] + kernel_img_mul_277[11] + 
                kernel_img_mul_277[12] + kernel_img_mul_277[13] + kernel_img_mul_277[14] + 
                kernel_img_mul_277[15] + kernel_img_mul_277[16] + kernel_img_mul_277[17] + 
                kernel_img_mul_277[18] + kernel_img_mul_277[19] + kernel_img_mul_277[20] + 
                kernel_img_mul_277[21] + kernel_img_mul_277[22] + kernel_img_mul_277[23] + 
                kernel_img_mul_277[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2223:2216] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2223:2216] <= kernel_img_sum_277[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2223:2216] <= 'd0;
end

wire  [39:0]  kernel_img_mul_278[0:24];
assign kernel_img_mul_278[0] = buffer_data_4[2215:2208] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_278[1] = buffer_data_4[2223:2216] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_278[2] = buffer_data_4[2231:2224] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_278[3] = buffer_data_4[2239:2232] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_278[4] = buffer_data_4[2247:2240] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_278[5] = buffer_data_3[2215:2208] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_278[6] = buffer_data_3[2223:2216] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_278[7] = buffer_data_3[2231:2224] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_278[8] = buffer_data_3[2239:2232] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_278[9] = buffer_data_3[2247:2240] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_278[10] = buffer_data_2[2215:2208] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_278[11] = buffer_data_2[2223:2216] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_278[12] = buffer_data_2[2231:2224] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_278[13] = buffer_data_2[2239:2232] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_278[14] = buffer_data_2[2247:2240] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_278[15] = buffer_data_1[2215:2208] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_278[16] = buffer_data_1[2223:2216] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_278[17] = buffer_data_1[2231:2224] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_278[18] = buffer_data_1[2239:2232] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_278[19] = buffer_data_1[2247:2240] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_278[20] = buffer_data_0[2215:2208] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_278[21] = buffer_data_0[2223:2216] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_278[22] = buffer_data_0[2231:2224] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_278[23] = buffer_data_0[2239:2232] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_278[24] = buffer_data_0[2247:2240] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_278 = kernel_img_mul_278[0] + kernel_img_mul_278[1] + kernel_img_mul_278[2] + 
                kernel_img_mul_278[3] + kernel_img_mul_278[4] + kernel_img_mul_278[5] + 
                kernel_img_mul_278[6] + kernel_img_mul_278[7] + kernel_img_mul_278[8] + 
                kernel_img_mul_278[9] + kernel_img_mul_278[10] + kernel_img_mul_278[11] + 
                kernel_img_mul_278[12] + kernel_img_mul_278[13] + kernel_img_mul_278[14] + 
                kernel_img_mul_278[15] + kernel_img_mul_278[16] + kernel_img_mul_278[17] + 
                kernel_img_mul_278[18] + kernel_img_mul_278[19] + kernel_img_mul_278[20] + 
                kernel_img_mul_278[21] + kernel_img_mul_278[22] + kernel_img_mul_278[23] + 
                kernel_img_mul_278[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2231:2224] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2231:2224] <= kernel_img_sum_278[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2231:2224] <= 'd0;
end

wire  [39:0]  kernel_img_mul_279[0:24];
assign kernel_img_mul_279[0] = buffer_data_4[2223:2216] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_279[1] = buffer_data_4[2231:2224] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_279[2] = buffer_data_4[2239:2232] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_279[3] = buffer_data_4[2247:2240] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_279[4] = buffer_data_4[2255:2248] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_279[5] = buffer_data_3[2223:2216] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_279[6] = buffer_data_3[2231:2224] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_279[7] = buffer_data_3[2239:2232] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_279[8] = buffer_data_3[2247:2240] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_279[9] = buffer_data_3[2255:2248] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_279[10] = buffer_data_2[2223:2216] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_279[11] = buffer_data_2[2231:2224] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_279[12] = buffer_data_2[2239:2232] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_279[13] = buffer_data_2[2247:2240] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_279[14] = buffer_data_2[2255:2248] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_279[15] = buffer_data_1[2223:2216] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_279[16] = buffer_data_1[2231:2224] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_279[17] = buffer_data_1[2239:2232] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_279[18] = buffer_data_1[2247:2240] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_279[19] = buffer_data_1[2255:2248] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_279[20] = buffer_data_0[2223:2216] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_279[21] = buffer_data_0[2231:2224] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_279[22] = buffer_data_0[2239:2232] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_279[23] = buffer_data_0[2247:2240] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_279[24] = buffer_data_0[2255:2248] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_279 = kernel_img_mul_279[0] + kernel_img_mul_279[1] + kernel_img_mul_279[2] + 
                kernel_img_mul_279[3] + kernel_img_mul_279[4] + kernel_img_mul_279[5] + 
                kernel_img_mul_279[6] + kernel_img_mul_279[7] + kernel_img_mul_279[8] + 
                kernel_img_mul_279[9] + kernel_img_mul_279[10] + kernel_img_mul_279[11] + 
                kernel_img_mul_279[12] + kernel_img_mul_279[13] + kernel_img_mul_279[14] + 
                kernel_img_mul_279[15] + kernel_img_mul_279[16] + kernel_img_mul_279[17] + 
                kernel_img_mul_279[18] + kernel_img_mul_279[19] + kernel_img_mul_279[20] + 
                kernel_img_mul_279[21] + kernel_img_mul_279[22] + kernel_img_mul_279[23] + 
                kernel_img_mul_279[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2239:2232] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2239:2232] <= kernel_img_sum_279[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2239:2232] <= 'd0;
end

wire  [39:0]  kernel_img_mul_280[0:24];
assign kernel_img_mul_280[0] = buffer_data_4[2231:2224] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_280[1] = buffer_data_4[2239:2232] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_280[2] = buffer_data_4[2247:2240] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_280[3] = buffer_data_4[2255:2248] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_280[4] = buffer_data_4[2263:2256] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_280[5] = buffer_data_3[2231:2224] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_280[6] = buffer_data_3[2239:2232] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_280[7] = buffer_data_3[2247:2240] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_280[8] = buffer_data_3[2255:2248] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_280[9] = buffer_data_3[2263:2256] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_280[10] = buffer_data_2[2231:2224] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_280[11] = buffer_data_2[2239:2232] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_280[12] = buffer_data_2[2247:2240] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_280[13] = buffer_data_2[2255:2248] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_280[14] = buffer_data_2[2263:2256] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_280[15] = buffer_data_1[2231:2224] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_280[16] = buffer_data_1[2239:2232] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_280[17] = buffer_data_1[2247:2240] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_280[18] = buffer_data_1[2255:2248] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_280[19] = buffer_data_1[2263:2256] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_280[20] = buffer_data_0[2231:2224] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_280[21] = buffer_data_0[2239:2232] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_280[22] = buffer_data_0[2247:2240] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_280[23] = buffer_data_0[2255:2248] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_280[24] = buffer_data_0[2263:2256] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_280 = kernel_img_mul_280[0] + kernel_img_mul_280[1] + kernel_img_mul_280[2] + 
                kernel_img_mul_280[3] + kernel_img_mul_280[4] + kernel_img_mul_280[5] + 
                kernel_img_mul_280[6] + kernel_img_mul_280[7] + kernel_img_mul_280[8] + 
                kernel_img_mul_280[9] + kernel_img_mul_280[10] + kernel_img_mul_280[11] + 
                kernel_img_mul_280[12] + kernel_img_mul_280[13] + kernel_img_mul_280[14] + 
                kernel_img_mul_280[15] + kernel_img_mul_280[16] + kernel_img_mul_280[17] + 
                kernel_img_mul_280[18] + kernel_img_mul_280[19] + kernel_img_mul_280[20] + 
                kernel_img_mul_280[21] + kernel_img_mul_280[22] + kernel_img_mul_280[23] + 
                kernel_img_mul_280[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2247:2240] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2247:2240] <= kernel_img_sum_280[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2247:2240] <= 'd0;
end

wire  [39:0]  kernel_img_mul_281[0:24];
assign kernel_img_mul_281[0] = buffer_data_4[2239:2232] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_281[1] = buffer_data_4[2247:2240] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_281[2] = buffer_data_4[2255:2248] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_281[3] = buffer_data_4[2263:2256] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_281[4] = buffer_data_4[2271:2264] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_281[5] = buffer_data_3[2239:2232] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_281[6] = buffer_data_3[2247:2240] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_281[7] = buffer_data_3[2255:2248] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_281[8] = buffer_data_3[2263:2256] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_281[9] = buffer_data_3[2271:2264] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_281[10] = buffer_data_2[2239:2232] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_281[11] = buffer_data_2[2247:2240] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_281[12] = buffer_data_2[2255:2248] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_281[13] = buffer_data_2[2263:2256] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_281[14] = buffer_data_2[2271:2264] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_281[15] = buffer_data_1[2239:2232] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_281[16] = buffer_data_1[2247:2240] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_281[17] = buffer_data_1[2255:2248] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_281[18] = buffer_data_1[2263:2256] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_281[19] = buffer_data_1[2271:2264] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_281[20] = buffer_data_0[2239:2232] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_281[21] = buffer_data_0[2247:2240] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_281[22] = buffer_data_0[2255:2248] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_281[23] = buffer_data_0[2263:2256] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_281[24] = buffer_data_0[2271:2264] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_281 = kernel_img_mul_281[0] + kernel_img_mul_281[1] + kernel_img_mul_281[2] + 
                kernel_img_mul_281[3] + kernel_img_mul_281[4] + kernel_img_mul_281[5] + 
                kernel_img_mul_281[6] + kernel_img_mul_281[7] + kernel_img_mul_281[8] + 
                kernel_img_mul_281[9] + kernel_img_mul_281[10] + kernel_img_mul_281[11] + 
                kernel_img_mul_281[12] + kernel_img_mul_281[13] + kernel_img_mul_281[14] + 
                kernel_img_mul_281[15] + kernel_img_mul_281[16] + kernel_img_mul_281[17] + 
                kernel_img_mul_281[18] + kernel_img_mul_281[19] + kernel_img_mul_281[20] + 
                kernel_img_mul_281[21] + kernel_img_mul_281[22] + kernel_img_mul_281[23] + 
                kernel_img_mul_281[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2255:2248] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2255:2248] <= kernel_img_sum_281[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2255:2248] <= 'd0;
end

wire  [39:0]  kernel_img_mul_282[0:24];
assign kernel_img_mul_282[0] = buffer_data_4[2247:2240] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_282[1] = buffer_data_4[2255:2248] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_282[2] = buffer_data_4[2263:2256] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_282[3] = buffer_data_4[2271:2264] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_282[4] = buffer_data_4[2279:2272] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_282[5] = buffer_data_3[2247:2240] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_282[6] = buffer_data_3[2255:2248] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_282[7] = buffer_data_3[2263:2256] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_282[8] = buffer_data_3[2271:2264] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_282[9] = buffer_data_3[2279:2272] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_282[10] = buffer_data_2[2247:2240] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_282[11] = buffer_data_2[2255:2248] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_282[12] = buffer_data_2[2263:2256] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_282[13] = buffer_data_2[2271:2264] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_282[14] = buffer_data_2[2279:2272] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_282[15] = buffer_data_1[2247:2240] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_282[16] = buffer_data_1[2255:2248] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_282[17] = buffer_data_1[2263:2256] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_282[18] = buffer_data_1[2271:2264] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_282[19] = buffer_data_1[2279:2272] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_282[20] = buffer_data_0[2247:2240] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_282[21] = buffer_data_0[2255:2248] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_282[22] = buffer_data_0[2263:2256] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_282[23] = buffer_data_0[2271:2264] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_282[24] = buffer_data_0[2279:2272] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_282 = kernel_img_mul_282[0] + kernel_img_mul_282[1] + kernel_img_mul_282[2] + 
                kernel_img_mul_282[3] + kernel_img_mul_282[4] + kernel_img_mul_282[5] + 
                kernel_img_mul_282[6] + kernel_img_mul_282[7] + kernel_img_mul_282[8] + 
                kernel_img_mul_282[9] + kernel_img_mul_282[10] + kernel_img_mul_282[11] + 
                kernel_img_mul_282[12] + kernel_img_mul_282[13] + kernel_img_mul_282[14] + 
                kernel_img_mul_282[15] + kernel_img_mul_282[16] + kernel_img_mul_282[17] + 
                kernel_img_mul_282[18] + kernel_img_mul_282[19] + kernel_img_mul_282[20] + 
                kernel_img_mul_282[21] + kernel_img_mul_282[22] + kernel_img_mul_282[23] + 
                kernel_img_mul_282[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2263:2256] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2263:2256] <= kernel_img_sum_282[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2263:2256] <= 'd0;
end

wire  [39:0]  kernel_img_mul_283[0:24];
assign kernel_img_mul_283[0] = buffer_data_4[2255:2248] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_283[1] = buffer_data_4[2263:2256] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_283[2] = buffer_data_4[2271:2264] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_283[3] = buffer_data_4[2279:2272] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_283[4] = buffer_data_4[2287:2280] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_283[5] = buffer_data_3[2255:2248] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_283[6] = buffer_data_3[2263:2256] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_283[7] = buffer_data_3[2271:2264] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_283[8] = buffer_data_3[2279:2272] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_283[9] = buffer_data_3[2287:2280] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_283[10] = buffer_data_2[2255:2248] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_283[11] = buffer_data_2[2263:2256] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_283[12] = buffer_data_2[2271:2264] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_283[13] = buffer_data_2[2279:2272] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_283[14] = buffer_data_2[2287:2280] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_283[15] = buffer_data_1[2255:2248] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_283[16] = buffer_data_1[2263:2256] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_283[17] = buffer_data_1[2271:2264] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_283[18] = buffer_data_1[2279:2272] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_283[19] = buffer_data_1[2287:2280] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_283[20] = buffer_data_0[2255:2248] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_283[21] = buffer_data_0[2263:2256] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_283[22] = buffer_data_0[2271:2264] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_283[23] = buffer_data_0[2279:2272] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_283[24] = buffer_data_0[2287:2280] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_283 = kernel_img_mul_283[0] + kernel_img_mul_283[1] + kernel_img_mul_283[2] + 
                kernel_img_mul_283[3] + kernel_img_mul_283[4] + kernel_img_mul_283[5] + 
                kernel_img_mul_283[6] + kernel_img_mul_283[7] + kernel_img_mul_283[8] + 
                kernel_img_mul_283[9] + kernel_img_mul_283[10] + kernel_img_mul_283[11] + 
                kernel_img_mul_283[12] + kernel_img_mul_283[13] + kernel_img_mul_283[14] + 
                kernel_img_mul_283[15] + kernel_img_mul_283[16] + kernel_img_mul_283[17] + 
                kernel_img_mul_283[18] + kernel_img_mul_283[19] + kernel_img_mul_283[20] + 
                kernel_img_mul_283[21] + kernel_img_mul_283[22] + kernel_img_mul_283[23] + 
                kernel_img_mul_283[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2271:2264] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2271:2264] <= kernel_img_sum_283[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2271:2264] <= 'd0;
end

wire  [39:0]  kernel_img_mul_284[0:24];
assign kernel_img_mul_284[0] = buffer_data_4[2263:2256] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_284[1] = buffer_data_4[2271:2264] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_284[2] = buffer_data_4[2279:2272] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_284[3] = buffer_data_4[2287:2280] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_284[4] = buffer_data_4[2295:2288] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_284[5] = buffer_data_3[2263:2256] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_284[6] = buffer_data_3[2271:2264] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_284[7] = buffer_data_3[2279:2272] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_284[8] = buffer_data_3[2287:2280] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_284[9] = buffer_data_3[2295:2288] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_284[10] = buffer_data_2[2263:2256] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_284[11] = buffer_data_2[2271:2264] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_284[12] = buffer_data_2[2279:2272] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_284[13] = buffer_data_2[2287:2280] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_284[14] = buffer_data_2[2295:2288] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_284[15] = buffer_data_1[2263:2256] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_284[16] = buffer_data_1[2271:2264] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_284[17] = buffer_data_1[2279:2272] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_284[18] = buffer_data_1[2287:2280] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_284[19] = buffer_data_1[2295:2288] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_284[20] = buffer_data_0[2263:2256] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_284[21] = buffer_data_0[2271:2264] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_284[22] = buffer_data_0[2279:2272] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_284[23] = buffer_data_0[2287:2280] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_284[24] = buffer_data_0[2295:2288] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_284 = kernel_img_mul_284[0] + kernel_img_mul_284[1] + kernel_img_mul_284[2] + 
                kernel_img_mul_284[3] + kernel_img_mul_284[4] + kernel_img_mul_284[5] + 
                kernel_img_mul_284[6] + kernel_img_mul_284[7] + kernel_img_mul_284[8] + 
                kernel_img_mul_284[9] + kernel_img_mul_284[10] + kernel_img_mul_284[11] + 
                kernel_img_mul_284[12] + kernel_img_mul_284[13] + kernel_img_mul_284[14] + 
                kernel_img_mul_284[15] + kernel_img_mul_284[16] + kernel_img_mul_284[17] + 
                kernel_img_mul_284[18] + kernel_img_mul_284[19] + kernel_img_mul_284[20] + 
                kernel_img_mul_284[21] + kernel_img_mul_284[22] + kernel_img_mul_284[23] + 
                kernel_img_mul_284[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2279:2272] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2279:2272] <= kernel_img_sum_284[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2279:2272] <= 'd0;
end

wire  [39:0]  kernel_img_mul_285[0:24];
assign kernel_img_mul_285[0] = buffer_data_4[2271:2264] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_285[1] = buffer_data_4[2279:2272] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_285[2] = buffer_data_4[2287:2280] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_285[3] = buffer_data_4[2295:2288] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_285[4] = buffer_data_4[2303:2296] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_285[5] = buffer_data_3[2271:2264] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_285[6] = buffer_data_3[2279:2272] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_285[7] = buffer_data_3[2287:2280] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_285[8] = buffer_data_3[2295:2288] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_285[9] = buffer_data_3[2303:2296] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_285[10] = buffer_data_2[2271:2264] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_285[11] = buffer_data_2[2279:2272] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_285[12] = buffer_data_2[2287:2280] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_285[13] = buffer_data_2[2295:2288] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_285[14] = buffer_data_2[2303:2296] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_285[15] = buffer_data_1[2271:2264] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_285[16] = buffer_data_1[2279:2272] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_285[17] = buffer_data_1[2287:2280] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_285[18] = buffer_data_1[2295:2288] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_285[19] = buffer_data_1[2303:2296] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_285[20] = buffer_data_0[2271:2264] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_285[21] = buffer_data_0[2279:2272] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_285[22] = buffer_data_0[2287:2280] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_285[23] = buffer_data_0[2295:2288] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_285[24] = buffer_data_0[2303:2296] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_285 = kernel_img_mul_285[0] + kernel_img_mul_285[1] + kernel_img_mul_285[2] + 
                kernel_img_mul_285[3] + kernel_img_mul_285[4] + kernel_img_mul_285[5] + 
                kernel_img_mul_285[6] + kernel_img_mul_285[7] + kernel_img_mul_285[8] + 
                kernel_img_mul_285[9] + kernel_img_mul_285[10] + kernel_img_mul_285[11] + 
                kernel_img_mul_285[12] + kernel_img_mul_285[13] + kernel_img_mul_285[14] + 
                kernel_img_mul_285[15] + kernel_img_mul_285[16] + kernel_img_mul_285[17] + 
                kernel_img_mul_285[18] + kernel_img_mul_285[19] + kernel_img_mul_285[20] + 
                kernel_img_mul_285[21] + kernel_img_mul_285[22] + kernel_img_mul_285[23] + 
                kernel_img_mul_285[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2287:2280] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2287:2280] <= kernel_img_sum_285[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2287:2280] <= 'd0;
end

wire  [39:0]  kernel_img_mul_286[0:24];
assign kernel_img_mul_286[0] = buffer_data_4[2279:2272] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_286[1] = buffer_data_4[2287:2280] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_286[2] = buffer_data_4[2295:2288] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_286[3] = buffer_data_4[2303:2296] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_286[4] = buffer_data_4[2311:2304] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_286[5] = buffer_data_3[2279:2272] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_286[6] = buffer_data_3[2287:2280] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_286[7] = buffer_data_3[2295:2288] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_286[8] = buffer_data_3[2303:2296] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_286[9] = buffer_data_3[2311:2304] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_286[10] = buffer_data_2[2279:2272] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_286[11] = buffer_data_2[2287:2280] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_286[12] = buffer_data_2[2295:2288] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_286[13] = buffer_data_2[2303:2296] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_286[14] = buffer_data_2[2311:2304] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_286[15] = buffer_data_1[2279:2272] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_286[16] = buffer_data_1[2287:2280] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_286[17] = buffer_data_1[2295:2288] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_286[18] = buffer_data_1[2303:2296] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_286[19] = buffer_data_1[2311:2304] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_286[20] = buffer_data_0[2279:2272] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_286[21] = buffer_data_0[2287:2280] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_286[22] = buffer_data_0[2295:2288] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_286[23] = buffer_data_0[2303:2296] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_286[24] = buffer_data_0[2311:2304] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_286 = kernel_img_mul_286[0] + kernel_img_mul_286[1] + kernel_img_mul_286[2] + 
                kernel_img_mul_286[3] + kernel_img_mul_286[4] + kernel_img_mul_286[5] + 
                kernel_img_mul_286[6] + kernel_img_mul_286[7] + kernel_img_mul_286[8] + 
                kernel_img_mul_286[9] + kernel_img_mul_286[10] + kernel_img_mul_286[11] + 
                kernel_img_mul_286[12] + kernel_img_mul_286[13] + kernel_img_mul_286[14] + 
                kernel_img_mul_286[15] + kernel_img_mul_286[16] + kernel_img_mul_286[17] + 
                kernel_img_mul_286[18] + kernel_img_mul_286[19] + kernel_img_mul_286[20] + 
                kernel_img_mul_286[21] + kernel_img_mul_286[22] + kernel_img_mul_286[23] + 
                kernel_img_mul_286[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2295:2288] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2295:2288] <= kernel_img_sum_286[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2295:2288] <= 'd0;
end

wire  [39:0]  kernel_img_mul_287[0:24];
assign kernel_img_mul_287[0] = buffer_data_4[2287:2280] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_287[1] = buffer_data_4[2295:2288] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_287[2] = buffer_data_4[2303:2296] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_287[3] = buffer_data_4[2311:2304] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_287[4] = buffer_data_4[2319:2312] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_287[5] = buffer_data_3[2287:2280] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_287[6] = buffer_data_3[2295:2288] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_287[7] = buffer_data_3[2303:2296] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_287[8] = buffer_data_3[2311:2304] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_287[9] = buffer_data_3[2319:2312] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_287[10] = buffer_data_2[2287:2280] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_287[11] = buffer_data_2[2295:2288] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_287[12] = buffer_data_2[2303:2296] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_287[13] = buffer_data_2[2311:2304] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_287[14] = buffer_data_2[2319:2312] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_287[15] = buffer_data_1[2287:2280] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_287[16] = buffer_data_1[2295:2288] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_287[17] = buffer_data_1[2303:2296] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_287[18] = buffer_data_1[2311:2304] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_287[19] = buffer_data_1[2319:2312] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_287[20] = buffer_data_0[2287:2280] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_287[21] = buffer_data_0[2295:2288] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_287[22] = buffer_data_0[2303:2296] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_287[23] = buffer_data_0[2311:2304] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_287[24] = buffer_data_0[2319:2312] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_287 = kernel_img_mul_287[0] + kernel_img_mul_287[1] + kernel_img_mul_287[2] + 
                kernel_img_mul_287[3] + kernel_img_mul_287[4] + kernel_img_mul_287[5] + 
                kernel_img_mul_287[6] + kernel_img_mul_287[7] + kernel_img_mul_287[8] + 
                kernel_img_mul_287[9] + kernel_img_mul_287[10] + kernel_img_mul_287[11] + 
                kernel_img_mul_287[12] + kernel_img_mul_287[13] + kernel_img_mul_287[14] + 
                kernel_img_mul_287[15] + kernel_img_mul_287[16] + kernel_img_mul_287[17] + 
                kernel_img_mul_287[18] + kernel_img_mul_287[19] + kernel_img_mul_287[20] + 
                kernel_img_mul_287[21] + kernel_img_mul_287[22] + kernel_img_mul_287[23] + 
                kernel_img_mul_287[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2303:2296] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2303:2296] <= kernel_img_sum_287[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2303:2296] <= 'd0;
end

wire  [39:0]  kernel_img_mul_288[0:24];
assign kernel_img_mul_288[0] = buffer_data_4[2295:2288] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_288[1] = buffer_data_4[2303:2296] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_288[2] = buffer_data_4[2311:2304] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_288[3] = buffer_data_4[2319:2312] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_288[4] = buffer_data_4[2327:2320] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_288[5] = buffer_data_3[2295:2288] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_288[6] = buffer_data_3[2303:2296] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_288[7] = buffer_data_3[2311:2304] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_288[8] = buffer_data_3[2319:2312] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_288[9] = buffer_data_3[2327:2320] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_288[10] = buffer_data_2[2295:2288] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_288[11] = buffer_data_2[2303:2296] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_288[12] = buffer_data_2[2311:2304] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_288[13] = buffer_data_2[2319:2312] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_288[14] = buffer_data_2[2327:2320] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_288[15] = buffer_data_1[2295:2288] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_288[16] = buffer_data_1[2303:2296] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_288[17] = buffer_data_1[2311:2304] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_288[18] = buffer_data_1[2319:2312] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_288[19] = buffer_data_1[2327:2320] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_288[20] = buffer_data_0[2295:2288] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_288[21] = buffer_data_0[2303:2296] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_288[22] = buffer_data_0[2311:2304] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_288[23] = buffer_data_0[2319:2312] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_288[24] = buffer_data_0[2327:2320] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_288 = kernel_img_mul_288[0] + kernel_img_mul_288[1] + kernel_img_mul_288[2] + 
                kernel_img_mul_288[3] + kernel_img_mul_288[4] + kernel_img_mul_288[5] + 
                kernel_img_mul_288[6] + kernel_img_mul_288[7] + kernel_img_mul_288[8] + 
                kernel_img_mul_288[9] + kernel_img_mul_288[10] + kernel_img_mul_288[11] + 
                kernel_img_mul_288[12] + kernel_img_mul_288[13] + kernel_img_mul_288[14] + 
                kernel_img_mul_288[15] + kernel_img_mul_288[16] + kernel_img_mul_288[17] + 
                kernel_img_mul_288[18] + kernel_img_mul_288[19] + kernel_img_mul_288[20] + 
                kernel_img_mul_288[21] + kernel_img_mul_288[22] + kernel_img_mul_288[23] + 
                kernel_img_mul_288[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2311:2304] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2311:2304] <= kernel_img_sum_288[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2311:2304] <= 'd0;
end

wire  [39:0]  kernel_img_mul_289[0:24];
assign kernel_img_mul_289[0] = buffer_data_4[2303:2296] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_289[1] = buffer_data_4[2311:2304] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_289[2] = buffer_data_4[2319:2312] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_289[3] = buffer_data_4[2327:2320] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_289[4] = buffer_data_4[2335:2328] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_289[5] = buffer_data_3[2303:2296] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_289[6] = buffer_data_3[2311:2304] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_289[7] = buffer_data_3[2319:2312] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_289[8] = buffer_data_3[2327:2320] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_289[9] = buffer_data_3[2335:2328] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_289[10] = buffer_data_2[2303:2296] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_289[11] = buffer_data_2[2311:2304] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_289[12] = buffer_data_2[2319:2312] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_289[13] = buffer_data_2[2327:2320] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_289[14] = buffer_data_2[2335:2328] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_289[15] = buffer_data_1[2303:2296] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_289[16] = buffer_data_1[2311:2304] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_289[17] = buffer_data_1[2319:2312] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_289[18] = buffer_data_1[2327:2320] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_289[19] = buffer_data_1[2335:2328] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_289[20] = buffer_data_0[2303:2296] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_289[21] = buffer_data_0[2311:2304] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_289[22] = buffer_data_0[2319:2312] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_289[23] = buffer_data_0[2327:2320] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_289[24] = buffer_data_0[2335:2328] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_289 = kernel_img_mul_289[0] + kernel_img_mul_289[1] + kernel_img_mul_289[2] + 
                kernel_img_mul_289[3] + kernel_img_mul_289[4] + kernel_img_mul_289[5] + 
                kernel_img_mul_289[6] + kernel_img_mul_289[7] + kernel_img_mul_289[8] + 
                kernel_img_mul_289[9] + kernel_img_mul_289[10] + kernel_img_mul_289[11] + 
                kernel_img_mul_289[12] + kernel_img_mul_289[13] + kernel_img_mul_289[14] + 
                kernel_img_mul_289[15] + kernel_img_mul_289[16] + kernel_img_mul_289[17] + 
                kernel_img_mul_289[18] + kernel_img_mul_289[19] + kernel_img_mul_289[20] + 
                kernel_img_mul_289[21] + kernel_img_mul_289[22] + kernel_img_mul_289[23] + 
                kernel_img_mul_289[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2319:2312] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2319:2312] <= kernel_img_sum_289[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2319:2312] <= 'd0;
end

wire  [39:0]  kernel_img_mul_290[0:24];
assign kernel_img_mul_290[0] = buffer_data_4[2311:2304] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_290[1] = buffer_data_4[2319:2312] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_290[2] = buffer_data_4[2327:2320] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_290[3] = buffer_data_4[2335:2328] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_290[4] = buffer_data_4[2343:2336] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_290[5] = buffer_data_3[2311:2304] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_290[6] = buffer_data_3[2319:2312] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_290[7] = buffer_data_3[2327:2320] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_290[8] = buffer_data_3[2335:2328] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_290[9] = buffer_data_3[2343:2336] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_290[10] = buffer_data_2[2311:2304] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_290[11] = buffer_data_2[2319:2312] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_290[12] = buffer_data_2[2327:2320] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_290[13] = buffer_data_2[2335:2328] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_290[14] = buffer_data_2[2343:2336] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_290[15] = buffer_data_1[2311:2304] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_290[16] = buffer_data_1[2319:2312] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_290[17] = buffer_data_1[2327:2320] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_290[18] = buffer_data_1[2335:2328] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_290[19] = buffer_data_1[2343:2336] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_290[20] = buffer_data_0[2311:2304] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_290[21] = buffer_data_0[2319:2312] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_290[22] = buffer_data_0[2327:2320] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_290[23] = buffer_data_0[2335:2328] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_290[24] = buffer_data_0[2343:2336] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_290 = kernel_img_mul_290[0] + kernel_img_mul_290[1] + kernel_img_mul_290[2] + 
                kernel_img_mul_290[3] + kernel_img_mul_290[4] + kernel_img_mul_290[5] + 
                kernel_img_mul_290[6] + kernel_img_mul_290[7] + kernel_img_mul_290[8] + 
                kernel_img_mul_290[9] + kernel_img_mul_290[10] + kernel_img_mul_290[11] + 
                kernel_img_mul_290[12] + kernel_img_mul_290[13] + kernel_img_mul_290[14] + 
                kernel_img_mul_290[15] + kernel_img_mul_290[16] + kernel_img_mul_290[17] + 
                kernel_img_mul_290[18] + kernel_img_mul_290[19] + kernel_img_mul_290[20] + 
                kernel_img_mul_290[21] + kernel_img_mul_290[22] + kernel_img_mul_290[23] + 
                kernel_img_mul_290[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2327:2320] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2327:2320] <= kernel_img_sum_290[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2327:2320] <= 'd0;
end

wire  [39:0]  kernel_img_mul_291[0:24];
assign kernel_img_mul_291[0] = buffer_data_4[2319:2312] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_291[1] = buffer_data_4[2327:2320] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_291[2] = buffer_data_4[2335:2328] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_291[3] = buffer_data_4[2343:2336] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_291[4] = buffer_data_4[2351:2344] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_291[5] = buffer_data_3[2319:2312] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_291[6] = buffer_data_3[2327:2320] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_291[7] = buffer_data_3[2335:2328] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_291[8] = buffer_data_3[2343:2336] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_291[9] = buffer_data_3[2351:2344] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_291[10] = buffer_data_2[2319:2312] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_291[11] = buffer_data_2[2327:2320] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_291[12] = buffer_data_2[2335:2328] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_291[13] = buffer_data_2[2343:2336] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_291[14] = buffer_data_2[2351:2344] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_291[15] = buffer_data_1[2319:2312] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_291[16] = buffer_data_1[2327:2320] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_291[17] = buffer_data_1[2335:2328] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_291[18] = buffer_data_1[2343:2336] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_291[19] = buffer_data_1[2351:2344] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_291[20] = buffer_data_0[2319:2312] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_291[21] = buffer_data_0[2327:2320] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_291[22] = buffer_data_0[2335:2328] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_291[23] = buffer_data_0[2343:2336] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_291[24] = buffer_data_0[2351:2344] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_291 = kernel_img_mul_291[0] + kernel_img_mul_291[1] + kernel_img_mul_291[2] + 
                kernel_img_mul_291[3] + kernel_img_mul_291[4] + kernel_img_mul_291[5] + 
                kernel_img_mul_291[6] + kernel_img_mul_291[7] + kernel_img_mul_291[8] + 
                kernel_img_mul_291[9] + kernel_img_mul_291[10] + kernel_img_mul_291[11] + 
                kernel_img_mul_291[12] + kernel_img_mul_291[13] + kernel_img_mul_291[14] + 
                kernel_img_mul_291[15] + kernel_img_mul_291[16] + kernel_img_mul_291[17] + 
                kernel_img_mul_291[18] + kernel_img_mul_291[19] + kernel_img_mul_291[20] + 
                kernel_img_mul_291[21] + kernel_img_mul_291[22] + kernel_img_mul_291[23] + 
                kernel_img_mul_291[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2335:2328] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2335:2328] <= kernel_img_sum_291[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2335:2328] <= 'd0;
end

wire  [39:0]  kernel_img_mul_292[0:24];
assign kernel_img_mul_292[0] = buffer_data_4[2327:2320] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_292[1] = buffer_data_4[2335:2328] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_292[2] = buffer_data_4[2343:2336] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_292[3] = buffer_data_4[2351:2344] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_292[4] = buffer_data_4[2359:2352] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_292[5] = buffer_data_3[2327:2320] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_292[6] = buffer_data_3[2335:2328] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_292[7] = buffer_data_3[2343:2336] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_292[8] = buffer_data_3[2351:2344] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_292[9] = buffer_data_3[2359:2352] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_292[10] = buffer_data_2[2327:2320] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_292[11] = buffer_data_2[2335:2328] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_292[12] = buffer_data_2[2343:2336] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_292[13] = buffer_data_2[2351:2344] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_292[14] = buffer_data_2[2359:2352] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_292[15] = buffer_data_1[2327:2320] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_292[16] = buffer_data_1[2335:2328] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_292[17] = buffer_data_1[2343:2336] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_292[18] = buffer_data_1[2351:2344] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_292[19] = buffer_data_1[2359:2352] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_292[20] = buffer_data_0[2327:2320] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_292[21] = buffer_data_0[2335:2328] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_292[22] = buffer_data_0[2343:2336] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_292[23] = buffer_data_0[2351:2344] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_292[24] = buffer_data_0[2359:2352] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_292 = kernel_img_mul_292[0] + kernel_img_mul_292[1] + kernel_img_mul_292[2] + 
                kernel_img_mul_292[3] + kernel_img_mul_292[4] + kernel_img_mul_292[5] + 
                kernel_img_mul_292[6] + kernel_img_mul_292[7] + kernel_img_mul_292[8] + 
                kernel_img_mul_292[9] + kernel_img_mul_292[10] + kernel_img_mul_292[11] + 
                kernel_img_mul_292[12] + kernel_img_mul_292[13] + kernel_img_mul_292[14] + 
                kernel_img_mul_292[15] + kernel_img_mul_292[16] + kernel_img_mul_292[17] + 
                kernel_img_mul_292[18] + kernel_img_mul_292[19] + kernel_img_mul_292[20] + 
                kernel_img_mul_292[21] + kernel_img_mul_292[22] + kernel_img_mul_292[23] + 
                kernel_img_mul_292[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2343:2336] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2343:2336] <= kernel_img_sum_292[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2343:2336] <= 'd0;
end

wire  [39:0]  kernel_img_mul_293[0:24];
assign kernel_img_mul_293[0] = buffer_data_4[2335:2328] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_293[1] = buffer_data_4[2343:2336] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_293[2] = buffer_data_4[2351:2344] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_293[3] = buffer_data_4[2359:2352] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_293[4] = buffer_data_4[2367:2360] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_293[5] = buffer_data_3[2335:2328] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_293[6] = buffer_data_3[2343:2336] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_293[7] = buffer_data_3[2351:2344] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_293[8] = buffer_data_3[2359:2352] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_293[9] = buffer_data_3[2367:2360] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_293[10] = buffer_data_2[2335:2328] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_293[11] = buffer_data_2[2343:2336] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_293[12] = buffer_data_2[2351:2344] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_293[13] = buffer_data_2[2359:2352] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_293[14] = buffer_data_2[2367:2360] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_293[15] = buffer_data_1[2335:2328] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_293[16] = buffer_data_1[2343:2336] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_293[17] = buffer_data_1[2351:2344] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_293[18] = buffer_data_1[2359:2352] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_293[19] = buffer_data_1[2367:2360] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_293[20] = buffer_data_0[2335:2328] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_293[21] = buffer_data_0[2343:2336] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_293[22] = buffer_data_0[2351:2344] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_293[23] = buffer_data_0[2359:2352] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_293[24] = buffer_data_0[2367:2360] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_293 = kernel_img_mul_293[0] + kernel_img_mul_293[1] + kernel_img_mul_293[2] + 
                kernel_img_mul_293[3] + kernel_img_mul_293[4] + kernel_img_mul_293[5] + 
                kernel_img_mul_293[6] + kernel_img_mul_293[7] + kernel_img_mul_293[8] + 
                kernel_img_mul_293[9] + kernel_img_mul_293[10] + kernel_img_mul_293[11] + 
                kernel_img_mul_293[12] + kernel_img_mul_293[13] + kernel_img_mul_293[14] + 
                kernel_img_mul_293[15] + kernel_img_mul_293[16] + kernel_img_mul_293[17] + 
                kernel_img_mul_293[18] + kernel_img_mul_293[19] + kernel_img_mul_293[20] + 
                kernel_img_mul_293[21] + kernel_img_mul_293[22] + kernel_img_mul_293[23] + 
                kernel_img_mul_293[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2351:2344] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2351:2344] <= kernel_img_sum_293[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2351:2344] <= 'd0;
end

wire  [39:0]  kernel_img_mul_294[0:24];
assign kernel_img_mul_294[0] = buffer_data_4[2343:2336] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_294[1] = buffer_data_4[2351:2344] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_294[2] = buffer_data_4[2359:2352] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_294[3] = buffer_data_4[2367:2360] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_294[4] = buffer_data_4[2375:2368] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_294[5] = buffer_data_3[2343:2336] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_294[6] = buffer_data_3[2351:2344] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_294[7] = buffer_data_3[2359:2352] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_294[8] = buffer_data_3[2367:2360] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_294[9] = buffer_data_3[2375:2368] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_294[10] = buffer_data_2[2343:2336] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_294[11] = buffer_data_2[2351:2344] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_294[12] = buffer_data_2[2359:2352] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_294[13] = buffer_data_2[2367:2360] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_294[14] = buffer_data_2[2375:2368] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_294[15] = buffer_data_1[2343:2336] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_294[16] = buffer_data_1[2351:2344] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_294[17] = buffer_data_1[2359:2352] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_294[18] = buffer_data_1[2367:2360] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_294[19] = buffer_data_1[2375:2368] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_294[20] = buffer_data_0[2343:2336] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_294[21] = buffer_data_0[2351:2344] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_294[22] = buffer_data_0[2359:2352] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_294[23] = buffer_data_0[2367:2360] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_294[24] = buffer_data_0[2375:2368] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_294 = kernel_img_mul_294[0] + kernel_img_mul_294[1] + kernel_img_mul_294[2] + 
                kernel_img_mul_294[3] + kernel_img_mul_294[4] + kernel_img_mul_294[5] + 
                kernel_img_mul_294[6] + kernel_img_mul_294[7] + kernel_img_mul_294[8] + 
                kernel_img_mul_294[9] + kernel_img_mul_294[10] + kernel_img_mul_294[11] + 
                kernel_img_mul_294[12] + kernel_img_mul_294[13] + kernel_img_mul_294[14] + 
                kernel_img_mul_294[15] + kernel_img_mul_294[16] + kernel_img_mul_294[17] + 
                kernel_img_mul_294[18] + kernel_img_mul_294[19] + kernel_img_mul_294[20] + 
                kernel_img_mul_294[21] + kernel_img_mul_294[22] + kernel_img_mul_294[23] + 
                kernel_img_mul_294[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2359:2352] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2359:2352] <= kernel_img_sum_294[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2359:2352] <= 'd0;
end

wire  [39:0]  kernel_img_mul_295[0:24];
assign kernel_img_mul_295[0] = buffer_data_4[2351:2344] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_295[1] = buffer_data_4[2359:2352] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_295[2] = buffer_data_4[2367:2360] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_295[3] = buffer_data_4[2375:2368] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_295[4] = buffer_data_4[2383:2376] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_295[5] = buffer_data_3[2351:2344] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_295[6] = buffer_data_3[2359:2352] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_295[7] = buffer_data_3[2367:2360] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_295[8] = buffer_data_3[2375:2368] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_295[9] = buffer_data_3[2383:2376] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_295[10] = buffer_data_2[2351:2344] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_295[11] = buffer_data_2[2359:2352] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_295[12] = buffer_data_2[2367:2360] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_295[13] = buffer_data_2[2375:2368] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_295[14] = buffer_data_2[2383:2376] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_295[15] = buffer_data_1[2351:2344] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_295[16] = buffer_data_1[2359:2352] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_295[17] = buffer_data_1[2367:2360] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_295[18] = buffer_data_1[2375:2368] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_295[19] = buffer_data_1[2383:2376] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_295[20] = buffer_data_0[2351:2344] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_295[21] = buffer_data_0[2359:2352] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_295[22] = buffer_data_0[2367:2360] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_295[23] = buffer_data_0[2375:2368] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_295[24] = buffer_data_0[2383:2376] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_295 = kernel_img_mul_295[0] + kernel_img_mul_295[1] + kernel_img_mul_295[2] + 
                kernel_img_mul_295[3] + kernel_img_mul_295[4] + kernel_img_mul_295[5] + 
                kernel_img_mul_295[6] + kernel_img_mul_295[7] + kernel_img_mul_295[8] + 
                kernel_img_mul_295[9] + kernel_img_mul_295[10] + kernel_img_mul_295[11] + 
                kernel_img_mul_295[12] + kernel_img_mul_295[13] + kernel_img_mul_295[14] + 
                kernel_img_mul_295[15] + kernel_img_mul_295[16] + kernel_img_mul_295[17] + 
                kernel_img_mul_295[18] + kernel_img_mul_295[19] + kernel_img_mul_295[20] + 
                kernel_img_mul_295[21] + kernel_img_mul_295[22] + kernel_img_mul_295[23] + 
                kernel_img_mul_295[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2367:2360] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2367:2360] <= kernel_img_sum_295[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2367:2360] <= 'd0;
end

wire  [39:0]  kernel_img_mul_296[0:24];
assign kernel_img_mul_296[0] = buffer_data_4[2359:2352] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_296[1] = buffer_data_4[2367:2360] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_296[2] = buffer_data_4[2375:2368] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_296[3] = buffer_data_4[2383:2376] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_296[4] = buffer_data_4[2391:2384] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_296[5] = buffer_data_3[2359:2352] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_296[6] = buffer_data_3[2367:2360] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_296[7] = buffer_data_3[2375:2368] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_296[8] = buffer_data_3[2383:2376] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_296[9] = buffer_data_3[2391:2384] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_296[10] = buffer_data_2[2359:2352] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_296[11] = buffer_data_2[2367:2360] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_296[12] = buffer_data_2[2375:2368] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_296[13] = buffer_data_2[2383:2376] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_296[14] = buffer_data_2[2391:2384] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_296[15] = buffer_data_1[2359:2352] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_296[16] = buffer_data_1[2367:2360] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_296[17] = buffer_data_1[2375:2368] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_296[18] = buffer_data_1[2383:2376] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_296[19] = buffer_data_1[2391:2384] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_296[20] = buffer_data_0[2359:2352] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_296[21] = buffer_data_0[2367:2360] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_296[22] = buffer_data_0[2375:2368] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_296[23] = buffer_data_0[2383:2376] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_296[24] = buffer_data_0[2391:2384] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_296 = kernel_img_mul_296[0] + kernel_img_mul_296[1] + kernel_img_mul_296[2] + 
                kernel_img_mul_296[3] + kernel_img_mul_296[4] + kernel_img_mul_296[5] + 
                kernel_img_mul_296[6] + kernel_img_mul_296[7] + kernel_img_mul_296[8] + 
                kernel_img_mul_296[9] + kernel_img_mul_296[10] + kernel_img_mul_296[11] + 
                kernel_img_mul_296[12] + kernel_img_mul_296[13] + kernel_img_mul_296[14] + 
                kernel_img_mul_296[15] + kernel_img_mul_296[16] + kernel_img_mul_296[17] + 
                kernel_img_mul_296[18] + kernel_img_mul_296[19] + kernel_img_mul_296[20] + 
                kernel_img_mul_296[21] + kernel_img_mul_296[22] + kernel_img_mul_296[23] + 
                kernel_img_mul_296[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2375:2368] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2375:2368] <= kernel_img_sum_296[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2375:2368] <= 'd0;
end

wire  [39:0]  kernel_img_mul_297[0:24];
assign kernel_img_mul_297[0] = buffer_data_4[2367:2360] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_297[1] = buffer_data_4[2375:2368] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_297[2] = buffer_data_4[2383:2376] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_297[3] = buffer_data_4[2391:2384] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_297[4] = buffer_data_4[2399:2392] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_297[5] = buffer_data_3[2367:2360] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_297[6] = buffer_data_3[2375:2368] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_297[7] = buffer_data_3[2383:2376] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_297[8] = buffer_data_3[2391:2384] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_297[9] = buffer_data_3[2399:2392] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_297[10] = buffer_data_2[2367:2360] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_297[11] = buffer_data_2[2375:2368] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_297[12] = buffer_data_2[2383:2376] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_297[13] = buffer_data_2[2391:2384] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_297[14] = buffer_data_2[2399:2392] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_297[15] = buffer_data_1[2367:2360] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_297[16] = buffer_data_1[2375:2368] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_297[17] = buffer_data_1[2383:2376] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_297[18] = buffer_data_1[2391:2384] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_297[19] = buffer_data_1[2399:2392] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_297[20] = buffer_data_0[2367:2360] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_297[21] = buffer_data_0[2375:2368] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_297[22] = buffer_data_0[2383:2376] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_297[23] = buffer_data_0[2391:2384] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_297[24] = buffer_data_0[2399:2392] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_297 = kernel_img_mul_297[0] + kernel_img_mul_297[1] + kernel_img_mul_297[2] + 
                kernel_img_mul_297[3] + kernel_img_mul_297[4] + kernel_img_mul_297[5] + 
                kernel_img_mul_297[6] + kernel_img_mul_297[7] + kernel_img_mul_297[8] + 
                kernel_img_mul_297[9] + kernel_img_mul_297[10] + kernel_img_mul_297[11] + 
                kernel_img_mul_297[12] + kernel_img_mul_297[13] + kernel_img_mul_297[14] + 
                kernel_img_mul_297[15] + kernel_img_mul_297[16] + kernel_img_mul_297[17] + 
                kernel_img_mul_297[18] + kernel_img_mul_297[19] + kernel_img_mul_297[20] + 
                kernel_img_mul_297[21] + kernel_img_mul_297[22] + kernel_img_mul_297[23] + 
                kernel_img_mul_297[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2383:2376] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2383:2376] <= kernel_img_sum_297[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2383:2376] <= 'd0;
end

wire  [39:0]  kernel_img_mul_298[0:24];
assign kernel_img_mul_298[0] = buffer_data_4[2375:2368] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_298[1] = buffer_data_4[2383:2376] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_298[2] = buffer_data_4[2391:2384] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_298[3] = buffer_data_4[2399:2392] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_298[4] = buffer_data_4[2407:2400] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_298[5] = buffer_data_3[2375:2368] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_298[6] = buffer_data_3[2383:2376] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_298[7] = buffer_data_3[2391:2384] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_298[8] = buffer_data_3[2399:2392] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_298[9] = buffer_data_3[2407:2400] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_298[10] = buffer_data_2[2375:2368] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_298[11] = buffer_data_2[2383:2376] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_298[12] = buffer_data_2[2391:2384] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_298[13] = buffer_data_2[2399:2392] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_298[14] = buffer_data_2[2407:2400] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_298[15] = buffer_data_1[2375:2368] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_298[16] = buffer_data_1[2383:2376] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_298[17] = buffer_data_1[2391:2384] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_298[18] = buffer_data_1[2399:2392] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_298[19] = buffer_data_1[2407:2400] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_298[20] = buffer_data_0[2375:2368] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_298[21] = buffer_data_0[2383:2376] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_298[22] = buffer_data_0[2391:2384] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_298[23] = buffer_data_0[2399:2392] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_298[24] = buffer_data_0[2407:2400] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_298 = kernel_img_mul_298[0] + kernel_img_mul_298[1] + kernel_img_mul_298[2] + 
                kernel_img_mul_298[3] + kernel_img_mul_298[4] + kernel_img_mul_298[5] + 
                kernel_img_mul_298[6] + kernel_img_mul_298[7] + kernel_img_mul_298[8] + 
                kernel_img_mul_298[9] + kernel_img_mul_298[10] + kernel_img_mul_298[11] + 
                kernel_img_mul_298[12] + kernel_img_mul_298[13] + kernel_img_mul_298[14] + 
                kernel_img_mul_298[15] + kernel_img_mul_298[16] + kernel_img_mul_298[17] + 
                kernel_img_mul_298[18] + kernel_img_mul_298[19] + kernel_img_mul_298[20] + 
                kernel_img_mul_298[21] + kernel_img_mul_298[22] + kernel_img_mul_298[23] + 
                kernel_img_mul_298[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2391:2384] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2391:2384] <= kernel_img_sum_298[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2391:2384] <= 'd0;
end

wire  [39:0]  kernel_img_mul_299[0:24];
assign kernel_img_mul_299[0] = buffer_data_4[2383:2376] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_299[1] = buffer_data_4[2391:2384] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_299[2] = buffer_data_4[2399:2392] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_299[3] = buffer_data_4[2407:2400] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_299[4] = buffer_data_4[2415:2408] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_299[5] = buffer_data_3[2383:2376] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_299[6] = buffer_data_3[2391:2384] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_299[7] = buffer_data_3[2399:2392] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_299[8] = buffer_data_3[2407:2400] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_299[9] = buffer_data_3[2415:2408] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_299[10] = buffer_data_2[2383:2376] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_299[11] = buffer_data_2[2391:2384] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_299[12] = buffer_data_2[2399:2392] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_299[13] = buffer_data_2[2407:2400] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_299[14] = buffer_data_2[2415:2408] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_299[15] = buffer_data_1[2383:2376] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_299[16] = buffer_data_1[2391:2384] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_299[17] = buffer_data_1[2399:2392] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_299[18] = buffer_data_1[2407:2400] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_299[19] = buffer_data_1[2415:2408] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_299[20] = buffer_data_0[2383:2376] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_299[21] = buffer_data_0[2391:2384] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_299[22] = buffer_data_0[2399:2392] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_299[23] = buffer_data_0[2407:2400] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_299[24] = buffer_data_0[2415:2408] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_299 = kernel_img_mul_299[0] + kernel_img_mul_299[1] + kernel_img_mul_299[2] + 
                kernel_img_mul_299[3] + kernel_img_mul_299[4] + kernel_img_mul_299[5] + 
                kernel_img_mul_299[6] + kernel_img_mul_299[7] + kernel_img_mul_299[8] + 
                kernel_img_mul_299[9] + kernel_img_mul_299[10] + kernel_img_mul_299[11] + 
                kernel_img_mul_299[12] + kernel_img_mul_299[13] + kernel_img_mul_299[14] + 
                kernel_img_mul_299[15] + kernel_img_mul_299[16] + kernel_img_mul_299[17] + 
                kernel_img_mul_299[18] + kernel_img_mul_299[19] + kernel_img_mul_299[20] + 
                kernel_img_mul_299[21] + kernel_img_mul_299[22] + kernel_img_mul_299[23] + 
                kernel_img_mul_299[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2399:2392] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2399:2392] <= kernel_img_sum_299[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2399:2392] <= 'd0;
end

wire  [39:0]  kernel_img_mul_300[0:24];
assign kernel_img_mul_300[0] = buffer_data_4[2391:2384] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_300[1] = buffer_data_4[2399:2392] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_300[2] = buffer_data_4[2407:2400] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_300[3] = buffer_data_4[2415:2408] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_300[4] = buffer_data_4[2423:2416] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_300[5] = buffer_data_3[2391:2384] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_300[6] = buffer_data_3[2399:2392] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_300[7] = buffer_data_3[2407:2400] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_300[8] = buffer_data_3[2415:2408] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_300[9] = buffer_data_3[2423:2416] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_300[10] = buffer_data_2[2391:2384] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_300[11] = buffer_data_2[2399:2392] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_300[12] = buffer_data_2[2407:2400] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_300[13] = buffer_data_2[2415:2408] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_300[14] = buffer_data_2[2423:2416] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_300[15] = buffer_data_1[2391:2384] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_300[16] = buffer_data_1[2399:2392] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_300[17] = buffer_data_1[2407:2400] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_300[18] = buffer_data_1[2415:2408] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_300[19] = buffer_data_1[2423:2416] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_300[20] = buffer_data_0[2391:2384] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_300[21] = buffer_data_0[2399:2392] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_300[22] = buffer_data_0[2407:2400] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_300[23] = buffer_data_0[2415:2408] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_300[24] = buffer_data_0[2423:2416] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_300 = kernel_img_mul_300[0] + kernel_img_mul_300[1] + kernel_img_mul_300[2] + 
                kernel_img_mul_300[3] + kernel_img_mul_300[4] + kernel_img_mul_300[5] + 
                kernel_img_mul_300[6] + kernel_img_mul_300[7] + kernel_img_mul_300[8] + 
                kernel_img_mul_300[9] + kernel_img_mul_300[10] + kernel_img_mul_300[11] + 
                kernel_img_mul_300[12] + kernel_img_mul_300[13] + kernel_img_mul_300[14] + 
                kernel_img_mul_300[15] + kernel_img_mul_300[16] + kernel_img_mul_300[17] + 
                kernel_img_mul_300[18] + kernel_img_mul_300[19] + kernel_img_mul_300[20] + 
                kernel_img_mul_300[21] + kernel_img_mul_300[22] + kernel_img_mul_300[23] + 
                kernel_img_mul_300[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2407:2400] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2407:2400] <= kernel_img_sum_300[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2407:2400] <= 'd0;
end

wire  [39:0]  kernel_img_mul_301[0:24];
assign kernel_img_mul_301[0] = buffer_data_4[2399:2392] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_301[1] = buffer_data_4[2407:2400] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_301[2] = buffer_data_4[2415:2408] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_301[3] = buffer_data_4[2423:2416] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_301[4] = buffer_data_4[2431:2424] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_301[5] = buffer_data_3[2399:2392] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_301[6] = buffer_data_3[2407:2400] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_301[7] = buffer_data_3[2415:2408] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_301[8] = buffer_data_3[2423:2416] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_301[9] = buffer_data_3[2431:2424] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_301[10] = buffer_data_2[2399:2392] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_301[11] = buffer_data_2[2407:2400] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_301[12] = buffer_data_2[2415:2408] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_301[13] = buffer_data_2[2423:2416] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_301[14] = buffer_data_2[2431:2424] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_301[15] = buffer_data_1[2399:2392] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_301[16] = buffer_data_1[2407:2400] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_301[17] = buffer_data_1[2415:2408] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_301[18] = buffer_data_1[2423:2416] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_301[19] = buffer_data_1[2431:2424] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_301[20] = buffer_data_0[2399:2392] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_301[21] = buffer_data_0[2407:2400] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_301[22] = buffer_data_0[2415:2408] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_301[23] = buffer_data_0[2423:2416] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_301[24] = buffer_data_0[2431:2424] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_301 = kernel_img_mul_301[0] + kernel_img_mul_301[1] + kernel_img_mul_301[2] + 
                kernel_img_mul_301[3] + kernel_img_mul_301[4] + kernel_img_mul_301[5] + 
                kernel_img_mul_301[6] + kernel_img_mul_301[7] + kernel_img_mul_301[8] + 
                kernel_img_mul_301[9] + kernel_img_mul_301[10] + kernel_img_mul_301[11] + 
                kernel_img_mul_301[12] + kernel_img_mul_301[13] + kernel_img_mul_301[14] + 
                kernel_img_mul_301[15] + kernel_img_mul_301[16] + kernel_img_mul_301[17] + 
                kernel_img_mul_301[18] + kernel_img_mul_301[19] + kernel_img_mul_301[20] + 
                kernel_img_mul_301[21] + kernel_img_mul_301[22] + kernel_img_mul_301[23] + 
                kernel_img_mul_301[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2415:2408] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2415:2408] <= kernel_img_sum_301[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2415:2408] <= 'd0;
end

wire  [39:0]  kernel_img_mul_302[0:24];
assign kernel_img_mul_302[0] = buffer_data_4[2407:2400] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_302[1] = buffer_data_4[2415:2408] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_302[2] = buffer_data_4[2423:2416] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_302[3] = buffer_data_4[2431:2424] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_302[4] = buffer_data_4[2439:2432] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_302[5] = buffer_data_3[2407:2400] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_302[6] = buffer_data_3[2415:2408] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_302[7] = buffer_data_3[2423:2416] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_302[8] = buffer_data_3[2431:2424] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_302[9] = buffer_data_3[2439:2432] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_302[10] = buffer_data_2[2407:2400] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_302[11] = buffer_data_2[2415:2408] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_302[12] = buffer_data_2[2423:2416] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_302[13] = buffer_data_2[2431:2424] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_302[14] = buffer_data_2[2439:2432] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_302[15] = buffer_data_1[2407:2400] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_302[16] = buffer_data_1[2415:2408] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_302[17] = buffer_data_1[2423:2416] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_302[18] = buffer_data_1[2431:2424] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_302[19] = buffer_data_1[2439:2432] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_302[20] = buffer_data_0[2407:2400] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_302[21] = buffer_data_0[2415:2408] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_302[22] = buffer_data_0[2423:2416] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_302[23] = buffer_data_0[2431:2424] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_302[24] = buffer_data_0[2439:2432] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_302 = kernel_img_mul_302[0] + kernel_img_mul_302[1] + kernel_img_mul_302[2] + 
                kernel_img_mul_302[3] + kernel_img_mul_302[4] + kernel_img_mul_302[5] + 
                kernel_img_mul_302[6] + kernel_img_mul_302[7] + kernel_img_mul_302[8] + 
                kernel_img_mul_302[9] + kernel_img_mul_302[10] + kernel_img_mul_302[11] + 
                kernel_img_mul_302[12] + kernel_img_mul_302[13] + kernel_img_mul_302[14] + 
                kernel_img_mul_302[15] + kernel_img_mul_302[16] + kernel_img_mul_302[17] + 
                kernel_img_mul_302[18] + kernel_img_mul_302[19] + kernel_img_mul_302[20] + 
                kernel_img_mul_302[21] + kernel_img_mul_302[22] + kernel_img_mul_302[23] + 
                kernel_img_mul_302[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2423:2416] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2423:2416] <= kernel_img_sum_302[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2423:2416] <= 'd0;
end

wire  [39:0]  kernel_img_mul_303[0:24];
assign kernel_img_mul_303[0] = buffer_data_4[2415:2408] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_303[1] = buffer_data_4[2423:2416] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_303[2] = buffer_data_4[2431:2424] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_303[3] = buffer_data_4[2439:2432] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_303[4] = buffer_data_4[2447:2440] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_303[5] = buffer_data_3[2415:2408] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_303[6] = buffer_data_3[2423:2416] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_303[7] = buffer_data_3[2431:2424] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_303[8] = buffer_data_3[2439:2432] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_303[9] = buffer_data_3[2447:2440] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_303[10] = buffer_data_2[2415:2408] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_303[11] = buffer_data_2[2423:2416] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_303[12] = buffer_data_2[2431:2424] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_303[13] = buffer_data_2[2439:2432] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_303[14] = buffer_data_2[2447:2440] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_303[15] = buffer_data_1[2415:2408] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_303[16] = buffer_data_1[2423:2416] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_303[17] = buffer_data_1[2431:2424] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_303[18] = buffer_data_1[2439:2432] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_303[19] = buffer_data_1[2447:2440] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_303[20] = buffer_data_0[2415:2408] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_303[21] = buffer_data_0[2423:2416] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_303[22] = buffer_data_0[2431:2424] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_303[23] = buffer_data_0[2439:2432] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_303[24] = buffer_data_0[2447:2440] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_303 = kernel_img_mul_303[0] + kernel_img_mul_303[1] + kernel_img_mul_303[2] + 
                kernel_img_mul_303[3] + kernel_img_mul_303[4] + kernel_img_mul_303[5] + 
                kernel_img_mul_303[6] + kernel_img_mul_303[7] + kernel_img_mul_303[8] + 
                kernel_img_mul_303[9] + kernel_img_mul_303[10] + kernel_img_mul_303[11] + 
                kernel_img_mul_303[12] + kernel_img_mul_303[13] + kernel_img_mul_303[14] + 
                kernel_img_mul_303[15] + kernel_img_mul_303[16] + kernel_img_mul_303[17] + 
                kernel_img_mul_303[18] + kernel_img_mul_303[19] + kernel_img_mul_303[20] + 
                kernel_img_mul_303[21] + kernel_img_mul_303[22] + kernel_img_mul_303[23] + 
                kernel_img_mul_303[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2431:2424] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2431:2424] <= kernel_img_sum_303[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2431:2424] <= 'd0;
end

wire  [39:0]  kernel_img_mul_304[0:24];
assign kernel_img_mul_304[0] = buffer_data_4[2423:2416] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_304[1] = buffer_data_4[2431:2424] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_304[2] = buffer_data_4[2439:2432] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_304[3] = buffer_data_4[2447:2440] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_304[4] = buffer_data_4[2455:2448] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_304[5] = buffer_data_3[2423:2416] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_304[6] = buffer_data_3[2431:2424] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_304[7] = buffer_data_3[2439:2432] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_304[8] = buffer_data_3[2447:2440] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_304[9] = buffer_data_3[2455:2448] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_304[10] = buffer_data_2[2423:2416] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_304[11] = buffer_data_2[2431:2424] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_304[12] = buffer_data_2[2439:2432] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_304[13] = buffer_data_2[2447:2440] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_304[14] = buffer_data_2[2455:2448] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_304[15] = buffer_data_1[2423:2416] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_304[16] = buffer_data_1[2431:2424] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_304[17] = buffer_data_1[2439:2432] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_304[18] = buffer_data_1[2447:2440] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_304[19] = buffer_data_1[2455:2448] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_304[20] = buffer_data_0[2423:2416] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_304[21] = buffer_data_0[2431:2424] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_304[22] = buffer_data_0[2439:2432] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_304[23] = buffer_data_0[2447:2440] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_304[24] = buffer_data_0[2455:2448] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_304 = kernel_img_mul_304[0] + kernel_img_mul_304[1] + kernel_img_mul_304[2] + 
                kernel_img_mul_304[3] + kernel_img_mul_304[4] + kernel_img_mul_304[5] + 
                kernel_img_mul_304[6] + kernel_img_mul_304[7] + kernel_img_mul_304[8] + 
                kernel_img_mul_304[9] + kernel_img_mul_304[10] + kernel_img_mul_304[11] + 
                kernel_img_mul_304[12] + kernel_img_mul_304[13] + kernel_img_mul_304[14] + 
                kernel_img_mul_304[15] + kernel_img_mul_304[16] + kernel_img_mul_304[17] + 
                kernel_img_mul_304[18] + kernel_img_mul_304[19] + kernel_img_mul_304[20] + 
                kernel_img_mul_304[21] + kernel_img_mul_304[22] + kernel_img_mul_304[23] + 
                kernel_img_mul_304[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2439:2432] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2439:2432] <= kernel_img_sum_304[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2439:2432] <= 'd0;
end

wire  [39:0]  kernel_img_mul_305[0:24];
assign kernel_img_mul_305[0] = buffer_data_4[2431:2424] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_305[1] = buffer_data_4[2439:2432] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_305[2] = buffer_data_4[2447:2440] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_305[3] = buffer_data_4[2455:2448] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_305[4] = buffer_data_4[2463:2456] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_305[5] = buffer_data_3[2431:2424] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_305[6] = buffer_data_3[2439:2432] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_305[7] = buffer_data_3[2447:2440] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_305[8] = buffer_data_3[2455:2448] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_305[9] = buffer_data_3[2463:2456] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_305[10] = buffer_data_2[2431:2424] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_305[11] = buffer_data_2[2439:2432] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_305[12] = buffer_data_2[2447:2440] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_305[13] = buffer_data_2[2455:2448] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_305[14] = buffer_data_2[2463:2456] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_305[15] = buffer_data_1[2431:2424] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_305[16] = buffer_data_1[2439:2432] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_305[17] = buffer_data_1[2447:2440] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_305[18] = buffer_data_1[2455:2448] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_305[19] = buffer_data_1[2463:2456] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_305[20] = buffer_data_0[2431:2424] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_305[21] = buffer_data_0[2439:2432] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_305[22] = buffer_data_0[2447:2440] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_305[23] = buffer_data_0[2455:2448] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_305[24] = buffer_data_0[2463:2456] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_305 = kernel_img_mul_305[0] + kernel_img_mul_305[1] + kernel_img_mul_305[2] + 
                kernel_img_mul_305[3] + kernel_img_mul_305[4] + kernel_img_mul_305[5] + 
                kernel_img_mul_305[6] + kernel_img_mul_305[7] + kernel_img_mul_305[8] + 
                kernel_img_mul_305[9] + kernel_img_mul_305[10] + kernel_img_mul_305[11] + 
                kernel_img_mul_305[12] + kernel_img_mul_305[13] + kernel_img_mul_305[14] + 
                kernel_img_mul_305[15] + kernel_img_mul_305[16] + kernel_img_mul_305[17] + 
                kernel_img_mul_305[18] + kernel_img_mul_305[19] + kernel_img_mul_305[20] + 
                kernel_img_mul_305[21] + kernel_img_mul_305[22] + kernel_img_mul_305[23] + 
                kernel_img_mul_305[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2447:2440] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2447:2440] <= kernel_img_sum_305[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2447:2440] <= 'd0;
end

wire  [39:0]  kernel_img_mul_306[0:24];
assign kernel_img_mul_306[0] = buffer_data_4[2439:2432] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_306[1] = buffer_data_4[2447:2440] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_306[2] = buffer_data_4[2455:2448] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_306[3] = buffer_data_4[2463:2456] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_306[4] = buffer_data_4[2471:2464] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_306[5] = buffer_data_3[2439:2432] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_306[6] = buffer_data_3[2447:2440] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_306[7] = buffer_data_3[2455:2448] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_306[8] = buffer_data_3[2463:2456] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_306[9] = buffer_data_3[2471:2464] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_306[10] = buffer_data_2[2439:2432] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_306[11] = buffer_data_2[2447:2440] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_306[12] = buffer_data_2[2455:2448] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_306[13] = buffer_data_2[2463:2456] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_306[14] = buffer_data_2[2471:2464] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_306[15] = buffer_data_1[2439:2432] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_306[16] = buffer_data_1[2447:2440] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_306[17] = buffer_data_1[2455:2448] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_306[18] = buffer_data_1[2463:2456] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_306[19] = buffer_data_1[2471:2464] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_306[20] = buffer_data_0[2439:2432] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_306[21] = buffer_data_0[2447:2440] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_306[22] = buffer_data_0[2455:2448] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_306[23] = buffer_data_0[2463:2456] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_306[24] = buffer_data_0[2471:2464] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_306 = kernel_img_mul_306[0] + kernel_img_mul_306[1] + kernel_img_mul_306[2] + 
                kernel_img_mul_306[3] + kernel_img_mul_306[4] + kernel_img_mul_306[5] + 
                kernel_img_mul_306[6] + kernel_img_mul_306[7] + kernel_img_mul_306[8] + 
                kernel_img_mul_306[9] + kernel_img_mul_306[10] + kernel_img_mul_306[11] + 
                kernel_img_mul_306[12] + kernel_img_mul_306[13] + kernel_img_mul_306[14] + 
                kernel_img_mul_306[15] + kernel_img_mul_306[16] + kernel_img_mul_306[17] + 
                kernel_img_mul_306[18] + kernel_img_mul_306[19] + kernel_img_mul_306[20] + 
                kernel_img_mul_306[21] + kernel_img_mul_306[22] + kernel_img_mul_306[23] + 
                kernel_img_mul_306[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2455:2448] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2455:2448] <= kernel_img_sum_306[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2455:2448] <= 'd0;
end

wire  [39:0]  kernel_img_mul_307[0:24];
assign kernel_img_mul_307[0] = buffer_data_4[2447:2440] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_307[1] = buffer_data_4[2455:2448] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_307[2] = buffer_data_4[2463:2456] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_307[3] = buffer_data_4[2471:2464] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_307[4] = buffer_data_4[2479:2472] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_307[5] = buffer_data_3[2447:2440] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_307[6] = buffer_data_3[2455:2448] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_307[7] = buffer_data_3[2463:2456] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_307[8] = buffer_data_3[2471:2464] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_307[9] = buffer_data_3[2479:2472] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_307[10] = buffer_data_2[2447:2440] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_307[11] = buffer_data_2[2455:2448] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_307[12] = buffer_data_2[2463:2456] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_307[13] = buffer_data_2[2471:2464] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_307[14] = buffer_data_2[2479:2472] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_307[15] = buffer_data_1[2447:2440] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_307[16] = buffer_data_1[2455:2448] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_307[17] = buffer_data_1[2463:2456] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_307[18] = buffer_data_1[2471:2464] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_307[19] = buffer_data_1[2479:2472] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_307[20] = buffer_data_0[2447:2440] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_307[21] = buffer_data_0[2455:2448] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_307[22] = buffer_data_0[2463:2456] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_307[23] = buffer_data_0[2471:2464] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_307[24] = buffer_data_0[2479:2472] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_307 = kernel_img_mul_307[0] + kernel_img_mul_307[1] + kernel_img_mul_307[2] + 
                kernel_img_mul_307[3] + kernel_img_mul_307[4] + kernel_img_mul_307[5] + 
                kernel_img_mul_307[6] + kernel_img_mul_307[7] + kernel_img_mul_307[8] + 
                kernel_img_mul_307[9] + kernel_img_mul_307[10] + kernel_img_mul_307[11] + 
                kernel_img_mul_307[12] + kernel_img_mul_307[13] + kernel_img_mul_307[14] + 
                kernel_img_mul_307[15] + kernel_img_mul_307[16] + kernel_img_mul_307[17] + 
                kernel_img_mul_307[18] + kernel_img_mul_307[19] + kernel_img_mul_307[20] + 
                kernel_img_mul_307[21] + kernel_img_mul_307[22] + kernel_img_mul_307[23] + 
                kernel_img_mul_307[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2463:2456] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2463:2456] <= kernel_img_sum_307[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2463:2456] <= 'd0;
end

wire  [39:0]  kernel_img_mul_308[0:24];
assign kernel_img_mul_308[0] = buffer_data_4[2455:2448] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_308[1] = buffer_data_4[2463:2456] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_308[2] = buffer_data_4[2471:2464] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_308[3] = buffer_data_4[2479:2472] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_308[4] = buffer_data_4[2487:2480] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_308[5] = buffer_data_3[2455:2448] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_308[6] = buffer_data_3[2463:2456] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_308[7] = buffer_data_3[2471:2464] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_308[8] = buffer_data_3[2479:2472] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_308[9] = buffer_data_3[2487:2480] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_308[10] = buffer_data_2[2455:2448] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_308[11] = buffer_data_2[2463:2456] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_308[12] = buffer_data_2[2471:2464] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_308[13] = buffer_data_2[2479:2472] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_308[14] = buffer_data_2[2487:2480] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_308[15] = buffer_data_1[2455:2448] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_308[16] = buffer_data_1[2463:2456] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_308[17] = buffer_data_1[2471:2464] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_308[18] = buffer_data_1[2479:2472] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_308[19] = buffer_data_1[2487:2480] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_308[20] = buffer_data_0[2455:2448] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_308[21] = buffer_data_0[2463:2456] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_308[22] = buffer_data_0[2471:2464] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_308[23] = buffer_data_0[2479:2472] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_308[24] = buffer_data_0[2487:2480] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_308 = kernel_img_mul_308[0] + kernel_img_mul_308[1] + kernel_img_mul_308[2] + 
                kernel_img_mul_308[3] + kernel_img_mul_308[4] + kernel_img_mul_308[5] + 
                kernel_img_mul_308[6] + kernel_img_mul_308[7] + kernel_img_mul_308[8] + 
                kernel_img_mul_308[9] + kernel_img_mul_308[10] + kernel_img_mul_308[11] + 
                kernel_img_mul_308[12] + kernel_img_mul_308[13] + kernel_img_mul_308[14] + 
                kernel_img_mul_308[15] + kernel_img_mul_308[16] + kernel_img_mul_308[17] + 
                kernel_img_mul_308[18] + kernel_img_mul_308[19] + kernel_img_mul_308[20] + 
                kernel_img_mul_308[21] + kernel_img_mul_308[22] + kernel_img_mul_308[23] + 
                kernel_img_mul_308[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2471:2464] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2471:2464] <= kernel_img_sum_308[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2471:2464] <= 'd0;
end

wire  [39:0]  kernel_img_mul_309[0:24];
assign kernel_img_mul_309[0] = buffer_data_4[2463:2456] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_309[1] = buffer_data_4[2471:2464] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_309[2] = buffer_data_4[2479:2472] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_309[3] = buffer_data_4[2487:2480] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_309[4] = buffer_data_4[2495:2488] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_309[5] = buffer_data_3[2463:2456] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_309[6] = buffer_data_3[2471:2464] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_309[7] = buffer_data_3[2479:2472] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_309[8] = buffer_data_3[2487:2480] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_309[9] = buffer_data_3[2495:2488] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_309[10] = buffer_data_2[2463:2456] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_309[11] = buffer_data_2[2471:2464] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_309[12] = buffer_data_2[2479:2472] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_309[13] = buffer_data_2[2487:2480] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_309[14] = buffer_data_2[2495:2488] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_309[15] = buffer_data_1[2463:2456] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_309[16] = buffer_data_1[2471:2464] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_309[17] = buffer_data_1[2479:2472] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_309[18] = buffer_data_1[2487:2480] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_309[19] = buffer_data_1[2495:2488] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_309[20] = buffer_data_0[2463:2456] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_309[21] = buffer_data_0[2471:2464] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_309[22] = buffer_data_0[2479:2472] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_309[23] = buffer_data_0[2487:2480] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_309[24] = buffer_data_0[2495:2488] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_309 = kernel_img_mul_309[0] + kernel_img_mul_309[1] + kernel_img_mul_309[2] + 
                kernel_img_mul_309[3] + kernel_img_mul_309[4] + kernel_img_mul_309[5] + 
                kernel_img_mul_309[6] + kernel_img_mul_309[7] + kernel_img_mul_309[8] + 
                kernel_img_mul_309[9] + kernel_img_mul_309[10] + kernel_img_mul_309[11] + 
                kernel_img_mul_309[12] + kernel_img_mul_309[13] + kernel_img_mul_309[14] + 
                kernel_img_mul_309[15] + kernel_img_mul_309[16] + kernel_img_mul_309[17] + 
                kernel_img_mul_309[18] + kernel_img_mul_309[19] + kernel_img_mul_309[20] + 
                kernel_img_mul_309[21] + kernel_img_mul_309[22] + kernel_img_mul_309[23] + 
                kernel_img_mul_309[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2479:2472] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2479:2472] <= kernel_img_sum_309[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2479:2472] <= 'd0;
end

wire  [39:0]  kernel_img_mul_310[0:24];
assign kernel_img_mul_310[0] = buffer_data_4[2471:2464] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_310[1] = buffer_data_4[2479:2472] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_310[2] = buffer_data_4[2487:2480] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_310[3] = buffer_data_4[2495:2488] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_310[4] = buffer_data_4[2503:2496] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_310[5] = buffer_data_3[2471:2464] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_310[6] = buffer_data_3[2479:2472] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_310[7] = buffer_data_3[2487:2480] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_310[8] = buffer_data_3[2495:2488] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_310[9] = buffer_data_3[2503:2496] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_310[10] = buffer_data_2[2471:2464] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_310[11] = buffer_data_2[2479:2472] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_310[12] = buffer_data_2[2487:2480] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_310[13] = buffer_data_2[2495:2488] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_310[14] = buffer_data_2[2503:2496] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_310[15] = buffer_data_1[2471:2464] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_310[16] = buffer_data_1[2479:2472] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_310[17] = buffer_data_1[2487:2480] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_310[18] = buffer_data_1[2495:2488] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_310[19] = buffer_data_1[2503:2496] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_310[20] = buffer_data_0[2471:2464] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_310[21] = buffer_data_0[2479:2472] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_310[22] = buffer_data_0[2487:2480] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_310[23] = buffer_data_0[2495:2488] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_310[24] = buffer_data_0[2503:2496] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_310 = kernel_img_mul_310[0] + kernel_img_mul_310[1] + kernel_img_mul_310[2] + 
                kernel_img_mul_310[3] + kernel_img_mul_310[4] + kernel_img_mul_310[5] + 
                kernel_img_mul_310[6] + kernel_img_mul_310[7] + kernel_img_mul_310[8] + 
                kernel_img_mul_310[9] + kernel_img_mul_310[10] + kernel_img_mul_310[11] + 
                kernel_img_mul_310[12] + kernel_img_mul_310[13] + kernel_img_mul_310[14] + 
                kernel_img_mul_310[15] + kernel_img_mul_310[16] + kernel_img_mul_310[17] + 
                kernel_img_mul_310[18] + kernel_img_mul_310[19] + kernel_img_mul_310[20] + 
                kernel_img_mul_310[21] + kernel_img_mul_310[22] + kernel_img_mul_310[23] + 
                kernel_img_mul_310[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2487:2480] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2487:2480] <= kernel_img_sum_310[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2487:2480] <= 'd0;
end

wire  [39:0]  kernel_img_mul_311[0:24];
assign kernel_img_mul_311[0] = buffer_data_4[2479:2472] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_311[1] = buffer_data_4[2487:2480] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_311[2] = buffer_data_4[2495:2488] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_311[3] = buffer_data_4[2503:2496] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_311[4] = buffer_data_4[2511:2504] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_311[5] = buffer_data_3[2479:2472] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_311[6] = buffer_data_3[2487:2480] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_311[7] = buffer_data_3[2495:2488] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_311[8] = buffer_data_3[2503:2496] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_311[9] = buffer_data_3[2511:2504] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_311[10] = buffer_data_2[2479:2472] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_311[11] = buffer_data_2[2487:2480] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_311[12] = buffer_data_2[2495:2488] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_311[13] = buffer_data_2[2503:2496] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_311[14] = buffer_data_2[2511:2504] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_311[15] = buffer_data_1[2479:2472] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_311[16] = buffer_data_1[2487:2480] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_311[17] = buffer_data_1[2495:2488] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_311[18] = buffer_data_1[2503:2496] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_311[19] = buffer_data_1[2511:2504] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_311[20] = buffer_data_0[2479:2472] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_311[21] = buffer_data_0[2487:2480] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_311[22] = buffer_data_0[2495:2488] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_311[23] = buffer_data_0[2503:2496] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_311[24] = buffer_data_0[2511:2504] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_311 = kernel_img_mul_311[0] + kernel_img_mul_311[1] + kernel_img_mul_311[2] + 
                kernel_img_mul_311[3] + kernel_img_mul_311[4] + kernel_img_mul_311[5] + 
                kernel_img_mul_311[6] + kernel_img_mul_311[7] + kernel_img_mul_311[8] + 
                kernel_img_mul_311[9] + kernel_img_mul_311[10] + kernel_img_mul_311[11] + 
                kernel_img_mul_311[12] + kernel_img_mul_311[13] + kernel_img_mul_311[14] + 
                kernel_img_mul_311[15] + kernel_img_mul_311[16] + kernel_img_mul_311[17] + 
                kernel_img_mul_311[18] + kernel_img_mul_311[19] + kernel_img_mul_311[20] + 
                kernel_img_mul_311[21] + kernel_img_mul_311[22] + kernel_img_mul_311[23] + 
                kernel_img_mul_311[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2495:2488] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2495:2488] <= kernel_img_sum_311[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2495:2488] <= 'd0;
end

wire  [39:0]  kernel_img_mul_312[0:24];
assign kernel_img_mul_312[0] = buffer_data_4[2487:2480] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_312[1] = buffer_data_4[2495:2488] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_312[2] = buffer_data_4[2503:2496] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_312[3] = buffer_data_4[2511:2504] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_312[4] = buffer_data_4[2519:2512] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_312[5] = buffer_data_3[2487:2480] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_312[6] = buffer_data_3[2495:2488] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_312[7] = buffer_data_3[2503:2496] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_312[8] = buffer_data_3[2511:2504] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_312[9] = buffer_data_3[2519:2512] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_312[10] = buffer_data_2[2487:2480] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_312[11] = buffer_data_2[2495:2488] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_312[12] = buffer_data_2[2503:2496] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_312[13] = buffer_data_2[2511:2504] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_312[14] = buffer_data_2[2519:2512] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_312[15] = buffer_data_1[2487:2480] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_312[16] = buffer_data_1[2495:2488] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_312[17] = buffer_data_1[2503:2496] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_312[18] = buffer_data_1[2511:2504] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_312[19] = buffer_data_1[2519:2512] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_312[20] = buffer_data_0[2487:2480] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_312[21] = buffer_data_0[2495:2488] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_312[22] = buffer_data_0[2503:2496] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_312[23] = buffer_data_0[2511:2504] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_312[24] = buffer_data_0[2519:2512] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_312 = kernel_img_mul_312[0] + kernel_img_mul_312[1] + kernel_img_mul_312[2] + 
                kernel_img_mul_312[3] + kernel_img_mul_312[4] + kernel_img_mul_312[5] + 
                kernel_img_mul_312[6] + kernel_img_mul_312[7] + kernel_img_mul_312[8] + 
                kernel_img_mul_312[9] + kernel_img_mul_312[10] + kernel_img_mul_312[11] + 
                kernel_img_mul_312[12] + kernel_img_mul_312[13] + kernel_img_mul_312[14] + 
                kernel_img_mul_312[15] + kernel_img_mul_312[16] + kernel_img_mul_312[17] + 
                kernel_img_mul_312[18] + kernel_img_mul_312[19] + kernel_img_mul_312[20] + 
                kernel_img_mul_312[21] + kernel_img_mul_312[22] + kernel_img_mul_312[23] + 
                kernel_img_mul_312[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2503:2496] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2503:2496] <= kernel_img_sum_312[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2503:2496] <= 'd0;
end

wire  [39:0]  kernel_img_mul_313[0:24];
assign kernel_img_mul_313[0] = buffer_data_4[2495:2488] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_313[1] = buffer_data_4[2503:2496] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_313[2] = buffer_data_4[2511:2504] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_313[3] = buffer_data_4[2519:2512] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_313[4] = buffer_data_4[2527:2520] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_313[5] = buffer_data_3[2495:2488] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_313[6] = buffer_data_3[2503:2496] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_313[7] = buffer_data_3[2511:2504] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_313[8] = buffer_data_3[2519:2512] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_313[9] = buffer_data_3[2527:2520] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_313[10] = buffer_data_2[2495:2488] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_313[11] = buffer_data_2[2503:2496] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_313[12] = buffer_data_2[2511:2504] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_313[13] = buffer_data_2[2519:2512] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_313[14] = buffer_data_2[2527:2520] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_313[15] = buffer_data_1[2495:2488] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_313[16] = buffer_data_1[2503:2496] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_313[17] = buffer_data_1[2511:2504] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_313[18] = buffer_data_1[2519:2512] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_313[19] = buffer_data_1[2527:2520] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_313[20] = buffer_data_0[2495:2488] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_313[21] = buffer_data_0[2503:2496] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_313[22] = buffer_data_0[2511:2504] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_313[23] = buffer_data_0[2519:2512] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_313[24] = buffer_data_0[2527:2520] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_313 = kernel_img_mul_313[0] + kernel_img_mul_313[1] + kernel_img_mul_313[2] + 
                kernel_img_mul_313[3] + kernel_img_mul_313[4] + kernel_img_mul_313[5] + 
                kernel_img_mul_313[6] + kernel_img_mul_313[7] + kernel_img_mul_313[8] + 
                kernel_img_mul_313[9] + kernel_img_mul_313[10] + kernel_img_mul_313[11] + 
                kernel_img_mul_313[12] + kernel_img_mul_313[13] + kernel_img_mul_313[14] + 
                kernel_img_mul_313[15] + kernel_img_mul_313[16] + kernel_img_mul_313[17] + 
                kernel_img_mul_313[18] + kernel_img_mul_313[19] + kernel_img_mul_313[20] + 
                kernel_img_mul_313[21] + kernel_img_mul_313[22] + kernel_img_mul_313[23] + 
                kernel_img_mul_313[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2511:2504] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2511:2504] <= kernel_img_sum_313[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2511:2504] <= 'd0;
end

wire  [39:0]  kernel_img_mul_314[0:24];
assign kernel_img_mul_314[0] = buffer_data_4[2503:2496] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_314[1] = buffer_data_4[2511:2504] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_314[2] = buffer_data_4[2519:2512] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_314[3] = buffer_data_4[2527:2520] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_314[4] = buffer_data_4[2535:2528] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_314[5] = buffer_data_3[2503:2496] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_314[6] = buffer_data_3[2511:2504] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_314[7] = buffer_data_3[2519:2512] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_314[8] = buffer_data_3[2527:2520] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_314[9] = buffer_data_3[2535:2528] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_314[10] = buffer_data_2[2503:2496] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_314[11] = buffer_data_2[2511:2504] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_314[12] = buffer_data_2[2519:2512] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_314[13] = buffer_data_2[2527:2520] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_314[14] = buffer_data_2[2535:2528] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_314[15] = buffer_data_1[2503:2496] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_314[16] = buffer_data_1[2511:2504] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_314[17] = buffer_data_1[2519:2512] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_314[18] = buffer_data_1[2527:2520] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_314[19] = buffer_data_1[2535:2528] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_314[20] = buffer_data_0[2503:2496] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_314[21] = buffer_data_0[2511:2504] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_314[22] = buffer_data_0[2519:2512] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_314[23] = buffer_data_0[2527:2520] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_314[24] = buffer_data_0[2535:2528] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_314 = kernel_img_mul_314[0] + kernel_img_mul_314[1] + kernel_img_mul_314[2] + 
                kernel_img_mul_314[3] + kernel_img_mul_314[4] + kernel_img_mul_314[5] + 
                kernel_img_mul_314[6] + kernel_img_mul_314[7] + kernel_img_mul_314[8] + 
                kernel_img_mul_314[9] + kernel_img_mul_314[10] + kernel_img_mul_314[11] + 
                kernel_img_mul_314[12] + kernel_img_mul_314[13] + kernel_img_mul_314[14] + 
                kernel_img_mul_314[15] + kernel_img_mul_314[16] + kernel_img_mul_314[17] + 
                kernel_img_mul_314[18] + kernel_img_mul_314[19] + kernel_img_mul_314[20] + 
                kernel_img_mul_314[21] + kernel_img_mul_314[22] + kernel_img_mul_314[23] + 
                kernel_img_mul_314[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2519:2512] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2519:2512] <= kernel_img_sum_314[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2519:2512] <= 'd0;
end

wire  [39:0]  kernel_img_mul_315[0:24];
assign kernel_img_mul_315[0] = buffer_data_4[2511:2504] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_315[1] = buffer_data_4[2519:2512] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_315[2] = buffer_data_4[2527:2520] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_315[3] = buffer_data_4[2535:2528] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_315[4] = buffer_data_4[2543:2536] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_315[5] = buffer_data_3[2511:2504] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_315[6] = buffer_data_3[2519:2512] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_315[7] = buffer_data_3[2527:2520] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_315[8] = buffer_data_3[2535:2528] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_315[9] = buffer_data_3[2543:2536] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_315[10] = buffer_data_2[2511:2504] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_315[11] = buffer_data_2[2519:2512] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_315[12] = buffer_data_2[2527:2520] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_315[13] = buffer_data_2[2535:2528] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_315[14] = buffer_data_2[2543:2536] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_315[15] = buffer_data_1[2511:2504] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_315[16] = buffer_data_1[2519:2512] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_315[17] = buffer_data_1[2527:2520] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_315[18] = buffer_data_1[2535:2528] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_315[19] = buffer_data_1[2543:2536] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_315[20] = buffer_data_0[2511:2504] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_315[21] = buffer_data_0[2519:2512] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_315[22] = buffer_data_0[2527:2520] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_315[23] = buffer_data_0[2535:2528] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_315[24] = buffer_data_0[2543:2536] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_315 = kernel_img_mul_315[0] + kernel_img_mul_315[1] + kernel_img_mul_315[2] + 
                kernel_img_mul_315[3] + kernel_img_mul_315[4] + kernel_img_mul_315[5] + 
                kernel_img_mul_315[6] + kernel_img_mul_315[7] + kernel_img_mul_315[8] + 
                kernel_img_mul_315[9] + kernel_img_mul_315[10] + kernel_img_mul_315[11] + 
                kernel_img_mul_315[12] + kernel_img_mul_315[13] + kernel_img_mul_315[14] + 
                kernel_img_mul_315[15] + kernel_img_mul_315[16] + kernel_img_mul_315[17] + 
                kernel_img_mul_315[18] + kernel_img_mul_315[19] + kernel_img_mul_315[20] + 
                kernel_img_mul_315[21] + kernel_img_mul_315[22] + kernel_img_mul_315[23] + 
                kernel_img_mul_315[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2527:2520] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2527:2520] <= kernel_img_sum_315[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2527:2520] <= 'd0;
end

wire  [39:0]  kernel_img_mul_316[0:24];
assign kernel_img_mul_316[0] = buffer_data_4[2519:2512] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_316[1] = buffer_data_4[2527:2520] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_316[2] = buffer_data_4[2535:2528] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_316[3] = buffer_data_4[2543:2536] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_316[4] = buffer_data_4[2551:2544] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_316[5] = buffer_data_3[2519:2512] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_316[6] = buffer_data_3[2527:2520] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_316[7] = buffer_data_3[2535:2528] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_316[8] = buffer_data_3[2543:2536] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_316[9] = buffer_data_3[2551:2544] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_316[10] = buffer_data_2[2519:2512] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_316[11] = buffer_data_2[2527:2520] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_316[12] = buffer_data_2[2535:2528] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_316[13] = buffer_data_2[2543:2536] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_316[14] = buffer_data_2[2551:2544] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_316[15] = buffer_data_1[2519:2512] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_316[16] = buffer_data_1[2527:2520] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_316[17] = buffer_data_1[2535:2528] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_316[18] = buffer_data_1[2543:2536] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_316[19] = buffer_data_1[2551:2544] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_316[20] = buffer_data_0[2519:2512] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_316[21] = buffer_data_0[2527:2520] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_316[22] = buffer_data_0[2535:2528] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_316[23] = buffer_data_0[2543:2536] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_316[24] = buffer_data_0[2551:2544] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_316 = kernel_img_mul_316[0] + kernel_img_mul_316[1] + kernel_img_mul_316[2] + 
                kernel_img_mul_316[3] + kernel_img_mul_316[4] + kernel_img_mul_316[5] + 
                kernel_img_mul_316[6] + kernel_img_mul_316[7] + kernel_img_mul_316[8] + 
                kernel_img_mul_316[9] + kernel_img_mul_316[10] + kernel_img_mul_316[11] + 
                kernel_img_mul_316[12] + kernel_img_mul_316[13] + kernel_img_mul_316[14] + 
                kernel_img_mul_316[15] + kernel_img_mul_316[16] + kernel_img_mul_316[17] + 
                kernel_img_mul_316[18] + kernel_img_mul_316[19] + kernel_img_mul_316[20] + 
                kernel_img_mul_316[21] + kernel_img_mul_316[22] + kernel_img_mul_316[23] + 
                kernel_img_mul_316[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2535:2528] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2535:2528] <= kernel_img_sum_316[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2535:2528] <= 'd0;
end

wire  [39:0]  kernel_img_mul_317[0:24];
assign kernel_img_mul_317[0] = buffer_data_4[2527:2520] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_317[1] = buffer_data_4[2535:2528] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_317[2] = buffer_data_4[2543:2536] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_317[3] = buffer_data_4[2551:2544] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_317[4] = buffer_data_4[2559:2552] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_317[5] = buffer_data_3[2527:2520] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_317[6] = buffer_data_3[2535:2528] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_317[7] = buffer_data_3[2543:2536] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_317[8] = buffer_data_3[2551:2544] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_317[9] = buffer_data_3[2559:2552] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_317[10] = buffer_data_2[2527:2520] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_317[11] = buffer_data_2[2535:2528] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_317[12] = buffer_data_2[2543:2536] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_317[13] = buffer_data_2[2551:2544] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_317[14] = buffer_data_2[2559:2552] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_317[15] = buffer_data_1[2527:2520] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_317[16] = buffer_data_1[2535:2528] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_317[17] = buffer_data_1[2543:2536] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_317[18] = buffer_data_1[2551:2544] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_317[19] = buffer_data_1[2559:2552] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_317[20] = buffer_data_0[2527:2520] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_317[21] = buffer_data_0[2535:2528] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_317[22] = buffer_data_0[2543:2536] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_317[23] = buffer_data_0[2551:2544] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_317[24] = buffer_data_0[2559:2552] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_317 = kernel_img_mul_317[0] + kernel_img_mul_317[1] + kernel_img_mul_317[2] + 
                kernel_img_mul_317[3] + kernel_img_mul_317[4] + kernel_img_mul_317[5] + 
                kernel_img_mul_317[6] + kernel_img_mul_317[7] + kernel_img_mul_317[8] + 
                kernel_img_mul_317[9] + kernel_img_mul_317[10] + kernel_img_mul_317[11] + 
                kernel_img_mul_317[12] + kernel_img_mul_317[13] + kernel_img_mul_317[14] + 
                kernel_img_mul_317[15] + kernel_img_mul_317[16] + kernel_img_mul_317[17] + 
                kernel_img_mul_317[18] + kernel_img_mul_317[19] + kernel_img_mul_317[20] + 
                kernel_img_mul_317[21] + kernel_img_mul_317[22] + kernel_img_mul_317[23] + 
                kernel_img_mul_317[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2543:2536] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2543:2536] <= kernel_img_sum_317[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2543:2536] <= 'd0;
end

wire  [39:0]  kernel_img_mul_318[0:24];
assign kernel_img_mul_318[0] = buffer_data_4[2535:2528] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_318[1] = buffer_data_4[2543:2536] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_318[2] = buffer_data_4[2551:2544] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_318[3] = buffer_data_4[2559:2552] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_318[4] = buffer_data_4[2567:2560] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_318[5] = buffer_data_3[2535:2528] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_318[6] = buffer_data_3[2543:2536] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_318[7] = buffer_data_3[2551:2544] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_318[8] = buffer_data_3[2559:2552] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_318[9] = buffer_data_3[2567:2560] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_318[10] = buffer_data_2[2535:2528] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_318[11] = buffer_data_2[2543:2536] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_318[12] = buffer_data_2[2551:2544] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_318[13] = buffer_data_2[2559:2552] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_318[14] = buffer_data_2[2567:2560] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_318[15] = buffer_data_1[2535:2528] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_318[16] = buffer_data_1[2543:2536] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_318[17] = buffer_data_1[2551:2544] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_318[18] = buffer_data_1[2559:2552] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_318[19] = buffer_data_1[2567:2560] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_318[20] = buffer_data_0[2535:2528] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_318[21] = buffer_data_0[2543:2536] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_318[22] = buffer_data_0[2551:2544] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_318[23] = buffer_data_0[2559:2552] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_318[24] = buffer_data_0[2567:2560] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_318 = kernel_img_mul_318[0] + kernel_img_mul_318[1] + kernel_img_mul_318[2] + 
                kernel_img_mul_318[3] + kernel_img_mul_318[4] + kernel_img_mul_318[5] + 
                kernel_img_mul_318[6] + kernel_img_mul_318[7] + kernel_img_mul_318[8] + 
                kernel_img_mul_318[9] + kernel_img_mul_318[10] + kernel_img_mul_318[11] + 
                kernel_img_mul_318[12] + kernel_img_mul_318[13] + kernel_img_mul_318[14] + 
                kernel_img_mul_318[15] + kernel_img_mul_318[16] + kernel_img_mul_318[17] + 
                kernel_img_mul_318[18] + kernel_img_mul_318[19] + kernel_img_mul_318[20] + 
                kernel_img_mul_318[21] + kernel_img_mul_318[22] + kernel_img_mul_318[23] + 
                kernel_img_mul_318[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2551:2544] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2551:2544] <= kernel_img_sum_318[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2551:2544] <= 'd0;
end

wire  [39:0]  kernel_img_mul_319[0:24];
assign kernel_img_mul_319[0] = buffer_data_4[2543:2536] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_319[1] = buffer_data_4[2551:2544] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_319[2] = buffer_data_4[2559:2552] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_319[3] = buffer_data_4[2567:2560] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_319[4] = buffer_data_4[2575:2568] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_319[5] = buffer_data_3[2543:2536] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_319[6] = buffer_data_3[2551:2544] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_319[7] = buffer_data_3[2559:2552] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_319[8] = buffer_data_3[2567:2560] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_319[9] = buffer_data_3[2575:2568] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_319[10] = buffer_data_2[2543:2536] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_319[11] = buffer_data_2[2551:2544] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_319[12] = buffer_data_2[2559:2552] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_319[13] = buffer_data_2[2567:2560] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_319[14] = buffer_data_2[2575:2568] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_319[15] = buffer_data_1[2543:2536] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_319[16] = buffer_data_1[2551:2544] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_319[17] = buffer_data_1[2559:2552] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_319[18] = buffer_data_1[2567:2560] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_319[19] = buffer_data_1[2575:2568] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_319[20] = buffer_data_0[2543:2536] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_319[21] = buffer_data_0[2551:2544] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_319[22] = buffer_data_0[2559:2552] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_319[23] = buffer_data_0[2567:2560] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_319[24] = buffer_data_0[2575:2568] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_319 = kernel_img_mul_319[0] + kernel_img_mul_319[1] + kernel_img_mul_319[2] + 
                kernel_img_mul_319[3] + kernel_img_mul_319[4] + kernel_img_mul_319[5] + 
                kernel_img_mul_319[6] + kernel_img_mul_319[7] + kernel_img_mul_319[8] + 
                kernel_img_mul_319[9] + kernel_img_mul_319[10] + kernel_img_mul_319[11] + 
                kernel_img_mul_319[12] + kernel_img_mul_319[13] + kernel_img_mul_319[14] + 
                kernel_img_mul_319[15] + kernel_img_mul_319[16] + kernel_img_mul_319[17] + 
                kernel_img_mul_319[18] + kernel_img_mul_319[19] + kernel_img_mul_319[20] + 
                kernel_img_mul_319[21] + kernel_img_mul_319[22] + kernel_img_mul_319[23] + 
                kernel_img_mul_319[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2559:2552] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2559:2552] <= kernel_img_sum_319[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2559:2552] <= 'd0;
end

wire  [39:0]  kernel_img_mul_320[0:24];
assign kernel_img_mul_320[0] = buffer_data_4[2551:2544] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_320[1] = buffer_data_4[2559:2552] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_320[2] = buffer_data_4[2567:2560] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_320[3] = buffer_data_4[2575:2568] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_320[4] = buffer_data_4[2583:2576] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_320[5] = buffer_data_3[2551:2544] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_320[6] = buffer_data_3[2559:2552] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_320[7] = buffer_data_3[2567:2560] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_320[8] = buffer_data_3[2575:2568] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_320[9] = buffer_data_3[2583:2576] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_320[10] = buffer_data_2[2551:2544] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_320[11] = buffer_data_2[2559:2552] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_320[12] = buffer_data_2[2567:2560] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_320[13] = buffer_data_2[2575:2568] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_320[14] = buffer_data_2[2583:2576] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_320[15] = buffer_data_1[2551:2544] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_320[16] = buffer_data_1[2559:2552] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_320[17] = buffer_data_1[2567:2560] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_320[18] = buffer_data_1[2575:2568] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_320[19] = buffer_data_1[2583:2576] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_320[20] = buffer_data_0[2551:2544] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_320[21] = buffer_data_0[2559:2552] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_320[22] = buffer_data_0[2567:2560] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_320[23] = buffer_data_0[2575:2568] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_320[24] = buffer_data_0[2583:2576] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_320 = kernel_img_mul_320[0] + kernel_img_mul_320[1] + kernel_img_mul_320[2] + 
                kernel_img_mul_320[3] + kernel_img_mul_320[4] + kernel_img_mul_320[5] + 
                kernel_img_mul_320[6] + kernel_img_mul_320[7] + kernel_img_mul_320[8] + 
                kernel_img_mul_320[9] + kernel_img_mul_320[10] + kernel_img_mul_320[11] + 
                kernel_img_mul_320[12] + kernel_img_mul_320[13] + kernel_img_mul_320[14] + 
                kernel_img_mul_320[15] + kernel_img_mul_320[16] + kernel_img_mul_320[17] + 
                kernel_img_mul_320[18] + kernel_img_mul_320[19] + kernel_img_mul_320[20] + 
                kernel_img_mul_320[21] + kernel_img_mul_320[22] + kernel_img_mul_320[23] + 
                kernel_img_mul_320[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2567:2560] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2567:2560] <= kernel_img_sum_320[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2567:2560] <= 'd0;
end

wire  [39:0]  kernel_img_mul_321[0:24];
assign kernel_img_mul_321[0] = buffer_data_4[2559:2552] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_321[1] = buffer_data_4[2567:2560] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_321[2] = buffer_data_4[2575:2568] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_321[3] = buffer_data_4[2583:2576] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_321[4] = buffer_data_4[2591:2584] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_321[5] = buffer_data_3[2559:2552] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_321[6] = buffer_data_3[2567:2560] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_321[7] = buffer_data_3[2575:2568] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_321[8] = buffer_data_3[2583:2576] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_321[9] = buffer_data_3[2591:2584] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_321[10] = buffer_data_2[2559:2552] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_321[11] = buffer_data_2[2567:2560] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_321[12] = buffer_data_2[2575:2568] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_321[13] = buffer_data_2[2583:2576] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_321[14] = buffer_data_2[2591:2584] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_321[15] = buffer_data_1[2559:2552] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_321[16] = buffer_data_1[2567:2560] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_321[17] = buffer_data_1[2575:2568] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_321[18] = buffer_data_1[2583:2576] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_321[19] = buffer_data_1[2591:2584] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_321[20] = buffer_data_0[2559:2552] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_321[21] = buffer_data_0[2567:2560] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_321[22] = buffer_data_0[2575:2568] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_321[23] = buffer_data_0[2583:2576] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_321[24] = buffer_data_0[2591:2584] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_321 = kernel_img_mul_321[0] + kernel_img_mul_321[1] + kernel_img_mul_321[2] + 
                kernel_img_mul_321[3] + kernel_img_mul_321[4] + kernel_img_mul_321[5] + 
                kernel_img_mul_321[6] + kernel_img_mul_321[7] + kernel_img_mul_321[8] + 
                kernel_img_mul_321[9] + kernel_img_mul_321[10] + kernel_img_mul_321[11] + 
                kernel_img_mul_321[12] + kernel_img_mul_321[13] + kernel_img_mul_321[14] + 
                kernel_img_mul_321[15] + kernel_img_mul_321[16] + kernel_img_mul_321[17] + 
                kernel_img_mul_321[18] + kernel_img_mul_321[19] + kernel_img_mul_321[20] + 
                kernel_img_mul_321[21] + kernel_img_mul_321[22] + kernel_img_mul_321[23] + 
                kernel_img_mul_321[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2575:2568] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2575:2568] <= kernel_img_sum_321[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2575:2568] <= 'd0;
end

wire  [39:0]  kernel_img_mul_322[0:24];
assign kernel_img_mul_322[0] = buffer_data_4[2567:2560] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_322[1] = buffer_data_4[2575:2568] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_322[2] = buffer_data_4[2583:2576] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_322[3] = buffer_data_4[2591:2584] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_322[4] = buffer_data_4[2599:2592] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_322[5] = buffer_data_3[2567:2560] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_322[6] = buffer_data_3[2575:2568] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_322[7] = buffer_data_3[2583:2576] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_322[8] = buffer_data_3[2591:2584] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_322[9] = buffer_data_3[2599:2592] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_322[10] = buffer_data_2[2567:2560] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_322[11] = buffer_data_2[2575:2568] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_322[12] = buffer_data_2[2583:2576] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_322[13] = buffer_data_2[2591:2584] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_322[14] = buffer_data_2[2599:2592] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_322[15] = buffer_data_1[2567:2560] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_322[16] = buffer_data_1[2575:2568] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_322[17] = buffer_data_1[2583:2576] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_322[18] = buffer_data_1[2591:2584] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_322[19] = buffer_data_1[2599:2592] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_322[20] = buffer_data_0[2567:2560] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_322[21] = buffer_data_0[2575:2568] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_322[22] = buffer_data_0[2583:2576] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_322[23] = buffer_data_0[2591:2584] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_322[24] = buffer_data_0[2599:2592] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_322 = kernel_img_mul_322[0] + kernel_img_mul_322[1] + kernel_img_mul_322[2] + 
                kernel_img_mul_322[3] + kernel_img_mul_322[4] + kernel_img_mul_322[5] + 
                kernel_img_mul_322[6] + kernel_img_mul_322[7] + kernel_img_mul_322[8] + 
                kernel_img_mul_322[9] + kernel_img_mul_322[10] + kernel_img_mul_322[11] + 
                kernel_img_mul_322[12] + kernel_img_mul_322[13] + kernel_img_mul_322[14] + 
                kernel_img_mul_322[15] + kernel_img_mul_322[16] + kernel_img_mul_322[17] + 
                kernel_img_mul_322[18] + kernel_img_mul_322[19] + kernel_img_mul_322[20] + 
                kernel_img_mul_322[21] + kernel_img_mul_322[22] + kernel_img_mul_322[23] + 
                kernel_img_mul_322[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2583:2576] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2583:2576] <= kernel_img_sum_322[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2583:2576] <= 'd0;
end

wire  [39:0]  kernel_img_mul_323[0:24];
assign kernel_img_mul_323[0] = buffer_data_4[2575:2568] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_323[1] = buffer_data_4[2583:2576] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_323[2] = buffer_data_4[2591:2584] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_323[3] = buffer_data_4[2599:2592] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_323[4] = buffer_data_4[2607:2600] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_323[5] = buffer_data_3[2575:2568] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_323[6] = buffer_data_3[2583:2576] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_323[7] = buffer_data_3[2591:2584] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_323[8] = buffer_data_3[2599:2592] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_323[9] = buffer_data_3[2607:2600] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_323[10] = buffer_data_2[2575:2568] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_323[11] = buffer_data_2[2583:2576] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_323[12] = buffer_data_2[2591:2584] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_323[13] = buffer_data_2[2599:2592] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_323[14] = buffer_data_2[2607:2600] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_323[15] = buffer_data_1[2575:2568] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_323[16] = buffer_data_1[2583:2576] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_323[17] = buffer_data_1[2591:2584] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_323[18] = buffer_data_1[2599:2592] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_323[19] = buffer_data_1[2607:2600] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_323[20] = buffer_data_0[2575:2568] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_323[21] = buffer_data_0[2583:2576] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_323[22] = buffer_data_0[2591:2584] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_323[23] = buffer_data_0[2599:2592] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_323[24] = buffer_data_0[2607:2600] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_323 = kernel_img_mul_323[0] + kernel_img_mul_323[1] + kernel_img_mul_323[2] + 
                kernel_img_mul_323[3] + kernel_img_mul_323[4] + kernel_img_mul_323[5] + 
                kernel_img_mul_323[6] + kernel_img_mul_323[7] + kernel_img_mul_323[8] + 
                kernel_img_mul_323[9] + kernel_img_mul_323[10] + kernel_img_mul_323[11] + 
                kernel_img_mul_323[12] + kernel_img_mul_323[13] + kernel_img_mul_323[14] + 
                kernel_img_mul_323[15] + kernel_img_mul_323[16] + kernel_img_mul_323[17] + 
                kernel_img_mul_323[18] + kernel_img_mul_323[19] + kernel_img_mul_323[20] + 
                kernel_img_mul_323[21] + kernel_img_mul_323[22] + kernel_img_mul_323[23] + 
                kernel_img_mul_323[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2591:2584] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2591:2584] <= kernel_img_sum_323[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2591:2584] <= 'd0;
end

wire  [39:0]  kernel_img_mul_324[0:24];
assign kernel_img_mul_324[0] = buffer_data_4[2583:2576] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_324[1] = buffer_data_4[2591:2584] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_324[2] = buffer_data_4[2599:2592] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_324[3] = buffer_data_4[2607:2600] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_324[4] = buffer_data_4[2615:2608] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_324[5] = buffer_data_3[2583:2576] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_324[6] = buffer_data_3[2591:2584] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_324[7] = buffer_data_3[2599:2592] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_324[8] = buffer_data_3[2607:2600] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_324[9] = buffer_data_3[2615:2608] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_324[10] = buffer_data_2[2583:2576] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_324[11] = buffer_data_2[2591:2584] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_324[12] = buffer_data_2[2599:2592] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_324[13] = buffer_data_2[2607:2600] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_324[14] = buffer_data_2[2615:2608] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_324[15] = buffer_data_1[2583:2576] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_324[16] = buffer_data_1[2591:2584] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_324[17] = buffer_data_1[2599:2592] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_324[18] = buffer_data_1[2607:2600] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_324[19] = buffer_data_1[2615:2608] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_324[20] = buffer_data_0[2583:2576] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_324[21] = buffer_data_0[2591:2584] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_324[22] = buffer_data_0[2599:2592] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_324[23] = buffer_data_0[2607:2600] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_324[24] = buffer_data_0[2615:2608] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_324 = kernel_img_mul_324[0] + kernel_img_mul_324[1] + kernel_img_mul_324[2] + 
                kernel_img_mul_324[3] + kernel_img_mul_324[4] + kernel_img_mul_324[5] + 
                kernel_img_mul_324[6] + kernel_img_mul_324[7] + kernel_img_mul_324[8] + 
                kernel_img_mul_324[9] + kernel_img_mul_324[10] + kernel_img_mul_324[11] + 
                kernel_img_mul_324[12] + kernel_img_mul_324[13] + kernel_img_mul_324[14] + 
                kernel_img_mul_324[15] + kernel_img_mul_324[16] + kernel_img_mul_324[17] + 
                kernel_img_mul_324[18] + kernel_img_mul_324[19] + kernel_img_mul_324[20] + 
                kernel_img_mul_324[21] + kernel_img_mul_324[22] + kernel_img_mul_324[23] + 
                kernel_img_mul_324[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2599:2592] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2599:2592] <= kernel_img_sum_324[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2599:2592] <= 'd0;
end

wire  [39:0]  kernel_img_mul_325[0:24];
assign kernel_img_mul_325[0] = buffer_data_4[2591:2584] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_325[1] = buffer_data_4[2599:2592] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_325[2] = buffer_data_4[2607:2600] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_325[3] = buffer_data_4[2615:2608] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_325[4] = buffer_data_4[2623:2616] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_325[5] = buffer_data_3[2591:2584] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_325[6] = buffer_data_3[2599:2592] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_325[7] = buffer_data_3[2607:2600] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_325[8] = buffer_data_3[2615:2608] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_325[9] = buffer_data_3[2623:2616] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_325[10] = buffer_data_2[2591:2584] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_325[11] = buffer_data_2[2599:2592] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_325[12] = buffer_data_2[2607:2600] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_325[13] = buffer_data_2[2615:2608] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_325[14] = buffer_data_2[2623:2616] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_325[15] = buffer_data_1[2591:2584] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_325[16] = buffer_data_1[2599:2592] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_325[17] = buffer_data_1[2607:2600] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_325[18] = buffer_data_1[2615:2608] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_325[19] = buffer_data_1[2623:2616] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_325[20] = buffer_data_0[2591:2584] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_325[21] = buffer_data_0[2599:2592] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_325[22] = buffer_data_0[2607:2600] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_325[23] = buffer_data_0[2615:2608] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_325[24] = buffer_data_0[2623:2616] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_325 = kernel_img_mul_325[0] + kernel_img_mul_325[1] + kernel_img_mul_325[2] + 
                kernel_img_mul_325[3] + kernel_img_mul_325[4] + kernel_img_mul_325[5] + 
                kernel_img_mul_325[6] + kernel_img_mul_325[7] + kernel_img_mul_325[8] + 
                kernel_img_mul_325[9] + kernel_img_mul_325[10] + kernel_img_mul_325[11] + 
                kernel_img_mul_325[12] + kernel_img_mul_325[13] + kernel_img_mul_325[14] + 
                kernel_img_mul_325[15] + kernel_img_mul_325[16] + kernel_img_mul_325[17] + 
                kernel_img_mul_325[18] + kernel_img_mul_325[19] + kernel_img_mul_325[20] + 
                kernel_img_mul_325[21] + kernel_img_mul_325[22] + kernel_img_mul_325[23] + 
                kernel_img_mul_325[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2607:2600] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2607:2600] <= kernel_img_sum_325[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2607:2600] <= 'd0;
end

wire  [39:0]  kernel_img_mul_326[0:24];
assign kernel_img_mul_326[0] = buffer_data_4[2599:2592] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_326[1] = buffer_data_4[2607:2600] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_326[2] = buffer_data_4[2615:2608] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_326[3] = buffer_data_4[2623:2616] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_326[4] = buffer_data_4[2631:2624] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_326[5] = buffer_data_3[2599:2592] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_326[6] = buffer_data_3[2607:2600] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_326[7] = buffer_data_3[2615:2608] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_326[8] = buffer_data_3[2623:2616] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_326[9] = buffer_data_3[2631:2624] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_326[10] = buffer_data_2[2599:2592] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_326[11] = buffer_data_2[2607:2600] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_326[12] = buffer_data_2[2615:2608] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_326[13] = buffer_data_2[2623:2616] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_326[14] = buffer_data_2[2631:2624] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_326[15] = buffer_data_1[2599:2592] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_326[16] = buffer_data_1[2607:2600] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_326[17] = buffer_data_1[2615:2608] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_326[18] = buffer_data_1[2623:2616] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_326[19] = buffer_data_1[2631:2624] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_326[20] = buffer_data_0[2599:2592] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_326[21] = buffer_data_0[2607:2600] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_326[22] = buffer_data_0[2615:2608] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_326[23] = buffer_data_0[2623:2616] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_326[24] = buffer_data_0[2631:2624] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_326 = kernel_img_mul_326[0] + kernel_img_mul_326[1] + kernel_img_mul_326[2] + 
                kernel_img_mul_326[3] + kernel_img_mul_326[4] + kernel_img_mul_326[5] + 
                kernel_img_mul_326[6] + kernel_img_mul_326[7] + kernel_img_mul_326[8] + 
                kernel_img_mul_326[9] + kernel_img_mul_326[10] + kernel_img_mul_326[11] + 
                kernel_img_mul_326[12] + kernel_img_mul_326[13] + kernel_img_mul_326[14] + 
                kernel_img_mul_326[15] + kernel_img_mul_326[16] + kernel_img_mul_326[17] + 
                kernel_img_mul_326[18] + kernel_img_mul_326[19] + kernel_img_mul_326[20] + 
                kernel_img_mul_326[21] + kernel_img_mul_326[22] + kernel_img_mul_326[23] + 
                kernel_img_mul_326[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2615:2608] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2615:2608] <= kernel_img_sum_326[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2615:2608] <= 'd0;
end

wire  [39:0]  kernel_img_mul_327[0:24];
assign kernel_img_mul_327[0] = buffer_data_4[2607:2600] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_327[1] = buffer_data_4[2615:2608] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_327[2] = buffer_data_4[2623:2616] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_327[3] = buffer_data_4[2631:2624] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_327[4] = buffer_data_4[2639:2632] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_327[5] = buffer_data_3[2607:2600] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_327[6] = buffer_data_3[2615:2608] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_327[7] = buffer_data_3[2623:2616] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_327[8] = buffer_data_3[2631:2624] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_327[9] = buffer_data_3[2639:2632] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_327[10] = buffer_data_2[2607:2600] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_327[11] = buffer_data_2[2615:2608] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_327[12] = buffer_data_2[2623:2616] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_327[13] = buffer_data_2[2631:2624] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_327[14] = buffer_data_2[2639:2632] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_327[15] = buffer_data_1[2607:2600] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_327[16] = buffer_data_1[2615:2608] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_327[17] = buffer_data_1[2623:2616] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_327[18] = buffer_data_1[2631:2624] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_327[19] = buffer_data_1[2639:2632] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_327[20] = buffer_data_0[2607:2600] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_327[21] = buffer_data_0[2615:2608] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_327[22] = buffer_data_0[2623:2616] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_327[23] = buffer_data_0[2631:2624] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_327[24] = buffer_data_0[2639:2632] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_327 = kernel_img_mul_327[0] + kernel_img_mul_327[1] + kernel_img_mul_327[2] + 
                kernel_img_mul_327[3] + kernel_img_mul_327[4] + kernel_img_mul_327[5] + 
                kernel_img_mul_327[6] + kernel_img_mul_327[7] + kernel_img_mul_327[8] + 
                kernel_img_mul_327[9] + kernel_img_mul_327[10] + kernel_img_mul_327[11] + 
                kernel_img_mul_327[12] + kernel_img_mul_327[13] + kernel_img_mul_327[14] + 
                kernel_img_mul_327[15] + kernel_img_mul_327[16] + kernel_img_mul_327[17] + 
                kernel_img_mul_327[18] + kernel_img_mul_327[19] + kernel_img_mul_327[20] + 
                kernel_img_mul_327[21] + kernel_img_mul_327[22] + kernel_img_mul_327[23] + 
                kernel_img_mul_327[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2623:2616] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2623:2616] <= kernel_img_sum_327[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2623:2616] <= 'd0;
end

wire  [39:0]  kernel_img_mul_328[0:24];
assign kernel_img_mul_328[0] = buffer_data_4[2615:2608] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_328[1] = buffer_data_4[2623:2616] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_328[2] = buffer_data_4[2631:2624] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_328[3] = buffer_data_4[2639:2632] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_328[4] = buffer_data_4[2647:2640] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_328[5] = buffer_data_3[2615:2608] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_328[6] = buffer_data_3[2623:2616] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_328[7] = buffer_data_3[2631:2624] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_328[8] = buffer_data_3[2639:2632] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_328[9] = buffer_data_3[2647:2640] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_328[10] = buffer_data_2[2615:2608] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_328[11] = buffer_data_2[2623:2616] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_328[12] = buffer_data_2[2631:2624] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_328[13] = buffer_data_2[2639:2632] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_328[14] = buffer_data_2[2647:2640] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_328[15] = buffer_data_1[2615:2608] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_328[16] = buffer_data_1[2623:2616] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_328[17] = buffer_data_1[2631:2624] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_328[18] = buffer_data_1[2639:2632] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_328[19] = buffer_data_1[2647:2640] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_328[20] = buffer_data_0[2615:2608] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_328[21] = buffer_data_0[2623:2616] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_328[22] = buffer_data_0[2631:2624] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_328[23] = buffer_data_0[2639:2632] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_328[24] = buffer_data_0[2647:2640] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_328 = kernel_img_mul_328[0] + kernel_img_mul_328[1] + kernel_img_mul_328[2] + 
                kernel_img_mul_328[3] + kernel_img_mul_328[4] + kernel_img_mul_328[5] + 
                kernel_img_mul_328[6] + kernel_img_mul_328[7] + kernel_img_mul_328[8] + 
                kernel_img_mul_328[9] + kernel_img_mul_328[10] + kernel_img_mul_328[11] + 
                kernel_img_mul_328[12] + kernel_img_mul_328[13] + kernel_img_mul_328[14] + 
                kernel_img_mul_328[15] + kernel_img_mul_328[16] + kernel_img_mul_328[17] + 
                kernel_img_mul_328[18] + kernel_img_mul_328[19] + kernel_img_mul_328[20] + 
                kernel_img_mul_328[21] + kernel_img_mul_328[22] + kernel_img_mul_328[23] + 
                kernel_img_mul_328[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2631:2624] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2631:2624] <= kernel_img_sum_328[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2631:2624] <= 'd0;
end

wire  [39:0]  kernel_img_mul_329[0:24];
assign kernel_img_mul_329[0] = buffer_data_4[2623:2616] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_329[1] = buffer_data_4[2631:2624] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_329[2] = buffer_data_4[2639:2632] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_329[3] = buffer_data_4[2647:2640] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_329[4] = buffer_data_4[2655:2648] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_329[5] = buffer_data_3[2623:2616] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_329[6] = buffer_data_3[2631:2624] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_329[7] = buffer_data_3[2639:2632] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_329[8] = buffer_data_3[2647:2640] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_329[9] = buffer_data_3[2655:2648] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_329[10] = buffer_data_2[2623:2616] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_329[11] = buffer_data_2[2631:2624] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_329[12] = buffer_data_2[2639:2632] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_329[13] = buffer_data_2[2647:2640] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_329[14] = buffer_data_2[2655:2648] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_329[15] = buffer_data_1[2623:2616] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_329[16] = buffer_data_1[2631:2624] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_329[17] = buffer_data_1[2639:2632] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_329[18] = buffer_data_1[2647:2640] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_329[19] = buffer_data_1[2655:2648] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_329[20] = buffer_data_0[2623:2616] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_329[21] = buffer_data_0[2631:2624] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_329[22] = buffer_data_0[2639:2632] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_329[23] = buffer_data_0[2647:2640] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_329[24] = buffer_data_0[2655:2648] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_329 = kernel_img_mul_329[0] + kernel_img_mul_329[1] + kernel_img_mul_329[2] + 
                kernel_img_mul_329[3] + kernel_img_mul_329[4] + kernel_img_mul_329[5] + 
                kernel_img_mul_329[6] + kernel_img_mul_329[7] + kernel_img_mul_329[8] + 
                kernel_img_mul_329[9] + kernel_img_mul_329[10] + kernel_img_mul_329[11] + 
                kernel_img_mul_329[12] + kernel_img_mul_329[13] + kernel_img_mul_329[14] + 
                kernel_img_mul_329[15] + kernel_img_mul_329[16] + kernel_img_mul_329[17] + 
                kernel_img_mul_329[18] + kernel_img_mul_329[19] + kernel_img_mul_329[20] + 
                kernel_img_mul_329[21] + kernel_img_mul_329[22] + kernel_img_mul_329[23] + 
                kernel_img_mul_329[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2639:2632] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2639:2632] <= kernel_img_sum_329[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2639:2632] <= 'd0;
end

wire  [39:0]  kernel_img_mul_330[0:24];
assign kernel_img_mul_330[0] = buffer_data_4[2631:2624] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_330[1] = buffer_data_4[2639:2632] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_330[2] = buffer_data_4[2647:2640] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_330[3] = buffer_data_4[2655:2648] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_330[4] = buffer_data_4[2663:2656] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_330[5] = buffer_data_3[2631:2624] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_330[6] = buffer_data_3[2639:2632] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_330[7] = buffer_data_3[2647:2640] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_330[8] = buffer_data_3[2655:2648] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_330[9] = buffer_data_3[2663:2656] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_330[10] = buffer_data_2[2631:2624] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_330[11] = buffer_data_2[2639:2632] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_330[12] = buffer_data_2[2647:2640] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_330[13] = buffer_data_2[2655:2648] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_330[14] = buffer_data_2[2663:2656] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_330[15] = buffer_data_1[2631:2624] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_330[16] = buffer_data_1[2639:2632] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_330[17] = buffer_data_1[2647:2640] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_330[18] = buffer_data_1[2655:2648] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_330[19] = buffer_data_1[2663:2656] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_330[20] = buffer_data_0[2631:2624] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_330[21] = buffer_data_0[2639:2632] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_330[22] = buffer_data_0[2647:2640] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_330[23] = buffer_data_0[2655:2648] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_330[24] = buffer_data_0[2663:2656] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_330 = kernel_img_mul_330[0] + kernel_img_mul_330[1] + kernel_img_mul_330[2] + 
                kernel_img_mul_330[3] + kernel_img_mul_330[4] + kernel_img_mul_330[5] + 
                kernel_img_mul_330[6] + kernel_img_mul_330[7] + kernel_img_mul_330[8] + 
                kernel_img_mul_330[9] + kernel_img_mul_330[10] + kernel_img_mul_330[11] + 
                kernel_img_mul_330[12] + kernel_img_mul_330[13] + kernel_img_mul_330[14] + 
                kernel_img_mul_330[15] + kernel_img_mul_330[16] + kernel_img_mul_330[17] + 
                kernel_img_mul_330[18] + kernel_img_mul_330[19] + kernel_img_mul_330[20] + 
                kernel_img_mul_330[21] + kernel_img_mul_330[22] + kernel_img_mul_330[23] + 
                kernel_img_mul_330[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2647:2640] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2647:2640] <= kernel_img_sum_330[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2647:2640] <= 'd0;
end

wire  [39:0]  kernel_img_mul_331[0:24];
assign kernel_img_mul_331[0] = buffer_data_4[2639:2632] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_331[1] = buffer_data_4[2647:2640] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_331[2] = buffer_data_4[2655:2648] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_331[3] = buffer_data_4[2663:2656] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_331[4] = buffer_data_4[2671:2664] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_331[5] = buffer_data_3[2639:2632] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_331[6] = buffer_data_3[2647:2640] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_331[7] = buffer_data_3[2655:2648] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_331[8] = buffer_data_3[2663:2656] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_331[9] = buffer_data_3[2671:2664] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_331[10] = buffer_data_2[2639:2632] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_331[11] = buffer_data_2[2647:2640] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_331[12] = buffer_data_2[2655:2648] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_331[13] = buffer_data_2[2663:2656] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_331[14] = buffer_data_2[2671:2664] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_331[15] = buffer_data_1[2639:2632] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_331[16] = buffer_data_1[2647:2640] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_331[17] = buffer_data_1[2655:2648] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_331[18] = buffer_data_1[2663:2656] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_331[19] = buffer_data_1[2671:2664] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_331[20] = buffer_data_0[2639:2632] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_331[21] = buffer_data_0[2647:2640] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_331[22] = buffer_data_0[2655:2648] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_331[23] = buffer_data_0[2663:2656] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_331[24] = buffer_data_0[2671:2664] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_331 = kernel_img_mul_331[0] + kernel_img_mul_331[1] + kernel_img_mul_331[2] + 
                kernel_img_mul_331[3] + kernel_img_mul_331[4] + kernel_img_mul_331[5] + 
                kernel_img_mul_331[6] + kernel_img_mul_331[7] + kernel_img_mul_331[8] + 
                kernel_img_mul_331[9] + kernel_img_mul_331[10] + kernel_img_mul_331[11] + 
                kernel_img_mul_331[12] + kernel_img_mul_331[13] + kernel_img_mul_331[14] + 
                kernel_img_mul_331[15] + kernel_img_mul_331[16] + kernel_img_mul_331[17] + 
                kernel_img_mul_331[18] + kernel_img_mul_331[19] + kernel_img_mul_331[20] + 
                kernel_img_mul_331[21] + kernel_img_mul_331[22] + kernel_img_mul_331[23] + 
                kernel_img_mul_331[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2655:2648] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2655:2648] <= kernel_img_sum_331[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2655:2648] <= 'd0;
end

wire  [39:0]  kernel_img_mul_332[0:24];
assign kernel_img_mul_332[0] = buffer_data_4[2647:2640] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_332[1] = buffer_data_4[2655:2648] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_332[2] = buffer_data_4[2663:2656] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_332[3] = buffer_data_4[2671:2664] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_332[4] = buffer_data_4[2679:2672] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_332[5] = buffer_data_3[2647:2640] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_332[6] = buffer_data_3[2655:2648] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_332[7] = buffer_data_3[2663:2656] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_332[8] = buffer_data_3[2671:2664] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_332[9] = buffer_data_3[2679:2672] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_332[10] = buffer_data_2[2647:2640] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_332[11] = buffer_data_2[2655:2648] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_332[12] = buffer_data_2[2663:2656] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_332[13] = buffer_data_2[2671:2664] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_332[14] = buffer_data_2[2679:2672] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_332[15] = buffer_data_1[2647:2640] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_332[16] = buffer_data_1[2655:2648] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_332[17] = buffer_data_1[2663:2656] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_332[18] = buffer_data_1[2671:2664] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_332[19] = buffer_data_1[2679:2672] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_332[20] = buffer_data_0[2647:2640] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_332[21] = buffer_data_0[2655:2648] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_332[22] = buffer_data_0[2663:2656] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_332[23] = buffer_data_0[2671:2664] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_332[24] = buffer_data_0[2679:2672] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_332 = kernel_img_mul_332[0] + kernel_img_mul_332[1] + kernel_img_mul_332[2] + 
                kernel_img_mul_332[3] + kernel_img_mul_332[4] + kernel_img_mul_332[5] + 
                kernel_img_mul_332[6] + kernel_img_mul_332[7] + kernel_img_mul_332[8] + 
                kernel_img_mul_332[9] + kernel_img_mul_332[10] + kernel_img_mul_332[11] + 
                kernel_img_mul_332[12] + kernel_img_mul_332[13] + kernel_img_mul_332[14] + 
                kernel_img_mul_332[15] + kernel_img_mul_332[16] + kernel_img_mul_332[17] + 
                kernel_img_mul_332[18] + kernel_img_mul_332[19] + kernel_img_mul_332[20] + 
                kernel_img_mul_332[21] + kernel_img_mul_332[22] + kernel_img_mul_332[23] + 
                kernel_img_mul_332[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2663:2656] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2663:2656] <= kernel_img_sum_332[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2663:2656] <= 'd0;
end

wire  [39:0]  kernel_img_mul_333[0:24];
assign kernel_img_mul_333[0] = buffer_data_4[2655:2648] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_333[1] = buffer_data_4[2663:2656] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_333[2] = buffer_data_4[2671:2664] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_333[3] = buffer_data_4[2679:2672] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_333[4] = buffer_data_4[2687:2680] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_333[5] = buffer_data_3[2655:2648] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_333[6] = buffer_data_3[2663:2656] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_333[7] = buffer_data_3[2671:2664] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_333[8] = buffer_data_3[2679:2672] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_333[9] = buffer_data_3[2687:2680] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_333[10] = buffer_data_2[2655:2648] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_333[11] = buffer_data_2[2663:2656] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_333[12] = buffer_data_2[2671:2664] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_333[13] = buffer_data_2[2679:2672] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_333[14] = buffer_data_2[2687:2680] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_333[15] = buffer_data_1[2655:2648] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_333[16] = buffer_data_1[2663:2656] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_333[17] = buffer_data_1[2671:2664] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_333[18] = buffer_data_1[2679:2672] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_333[19] = buffer_data_1[2687:2680] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_333[20] = buffer_data_0[2655:2648] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_333[21] = buffer_data_0[2663:2656] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_333[22] = buffer_data_0[2671:2664] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_333[23] = buffer_data_0[2679:2672] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_333[24] = buffer_data_0[2687:2680] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_333 = kernel_img_mul_333[0] + kernel_img_mul_333[1] + kernel_img_mul_333[2] + 
                kernel_img_mul_333[3] + kernel_img_mul_333[4] + kernel_img_mul_333[5] + 
                kernel_img_mul_333[6] + kernel_img_mul_333[7] + kernel_img_mul_333[8] + 
                kernel_img_mul_333[9] + kernel_img_mul_333[10] + kernel_img_mul_333[11] + 
                kernel_img_mul_333[12] + kernel_img_mul_333[13] + kernel_img_mul_333[14] + 
                kernel_img_mul_333[15] + kernel_img_mul_333[16] + kernel_img_mul_333[17] + 
                kernel_img_mul_333[18] + kernel_img_mul_333[19] + kernel_img_mul_333[20] + 
                kernel_img_mul_333[21] + kernel_img_mul_333[22] + kernel_img_mul_333[23] + 
                kernel_img_mul_333[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2671:2664] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2671:2664] <= kernel_img_sum_333[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2671:2664] <= 'd0;
end

wire  [39:0]  kernel_img_mul_334[0:24];
assign kernel_img_mul_334[0] = buffer_data_4[2663:2656] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_334[1] = buffer_data_4[2671:2664] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_334[2] = buffer_data_4[2679:2672] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_334[3] = buffer_data_4[2687:2680] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_334[4] = buffer_data_4[2695:2688] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_334[5] = buffer_data_3[2663:2656] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_334[6] = buffer_data_3[2671:2664] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_334[7] = buffer_data_3[2679:2672] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_334[8] = buffer_data_3[2687:2680] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_334[9] = buffer_data_3[2695:2688] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_334[10] = buffer_data_2[2663:2656] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_334[11] = buffer_data_2[2671:2664] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_334[12] = buffer_data_2[2679:2672] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_334[13] = buffer_data_2[2687:2680] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_334[14] = buffer_data_2[2695:2688] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_334[15] = buffer_data_1[2663:2656] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_334[16] = buffer_data_1[2671:2664] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_334[17] = buffer_data_1[2679:2672] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_334[18] = buffer_data_1[2687:2680] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_334[19] = buffer_data_1[2695:2688] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_334[20] = buffer_data_0[2663:2656] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_334[21] = buffer_data_0[2671:2664] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_334[22] = buffer_data_0[2679:2672] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_334[23] = buffer_data_0[2687:2680] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_334[24] = buffer_data_0[2695:2688] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_334 = kernel_img_mul_334[0] + kernel_img_mul_334[1] + kernel_img_mul_334[2] + 
                kernel_img_mul_334[3] + kernel_img_mul_334[4] + kernel_img_mul_334[5] + 
                kernel_img_mul_334[6] + kernel_img_mul_334[7] + kernel_img_mul_334[8] + 
                kernel_img_mul_334[9] + kernel_img_mul_334[10] + kernel_img_mul_334[11] + 
                kernel_img_mul_334[12] + kernel_img_mul_334[13] + kernel_img_mul_334[14] + 
                kernel_img_mul_334[15] + kernel_img_mul_334[16] + kernel_img_mul_334[17] + 
                kernel_img_mul_334[18] + kernel_img_mul_334[19] + kernel_img_mul_334[20] + 
                kernel_img_mul_334[21] + kernel_img_mul_334[22] + kernel_img_mul_334[23] + 
                kernel_img_mul_334[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2679:2672] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2679:2672] <= kernel_img_sum_334[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2679:2672] <= 'd0;
end

wire  [39:0]  kernel_img_mul_335[0:24];
assign kernel_img_mul_335[0] = buffer_data_4[2671:2664] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_335[1] = buffer_data_4[2679:2672] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_335[2] = buffer_data_4[2687:2680] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_335[3] = buffer_data_4[2695:2688] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_335[4] = buffer_data_4[2703:2696] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_335[5] = buffer_data_3[2671:2664] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_335[6] = buffer_data_3[2679:2672] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_335[7] = buffer_data_3[2687:2680] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_335[8] = buffer_data_3[2695:2688] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_335[9] = buffer_data_3[2703:2696] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_335[10] = buffer_data_2[2671:2664] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_335[11] = buffer_data_2[2679:2672] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_335[12] = buffer_data_2[2687:2680] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_335[13] = buffer_data_2[2695:2688] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_335[14] = buffer_data_2[2703:2696] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_335[15] = buffer_data_1[2671:2664] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_335[16] = buffer_data_1[2679:2672] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_335[17] = buffer_data_1[2687:2680] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_335[18] = buffer_data_1[2695:2688] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_335[19] = buffer_data_1[2703:2696] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_335[20] = buffer_data_0[2671:2664] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_335[21] = buffer_data_0[2679:2672] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_335[22] = buffer_data_0[2687:2680] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_335[23] = buffer_data_0[2695:2688] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_335[24] = buffer_data_0[2703:2696] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_335 = kernel_img_mul_335[0] + kernel_img_mul_335[1] + kernel_img_mul_335[2] + 
                kernel_img_mul_335[3] + kernel_img_mul_335[4] + kernel_img_mul_335[5] + 
                kernel_img_mul_335[6] + kernel_img_mul_335[7] + kernel_img_mul_335[8] + 
                kernel_img_mul_335[9] + kernel_img_mul_335[10] + kernel_img_mul_335[11] + 
                kernel_img_mul_335[12] + kernel_img_mul_335[13] + kernel_img_mul_335[14] + 
                kernel_img_mul_335[15] + kernel_img_mul_335[16] + kernel_img_mul_335[17] + 
                kernel_img_mul_335[18] + kernel_img_mul_335[19] + kernel_img_mul_335[20] + 
                kernel_img_mul_335[21] + kernel_img_mul_335[22] + kernel_img_mul_335[23] + 
                kernel_img_mul_335[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2687:2680] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2687:2680] <= kernel_img_sum_335[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2687:2680] <= 'd0;
end

wire  [39:0]  kernel_img_mul_336[0:24];
assign kernel_img_mul_336[0] = buffer_data_4[2679:2672] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_336[1] = buffer_data_4[2687:2680] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_336[2] = buffer_data_4[2695:2688] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_336[3] = buffer_data_4[2703:2696] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_336[4] = buffer_data_4[2711:2704] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_336[5] = buffer_data_3[2679:2672] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_336[6] = buffer_data_3[2687:2680] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_336[7] = buffer_data_3[2695:2688] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_336[8] = buffer_data_3[2703:2696] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_336[9] = buffer_data_3[2711:2704] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_336[10] = buffer_data_2[2679:2672] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_336[11] = buffer_data_2[2687:2680] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_336[12] = buffer_data_2[2695:2688] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_336[13] = buffer_data_2[2703:2696] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_336[14] = buffer_data_2[2711:2704] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_336[15] = buffer_data_1[2679:2672] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_336[16] = buffer_data_1[2687:2680] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_336[17] = buffer_data_1[2695:2688] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_336[18] = buffer_data_1[2703:2696] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_336[19] = buffer_data_1[2711:2704] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_336[20] = buffer_data_0[2679:2672] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_336[21] = buffer_data_0[2687:2680] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_336[22] = buffer_data_0[2695:2688] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_336[23] = buffer_data_0[2703:2696] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_336[24] = buffer_data_0[2711:2704] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_336 = kernel_img_mul_336[0] + kernel_img_mul_336[1] + kernel_img_mul_336[2] + 
                kernel_img_mul_336[3] + kernel_img_mul_336[4] + kernel_img_mul_336[5] + 
                kernel_img_mul_336[6] + kernel_img_mul_336[7] + kernel_img_mul_336[8] + 
                kernel_img_mul_336[9] + kernel_img_mul_336[10] + kernel_img_mul_336[11] + 
                kernel_img_mul_336[12] + kernel_img_mul_336[13] + kernel_img_mul_336[14] + 
                kernel_img_mul_336[15] + kernel_img_mul_336[16] + kernel_img_mul_336[17] + 
                kernel_img_mul_336[18] + kernel_img_mul_336[19] + kernel_img_mul_336[20] + 
                kernel_img_mul_336[21] + kernel_img_mul_336[22] + kernel_img_mul_336[23] + 
                kernel_img_mul_336[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2695:2688] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2695:2688] <= kernel_img_sum_336[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2695:2688] <= 'd0;
end

wire  [39:0]  kernel_img_mul_337[0:24];
assign kernel_img_mul_337[0] = buffer_data_4[2687:2680] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_337[1] = buffer_data_4[2695:2688] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_337[2] = buffer_data_4[2703:2696] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_337[3] = buffer_data_4[2711:2704] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_337[4] = buffer_data_4[2719:2712] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_337[5] = buffer_data_3[2687:2680] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_337[6] = buffer_data_3[2695:2688] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_337[7] = buffer_data_3[2703:2696] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_337[8] = buffer_data_3[2711:2704] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_337[9] = buffer_data_3[2719:2712] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_337[10] = buffer_data_2[2687:2680] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_337[11] = buffer_data_2[2695:2688] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_337[12] = buffer_data_2[2703:2696] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_337[13] = buffer_data_2[2711:2704] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_337[14] = buffer_data_2[2719:2712] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_337[15] = buffer_data_1[2687:2680] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_337[16] = buffer_data_1[2695:2688] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_337[17] = buffer_data_1[2703:2696] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_337[18] = buffer_data_1[2711:2704] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_337[19] = buffer_data_1[2719:2712] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_337[20] = buffer_data_0[2687:2680] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_337[21] = buffer_data_0[2695:2688] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_337[22] = buffer_data_0[2703:2696] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_337[23] = buffer_data_0[2711:2704] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_337[24] = buffer_data_0[2719:2712] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_337 = kernel_img_mul_337[0] + kernel_img_mul_337[1] + kernel_img_mul_337[2] + 
                kernel_img_mul_337[3] + kernel_img_mul_337[4] + kernel_img_mul_337[5] + 
                kernel_img_mul_337[6] + kernel_img_mul_337[7] + kernel_img_mul_337[8] + 
                kernel_img_mul_337[9] + kernel_img_mul_337[10] + kernel_img_mul_337[11] + 
                kernel_img_mul_337[12] + kernel_img_mul_337[13] + kernel_img_mul_337[14] + 
                kernel_img_mul_337[15] + kernel_img_mul_337[16] + kernel_img_mul_337[17] + 
                kernel_img_mul_337[18] + kernel_img_mul_337[19] + kernel_img_mul_337[20] + 
                kernel_img_mul_337[21] + kernel_img_mul_337[22] + kernel_img_mul_337[23] + 
                kernel_img_mul_337[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2703:2696] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2703:2696] <= kernel_img_sum_337[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2703:2696] <= 'd0;
end

wire  [39:0]  kernel_img_mul_338[0:24];
assign kernel_img_mul_338[0] = buffer_data_4[2695:2688] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_338[1] = buffer_data_4[2703:2696] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_338[2] = buffer_data_4[2711:2704] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_338[3] = buffer_data_4[2719:2712] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_338[4] = buffer_data_4[2727:2720] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_338[5] = buffer_data_3[2695:2688] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_338[6] = buffer_data_3[2703:2696] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_338[7] = buffer_data_3[2711:2704] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_338[8] = buffer_data_3[2719:2712] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_338[9] = buffer_data_3[2727:2720] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_338[10] = buffer_data_2[2695:2688] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_338[11] = buffer_data_2[2703:2696] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_338[12] = buffer_data_2[2711:2704] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_338[13] = buffer_data_2[2719:2712] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_338[14] = buffer_data_2[2727:2720] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_338[15] = buffer_data_1[2695:2688] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_338[16] = buffer_data_1[2703:2696] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_338[17] = buffer_data_1[2711:2704] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_338[18] = buffer_data_1[2719:2712] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_338[19] = buffer_data_1[2727:2720] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_338[20] = buffer_data_0[2695:2688] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_338[21] = buffer_data_0[2703:2696] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_338[22] = buffer_data_0[2711:2704] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_338[23] = buffer_data_0[2719:2712] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_338[24] = buffer_data_0[2727:2720] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_338 = kernel_img_mul_338[0] + kernel_img_mul_338[1] + kernel_img_mul_338[2] + 
                kernel_img_mul_338[3] + kernel_img_mul_338[4] + kernel_img_mul_338[5] + 
                kernel_img_mul_338[6] + kernel_img_mul_338[7] + kernel_img_mul_338[8] + 
                kernel_img_mul_338[9] + kernel_img_mul_338[10] + kernel_img_mul_338[11] + 
                kernel_img_mul_338[12] + kernel_img_mul_338[13] + kernel_img_mul_338[14] + 
                kernel_img_mul_338[15] + kernel_img_mul_338[16] + kernel_img_mul_338[17] + 
                kernel_img_mul_338[18] + kernel_img_mul_338[19] + kernel_img_mul_338[20] + 
                kernel_img_mul_338[21] + kernel_img_mul_338[22] + kernel_img_mul_338[23] + 
                kernel_img_mul_338[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2711:2704] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2711:2704] <= kernel_img_sum_338[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2711:2704] <= 'd0;
end

wire  [39:0]  kernel_img_mul_339[0:24];
assign kernel_img_mul_339[0] = buffer_data_4[2703:2696] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_339[1] = buffer_data_4[2711:2704] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_339[2] = buffer_data_4[2719:2712] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_339[3] = buffer_data_4[2727:2720] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_339[4] = buffer_data_4[2735:2728] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_339[5] = buffer_data_3[2703:2696] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_339[6] = buffer_data_3[2711:2704] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_339[7] = buffer_data_3[2719:2712] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_339[8] = buffer_data_3[2727:2720] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_339[9] = buffer_data_3[2735:2728] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_339[10] = buffer_data_2[2703:2696] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_339[11] = buffer_data_2[2711:2704] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_339[12] = buffer_data_2[2719:2712] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_339[13] = buffer_data_2[2727:2720] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_339[14] = buffer_data_2[2735:2728] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_339[15] = buffer_data_1[2703:2696] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_339[16] = buffer_data_1[2711:2704] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_339[17] = buffer_data_1[2719:2712] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_339[18] = buffer_data_1[2727:2720] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_339[19] = buffer_data_1[2735:2728] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_339[20] = buffer_data_0[2703:2696] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_339[21] = buffer_data_0[2711:2704] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_339[22] = buffer_data_0[2719:2712] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_339[23] = buffer_data_0[2727:2720] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_339[24] = buffer_data_0[2735:2728] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_339 = kernel_img_mul_339[0] + kernel_img_mul_339[1] + kernel_img_mul_339[2] + 
                kernel_img_mul_339[3] + kernel_img_mul_339[4] + kernel_img_mul_339[5] + 
                kernel_img_mul_339[6] + kernel_img_mul_339[7] + kernel_img_mul_339[8] + 
                kernel_img_mul_339[9] + kernel_img_mul_339[10] + kernel_img_mul_339[11] + 
                kernel_img_mul_339[12] + kernel_img_mul_339[13] + kernel_img_mul_339[14] + 
                kernel_img_mul_339[15] + kernel_img_mul_339[16] + kernel_img_mul_339[17] + 
                kernel_img_mul_339[18] + kernel_img_mul_339[19] + kernel_img_mul_339[20] + 
                kernel_img_mul_339[21] + kernel_img_mul_339[22] + kernel_img_mul_339[23] + 
                kernel_img_mul_339[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2719:2712] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2719:2712] <= kernel_img_sum_339[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2719:2712] <= 'd0;
end

wire  [39:0]  kernel_img_mul_340[0:24];
assign kernel_img_mul_340[0] = buffer_data_4[2711:2704] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_340[1] = buffer_data_4[2719:2712] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_340[2] = buffer_data_4[2727:2720] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_340[3] = buffer_data_4[2735:2728] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_340[4] = buffer_data_4[2743:2736] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_340[5] = buffer_data_3[2711:2704] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_340[6] = buffer_data_3[2719:2712] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_340[7] = buffer_data_3[2727:2720] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_340[8] = buffer_data_3[2735:2728] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_340[9] = buffer_data_3[2743:2736] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_340[10] = buffer_data_2[2711:2704] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_340[11] = buffer_data_2[2719:2712] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_340[12] = buffer_data_2[2727:2720] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_340[13] = buffer_data_2[2735:2728] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_340[14] = buffer_data_2[2743:2736] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_340[15] = buffer_data_1[2711:2704] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_340[16] = buffer_data_1[2719:2712] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_340[17] = buffer_data_1[2727:2720] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_340[18] = buffer_data_1[2735:2728] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_340[19] = buffer_data_1[2743:2736] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_340[20] = buffer_data_0[2711:2704] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_340[21] = buffer_data_0[2719:2712] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_340[22] = buffer_data_0[2727:2720] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_340[23] = buffer_data_0[2735:2728] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_340[24] = buffer_data_0[2743:2736] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_340 = kernel_img_mul_340[0] + kernel_img_mul_340[1] + kernel_img_mul_340[2] + 
                kernel_img_mul_340[3] + kernel_img_mul_340[4] + kernel_img_mul_340[5] + 
                kernel_img_mul_340[6] + kernel_img_mul_340[7] + kernel_img_mul_340[8] + 
                kernel_img_mul_340[9] + kernel_img_mul_340[10] + kernel_img_mul_340[11] + 
                kernel_img_mul_340[12] + kernel_img_mul_340[13] + kernel_img_mul_340[14] + 
                kernel_img_mul_340[15] + kernel_img_mul_340[16] + kernel_img_mul_340[17] + 
                kernel_img_mul_340[18] + kernel_img_mul_340[19] + kernel_img_mul_340[20] + 
                kernel_img_mul_340[21] + kernel_img_mul_340[22] + kernel_img_mul_340[23] + 
                kernel_img_mul_340[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2727:2720] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2727:2720] <= kernel_img_sum_340[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2727:2720] <= 'd0;
end

wire  [39:0]  kernel_img_mul_341[0:24];
assign kernel_img_mul_341[0] = buffer_data_4[2719:2712] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_341[1] = buffer_data_4[2727:2720] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_341[2] = buffer_data_4[2735:2728] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_341[3] = buffer_data_4[2743:2736] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_341[4] = buffer_data_4[2751:2744] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_341[5] = buffer_data_3[2719:2712] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_341[6] = buffer_data_3[2727:2720] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_341[7] = buffer_data_3[2735:2728] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_341[8] = buffer_data_3[2743:2736] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_341[9] = buffer_data_3[2751:2744] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_341[10] = buffer_data_2[2719:2712] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_341[11] = buffer_data_2[2727:2720] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_341[12] = buffer_data_2[2735:2728] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_341[13] = buffer_data_2[2743:2736] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_341[14] = buffer_data_2[2751:2744] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_341[15] = buffer_data_1[2719:2712] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_341[16] = buffer_data_1[2727:2720] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_341[17] = buffer_data_1[2735:2728] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_341[18] = buffer_data_1[2743:2736] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_341[19] = buffer_data_1[2751:2744] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_341[20] = buffer_data_0[2719:2712] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_341[21] = buffer_data_0[2727:2720] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_341[22] = buffer_data_0[2735:2728] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_341[23] = buffer_data_0[2743:2736] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_341[24] = buffer_data_0[2751:2744] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_341 = kernel_img_mul_341[0] + kernel_img_mul_341[1] + kernel_img_mul_341[2] + 
                kernel_img_mul_341[3] + kernel_img_mul_341[4] + kernel_img_mul_341[5] + 
                kernel_img_mul_341[6] + kernel_img_mul_341[7] + kernel_img_mul_341[8] + 
                kernel_img_mul_341[9] + kernel_img_mul_341[10] + kernel_img_mul_341[11] + 
                kernel_img_mul_341[12] + kernel_img_mul_341[13] + kernel_img_mul_341[14] + 
                kernel_img_mul_341[15] + kernel_img_mul_341[16] + kernel_img_mul_341[17] + 
                kernel_img_mul_341[18] + kernel_img_mul_341[19] + kernel_img_mul_341[20] + 
                kernel_img_mul_341[21] + kernel_img_mul_341[22] + kernel_img_mul_341[23] + 
                kernel_img_mul_341[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2735:2728] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2735:2728] <= kernel_img_sum_341[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2735:2728] <= 'd0;
end

wire  [39:0]  kernel_img_mul_342[0:24];
assign kernel_img_mul_342[0] = buffer_data_4[2727:2720] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_342[1] = buffer_data_4[2735:2728] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_342[2] = buffer_data_4[2743:2736] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_342[3] = buffer_data_4[2751:2744] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_342[4] = buffer_data_4[2759:2752] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_342[5] = buffer_data_3[2727:2720] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_342[6] = buffer_data_3[2735:2728] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_342[7] = buffer_data_3[2743:2736] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_342[8] = buffer_data_3[2751:2744] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_342[9] = buffer_data_3[2759:2752] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_342[10] = buffer_data_2[2727:2720] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_342[11] = buffer_data_2[2735:2728] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_342[12] = buffer_data_2[2743:2736] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_342[13] = buffer_data_2[2751:2744] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_342[14] = buffer_data_2[2759:2752] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_342[15] = buffer_data_1[2727:2720] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_342[16] = buffer_data_1[2735:2728] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_342[17] = buffer_data_1[2743:2736] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_342[18] = buffer_data_1[2751:2744] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_342[19] = buffer_data_1[2759:2752] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_342[20] = buffer_data_0[2727:2720] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_342[21] = buffer_data_0[2735:2728] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_342[22] = buffer_data_0[2743:2736] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_342[23] = buffer_data_0[2751:2744] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_342[24] = buffer_data_0[2759:2752] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_342 = kernel_img_mul_342[0] + kernel_img_mul_342[1] + kernel_img_mul_342[2] + 
                kernel_img_mul_342[3] + kernel_img_mul_342[4] + kernel_img_mul_342[5] + 
                kernel_img_mul_342[6] + kernel_img_mul_342[7] + kernel_img_mul_342[8] + 
                kernel_img_mul_342[9] + kernel_img_mul_342[10] + kernel_img_mul_342[11] + 
                kernel_img_mul_342[12] + kernel_img_mul_342[13] + kernel_img_mul_342[14] + 
                kernel_img_mul_342[15] + kernel_img_mul_342[16] + kernel_img_mul_342[17] + 
                kernel_img_mul_342[18] + kernel_img_mul_342[19] + kernel_img_mul_342[20] + 
                kernel_img_mul_342[21] + kernel_img_mul_342[22] + kernel_img_mul_342[23] + 
                kernel_img_mul_342[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2743:2736] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2743:2736] <= kernel_img_sum_342[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2743:2736] <= 'd0;
end

wire  [39:0]  kernel_img_mul_343[0:24];
assign kernel_img_mul_343[0] = buffer_data_4[2735:2728] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_343[1] = buffer_data_4[2743:2736] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_343[2] = buffer_data_4[2751:2744] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_343[3] = buffer_data_4[2759:2752] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_343[4] = buffer_data_4[2767:2760] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_343[5] = buffer_data_3[2735:2728] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_343[6] = buffer_data_3[2743:2736] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_343[7] = buffer_data_3[2751:2744] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_343[8] = buffer_data_3[2759:2752] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_343[9] = buffer_data_3[2767:2760] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_343[10] = buffer_data_2[2735:2728] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_343[11] = buffer_data_2[2743:2736] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_343[12] = buffer_data_2[2751:2744] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_343[13] = buffer_data_2[2759:2752] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_343[14] = buffer_data_2[2767:2760] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_343[15] = buffer_data_1[2735:2728] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_343[16] = buffer_data_1[2743:2736] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_343[17] = buffer_data_1[2751:2744] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_343[18] = buffer_data_1[2759:2752] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_343[19] = buffer_data_1[2767:2760] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_343[20] = buffer_data_0[2735:2728] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_343[21] = buffer_data_0[2743:2736] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_343[22] = buffer_data_0[2751:2744] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_343[23] = buffer_data_0[2759:2752] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_343[24] = buffer_data_0[2767:2760] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_343 = kernel_img_mul_343[0] + kernel_img_mul_343[1] + kernel_img_mul_343[2] + 
                kernel_img_mul_343[3] + kernel_img_mul_343[4] + kernel_img_mul_343[5] + 
                kernel_img_mul_343[6] + kernel_img_mul_343[7] + kernel_img_mul_343[8] + 
                kernel_img_mul_343[9] + kernel_img_mul_343[10] + kernel_img_mul_343[11] + 
                kernel_img_mul_343[12] + kernel_img_mul_343[13] + kernel_img_mul_343[14] + 
                kernel_img_mul_343[15] + kernel_img_mul_343[16] + kernel_img_mul_343[17] + 
                kernel_img_mul_343[18] + kernel_img_mul_343[19] + kernel_img_mul_343[20] + 
                kernel_img_mul_343[21] + kernel_img_mul_343[22] + kernel_img_mul_343[23] + 
                kernel_img_mul_343[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2751:2744] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2751:2744] <= kernel_img_sum_343[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2751:2744] <= 'd0;
end

wire  [39:0]  kernel_img_mul_344[0:24];
assign kernel_img_mul_344[0] = buffer_data_4[2743:2736] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_344[1] = buffer_data_4[2751:2744] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_344[2] = buffer_data_4[2759:2752] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_344[3] = buffer_data_4[2767:2760] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_344[4] = buffer_data_4[2775:2768] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_344[5] = buffer_data_3[2743:2736] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_344[6] = buffer_data_3[2751:2744] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_344[7] = buffer_data_3[2759:2752] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_344[8] = buffer_data_3[2767:2760] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_344[9] = buffer_data_3[2775:2768] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_344[10] = buffer_data_2[2743:2736] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_344[11] = buffer_data_2[2751:2744] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_344[12] = buffer_data_2[2759:2752] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_344[13] = buffer_data_2[2767:2760] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_344[14] = buffer_data_2[2775:2768] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_344[15] = buffer_data_1[2743:2736] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_344[16] = buffer_data_1[2751:2744] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_344[17] = buffer_data_1[2759:2752] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_344[18] = buffer_data_1[2767:2760] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_344[19] = buffer_data_1[2775:2768] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_344[20] = buffer_data_0[2743:2736] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_344[21] = buffer_data_0[2751:2744] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_344[22] = buffer_data_0[2759:2752] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_344[23] = buffer_data_0[2767:2760] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_344[24] = buffer_data_0[2775:2768] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_344 = kernel_img_mul_344[0] + kernel_img_mul_344[1] + kernel_img_mul_344[2] + 
                kernel_img_mul_344[3] + kernel_img_mul_344[4] + kernel_img_mul_344[5] + 
                kernel_img_mul_344[6] + kernel_img_mul_344[7] + kernel_img_mul_344[8] + 
                kernel_img_mul_344[9] + kernel_img_mul_344[10] + kernel_img_mul_344[11] + 
                kernel_img_mul_344[12] + kernel_img_mul_344[13] + kernel_img_mul_344[14] + 
                kernel_img_mul_344[15] + kernel_img_mul_344[16] + kernel_img_mul_344[17] + 
                kernel_img_mul_344[18] + kernel_img_mul_344[19] + kernel_img_mul_344[20] + 
                kernel_img_mul_344[21] + kernel_img_mul_344[22] + kernel_img_mul_344[23] + 
                kernel_img_mul_344[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2759:2752] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2759:2752] <= kernel_img_sum_344[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2759:2752] <= 'd0;
end

wire  [39:0]  kernel_img_mul_345[0:24];
assign kernel_img_mul_345[0] = buffer_data_4[2751:2744] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_345[1] = buffer_data_4[2759:2752] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_345[2] = buffer_data_4[2767:2760] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_345[3] = buffer_data_4[2775:2768] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_345[4] = buffer_data_4[2783:2776] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_345[5] = buffer_data_3[2751:2744] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_345[6] = buffer_data_3[2759:2752] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_345[7] = buffer_data_3[2767:2760] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_345[8] = buffer_data_3[2775:2768] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_345[9] = buffer_data_3[2783:2776] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_345[10] = buffer_data_2[2751:2744] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_345[11] = buffer_data_2[2759:2752] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_345[12] = buffer_data_2[2767:2760] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_345[13] = buffer_data_2[2775:2768] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_345[14] = buffer_data_2[2783:2776] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_345[15] = buffer_data_1[2751:2744] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_345[16] = buffer_data_1[2759:2752] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_345[17] = buffer_data_1[2767:2760] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_345[18] = buffer_data_1[2775:2768] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_345[19] = buffer_data_1[2783:2776] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_345[20] = buffer_data_0[2751:2744] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_345[21] = buffer_data_0[2759:2752] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_345[22] = buffer_data_0[2767:2760] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_345[23] = buffer_data_0[2775:2768] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_345[24] = buffer_data_0[2783:2776] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_345 = kernel_img_mul_345[0] + kernel_img_mul_345[1] + kernel_img_mul_345[2] + 
                kernel_img_mul_345[3] + kernel_img_mul_345[4] + kernel_img_mul_345[5] + 
                kernel_img_mul_345[6] + kernel_img_mul_345[7] + kernel_img_mul_345[8] + 
                kernel_img_mul_345[9] + kernel_img_mul_345[10] + kernel_img_mul_345[11] + 
                kernel_img_mul_345[12] + kernel_img_mul_345[13] + kernel_img_mul_345[14] + 
                kernel_img_mul_345[15] + kernel_img_mul_345[16] + kernel_img_mul_345[17] + 
                kernel_img_mul_345[18] + kernel_img_mul_345[19] + kernel_img_mul_345[20] + 
                kernel_img_mul_345[21] + kernel_img_mul_345[22] + kernel_img_mul_345[23] + 
                kernel_img_mul_345[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2767:2760] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2767:2760] <= kernel_img_sum_345[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2767:2760] <= 'd0;
end

wire  [39:0]  kernel_img_mul_346[0:24];
assign kernel_img_mul_346[0] = buffer_data_4[2759:2752] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_346[1] = buffer_data_4[2767:2760] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_346[2] = buffer_data_4[2775:2768] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_346[3] = buffer_data_4[2783:2776] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_346[4] = buffer_data_4[2791:2784] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_346[5] = buffer_data_3[2759:2752] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_346[6] = buffer_data_3[2767:2760] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_346[7] = buffer_data_3[2775:2768] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_346[8] = buffer_data_3[2783:2776] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_346[9] = buffer_data_3[2791:2784] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_346[10] = buffer_data_2[2759:2752] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_346[11] = buffer_data_2[2767:2760] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_346[12] = buffer_data_2[2775:2768] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_346[13] = buffer_data_2[2783:2776] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_346[14] = buffer_data_2[2791:2784] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_346[15] = buffer_data_1[2759:2752] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_346[16] = buffer_data_1[2767:2760] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_346[17] = buffer_data_1[2775:2768] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_346[18] = buffer_data_1[2783:2776] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_346[19] = buffer_data_1[2791:2784] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_346[20] = buffer_data_0[2759:2752] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_346[21] = buffer_data_0[2767:2760] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_346[22] = buffer_data_0[2775:2768] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_346[23] = buffer_data_0[2783:2776] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_346[24] = buffer_data_0[2791:2784] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_346 = kernel_img_mul_346[0] + kernel_img_mul_346[1] + kernel_img_mul_346[2] + 
                kernel_img_mul_346[3] + kernel_img_mul_346[4] + kernel_img_mul_346[5] + 
                kernel_img_mul_346[6] + kernel_img_mul_346[7] + kernel_img_mul_346[8] + 
                kernel_img_mul_346[9] + kernel_img_mul_346[10] + kernel_img_mul_346[11] + 
                kernel_img_mul_346[12] + kernel_img_mul_346[13] + kernel_img_mul_346[14] + 
                kernel_img_mul_346[15] + kernel_img_mul_346[16] + kernel_img_mul_346[17] + 
                kernel_img_mul_346[18] + kernel_img_mul_346[19] + kernel_img_mul_346[20] + 
                kernel_img_mul_346[21] + kernel_img_mul_346[22] + kernel_img_mul_346[23] + 
                kernel_img_mul_346[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2775:2768] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2775:2768] <= kernel_img_sum_346[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2775:2768] <= 'd0;
end

wire  [39:0]  kernel_img_mul_347[0:24];
assign kernel_img_mul_347[0] = buffer_data_4[2767:2760] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_347[1] = buffer_data_4[2775:2768] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_347[2] = buffer_data_4[2783:2776] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_347[3] = buffer_data_4[2791:2784] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_347[4] = buffer_data_4[2799:2792] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_347[5] = buffer_data_3[2767:2760] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_347[6] = buffer_data_3[2775:2768] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_347[7] = buffer_data_3[2783:2776] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_347[8] = buffer_data_3[2791:2784] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_347[9] = buffer_data_3[2799:2792] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_347[10] = buffer_data_2[2767:2760] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_347[11] = buffer_data_2[2775:2768] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_347[12] = buffer_data_2[2783:2776] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_347[13] = buffer_data_2[2791:2784] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_347[14] = buffer_data_2[2799:2792] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_347[15] = buffer_data_1[2767:2760] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_347[16] = buffer_data_1[2775:2768] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_347[17] = buffer_data_1[2783:2776] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_347[18] = buffer_data_1[2791:2784] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_347[19] = buffer_data_1[2799:2792] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_347[20] = buffer_data_0[2767:2760] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_347[21] = buffer_data_0[2775:2768] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_347[22] = buffer_data_0[2783:2776] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_347[23] = buffer_data_0[2791:2784] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_347[24] = buffer_data_0[2799:2792] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_347 = kernel_img_mul_347[0] + kernel_img_mul_347[1] + kernel_img_mul_347[2] + 
                kernel_img_mul_347[3] + kernel_img_mul_347[4] + kernel_img_mul_347[5] + 
                kernel_img_mul_347[6] + kernel_img_mul_347[7] + kernel_img_mul_347[8] + 
                kernel_img_mul_347[9] + kernel_img_mul_347[10] + kernel_img_mul_347[11] + 
                kernel_img_mul_347[12] + kernel_img_mul_347[13] + kernel_img_mul_347[14] + 
                kernel_img_mul_347[15] + kernel_img_mul_347[16] + kernel_img_mul_347[17] + 
                kernel_img_mul_347[18] + kernel_img_mul_347[19] + kernel_img_mul_347[20] + 
                kernel_img_mul_347[21] + kernel_img_mul_347[22] + kernel_img_mul_347[23] + 
                kernel_img_mul_347[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2783:2776] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2783:2776] <= kernel_img_sum_347[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2783:2776] <= 'd0;
end

wire  [39:0]  kernel_img_mul_348[0:24];
assign kernel_img_mul_348[0] = buffer_data_4[2775:2768] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_348[1] = buffer_data_4[2783:2776] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_348[2] = buffer_data_4[2791:2784] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_348[3] = buffer_data_4[2799:2792] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_348[4] = buffer_data_4[2807:2800] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_348[5] = buffer_data_3[2775:2768] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_348[6] = buffer_data_3[2783:2776] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_348[7] = buffer_data_3[2791:2784] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_348[8] = buffer_data_3[2799:2792] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_348[9] = buffer_data_3[2807:2800] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_348[10] = buffer_data_2[2775:2768] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_348[11] = buffer_data_2[2783:2776] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_348[12] = buffer_data_2[2791:2784] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_348[13] = buffer_data_2[2799:2792] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_348[14] = buffer_data_2[2807:2800] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_348[15] = buffer_data_1[2775:2768] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_348[16] = buffer_data_1[2783:2776] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_348[17] = buffer_data_1[2791:2784] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_348[18] = buffer_data_1[2799:2792] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_348[19] = buffer_data_1[2807:2800] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_348[20] = buffer_data_0[2775:2768] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_348[21] = buffer_data_0[2783:2776] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_348[22] = buffer_data_0[2791:2784] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_348[23] = buffer_data_0[2799:2792] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_348[24] = buffer_data_0[2807:2800] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_348 = kernel_img_mul_348[0] + kernel_img_mul_348[1] + kernel_img_mul_348[2] + 
                kernel_img_mul_348[3] + kernel_img_mul_348[4] + kernel_img_mul_348[5] + 
                kernel_img_mul_348[6] + kernel_img_mul_348[7] + kernel_img_mul_348[8] + 
                kernel_img_mul_348[9] + kernel_img_mul_348[10] + kernel_img_mul_348[11] + 
                kernel_img_mul_348[12] + kernel_img_mul_348[13] + kernel_img_mul_348[14] + 
                kernel_img_mul_348[15] + kernel_img_mul_348[16] + kernel_img_mul_348[17] + 
                kernel_img_mul_348[18] + kernel_img_mul_348[19] + kernel_img_mul_348[20] + 
                kernel_img_mul_348[21] + kernel_img_mul_348[22] + kernel_img_mul_348[23] + 
                kernel_img_mul_348[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2791:2784] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2791:2784] <= kernel_img_sum_348[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2791:2784] <= 'd0;
end

wire  [39:0]  kernel_img_mul_349[0:24];
assign kernel_img_mul_349[0] = buffer_data_4[2783:2776] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_349[1] = buffer_data_4[2791:2784] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_349[2] = buffer_data_4[2799:2792] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_349[3] = buffer_data_4[2807:2800] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_349[4] = buffer_data_4[2815:2808] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_349[5] = buffer_data_3[2783:2776] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_349[6] = buffer_data_3[2791:2784] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_349[7] = buffer_data_3[2799:2792] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_349[8] = buffer_data_3[2807:2800] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_349[9] = buffer_data_3[2815:2808] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_349[10] = buffer_data_2[2783:2776] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_349[11] = buffer_data_2[2791:2784] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_349[12] = buffer_data_2[2799:2792] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_349[13] = buffer_data_2[2807:2800] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_349[14] = buffer_data_2[2815:2808] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_349[15] = buffer_data_1[2783:2776] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_349[16] = buffer_data_1[2791:2784] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_349[17] = buffer_data_1[2799:2792] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_349[18] = buffer_data_1[2807:2800] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_349[19] = buffer_data_1[2815:2808] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_349[20] = buffer_data_0[2783:2776] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_349[21] = buffer_data_0[2791:2784] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_349[22] = buffer_data_0[2799:2792] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_349[23] = buffer_data_0[2807:2800] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_349[24] = buffer_data_0[2815:2808] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_349 = kernel_img_mul_349[0] + kernel_img_mul_349[1] + kernel_img_mul_349[2] + 
                kernel_img_mul_349[3] + kernel_img_mul_349[4] + kernel_img_mul_349[5] + 
                kernel_img_mul_349[6] + kernel_img_mul_349[7] + kernel_img_mul_349[8] + 
                kernel_img_mul_349[9] + kernel_img_mul_349[10] + kernel_img_mul_349[11] + 
                kernel_img_mul_349[12] + kernel_img_mul_349[13] + kernel_img_mul_349[14] + 
                kernel_img_mul_349[15] + kernel_img_mul_349[16] + kernel_img_mul_349[17] + 
                kernel_img_mul_349[18] + kernel_img_mul_349[19] + kernel_img_mul_349[20] + 
                kernel_img_mul_349[21] + kernel_img_mul_349[22] + kernel_img_mul_349[23] + 
                kernel_img_mul_349[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2799:2792] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2799:2792] <= kernel_img_sum_349[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2799:2792] <= 'd0;
end

wire  [39:0]  kernel_img_mul_350[0:24];
assign kernel_img_mul_350[0] = buffer_data_4[2791:2784] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_350[1] = buffer_data_4[2799:2792] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_350[2] = buffer_data_4[2807:2800] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_350[3] = buffer_data_4[2815:2808] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_350[4] = buffer_data_4[2823:2816] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_350[5] = buffer_data_3[2791:2784] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_350[6] = buffer_data_3[2799:2792] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_350[7] = buffer_data_3[2807:2800] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_350[8] = buffer_data_3[2815:2808] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_350[9] = buffer_data_3[2823:2816] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_350[10] = buffer_data_2[2791:2784] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_350[11] = buffer_data_2[2799:2792] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_350[12] = buffer_data_2[2807:2800] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_350[13] = buffer_data_2[2815:2808] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_350[14] = buffer_data_2[2823:2816] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_350[15] = buffer_data_1[2791:2784] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_350[16] = buffer_data_1[2799:2792] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_350[17] = buffer_data_1[2807:2800] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_350[18] = buffer_data_1[2815:2808] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_350[19] = buffer_data_1[2823:2816] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_350[20] = buffer_data_0[2791:2784] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_350[21] = buffer_data_0[2799:2792] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_350[22] = buffer_data_0[2807:2800] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_350[23] = buffer_data_0[2815:2808] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_350[24] = buffer_data_0[2823:2816] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_350 = kernel_img_mul_350[0] + kernel_img_mul_350[1] + kernel_img_mul_350[2] + 
                kernel_img_mul_350[3] + kernel_img_mul_350[4] + kernel_img_mul_350[5] + 
                kernel_img_mul_350[6] + kernel_img_mul_350[7] + kernel_img_mul_350[8] + 
                kernel_img_mul_350[9] + kernel_img_mul_350[10] + kernel_img_mul_350[11] + 
                kernel_img_mul_350[12] + kernel_img_mul_350[13] + kernel_img_mul_350[14] + 
                kernel_img_mul_350[15] + kernel_img_mul_350[16] + kernel_img_mul_350[17] + 
                kernel_img_mul_350[18] + kernel_img_mul_350[19] + kernel_img_mul_350[20] + 
                kernel_img_mul_350[21] + kernel_img_mul_350[22] + kernel_img_mul_350[23] + 
                kernel_img_mul_350[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2807:2800] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2807:2800] <= kernel_img_sum_350[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2807:2800] <= 'd0;
end

wire  [39:0]  kernel_img_mul_351[0:24];
assign kernel_img_mul_351[0] = buffer_data_4[2799:2792] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_351[1] = buffer_data_4[2807:2800] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_351[2] = buffer_data_4[2815:2808] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_351[3] = buffer_data_4[2823:2816] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_351[4] = buffer_data_4[2831:2824] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_351[5] = buffer_data_3[2799:2792] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_351[6] = buffer_data_3[2807:2800] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_351[7] = buffer_data_3[2815:2808] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_351[8] = buffer_data_3[2823:2816] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_351[9] = buffer_data_3[2831:2824] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_351[10] = buffer_data_2[2799:2792] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_351[11] = buffer_data_2[2807:2800] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_351[12] = buffer_data_2[2815:2808] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_351[13] = buffer_data_2[2823:2816] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_351[14] = buffer_data_2[2831:2824] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_351[15] = buffer_data_1[2799:2792] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_351[16] = buffer_data_1[2807:2800] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_351[17] = buffer_data_1[2815:2808] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_351[18] = buffer_data_1[2823:2816] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_351[19] = buffer_data_1[2831:2824] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_351[20] = buffer_data_0[2799:2792] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_351[21] = buffer_data_0[2807:2800] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_351[22] = buffer_data_0[2815:2808] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_351[23] = buffer_data_0[2823:2816] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_351[24] = buffer_data_0[2831:2824] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_351 = kernel_img_mul_351[0] + kernel_img_mul_351[1] + kernel_img_mul_351[2] + 
                kernel_img_mul_351[3] + kernel_img_mul_351[4] + kernel_img_mul_351[5] + 
                kernel_img_mul_351[6] + kernel_img_mul_351[7] + kernel_img_mul_351[8] + 
                kernel_img_mul_351[9] + kernel_img_mul_351[10] + kernel_img_mul_351[11] + 
                kernel_img_mul_351[12] + kernel_img_mul_351[13] + kernel_img_mul_351[14] + 
                kernel_img_mul_351[15] + kernel_img_mul_351[16] + kernel_img_mul_351[17] + 
                kernel_img_mul_351[18] + kernel_img_mul_351[19] + kernel_img_mul_351[20] + 
                kernel_img_mul_351[21] + kernel_img_mul_351[22] + kernel_img_mul_351[23] + 
                kernel_img_mul_351[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2815:2808] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2815:2808] <= kernel_img_sum_351[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2815:2808] <= 'd0;
end

wire  [39:0]  kernel_img_mul_352[0:24];
assign kernel_img_mul_352[0] = buffer_data_4[2807:2800] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_352[1] = buffer_data_4[2815:2808] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_352[2] = buffer_data_4[2823:2816] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_352[3] = buffer_data_4[2831:2824] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_352[4] = buffer_data_4[2839:2832] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_352[5] = buffer_data_3[2807:2800] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_352[6] = buffer_data_3[2815:2808] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_352[7] = buffer_data_3[2823:2816] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_352[8] = buffer_data_3[2831:2824] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_352[9] = buffer_data_3[2839:2832] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_352[10] = buffer_data_2[2807:2800] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_352[11] = buffer_data_2[2815:2808] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_352[12] = buffer_data_2[2823:2816] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_352[13] = buffer_data_2[2831:2824] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_352[14] = buffer_data_2[2839:2832] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_352[15] = buffer_data_1[2807:2800] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_352[16] = buffer_data_1[2815:2808] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_352[17] = buffer_data_1[2823:2816] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_352[18] = buffer_data_1[2831:2824] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_352[19] = buffer_data_1[2839:2832] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_352[20] = buffer_data_0[2807:2800] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_352[21] = buffer_data_0[2815:2808] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_352[22] = buffer_data_0[2823:2816] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_352[23] = buffer_data_0[2831:2824] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_352[24] = buffer_data_0[2839:2832] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_352 = kernel_img_mul_352[0] + kernel_img_mul_352[1] + kernel_img_mul_352[2] + 
                kernel_img_mul_352[3] + kernel_img_mul_352[4] + kernel_img_mul_352[5] + 
                kernel_img_mul_352[6] + kernel_img_mul_352[7] + kernel_img_mul_352[8] + 
                kernel_img_mul_352[9] + kernel_img_mul_352[10] + kernel_img_mul_352[11] + 
                kernel_img_mul_352[12] + kernel_img_mul_352[13] + kernel_img_mul_352[14] + 
                kernel_img_mul_352[15] + kernel_img_mul_352[16] + kernel_img_mul_352[17] + 
                kernel_img_mul_352[18] + kernel_img_mul_352[19] + kernel_img_mul_352[20] + 
                kernel_img_mul_352[21] + kernel_img_mul_352[22] + kernel_img_mul_352[23] + 
                kernel_img_mul_352[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2823:2816] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2823:2816] <= kernel_img_sum_352[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2823:2816] <= 'd0;
end

wire  [39:0]  kernel_img_mul_353[0:24];
assign kernel_img_mul_353[0] = buffer_data_4[2815:2808] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_353[1] = buffer_data_4[2823:2816] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_353[2] = buffer_data_4[2831:2824] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_353[3] = buffer_data_4[2839:2832] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_353[4] = buffer_data_4[2847:2840] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_353[5] = buffer_data_3[2815:2808] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_353[6] = buffer_data_3[2823:2816] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_353[7] = buffer_data_3[2831:2824] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_353[8] = buffer_data_3[2839:2832] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_353[9] = buffer_data_3[2847:2840] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_353[10] = buffer_data_2[2815:2808] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_353[11] = buffer_data_2[2823:2816] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_353[12] = buffer_data_2[2831:2824] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_353[13] = buffer_data_2[2839:2832] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_353[14] = buffer_data_2[2847:2840] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_353[15] = buffer_data_1[2815:2808] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_353[16] = buffer_data_1[2823:2816] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_353[17] = buffer_data_1[2831:2824] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_353[18] = buffer_data_1[2839:2832] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_353[19] = buffer_data_1[2847:2840] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_353[20] = buffer_data_0[2815:2808] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_353[21] = buffer_data_0[2823:2816] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_353[22] = buffer_data_0[2831:2824] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_353[23] = buffer_data_0[2839:2832] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_353[24] = buffer_data_0[2847:2840] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_353 = kernel_img_mul_353[0] + kernel_img_mul_353[1] + kernel_img_mul_353[2] + 
                kernel_img_mul_353[3] + kernel_img_mul_353[4] + kernel_img_mul_353[5] + 
                kernel_img_mul_353[6] + kernel_img_mul_353[7] + kernel_img_mul_353[8] + 
                kernel_img_mul_353[9] + kernel_img_mul_353[10] + kernel_img_mul_353[11] + 
                kernel_img_mul_353[12] + kernel_img_mul_353[13] + kernel_img_mul_353[14] + 
                kernel_img_mul_353[15] + kernel_img_mul_353[16] + kernel_img_mul_353[17] + 
                kernel_img_mul_353[18] + kernel_img_mul_353[19] + kernel_img_mul_353[20] + 
                kernel_img_mul_353[21] + kernel_img_mul_353[22] + kernel_img_mul_353[23] + 
                kernel_img_mul_353[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2831:2824] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2831:2824] <= kernel_img_sum_353[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2831:2824] <= 'd0;
end

wire  [39:0]  kernel_img_mul_354[0:24];
assign kernel_img_mul_354[0] = buffer_data_4[2823:2816] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_354[1] = buffer_data_4[2831:2824] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_354[2] = buffer_data_4[2839:2832] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_354[3] = buffer_data_4[2847:2840] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_354[4] = buffer_data_4[2855:2848] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_354[5] = buffer_data_3[2823:2816] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_354[6] = buffer_data_3[2831:2824] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_354[7] = buffer_data_3[2839:2832] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_354[8] = buffer_data_3[2847:2840] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_354[9] = buffer_data_3[2855:2848] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_354[10] = buffer_data_2[2823:2816] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_354[11] = buffer_data_2[2831:2824] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_354[12] = buffer_data_2[2839:2832] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_354[13] = buffer_data_2[2847:2840] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_354[14] = buffer_data_2[2855:2848] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_354[15] = buffer_data_1[2823:2816] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_354[16] = buffer_data_1[2831:2824] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_354[17] = buffer_data_1[2839:2832] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_354[18] = buffer_data_1[2847:2840] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_354[19] = buffer_data_1[2855:2848] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_354[20] = buffer_data_0[2823:2816] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_354[21] = buffer_data_0[2831:2824] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_354[22] = buffer_data_0[2839:2832] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_354[23] = buffer_data_0[2847:2840] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_354[24] = buffer_data_0[2855:2848] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_354 = kernel_img_mul_354[0] + kernel_img_mul_354[1] + kernel_img_mul_354[2] + 
                kernel_img_mul_354[3] + kernel_img_mul_354[4] + kernel_img_mul_354[5] + 
                kernel_img_mul_354[6] + kernel_img_mul_354[7] + kernel_img_mul_354[8] + 
                kernel_img_mul_354[9] + kernel_img_mul_354[10] + kernel_img_mul_354[11] + 
                kernel_img_mul_354[12] + kernel_img_mul_354[13] + kernel_img_mul_354[14] + 
                kernel_img_mul_354[15] + kernel_img_mul_354[16] + kernel_img_mul_354[17] + 
                kernel_img_mul_354[18] + kernel_img_mul_354[19] + kernel_img_mul_354[20] + 
                kernel_img_mul_354[21] + kernel_img_mul_354[22] + kernel_img_mul_354[23] + 
                kernel_img_mul_354[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2839:2832] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2839:2832] <= kernel_img_sum_354[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2839:2832] <= 'd0;
end

wire  [39:0]  kernel_img_mul_355[0:24];
assign kernel_img_mul_355[0] = buffer_data_4[2831:2824] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_355[1] = buffer_data_4[2839:2832] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_355[2] = buffer_data_4[2847:2840] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_355[3] = buffer_data_4[2855:2848] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_355[4] = buffer_data_4[2863:2856] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_355[5] = buffer_data_3[2831:2824] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_355[6] = buffer_data_3[2839:2832] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_355[7] = buffer_data_3[2847:2840] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_355[8] = buffer_data_3[2855:2848] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_355[9] = buffer_data_3[2863:2856] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_355[10] = buffer_data_2[2831:2824] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_355[11] = buffer_data_2[2839:2832] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_355[12] = buffer_data_2[2847:2840] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_355[13] = buffer_data_2[2855:2848] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_355[14] = buffer_data_2[2863:2856] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_355[15] = buffer_data_1[2831:2824] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_355[16] = buffer_data_1[2839:2832] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_355[17] = buffer_data_1[2847:2840] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_355[18] = buffer_data_1[2855:2848] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_355[19] = buffer_data_1[2863:2856] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_355[20] = buffer_data_0[2831:2824] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_355[21] = buffer_data_0[2839:2832] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_355[22] = buffer_data_0[2847:2840] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_355[23] = buffer_data_0[2855:2848] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_355[24] = buffer_data_0[2863:2856] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_355 = kernel_img_mul_355[0] + kernel_img_mul_355[1] + kernel_img_mul_355[2] + 
                kernel_img_mul_355[3] + kernel_img_mul_355[4] + kernel_img_mul_355[5] + 
                kernel_img_mul_355[6] + kernel_img_mul_355[7] + kernel_img_mul_355[8] + 
                kernel_img_mul_355[9] + kernel_img_mul_355[10] + kernel_img_mul_355[11] + 
                kernel_img_mul_355[12] + kernel_img_mul_355[13] + kernel_img_mul_355[14] + 
                kernel_img_mul_355[15] + kernel_img_mul_355[16] + kernel_img_mul_355[17] + 
                kernel_img_mul_355[18] + kernel_img_mul_355[19] + kernel_img_mul_355[20] + 
                kernel_img_mul_355[21] + kernel_img_mul_355[22] + kernel_img_mul_355[23] + 
                kernel_img_mul_355[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2847:2840] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2847:2840] <= kernel_img_sum_355[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2847:2840] <= 'd0;
end

wire  [39:0]  kernel_img_mul_356[0:24];
assign kernel_img_mul_356[0] = buffer_data_4[2839:2832] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_356[1] = buffer_data_4[2847:2840] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_356[2] = buffer_data_4[2855:2848] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_356[3] = buffer_data_4[2863:2856] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_356[4] = buffer_data_4[2871:2864] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_356[5] = buffer_data_3[2839:2832] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_356[6] = buffer_data_3[2847:2840] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_356[7] = buffer_data_3[2855:2848] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_356[8] = buffer_data_3[2863:2856] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_356[9] = buffer_data_3[2871:2864] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_356[10] = buffer_data_2[2839:2832] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_356[11] = buffer_data_2[2847:2840] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_356[12] = buffer_data_2[2855:2848] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_356[13] = buffer_data_2[2863:2856] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_356[14] = buffer_data_2[2871:2864] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_356[15] = buffer_data_1[2839:2832] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_356[16] = buffer_data_1[2847:2840] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_356[17] = buffer_data_1[2855:2848] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_356[18] = buffer_data_1[2863:2856] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_356[19] = buffer_data_1[2871:2864] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_356[20] = buffer_data_0[2839:2832] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_356[21] = buffer_data_0[2847:2840] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_356[22] = buffer_data_0[2855:2848] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_356[23] = buffer_data_0[2863:2856] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_356[24] = buffer_data_0[2871:2864] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_356 = kernel_img_mul_356[0] + kernel_img_mul_356[1] + kernel_img_mul_356[2] + 
                kernel_img_mul_356[3] + kernel_img_mul_356[4] + kernel_img_mul_356[5] + 
                kernel_img_mul_356[6] + kernel_img_mul_356[7] + kernel_img_mul_356[8] + 
                kernel_img_mul_356[9] + kernel_img_mul_356[10] + kernel_img_mul_356[11] + 
                kernel_img_mul_356[12] + kernel_img_mul_356[13] + kernel_img_mul_356[14] + 
                kernel_img_mul_356[15] + kernel_img_mul_356[16] + kernel_img_mul_356[17] + 
                kernel_img_mul_356[18] + kernel_img_mul_356[19] + kernel_img_mul_356[20] + 
                kernel_img_mul_356[21] + kernel_img_mul_356[22] + kernel_img_mul_356[23] + 
                kernel_img_mul_356[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2855:2848] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2855:2848] <= kernel_img_sum_356[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2855:2848] <= 'd0;
end

wire  [39:0]  kernel_img_mul_357[0:24];
assign kernel_img_mul_357[0] = buffer_data_4[2847:2840] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_357[1] = buffer_data_4[2855:2848] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_357[2] = buffer_data_4[2863:2856] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_357[3] = buffer_data_4[2871:2864] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_357[4] = buffer_data_4[2879:2872] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_357[5] = buffer_data_3[2847:2840] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_357[6] = buffer_data_3[2855:2848] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_357[7] = buffer_data_3[2863:2856] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_357[8] = buffer_data_3[2871:2864] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_357[9] = buffer_data_3[2879:2872] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_357[10] = buffer_data_2[2847:2840] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_357[11] = buffer_data_2[2855:2848] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_357[12] = buffer_data_2[2863:2856] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_357[13] = buffer_data_2[2871:2864] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_357[14] = buffer_data_2[2879:2872] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_357[15] = buffer_data_1[2847:2840] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_357[16] = buffer_data_1[2855:2848] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_357[17] = buffer_data_1[2863:2856] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_357[18] = buffer_data_1[2871:2864] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_357[19] = buffer_data_1[2879:2872] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_357[20] = buffer_data_0[2847:2840] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_357[21] = buffer_data_0[2855:2848] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_357[22] = buffer_data_0[2863:2856] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_357[23] = buffer_data_0[2871:2864] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_357[24] = buffer_data_0[2879:2872] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_357 = kernel_img_mul_357[0] + kernel_img_mul_357[1] + kernel_img_mul_357[2] + 
                kernel_img_mul_357[3] + kernel_img_mul_357[4] + kernel_img_mul_357[5] + 
                kernel_img_mul_357[6] + kernel_img_mul_357[7] + kernel_img_mul_357[8] + 
                kernel_img_mul_357[9] + kernel_img_mul_357[10] + kernel_img_mul_357[11] + 
                kernel_img_mul_357[12] + kernel_img_mul_357[13] + kernel_img_mul_357[14] + 
                kernel_img_mul_357[15] + kernel_img_mul_357[16] + kernel_img_mul_357[17] + 
                kernel_img_mul_357[18] + kernel_img_mul_357[19] + kernel_img_mul_357[20] + 
                kernel_img_mul_357[21] + kernel_img_mul_357[22] + kernel_img_mul_357[23] + 
                kernel_img_mul_357[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2863:2856] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2863:2856] <= kernel_img_sum_357[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2863:2856] <= 'd0;
end

wire  [39:0]  kernel_img_mul_358[0:24];
assign kernel_img_mul_358[0] = buffer_data_4[2855:2848] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_358[1] = buffer_data_4[2863:2856] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_358[2] = buffer_data_4[2871:2864] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_358[3] = buffer_data_4[2879:2872] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_358[4] = buffer_data_4[2887:2880] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_358[5] = buffer_data_3[2855:2848] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_358[6] = buffer_data_3[2863:2856] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_358[7] = buffer_data_3[2871:2864] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_358[8] = buffer_data_3[2879:2872] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_358[9] = buffer_data_3[2887:2880] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_358[10] = buffer_data_2[2855:2848] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_358[11] = buffer_data_2[2863:2856] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_358[12] = buffer_data_2[2871:2864] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_358[13] = buffer_data_2[2879:2872] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_358[14] = buffer_data_2[2887:2880] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_358[15] = buffer_data_1[2855:2848] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_358[16] = buffer_data_1[2863:2856] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_358[17] = buffer_data_1[2871:2864] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_358[18] = buffer_data_1[2879:2872] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_358[19] = buffer_data_1[2887:2880] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_358[20] = buffer_data_0[2855:2848] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_358[21] = buffer_data_0[2863:2856] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_358[22] = buffer_data_0[2871:2864] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_358[23] = buffer_data_0[2879:2872] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_358[24] = buffer_data_0[2887:2880] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_358 = kernel_img_mul_358[0] + kernel_img_mul_358[1] + kernel_img_mul_358[2] + 
                kernel_img_mul_358[3] + kernel_img_mul_358[4] + kernel_img_mul_358[5] + 
                kernel_img_mul_358[6] + kernel_img_mul_358[7] + kernel_img_mul_358[8] + 
                kernel_img_mul_358[9] + kernel_img_mul_358[10] + kernel_img_mul_358[11] + 
                kernel_img_mul_358[12] + kernel_img_mul_358[13] + kernel_img_mul_358[14] + 
                kernel_img_mul_358[15] + kernel_img_mul_358[16] + kernel_img_mul_358[17] + 
                kernel_img_mul_358[18] + kernel_img_mul_358[19] + kernel_img_mul_358[20] + 
                kernel_img_mul_358[21] + kernel_img_mul_358[22] + kernel_img_mul_358[23] + 
                kernel_img_mul_358[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2871:2864] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2871:2864] <= kernel_img_sum_358[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2871:2864] <= 'd0;
end

wire  [39:0]  kernel_img_mul_359[0:24];
assign kernel_img_mul_359[0] = buffer_data_4[2863:2856] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_359[1] = buffer_data_4[2871:2864] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_359[2] = buffer_data_4[2879:2872] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_359[3] = buffer_data_4[2887:2880] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_359[4] = buffer_data_4[2895:2888] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_359[5] = buffer_data_3[2863:2856] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_359[6] = buffer_data_3[2871:2864] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_359[7] = buffer_data_3[2879:2872] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_359[8] = buffer_data_3[2887:2880] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_359[9] = buffer_data_3[2895:2888] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_359[10] = buffer_data_2[2863:2856] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_359[11] = buffer_data_2[2871:2864] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_359[12] = buffer_data_2[2879:2872] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_359[13] = buffer_data_2[2887:2880] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_359[14] = buffer_data_2[2895:2888] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_359[15] = buffer_data_1[2863:2856] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_359[16] = buffer_data_1[2871:2864] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_359[17] = buffer_data_1[2879:2872] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_359[18] = buffer_data_1[2887:2880] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_359[19] = buffer_data_1[2895:2888] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_359[20] = buffer_data_0[2863:2856] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_359[21] = buffer_data_0[2871:2864] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_359[22] = buffer_data_0[2879:2872] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_359[23] = buffer_data_0[2887:2880] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_359[24] = buffer_data_0[2895:2888] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_359 = kernel_img_mul_359[0] + kernel_img_mul_359[1] + kernel_img_mul_359[2] + 
                kernel_img_mul_359[3] + kernel_img_mul_359[4] + kernel_img_mul_359[5] + 
                kernel_img_mul_359[6] + kernel_img_mul_359[7] + kernel_img_mul_359[8] + 
                kernel_img_mul_359[9] + kernel_img_mul_359[10] + kernel_img_mul_359[11] + 
                kernel_img_mul_359[12] + kernel_img_mul_359[13] + kernel_img_mul_359[14] + 
                kernel_img_mul_359[15] + kernel_img_mul_359[16] + kernel_img_mul_359[17] + 
                kernel_img_mul_359[18] + kernel_img_mul_359[19] + kernel_img_mul_359[20] + 
                kernel_img_mul_359[21] + kernel_img_mul_359[22] + kernel_img_mul_359[23] + 
                kernel_img_mul_359[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2879:2872] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2879:2872] <= kernel_img_sum_359[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2879:2872] <= 'd0;
end

wire  [39:0]  kernel_img_mul_360[0:24];
assign kernel_img_mul_360[0] = buffer_data_4[2871:2864] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_360[1] = buffer_data_4[2879:2872] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_360[2] = buffer_data_4[2887:2880] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_360[3] = buffer_data_4[2895:2888] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_360[4] = buffer_data_4[2903:2896] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_360[5] = buffer_data_3[2871:2864] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_360[6] = buffer_data_3[2879:2872] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_360[7] = buffer_data_3[2887:2880] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_360[8] = buffer_data_3[2895:2888] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_360[9] = buffer_data_3[2903:2896] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_360[10] = buffer_data_2[2871:2864] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_360[11] = buffer_data_2[2879:2872] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_360[12] = buffer_data_2[2887:2880] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_360[13] = buffer_data_2[2895:2888] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_360[14] = buffer_data_2[2903:2896] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_360[15] = buffer_data_1[2871:2864] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_360[16] = buffer_data_1[2879:2872] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_360[17] = buffer_data_1[2887:2880] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_360[18] = buffer_data_1[2895:2888] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_360[19] = buffer_data_1[2903:2896] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_360[20] = buffer_data_0[2871:2864] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_360[21] = buffer_data_0[2879:2872] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_360[22] = buffer_data_0[2887:2880] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_360[23] = buffer_data_0[2895:2888] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_360[24] = buffer_data_0[2903:2896] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_360 = kernel_img_mul_360[0] + kernel_img_mul_360[1] + kernel_img_mul_360[2] + 
                kernel_img_mul_360[3] + kernel_img_mul_360[4] + kernel_img_mul_360[5] + 
                kernel_img_mul_360[6] + kernel_img_mul_360[7] + kernel_img_mul_360[8] + 
                kernel_img_mul_360[9] + kernel_img_mul_360[10] + kernel_img_mul_360[11] + 
                kernel_img_mul_360[12] + kernel_img_mul_360[13] + kernel_img_mul_360[14] + 
                kernel_img_mul_360[15] + kernel_img_mul_360[16] + kernel_img_mul_360[17] + 
                kernel_img_mul_360[18] + kernel_img_mul_360[19] + kernel_img_mul_360[20] + 
                kernel_img_mul_360[21] + kernel_img_mul_360[22] + kernel_img_mul_360[23] + 
                kernel_img_mul_360[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2887:2880] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2887:2880] <= kernel_img_sum_360[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2887:2880] <= 'd0;
end

wire  [39:0]  kernel_img_mul_361[0:24];
assign kernel_img_mul_361[0] = buffer_data_4[2879:2872] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_361[1] = buffer_data_4[2887:2880] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_361[2] = buffer_data_4[2895:2888] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_361[3] = buffer_data_4[2903:2896] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_361[4] = buffer_data_4[2911:2904] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_361[5] = buffer_data_3[2879:2872] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_361[6] = buffer_data_3[2887:2880] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_361[7] = buffer_data_3[2895:2888] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_361[8] = buffer_data_3[2903:2896] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_361[9] = buffer_data_3[2911:2904] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_361[10] = buffer_data_2[2879:2872] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_361[11] = buffer_data_2[2887:2880] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_361[12] = buffer_data_2[2895:2888] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_361[13] = buffer_data_2[2903:2896] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_361[14] = buffer_data_2[2911:2904] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_361[15] = buffer_data_1[2879:2872] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_361[16] = buffer_data_1[2887:2880] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_361[17] = buffer_data_1[2895:2888] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_361[18] = buffer_data_1[2903:2896] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_361[19] = buffer_data_1[2911:2904] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_361[20] = buffer_data_0[2879:2872] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_361[21] = buffer_data_0[2887:2880] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_361[22] = buffer_data_0[2895:2888] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_361[23] = buffer_data_0[2903:2896] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_361[24] = buffer_data_0[2911:2904] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_361 = kernel_img_mul_361[0] + kernel_img_mul_361[1] + kernel_img_mul_361[2] + 
                kernel_img_mul_361[3] + kernel_img_mul_361[4] + kernel_img_mul_361[5] + 
                kernel_img_mul_361[6] + kernel_img_mul_361[7] + kernel_img_mul_361[8] + 
                kernel_img_mul_361[9] + kernel_img_mul_361[10] + kernel_img_mul_361[11] + 
                kernel_img_mul_361[12] + kernel_img_mul_361[13] + kernel_img_mul_361[14] + 
                kernel_img_mul_361[15] + kernel_img_mul_361[16] + kernel_img_mul_361[17] + 
                kernel_img_mul_361[18] + kernel_img_mul_361[19] + kernel_img_mul_361[20] + 
                kernel_img_mul_361[21] + kernel_img_mul_361[22] + kernel_img_mul_361[23] + 
                kernel_img_mul_361[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2895:2888] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2895:2888] <= kernel_img_sum_361[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2895:2888] <= 'd0;
end

wire  [39:0]  kernel_img_mul_362[0:24];
assign kernel_img_mul_362[0] = buffer_data_4[2887:2880] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_362[1] = buffer_data_4[2895:2888] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_362[2] = buffer_data_4[2903:2896] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_362[3] = buffer_data_4[2911:2904] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_362[4] = buffer_data_4[2919:2912] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_362[5] = buffer_data_3[2887:2880] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_362[6] = buffer_data_3[2895:2888] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_362[7] = buffer_data_3[2903:2896] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_362[8] = buffer_data_3[2911:2904] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_362[9] = buffer_data_3[2919:2912] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_362[10] = buffer_data_2[2887:2880] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_362[11] = buffer_data_2[2895:2888] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_362[12] = buffer_data_2[2903:2896] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_362[13] = buffer_data_2[2911:2904] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_362[14] = buffer_data_2[2919:2912] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_362[15] = buffer_data_1[2887:2880] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_362[16] = buffer_data_1[2895:2888] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_362[17] = buffer_data_1[2903:2896] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_362[18] = buffer_data_1[2911:2904] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_362[19] = buffer_data_1[2919:2912] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_362[20] = buffer_data_0[2887:2880] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_362[21] = buffer_data_0[2895:2888] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_362[22] = buffer_data_0[2903:2896] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_362[23] = buffer_data_0[2911:2904] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_362[24] = buffer_data_0[2919:2912] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_362 = kernel_img_mul_362[0] + kernel_img_mul_362[1] + kernel_img_mul_362[2] + 
                kernel_img_mul_362[3] + kernel_img_mul_362[4] + kernel_img_mul_362[5] + 
                kernel_img_mul_362[6] + kernel_img_mul_362[7] + kernel_img_mul_362[8] + 
                kernel_img_mul_362[9] + kernel_img_mul_362[10] + kernel_img_mul_362[11] + 
                kernel_img_mul_362[12] + kernel_img_mul_362[13] + kernel_img_mul_362[14] + 
                kernel_img_mul_362[15] + kernel_img_mul_362[16] + kernel_img_mul_362[17] + 
                kernel_img_mul_362[18] + kernel_img_mul_362[19] + kernel_img_mul_362[20] + 
                kernel_img_mul_362[21] + kernel_img_mul_362[22] + kernel_img_mul_362[23] + 
                kernel_img_mul_362[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2903:2896] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2903:2896] <= kernel_img_sum_362[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2903:2896] <= 'd0;
end

wire  [39:0]  kernel_img_mul_363[0:24];
assign kernel_img_mul_363[0] = buffer_data_4[2895:2888] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_363[1] = buffer_data_4[2903:2896] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_363[2] = buffer_data_4[2911:2904] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_363[3] = buffer_data_4[2919:2912] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_363[4] = buffer_data_4[2927:2920] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_363[5] = buffer_data_3[2895:2888] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_363[6] = buffer_data_3[2903:2896] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_363[7] = buffer_data_3[2911:2904] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_363[8] = buffer_data_3[2919:2912] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_363[9] = buffer_data_3[2927:2920] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_363[10] = buffer_data_2[2895:2888] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_363[11] = buffer_data_2[2903:2896] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_363[12] = buffer_data_2[2911:2904] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_363[13] = buffer_data_2[2919:2912] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_363[14] = buffer_data_2[2927:2920] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_363[15] = buffer_data_1[2895:2888] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_363[16] = buffer_data_1[2903:2896] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_363[17] = buffer_data_1[2911:2904] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_363[18] = buffer_data_1[2919:2912] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_363[19] = buffer_data_1[2927:2920] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_363[20] = buffer_data_0[2895:2888] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_363[21] = buffer_data_0[2903:2896] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_363[22] = buffer_data_0[2911:2904] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_363[23] = buffer_data_0[2919:2912] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_363[24] = buffer_data_0[2927:2920] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_363 = kernel_img_mul_363[0] + kernel_img_mul_363[1] + kernel_img_mul_363[2] + 
                kernel_img_mul_363[3] + kernel_img_mul_363[4] + kernel_img_mul_363[5] + 
                kernel_img_mul_363[6] + kernel_img_mul_363[7] + kernel_img_mul_363[8] + 
                kernel_img_mul_363[9] + kernel_img_mul_363[10] + kernel_img_mul_363[11] + 
                kernel_img_mul_363[12] + kernel_img_mul_363[13] + kernel_img_mul_363[14] + 
                kernel_img_mul_363[15] + kernel_img_mul_363[16] + kernel_img_mul_363[17] + 
                kernel_img_mul_363[18] + kernel_img_mul_363[19] + kernel_img_mul_363[20] + 
                kernel_img_mul_363[21] + kernel_img_mul_363[22] + kernel_img_mul_363[23] + 
                kernel_img_mul_363[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2911:2904] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2911:2904] <= kernel_img_sum_363[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2911:2904] <= 'd0;
end

wire  [39:0]  kernel_img_mul_364[0:24];
assign kernel_img_mul_364[0] = buffer_data_4[2903:2896] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_364[1] = buffer_data_4[2911:2904] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_364[2] = buffer_data_4[2919:2912] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_364[3] = buffer_data_4[2927:2920] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_364[4] = buffer_data_4[2935:2928] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_364[5] = buffer_data_3[2903:2896] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_364[6] = buffer_data_3[2911:2904] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_364[7] = buffer_data_3[2919:2912] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_364[8] = buffer_data_3[2927:2920] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_364[9] = buffer_data_3[2935:2928] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_364[10] = buffer_data_2[2903:2896] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_364[11] = buffer_data_2[2911:2904] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_364[12] = buffer_data_2[2919:2912] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_364[13] = buffer_data_2[2927:2920] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_364[14] = buffer_data_2[2935:2928] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_364[15] = buffer_data_1[2903:2896] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_364[16] = buffer_data_1[2911:2904] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_364[17] = buffer_data_1[2919:2912] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_364[18] = buffer_data_1[2927:2920] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_364[19] = buffer_data_1[2935:2928] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_364[20] = buffer_data_0[2903:2896] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_364[21] = buffer_data_0[2911:2904] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_364[22] = buffer_data_0[2919:2912] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_364[23] = buffer_data_0[2927:2920] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_364[24] = buffer_data_0[2935:2928] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_364 = kernel_img_mul_364[0] + kernel_img_mul_364[1] + kernel_img_mul_364[2] + 
                kernel_img_mul_364[3] + kernel_img_mul_364[4] + kernel_img_mul_364[5] + 
                kernel_img_mul_364[6] + kernel_img_mul_364[7] + kernel_img_mul_364[8] + 
                kernel_img_mul_364[9] + kernel_img_mul_364[10] + kernel_img_mul_364[11] + 
                kernel_img_mul_364[12] + kernel_img_mul_364[13] + kernel_img_mul_364[14] + 
                kernel_img_mul_364[15] + kernel_img_mul_364[16] + kernel_img_mul_364[17] + 
                kernel_img_mul_364[18] + kernel_img_mul_364[19] + kernel_img_mul_364[20] + 
                kernel_img_mul_364[21] + kernel_img_mul_364[22] + kernel_img_mul_364[23] + 
                kernel_img_mul_364[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2919:2912] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2919:2912] <= kernel_img_sum_364[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2919:2912] <= 'd0;
end

wire  [39:0]  kernel_img_mul_365[0:24];
assign kernel_img_mul_365[0] = buffer_data_4[2911:2904] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_365[1] = buffer_data_4[2919:2912] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_365[2] = buffer_data_4[2927:2920] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_365[3] = buffer_data_4[2935:2928] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_365[4] = buffer_data_4[2943:2936] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_365[5] = buffer_data_3[2911:2904] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_365[6] = buffer_data_3[2919:2912] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_365[7] = buffer_data_3[2927:2920] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_365[8] = buffer_data_3[2935:2928] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_365[9] = buffer_data_3[2943:2936] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_365[10] = buffer_data_2[2911:2904] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_365[11] = buffer_data_2[2919:2912] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_365[12] = buffer_data_2[2927:2920] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_365[13] = buffer_data_2[2935:2928] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_365[14] = buffer_data_2[2943:2936] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_365[15] = buffer_data_1[2911:2904] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_365[16] = buffer_data_1[2919:2912] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_365[17] = buffer_data_1[2927:2920] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_365[18] = buffer_data_1[2935:2928] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_365[19] = buffer_data_1[2943:2936] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_365[20] = buffer_data_0[2911:2904] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_365[21] = buffer_data_0[2919:2912] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_365[22] = buffer_data_0[2927:2920] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_365[23] = buffer_data_0[2935:2928] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_365[24] = buffer_data_0[2943:2936] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_365 = kernel_img_mul_365[0] + kernel_img_mul_365[1] + kernel_img_mul_365[2] + 
                kernel_img_mul_365[3] + kernel_img_mul_365[4] + kernel_img_mul_365[5] + 
                kernel_img_mul_365[6] + kernel_img_mul_365[7] + kernel_img_mul_365[8] + 
                kernel_img_mul_365[9] + kernel_img_mul_365[10] + kernel_img_mul_365[11] + 
                kernel_img_mul_365[12] + kernel_img_mul_365[13] + kernel_img_mul_365[14] + 
                kernel_img_mul_365[15] + kernel_img_mul_365[16] + kernel_img_mul_365[17] + 
                kernel_img_mul_365[18] + kernel_img_mul_365[19] + kernel_img_mul_365[20] + 
                kernel_img_mul_365[21] + kernel_img_mul_365[22] + kernel_img_mul_365[23] + 
                kernel_img_mul_365[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2927:2920] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2927:2920] <= kernel_img_sum_365[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2927:2920] <= 'd0;
end

wire  [39:0]  kernel_img_mul_366[0:24];
assign kernel_img_mul_366[0] = buffer_data_4[2919:2912] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_366[1] = buffer_data_4[2927:2920] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_366[2] = buffer_data_4[2935:2928] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_366[3] = buffer_data_4[2943:2936] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_366[4] = buffer_data_4[2951:2944] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_366[5] = buffer_data_3[2919:2912] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_366[6] = buffer_data_3[2927:2920] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_366[7] = buffer_data_3[2935:2928] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_366[8] = buffer_data_3[2943:2936] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_366[9] = buffer_data_3[2951:2944] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_366[10] = buffer_data_2[2919:2912] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_366[11] = buffer_data_2[2927:2920] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_366[12] = buffer_data_2[2935:2928] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_366[13] = buffer_data_2[2943:2936] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_366[14] = buffer_data_2[2951:2944] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_366[15] = buffer_data_1[2919:2912] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_366[16] = buffer_data_1[2927:2920] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_366[17] = buffer_data_1[2935:2928] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_366[18] = buffer_data_1[2943:2936] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_366[19] = buffer_data_1[2951:2944] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_366[20] = buffer_data_0[2919:2912] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_366[21] = buffer_data_0[2927:2920] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_366[22] = buffer_data_0[2935:2928] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_366[23] = buffer_data_0[2943:2936] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_366[24] = buffer_data_0[2951:2944] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_366 = kernel_img_mul_366[0] + kernel_img_mul_366[1] + kernel_img_mul_366[2] + 
                kernel_img_mul_366[3] + kernel_img_mul_366[4] + kernel_img_mul_366[5] + 
                kernel_img_mul_366[6] + kernel_img_mul_366[7] + kernel_img_mul_366[8] + 
                kernel_img_mul_366[9] + kernel_img_mul_366[10] + kernel_img_mul_366[11] + 
                kernel_img_mul_366[12] + kernel_img_mul_366[13] + kernel_img_mul_366[14] + 
                kernel_img_mul_366[15] + kernel_img_mul_366[16] + kernel_img_mul_366[17] + 
                kernel_img_mul_366[18] + kernel_img_mul_366[19] + kernel_img_mul_366[20] + 
                kernel_img_mul_366[21] + kernel_img_mul_366[22] + kernel_img_mul_366[23] + 
                kernel_img_mul_366[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2935:2928] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2935:2928] <= kernel_img_sum_366[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2935:2928] <= 'd0;
end

wire  [39:0]  kernel_img_mul_367[0:24];
assign kernel_img_mul_367[0] = buffer_data_4[2927:2920] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_367[1] = buffer_data_4[2935:2928] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_367[2] = buffer_data_4[2943:2936] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_367[3] = buffer_data_4[2951:2944] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_367[4] = buffer_data_4[2959:2952] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_367[5] = buffer_data_3[2927:2920] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_367[6] = buffer_data_3[2935:2928] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_367[7] = buffer_data_3[2943:2936] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_367[8] = buffer_data_3[2951:2944] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_367[9] = buffer_data_3[2959:2952] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_367[10] = buffer_data_2[2927:2920] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_367[11] = buffer_data_2[2935:2928] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_367[12] = buffer_data_2[2943:2936] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_367[13] = buffer_data_2[2951:2944] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_367[14] = buffer_data_2[2959:2952] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_367[15] = buffer_data_1[2927:2920] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_367[16] = buffer_data_1[2935:2928] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_367[17] = buffer_data_1[2943:2936] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_367[18] = buffer_data_1[2951:2944] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_367[19] = buffer_data_1[2959:2952] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_367[20] = buffer_data_0[2927:2920] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_367[21] = buffer_data_0[2935:2928] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_367[22] = buffer_data_0[2943:2936] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_367[23] = buffer_data_0[2951:2944] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_367[24] = buffer_data_0[2959:2952] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_367 = kernel_img_mul_367[0] + kernel_img_mul_367[1] + kernel_img_mul_367[2] + 
                kernel_img_mul_367[3] + kernel_img_mul_367[4] + kernel_img_mul_367[5] + 
                kernel_img_mul_367[6] + kernel_img_mul_367[7] + kernel_img_mul_367[8] + 
                kernel_img_mul_367[9] + kernel_img_mul_367[10] + kernel_img_mul_367[11] + 
                kernel_img_mul_367[12] + kernel_img_mul_367[13] + kernel_img_mul_367[14] + 
                kernel_img_mul_367[15] + kernel_img_mul_367[16] + kernel_img_mul_367[17] + 
                kernel_img_mul_367[18] + kernel_img_mul_367[19] + kernel_img_mul_367[20] + 
                kernel_img_mul_367[21] + kernel_img_mul_367[22] + kernel_img_mul_367[23] + 
                kernel_img_mul_367[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2943:2936] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2943:2936] <= kernel_img_sum_367[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2943:2936] <= 'd0;
end

wire  [39:0]  kernel_img_mul_368[0:24];
assign kernel_img_mul_368[0] = buffer_data_4[2935:2928] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_368[1] = buffer_data_4[2943:2936] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_368[2] = buffer_data_4[2951:2944] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_368[3] = buffer_data_4[2959:2952] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_368[4] = buffer_data_4[2967:2960] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_368[5] = buffer_data_3[2935:2928] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_368[6] = buffer_data_3[2943:2936] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_368[7] = buffer_data_3[2951:2944] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_368[8] = buffer_data_3[2959:2952] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_368[9] = buffer_data_3[2967:2960] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_368[10] = buffer_data_2[2935:2928] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_368[11] = buffer_data_2[2943:2936] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_368[12] = buffer_data_2[2951:2944] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_368[13] = buffer_data_2[2959:2952] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_368[14] = buffer_data_2[2967:2960] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_368[15] = buffer_data_1[2935:2928] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_368[16] = buffer_data_1[2943:2936] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_368[17] = buffer_data_1[2951:2944] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_368[18] = buffer_data_1[2959:2952] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_368[19] = buffer_data_1[2967:2960] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_368[20] = buffer_data_0[2935:2928] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_368[21] = buffer_data_0[2943:2936] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_368[22] = buffer_data_0[2951:2944] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_368[23] = buffer_data_0[2959:2952] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_368[24] = buffer_data_0[2967:2960] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_368 = kernel_img_mul_368[0] + kernel_img_mul_368[1] + kernel_img_mul_368[2] + 
                kernel_img_mul_368[3] + kernel_img_mul_368[4] + kernel_img_mul_368[5] + 
                kernel_img_mul_368[6] + kernel_img_mul_368[7] + kernel_img_mul_368[8] + 
                kernel_img_mul_368[9] + kernel_img_mul_368[10] + kernel_img_mul_368[11] + 
                kernel_img_mul_368[12] + kernel_img_mul_368[13] + kernel_img_mul_368[14] + 
                kernel_img_mul_368[15] + kernel_img_mul_368[16] + kernel_img_mul_368[17] + 
                kernel_img_mul_368[18] + kernel_img_mul_368[19] + kernel_img_mul_368[20] + 
                kernel_img_mul_368[21] + kernel_img_mul_368[22] + kernel_img_mul_368[23] + 
                kernel_img_mul_368[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2951:2944] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2951:2944] <= kernel_img_sum_368[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2951:2944] <= 'd0;
end

wire  [39:0]  kernel_img_mul_369[0:24];
assign kernel_img_mul_369[0] = buffer_data_4[2943:2936] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_369[1] = buffer_data_4[2951:2944] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_369[2] = buffer_data_4[2959:2952] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_369[3] = buffer_data_4[2967:2960] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_369[4] = buffer_data_4[2975:2968] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_369[5] = buffer_data_3[2943:2936] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_369[6] = buffer_data_3[2951:2944] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_369[7] = buffer_data_3[2959:2952] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_369[8] = buffer_data_3[2967:2960] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_369[9] = buffer_data_3[2975:2968] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_369[10] = buffer_data_2[2943:2936] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_369[11] = buffer_data_2[2951:2944] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_369[12] = buffer_data_2[2959:2952] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_369[13] = buffer_data_2[2967:2960] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_369[14] = buffer_data_2[2975:2968] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_369[15] = buffer_data_1[2943:2936] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_369[16] = buffer_data_1[2951:2944] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_369[17] = buffer_data_1[2959:2952] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_369[18] = buffer_data_1[2967:2960] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_369[19] = buffer_data_1[2975:2968] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_369[20] = buffer_data_0[2943:2936] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_369[21] = buffer_data_0[2951:2944] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_369[22] = buffer_data_0[2959:2952] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_369[23] = buffer_data_0[2967:2960] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_369[24] = buffer_data_0[2975:2968] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_369 = kernel_img_mul_369[0] + kernel_img_mul_369[1] + kernel_img_mul_369[2] + 
                kernel_img_mul_369[3] + kernel_img_mul_369[4] + kernel_img_mul_369[5] + 
                kernel_img_mul_369[6] + kernel_img_mul_369[7] + kernel_img_mul_369[8] + 
                kernel_img_mul_369[9] + kernel_img_mul_369[10] + kernel_img_mul_369[11] + 
                kernel_img_mul_369[12] + kernel_img_mul_369[13] + kernel_img_mul_369[14] + 
                kernel_img_mul_369[15] + kernel_img_mul_369[16] + kernel_img_mul_369[17] + 
                kernel_img_mul_369[18] + kernel_img_mul_369[19] + kernel_img_mul_369[20] + 
                kernel_img_mul_369[21] + kernel_img_mul_369[22] + kernel_img_mul_369[23] + 
                kernel_img_mul_369[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2959:2952] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2959:2952] <= kernel_img_sum_369[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2959:2952] <= 'd0;
end

wire  [39:0]  kernel_img_mul_370[0:24];
assign kernel_img_mul_370[0] = buffer_data_4[2951:2944] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_370[1] = buffer_data_4[2959:2952] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_370[2] = buffer_data_4[2967:2960] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_370[3] = buffer_data_4[2975:2968] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_370[4] = buffer_data_4[2983:2976] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_370[5] = buffer_data_3[2951:2944] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_370[6] = buffer_data_3[2959:2952] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_370[7] = buffer_data_3[2967:2960] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_370[8] = buffer_data_3[2975:2968] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_370[9] = buffer_data_3[2983:2976] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_370[10] = buffer_data_2[2951:2944] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_370[11] = buffer_data_2[2959:2952] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_370[12] = buffer_data_2[2967:2960] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_370[13] = buffer_data_2[2975:2968] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_370[14] = buffer_data_2[2983:2976] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_370[15] = buffer_data_1[2951:2944] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_370[16] = buffer_data_1[2959:2952] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_370[17] = buffer_data_1[2967:2960] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_370[18] = buffer_data_1[2975:2968] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_370[19] = buffer_data_1[2983:2976] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_370[20] = buffer_data_0[2951:2944] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_370[21] = buffer_data_0[2959:2952] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_370[22] = buffer_data_0[2967:2960] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_370[23] = buffer_data_0[2975:2968] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_370[24] = buffer_data_0[2983:2976] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_370 = kernel_img_mul_370[0] + kernel_img_mul_370[1] + kernel_img_mul_370[2] + 
                kernel_img_mul_370[3] + kernel_img_mul_370[4] + kernel_img_mul_370[5] + 
                kernel_img_mul_370[6] + kernel_img_mul_370[7] + kernel_img_mul_370[8] + 
                kernel_img_mul_370[9] + kernel_img_mul_370[10] + kernel_img_mul_370[11] + 
                kernel_img_mul_370[12] + kernel_img_mul_370[13] + kernel_img_mul_370[14] + 
                kernel_img_mul_370[15] + kernel_img_mul_370[16] + kernel_img_mul_370[17] + 
                kernel_img_mul_370[18] + kernel_img_mul_370[19] + kernel_img_mul_370[20] + 
                kernel_img_mul_370[21] + kernel_img_mul_370[22] + kernel_img_mul_370[23] + 
                kernel_img_mul_370[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2967:2960] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2967:2960] <= kernel_img_sum_370[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2967:2960] <= 'd0;
end

wire  [39:0]  kernel_img_mul_371[0:24];
assign kernel_img_mul_371[0] = buffer_data_4[2959:2952] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_371[1] = buffer_data_4[2967:2960] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_371[2] = buffer_data_4[2975:2968] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_371[3] = buffer_data_4[2983:2976] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_371[4] = buffer_data_4[2991:2984] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_371[5] = buffer_data_3[2959:2952] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_371[6] = buffer_data_3[2967:2960] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_371[7] = buffer_data_3[2975:2968] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_371[8] = buffer_data_3[2983:2976] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_371[9] = buffer_data_3[2991:2984] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_371[10] = buffer_data_2[2959:2952] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_371[11] = buffer_data_2[2967:2960] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_371[12] = buffer_data_2[2975:2968] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_371[13] = buffer_data_2[2983:2976] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_371[14] = buffer_data_2[2991:2984] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_371[15] = buffer_data_1[2959:2952] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_371[16] = buffer_data_1[2967:2960] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_371[17] = buffer_data_1[2975:2968] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_371[18] = buffer_data_1[2983:2976] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_371[19] = buffer_data_1[2991:2984] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_371[20] = buffer_data_0[2959:2952] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_371[21] = buffer_data_0[2967:2960] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_371[22] = buffer_data_0[2975:2968] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_371[23] = buffer_data_0[2983:2976] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_371[24] = buffer_data_0[2991:2984] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_371 = kernel_img_mul_371[0] + kernel_img_mul_371[1] + kernel_img_mul_371[2] + 
                kernel_img_mul_371[3] + kernel_img_mul_371[4] + kernel_img_mul_371[5] + 
                kernel_img_mul_371[6] + kernel_img_mul_371[7] + kernel_img_mul_371[8] + 
                kernel_img_mul_371[9] + kernel_img_mul_371[10] + kernel_img_mul_371[11] + 
                kernel_img_mul_371[12] + kernel_img_mul_371[13] + kernel_img_mul_371[14] + 
                kernel_img_mul_371[15] + kernel_img_mul_371[16] + kernel_img_mul_371[17] + 
                kernel_img_mul_371[18] + kernel_img_mul_371[19] + kernel_img_mul_371[20] + 
                kernel_img_mul_371[21] + kernel_img_mul_371[22] + kernel_img_mul_371[23] + 
                kernel_img_mul_371[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2975:2968] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2975:2968] <= kernel_img_sum_371[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2975:2968] <= 'd0;
end

wire  [39:0]  kernel_img_mul_372[0:24];
assign kernel_img_mul_372[0] = buffer_data_4[2967:2960] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_372[1] = buffer_data_4[2975:2968] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_372[2] = buffer_data_4[2983:2976] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_372[3] = buffer_data_4[2991:2984] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_372[4] = buffer_data_4[2999:2992] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_372[5] = buffer_data_3[2967:2960] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_372[6] = buffer_data_3[2975:2968] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_372[7] = buffer_data_3[2983:2976] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_372[8] = buffer_data_3[2991:2984] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_372[9] = buffer_data_3[2999:2992] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_372[10] = buffer_data_2[2967:2960] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_372[11] = buffer_data_2[2975:2968] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_372[12] = buffer_data_2[2983:2976] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_372[13] = buffer_data_2[2991:2984] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_372[14] = buffer_data_2[2999:2992] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_372[15] = buffer_data_1[2967:2960] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_372[16] = buffer_data_1[2975:2968] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_372[17] = buffer_data_1[2983:2976] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_372[18] = buffer_data_1[2991:2984] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_372[19] = buffer_data_1[2999:2992] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_372[20] = buffer_data_0[2967:2960] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_372[21] = buffer_data_0[2975:2968] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_372[22] = buffer_data_0[2983:2976] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_372[23] = buffer_data_0[2991:2984] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_372[24] = buffer_data_0[2999:2992] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_372 = kernel_img_mul_372[0] + kernel_img_mul_372[1] + kernel_img_mul_372[2] + 
                kernel_img_mul_372[3] + kernel_img_mul_372[4] + kernel_img_mul_372[5] + 
                kernel_img_mul_372[6] + kernel_img_mul_372[7] + kernel_img_mul_372[8] + 
                kernel_img_mul_372[9] + kernel_img_mul_372[10] + kernel_img_mul_372[11] + 
                kernel_img_mul_372[12] + kernel_img_mul_372[13] + kernel_img_mul_372[14] + 
                kernel_img_mul_372[15] + kernel_img_mul_372[16] + kernel_img_mul_372[17] + 
                kernel_img_mul_372[18] + kernel_img_mul_372[19] + kernel_img_mul_372[20] + 
                kernel_img_mul_372[21] + kernel_img_mul_372[22] + kernel_img_mul_372[23] + 
                kernel_img_mul_372[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2983:2976] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2983:2976] <= kernel_img_sum_372[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2983:2976] <= 'd0;
end

wire  [39:0]  kernel_img_mul_373[0:24];
assign kernel_img_mul_373[0] = buffer_data_4[2975:2968] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_373[1] = buffer_data_4[2983:2976] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_373[2] = buffer_data_4[2991:2984] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_373[3] = buffer_data_4[2999:2992] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_373[4] = buffer_data_4[3007:3000] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_373[5] = buffer_data_3[2975:2968] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_373[6] = buffer_data_3[2983:2976] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_373[7] = buffer_data_3[2991:2984] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_373[8] = buffer_data_3[2999:2992] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_373[9] = buffer_data_3[3007:3000] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_373[10] = buffer_data_2[2975:2968] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_373[11] = buffer_data_2[2983:2976] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_373[12] = buffer_data_2[2991:2984] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_373[13] = buffer_data_2[2999:2992] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_373[14] = buffer_data_2[3007:3000] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_373[15] = buffer_data_1[2975:2968] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_373[16] = buffer_data_1[2983:2976] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_373[17] = buffer_data_1[2991:2984] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_373[18] = buffer_data_1[2999:2992] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_373[19] = buffer_data_1[3007:3000] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_373[20] = buffer_data_0[2975:2968] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_373[21] = buffer_data_0[2983:2976] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_373[22] = buffer_data_0[2991:2984] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_373[23] = buffer_data_0[2999:2992] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_373[24] = buffer_data_0[3007:3000] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_373 = kernel_img_mul_373[0] + kernel_img_mul_373[1] + kernel_img_mul_373[2] + 
                kernel_img_mul_373[3] + kernel_img_mul_373[4] + kernel_img_mul_373[5] + 
                kernel_img_mul_373[6] + kernel_img_mul_373[7] + kernel_img_mul_373[8] + 
                kernel_img_mul_373[9] + kernel_img_mul_373[10] + kernel_img_mul_373[11] + 
                kernel_img_mul_373[12] + kernel_img_mul_373[13] + kernel_img_mul_373[14] + 
                kernel_img_mul_373[15] + kernel_img_mul_373[16] + kernel_img_mul_373[17] + 
                kernel_img_mul_373[18] + kernel_img_mul_373[19] + kernel_img_mul_373[20] + 
                kernel_img_mul_373[21] + kernel_img_mul_373[22] + kernel_img_mul_373[23] + 
                kernel_img_mul_373[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2991:2984] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2991:2984] <= kernel_img_sum_373[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2991:2984] <= 'd0;
end

wire  [39:0]  kernel_img_mul_374[0:24];
assign kernel_img_mul_374[0] = buffer_data_4[2983:2976] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_374[1] = buffer_data_4[2991:2984] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_374[2] = buffer_data_4[2999:2992] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_374[3] = buffer_data_4[3007:3000] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_374[4] = buffer_data_4[3015:3008] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_374[5] = buffer_data_3[2983:2976] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_374[6] = buffer_data_3[2991:2984] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_374[7] = buffer_data_3[2999:2992] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_374[8] = buffer_data_3[3007:3000] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_374[9] = buffer_data_3[3015:3008] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_374[10] = buffer_data_2[2983:2976] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_374[11] = buffer_data_2[2991:2984] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_374[12] = buffer_data_2[2999:2992] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_374[13] = buffer_data_2[3007:3000] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_374[14] = buffer_data_2[3015:3008] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_374[15] = buffer_data_1[2983:2976] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_374[16] = buffer_data_1[2991:2984] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_374[17] = buffer_data_1[2999:2992] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_374[18] = buffer_data_1[3007:3000] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_374[19] = buffer_data_1[3015:3008] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_374[20] = buffer_data_0[2983:2976] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_374[21] = buffer_data_0[2991:2984] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_374[22] = buffer_data_0[2999:2992] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_374[23] = buffer_data_0[3007:3000] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_374[24] = buffer_data_0[3015:3008] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_374 = kernel_img_mul_374[0] + kernel_img_mul_374[1] + kernel_img_mul_374[2] + 
                kernel_img_mul_374[3] + kernel_img_mul_374[4] + kernel_img_mul_374[5] + 
                kernel_img_mul_374[6] + kernel_img_mul_374[7] + kernel_img_mul_374[8] + 
                kernel_img_mul_374[9] + kernel_img_mul_374[10] + kernel_img_mul_374[11] + 
                kernel_img_mul_374[12] + kernel_img_mul_374[13] + kernel_img_mul_374[14] + 
                kernel_img_mul_374[15] + kernel_img_mul_374[16] + kernel_img_mul_374[17] + 
                kernel_img_mul_374[18] + kernel_img_mul_374[19] + kernel_img_mul_374[20] + 
                kernel_img_mul_374[21] + kernel_img_mul_374[22] + kernel_img_mul_374[23] + 
                kernel_img_mul_374[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[2999:2992] <= 'd0;
  else if (current_state==ST_START)
    blur_din[2999:2992] <= kernel_img_sum_374[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2999:2992] <= 'd0;
end

wire  [39:0]  kernel_img_mul_375[0:24];
assign kernel_img_mul_375[0] = buffer_data_4[2991:2984] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_375[1] = buffer_data_4[2999:2992] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_375[2] = buffer_data_4[3007:3000] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_375[3] = buffer_data_4[3015:3008] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_375[4] = buffer_data_4[3023:3016] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_375[5] = buffer_data_3[2991:2984] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_375[6] = buffer_data_3[2999:2992] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_375[7] = buffer_data_3[3007:3000] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_375[8] = buffer_data_3[3015:3008] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_375[9] = buffer_data_3[3023:3016] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_375[10] = buffer_data_2[2991:2984] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_375[11] = buffer_data_2[2999:2992] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_375[12] = buffer_data_2[3007:3000] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_375[13] = buffer_data_2[3015:3008] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_375[14] = buffer_data_2[3023:3016] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_375[15] = buffer_data_1[2991:2984] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_375[16] = buffer_data_1[2999:2992] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_375[17] = buffer_data_1[3007:3000] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_375[18] = buffer_data_1[3015:3008] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_375[19] = buffer_data_1[3023:3016] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_375[20] = buffer_data_0[2991:2984] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_375[21] = buffer_data_0[2999:2992] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_375[22] = buffer_data_0[3007:3000] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_375[23] = buffer_data_0[3015:3008] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_375[24] = buffer_data_0[3023:3016] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_375 = kernel_img_mul_375[0] + kernel_img_mul_375[1] + kernel_img_mul_375[2] + 
                kernel_img_mul_375[3] + kernel_img_mul_375[4] + kernel_img_mul_375[5] + 
                kernel_img_mul_375[6] + kernel_img_mul_375[7] + kernel_img_mul_375[8] + 
                kernel_img_mul_375[9] + kernel_img_mul_375[10] + kernel_img_mul_375[11] + 
                kernel_img_mul_375[12] + kernel_img_mul_375[13] + kernel_img_mul_375[14] + 
                kernel_img_mul_375[15] + kernel_img_mul_375[16] + kernel_img_mul_375[17] + 
                kernel_img_mul_375[18] + kernel_img_mul_375[19] + kernel_img_mul_375[20] + 
                kernel_img_mul_375[21] + kernel_img_mul_375[22] + kernel_img_mul_375[23] + 
                kernel_img_mul_375[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3007:3000] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3007:3000] <= kernel_img_sum_375[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3007:3000] <= 'd0;
end

wire  [39:0]  kernel_img_mul_376[0:24];
assign kernel_img_mul_376[0] = buffer_data_4[2999:2992] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_376[1] = buffer_data_4[3007:3000] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_376[2] = buffer_data_4[3015:3008] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_376[3] = buffer_data_4[3023:3016] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_376[4] = buffer_data_4[3031:3024] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_376[5] = buffer_data_3[2999:2992] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_376[6] = buffer_data_3[3007:3000] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_376[7] = buffer_data_3[3015:3008] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_376[8] = buffer_data_3[3023:3016] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_376[9] = buffer_data_3[3031:3024] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_376[10] = buffer_data_2[2999:2992] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_376[11] = buffer_data_2[3007:3000] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_376[12] = buffer_data_2[3015:3008] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_376[13] = buffer_data_2[3023:3016] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_376[14] = buffer_data_2[3031:3024] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_376[15] = buffer_data_1[2999:2992] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_376[16] = buffer_data_1[3007:3000] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_376[17] = buffer_data_1[3015:3008] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_376[18] = buffer_data_1[3023:3016] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_376[19] = buffer_data_1[3031:3024] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_376[20] = buffer_data_0[2999:2992] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_376[21] = buffer_data_0[3007:3000] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_376[22] = buffer_data_0[3015:3008] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_376[23] = buffer_data_0[3023:3016] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_376[24] = buffer_data_0[3031:3024] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_376 = kernel_img_mul_376[0] + kernel_img_mul_376[1] + kernel_img_mul_376[2] + 
                kernel_img_mul_376[3] + kernel_img_mul_376[4] + kernel_img_mul_376[5] + 
                kernel_img_mul_376[6] + kernel_img_mul_376[7] + kernel_img_mul_376[8] + 
                kernel_img_mul_376[9] + kernel_img_mul_376[10] + kernel_img_mul_376[11] + 
                kernel_img_mul_376[12] + kernel_img_mul_376[13] + kernel_img_mul_376[14] + 
                kernel_img_mul_376[15] + kernel_img_mul_376[16] + kernel_img_mul_376[17] + 
                kernel_img_mul_376[18] + kernel_img_mul_376[19] + kernel_img_mul_376[20] + 
                kernel_img_mul_376[21] + kernel_img_mul_376[22] + kernel_img_mul_376[23] + 
                kernel_img_mul_376[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3015:3008] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3015:3008] <= kernel_img_sum_376[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3015:3008] <= 'd0;
end

wire  [39:0]  kernel_img_mul_377[0:24];
assign kernel_img_mul_377[0] = buffer_data_4[3007:3000] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_377[1] = buffer_data_4[3015:3008] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_377[2] = buffer_data_4[3023:3016] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_377[3] = buffer_data_4[3031:3024] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_377[4] = buffer_data_4[3039:3032] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_377[5] = buffer_data_3[3007:3000] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_377[6] = buffer_data_3[3015:3008] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_377[7] = buffer_data_3[3023:3016] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_377[8] = buffer_data_3[3031:3024] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_377[9] = buffer_data_3[3039:3032] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_377[10] = buffer_data_2[3007:3000] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_377[11] = buffer_data_2[3015:3008] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_377[12] = buffer_data_2[3023:3016] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_377[13] = buffer_data_2[3031:3024] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_377[14] = buffer_data_2[3039:3032] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_377[15] = buffer_data_1[3007:3000] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_377[16] = buffer_data_1[3015:3008] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_377[17] = buffer_data_1[3023:3016] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_377[18] = buffer_data_1[3031:3024] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_377[19] = buffer_data_1[3039:3032] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_377[20] = buffer_data_0[3007:3000] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_377[21] = buffer_data_0[3015:3008] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_377[22] = buffer_data_0[3023:3016] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_377[23] = buffer_data_0[3031:3024] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_377[24] = buffer_data_0[3039:3032] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_377 = kernel_img_mul_377[0] + kernel_img_mul_377[1] + kernel_img_mul_377[2] + 
                kernel_img_mul_377[3] + kernel_img_mul_377[4] + kernel_img_mul_377[5] + 
                kernel_img_mul_377[6] + kernel_img_mul_377[7] + kernel_img_mul_377[8] + 
                kernel_img_mul_377[9] + kernel_img_mul_377[10] + kernel_img_mul_377[11] + 
                kernel_img_mul_377[12] + kernel_img_mul_377[13] + kernel_img_mul_377[14] + 
                kernel_img_mul_377[15] + kernel_img_mul_377[16] + kernel_img_mul_377[17] + 
                kernel_img_mul_377[18] + kernel_img_mul_377[19] + kernel_img_mul_377[20] + 
                kernel_img_mul_377[21] + kernel_img_mul_377[22] + kernel_img_mul_377[23] + 
                kernel_img_mul_377[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3023:3016] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3023:3016] <= kernel_img_sum_377[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3023:3016] <= 'd0;
end

wire  [39:0]  kernel_img_mul_378[0:24];
assign kernel_img_mul_378[0] = buffer_data_4[3015:3008] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_378[1] = buffer_data_4[3023:3016] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_378[2] = buffer_data_4[3031:3024] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_378[3] = buffer_data_4[3039:3032] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_378[4] = buffer_data_4[3047:3040] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_378[5] = buffer_data_3[3015:3008] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_378[6] = buffer_data_3[3023:3016] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_378[7] = buffer_data_3[3031:3024] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_378[8] = buffer_data_3[3039:3032] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_378[9] = buffer_data_3[3047:3040] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_378[10] = buffer_data_2[3015:3008] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_378[11] = buffer_data_2[3023:3016] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_378[12] = buffer_data_2[3031:3024] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_378[13] = buffer_data_2[3039:3032] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_378[14] = buffer_data_2[3047:3040] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_378[15] = buffer_data_1[3015:3008] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_378[16] = buffer_data_1[3023:3016] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_378[17] = buffer_data_1[3031:3024] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_378[18] = buffer_data_1[3039:3032] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_378[19] = buffer_data_1[3047:3040] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_378[20] = buffer_data_0[3015:3008] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_378[21] = buffer_data_0[3023:3016] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_378[22] = buffer_data_0[3031:3024] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_378[23] = buffer_data_0[3039:3032] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_378[24] = buffer_data_0[3047:3040] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_378 = kernel_img_mul_378[0] + kernel_img_mul_378[1] + kernel_img_mul_378[2] + 
                kernel_img_mul_378[3] + kernel_img_mul_378[4] + kernel_img_mul_378[5] + 
                kernel_img_mul_378[6] + kernel_img_mul_378[7] + kernel_img_mul_378[8] + 
                kernel_img_mul_378[9] + kernel_img_mul_378[10] + kernel_img_mul_378[11] + 
                kernel_img_mul_378[12] + kernel_img_mul_378[13] + kernel_img_mul_378[14] + 
                kernel_img_mul_378[15] + kernel_img_mul_378[16] + kernel_img_mul_378[17] + 
                kernel_img_mul_378[18] + kernel_img_mul_378[19] + kernel_img_mul_378[20] + 
                kernel_img_mul_378[21] + kernel_img_mul_378[22] + kernel_img_mul_378[23] + 
                kernel_img_mul_378[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3031:3024] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3031:3024] <= kernel_img_sum_378[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3031:3024] <= 'd0;
end

wire  [39:0]  kernel_img_mul_379[0:24];
assign kernel_img_mul_379[0] = buffer_data_4[3023:3016] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_379[1] = buffer_data_4[3031:3024] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_379[2] = buffer_data_4[3039:3032] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_379[3] = buffer_data_4[3047:3040] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_379[4] = buffer_data_4[3055:3048] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_379[5] = buffer_data_3[3023:3016] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_379[6] = buffer_data_3[3031:3024] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_379[7] = buffer_data_3[3039:3032] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_379[8] = buffer_data_3[3047:3040] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_379[9] = buffer_data_3[3055:3048] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_379[10] = buffer_data_2[3023:3016] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_379[11] = buffer_data_2[3031:3024] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_379[12] = buffer_data_2[3039:3032] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_379[13] = buffer_data_2[3047:3040] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_379[14] = buffer_data_2[3055:3048] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_379[15] = buffer_data_1[3023:3016] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_379[16] = buffer_data_1[3031:3024] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_379[17] = buffer_data_1[3039:3032] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_379[18] = buffer_data_1[3047:3040] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_379[19] = buffer_data_1[3055:3048] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_379[20] = buffer_data_0[3023:3016] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_379[21] = buffer_data_0[3031:3024] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_379[22] = buffer_data_0[3039:3032] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_379[23] = buffer_data_0[3047:3040] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_379[24] = buffer_data_0[3055:3048] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_379 = kernel_img_mul_379[0] + kernel_img_mul_379[1] + kernel_img_mul_379[2] + 
                kernel_img_mul_379[3] + kernel_img_mul_379[4] + kernel_img_mul_379[5] + 
                kernel_img_mul_379[6] + kernel_img_mul_379[7] + kernel_img_mul_379[8] + 
                kernel_img_mul_379[9] + kernel_img_mul_379[10] + kernel_img_mul_379[11] + 
                kernel_img_mul_379[12] + kernel_img_mul_379[13] + kernel_img_mul_379[14] + 
                kernel_img_mul_379[15] + kernel_img_mul_379[16] + kernel_img_mul_379[17] + 
                kernel_img_mul_379[18] + kernel_img_mul_379[19] + kernel_img_mul_379[20] + 
                kernel_img_mul_379[21] + kernel_img_mul_379[22] + kernel_img_mul_379[23] + 
                kernel_img_mul_379[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3039:3032] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3039:3032] <= kernel_img_sum_379[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3039:3032] <= 'd0;
end

wire  [39:0]  kernel_img_mul_380[0:24];
assign kernel_img_mul_380[0] = buffer_data_4[3031:3024] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_380[1] = buffer_data_4[3039:3032] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_380[2] = buffer_data_4[3047:3040] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_380[3] = buffer_data_4[3055:3048] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_380[4] = buffer_data_4[3063:3056] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_380[5] = buffer_data_3[3031:3024] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_380[6] = buffer_data_3[3039:3032] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_380[7] = buffer_data_3[3047:3040] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_380[8] = buffer_data_3[3055:3048] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_380[9] = buffer_data_3[3063:3056] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_380[10] = buffer_data_2[3031:3024] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_380[11] = buffer_data_2[3039:3032] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_380[12] = buffer_data_2[3047:3040] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_380[13] = buffer_data_2[3055:3048] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_380[14] = buffer_data_2[3063:3056] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_380[15] = buffer_data_1[3031:3024] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_380[16] = buffer_data_1[3039:3032] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_380[17] = buffer_data_1[3047:3040] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_380[18] = buffer_data_1[3055:3048] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_380[19] = buffer_data_1[3063:3056] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_380[20] = buffer_data_0[3031:3024] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_380[21] = buffer_data_0[3039:3032] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_380[22] = buffer_data_0[3047:3040] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_380[23] = buffer_data_0[3055:3048] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_380[24] = buffer_data_0[3063:3056] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_380 = kernel_img_mul_380[0] + kernel_img_mul_380[1] + kernel_img_mul_380[2] + 
                kernel_img_mul_380[3] + kernel_img_mul_380[4] + kernel_img_mul_380[5] + 
                kernel_img_mul_380[6] + kernel_img_mul_380[7] + kernel_img_mul_380[8] + 
                kernel_img_mul_380[9] + kernel_img_mul_380[10] + kernel_img_mul_380[11] + 
                kernel_img_mul_380[12] + kernel_img_mul_380[13] + kernel_img_mul_380[14] + 
                kernel_img_mul_380[15] + kernel_img_mul_380[16] + kernel_img_mul_380[17] + 
                kernel_img_mul_380[18] + kernel_img_mul_380[19] + kernel_img_mul_380[20] + 
                kernel_img_mul_380[21] + kernel_img_mul_380[22] + kernel_img_mul_380[23] + 
                kernel_img_mul_380[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3047:3040] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3047:3040] <= kernel_img_sum_380[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3047:3040] <= 'd0;
end

wire  [39:0]  kernel_img_mul_381[0:24];
assign kernel_img_mul_381[0] = buffer_data_4[3039:3032] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_381[1] = buffer_data_4[3047:3040] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_381[2] = buffer_data_4[3055:3048] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_381[3] = buffer_data_4[3063:3056] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_381[4] = buffer_data_4[3071:3064] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_381[5] = buffer_data_3[3039:3032] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_381[6] = buffer_data_3[3047:3040] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_381[7] = buffer_data_3[3055:3048] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_381[8] = buffer_data_3[3063:3056] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_381[9] = buffer_data_3[3071:3064] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_381[10] = buffer_data_2[3039:3032] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_381[11] = buffer_data_2[3047:3040] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_381[12] = buffer_data_2[3055:3048] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_381[13] = buffer_data_2[3063:3056] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_381[14] = buffer_data_2[3071:3064] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_381[15] = buffer_data_1[3039:3032] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_381[16] = buffer_data_1[3047:3040] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_381[17] = buffer_data_1[3055:3048] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_381[18] = buffer_data_1[3063:3056] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_381[19] = buffer_data_1[3071:3064] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_381[20] = buffer_data_0[3039:3032] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_381[21] = buffer_data_0[3047:3040] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_381[22] = buffer_data_0[3055:3048] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_381[23] = buffer_data_0[3063:3056] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_381[24] = buffer_data_0[3071:3064] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_381 = kernel_img_mul_381[0] + kernel_img_mul_381[1] + kernel_img_mul_381[2] + 
                kernel_img_mul_381[3] + kernel_img_mul_381[4] + kernel_img_mul_381[5] + 
                kernel_img_mul_381[6] + kernel_img_mul_381[7] + kernel_img_mul_381[8] + 
                kernel_img_mul_381[9] + kernel_img_mul_381[10] + kernel_img_mul_381[11] + 
                kernel_img_mul_381[12] + kernel_img_mul_381[13] + kernel_img_mul_381[14] + 
                kernel_img_mul_381[15] + kernel_img_mul_381[16] + kernel_img_mul_381[17] + 
                kernel_img_mul_381[18] + kernel_img_mul_381[19] + kernel_img_mul_381[20] + 
                kernel_img_mul_381[21] + kernel_img_mul_381[22] + kernel_img_mul_381[23] + 
                kernel_img_mul_381[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3055:3048] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3055:3048] <= kernel_img_sum_381[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3055:3048] <= 'd0;
end

wire  [39:0]  kernel_img_mul_382[0:24];
assign kernel_img_mul_382[0] = buffer_data_4[3047:3040] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_382[1] = buffer_data_4[3055:3048] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_382[2] = buffer_data_4[3063:3056] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_382[3] = buffer_data_4[3071:3064] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_382[4] = buffer_data_4[3079:3072] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_382[5] = buffer_data_3[3047:3040] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_382[6] = buffer_data_3[3055:3048] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_382[7] = buffer_data_3[3063:3056] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_382[8] = buffer_data_3[3071:3064] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_382[9] = buffer_data_3[3079:3072] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_382[10] = buffer_data_2[3047:3040] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_382[11] = buffer_data_2[3055:3048] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_382[12] = buffer_data_2[3063:3056] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_382[13] = buffer_data_2[3071:3064] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_382[14] = buffer_data_2[3079:3072] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_382[15] = buffer_data_1[3047:3040] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_382[16] = buffer_data_1[3055:3048] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_382[17] = buffer_data_1[3063:3056] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_382[18] = buffer_data_1[3071:3064] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_382[19] = buffer_data_1[3079:3072] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_382[20] = buffer_data_0[3047:3040] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_382[21] = buffer_data_0[3055:3048] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_382[22] = buffer_data_0[3063:3056] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_382[23] = buffer_data_0[3071:3064] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_382[24] = buffer_data_0[3079:3072] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_382 = kernel_img_mul_382[0] + kernel_img_mul_382[1] + kernel_img_mul_382[2] + 
                kernel_img_mul_382[3] + kernel_img_mul_382[4] + kernel_img_mul_382[5] + 
                kernel_img_mul_382[6] + kernel_img_mul_382[7] + kernel_img_mul_382[8] + 
                kernel_img_mul_382[9] + kernel_img_mul_382[10] + kernel_img_mul_382[11] + 
                kernel_img_mul_382[12] + kernel_img_mul_382[13] + kernel_img_mul_382[14] + 
                kernel_img_mul_382[15] + kernel_img_mul_382[16] + kernel_img_mul_382[17] + 
                kernel_img_mul_382[18] + kernel_img_mul_382[19] + kernel_img_mul_382[20] + 
                kernel_img_mul_382[21] + kernel_img_mul_382[22] + kernel_img_mul_382[23] + 
                kernel_img_mul_382[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3063:3056] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3063:3056] <= kernel_img_sum_382[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3063:3056] <= 'd0;
end

wire  [39:0]  kernel_img_mul_383[0:24];
assign kernel_img_mul_383[0] = buffer_data_4[3055:3048] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_383[1] = buffer_data_4[3063:3056] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_383[2] = buffer_data_4[3071:3064] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_383[3] = buffer_data_4[3079:3072] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_383[4] = buffer_data_4[3087:3080] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_383[5] = buffer_data_3[3055:3048] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_383[6] = buffer_data_3[3063:3056] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_383[7] = buffer_data_3[3071:3064] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_383[8] = buffer_data_3[3079:3072] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_383[9] = buffer_data_3[3087:3080] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_383[10] = buffer_data_2[3055:3048] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_383[11] = buffer_data_2[3063:3056] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_383[12] = buffer_data_2[3071:3064] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_383[13] = buffer_data_2[3079:3072] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_383[14] = buffer_data_2[3087:3080] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_383[15] = buffer_data_1[3055:3048] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_383[16] = buffer_data_1[3063:3056] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_383[17] = buffer_data_1[3071:3064] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_383[18] = buffer_data_1[3079:3072] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_383[19] = buffer_data_1[3087:3080] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_383[20] = buffer_data_0[3055:3048] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_383[21] = buffer_data_0[3063:3056] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_383[22] = buffer_data_0[3071:3064] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_383[23] = buffer_data_0[3079:3072] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_383[24] = buffer_data_0[3087:3080] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_383 = kernel_img_mul_383[0] + kernel_img_mul_383[1] + kernel_img_mul_383[2] + 
                kernel_img_mul_383[3] + kernel_img_mul_383[4] + kernel_img_mul_383[5] + 
                kernel_img_mul_383[6] + kernel_img_mul_383[7] + kernel_img_mul_383[8] + 
                kernel_img_mul_383[9] + kernel_img_mul_383[10] + kernel_img_mul_383[11] + 
                kernel_img_mul_383[12] + kernel_img_mul_383[13] + kernel_img_mul_383[14] + 
                kernel_img_mul_383[15] + kernel_img_mul_383[16] + kernel_img_mul_383[17] + 
                kernel_img_mul_383[18] + kernel_img_mul_383[19] + kernel_img_mul_383[20] + 
                kernel_img_mul_383[21] + kernel_img_mul_383[22] + kernel_img_mul_383[23] + 
                kernel_img_mul_383[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3071:3064] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3071:3064] <= kernel_img_sum_383[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3071:3064] <= 'd0;
end

wire  [39:0]  kernel_img_mul_384[0:24];
assign kernel_img_mul_384[0] = buffer_data_4[3063:3056] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_384[1] = buffer_data_4[3071:3064] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_384[2] = buffer_data_4[3079:3072] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_384[3] = buffer_data_4[3087:3080] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_384[4] = buffer_data_4[3095:3088] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_384[5] = buffer_data_3[3063:3056] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_384[6] = buffer_data_3[3071:3064] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_384[7] = buffer_data_3[3079:3072] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_384[8] = buffer_data_3[3087:3080] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_384[9] = buffer_data_3[3095:3088] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_384[10] = buffer_data_2[3063:3056] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_384[11] = buffer_data_2[3071:3064] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_384[12] = buffer_data_2[3079:3072] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_384[13] = buffer_data_2[3087:3080] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_384[14] = buffer_data_2[3095:3088] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_384[15] = buffer_data_1[3063:3056] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_384[16] = buffer_data_1[3071:3064] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_384[17] = buffer_data_1[3079:3072] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_384[18] = buffer_data_1[3087:3080] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_384[19] = buffer_data_1[3095:3088] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_384[20] = buffer_data_0[3063:3056] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_384[21] = buffer_data_0[3071:3064] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_384[22] = buffer_data_0[3079:3072] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_384[23] = buffer_data_0[3087:3080] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_384[24] = buffer_data_0[3095:3088] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_384 = kernel_img_mul_384[0] + kernel_img_mul_384[1] + kernel_img_mul_384[2] + 
                kernel_img_mul_384[3] + kernel_img_mul_384[4] + kernel_img_mul_384[5] + 
                kernel_img_mul_384[6] + kernel_img_mul_384[7] + kernel_img_mul_384[8] + 
                kernel_img_mul_384[9] + kernel_img_mul_384[10] + kernel_img_mul_384[11] + 
                kernel_img_mul_384[12] + kernel_img_mul_384[13] + kernel_img_mul_384[14] + 
                kernel_img_mul_384[15] + kernel_img_mul_384[16] + kernel_img_mul_384[17] + 
                kernel_img_mul_384[18] + kernel_img_mul_384[19] + kernel_img_mul_384[20] + 
                kernel_img_mul_384[21] + kernel_img_mul_384[22] + kernel_img_mul_384[23] + 
                kernel_img_mul_384[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3079:3072] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3079:3072] <= kernel_img_sum_384[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3079:3072] <= 'd0;
end

wire  [39:0]  kernel_img_mul_385[0:24];
assign kernel_img_mul_385[0] = buffer_data_4[3071:3064] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_385[1] = buffer_data_4[3079:3072] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_385[2] = buffer_data_4[3087:3080] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_385[3] = buffer_data_4[3095:3088] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_385[4] = buffer_data_4[3103:3096] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_385[5] = buffer_data_3[3071:3064] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_385[6] = buffer_data_3[3079:3072] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_385[7] = buffer_data_3[3087:3080] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_385[8] = buffer_data_3[3095:3088] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_385[9] = buffer_data_3[3103:3096] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_385[10] = buffer_data_2[3071:3064] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_385[11] = buffer_data_2[3079:3072] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_385[12] = buffer_data_2[3087:3080] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_385[13] = buffer_data_2[3095:3088] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_385[14] = buffer_data_2[3103:3096] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_385[15] = buffer_data_1[3071:3064] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_385[16] = buffer_data_1[3079:3072] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_385[17] = buffer_data_1[3087:3080] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_385[18] = buffer_data_1[3095:3088] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_385[19] = buffer_data_1[3103:3096] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_385[20] = buffer_data_0[3071:3064] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_385[21] = buffer_data_0[3079:3072] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_385[22] = buffer_data_0[3087:3080] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_385[23] = buffer_data_0[3095:3088] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_385[24] = buffer_data_0[3103:3096] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_385 = kernel_img_mul_385[0] + kernel_img_mul_385[1] + kernel_img_mul_385[2] + 
                kernel_img_mul_385[3] + kernel_img_mul_385[4] + kernel_img_mul_385[5] + 
                kernel_img_mul_385[6] + kernel_img_mul_385[7] + kernel_img_mul_385[8] + 
                kernel_img_mul_385[9] + kernel_img_mul_385[10] + kernel_img_mul_385[11] + 
                kernel_img_mul_385[12] + kernel_img_mul_385[13] + kernel_img_mul_385[14] + 
                kernel_img_mul_385[15] + kernel_img_mul_385[16] + kernel_img_mul_385[17] + 
                kernel_img_mul_385[18] + kernel_img_mul_385[19] + kernel_img_mul_385[20] + 
                kernel_img_mul_385[21] + kernel_img_mul_385[22] + kernel_img_mul_385[23] + 
                kernel_img_mul_385[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3087:3080] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3087:3080] <= kernel_img_sum_385[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3087:3080] <= 'd0;
end

wire  [39:0]  kernel_img_mul_386[0:24];
assign kernel_img_mul_386[0] = buffer_data_4[3079:3072] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_386[1] = buffer_data_4[3087:3080] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_386[2] = buffer_data_4[3095:3088] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_386[3] = buffer_data_4[3103:3096] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_386[4] = buffer_data_4[3111:3104] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_386[5] = buffer_data_3[3079:3072] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_386[6] = buffer_data_3[3087:3080] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_386[7] = buffer_data_3[3095:3088] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_386[8] = buffer_data_3[3103:3096] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_386[9] = buffer_data_3[3111:3104] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_386[10] = buffer_data_2[3079:3072] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_386[11] = buffer_data_2[3087:3080] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_386[12] = buffer_data_2[3095:3088] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_386[13] = buffer_data_2[3103:3096] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_386[14] = buffer_data_2[3111:3104] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_386[15] = buffer_data_1[3079:3072] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_386[16] = buffer_data_1[3087:3080] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_386[17] = buffer_data_1[3095:3088] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_386[18] = buffer_data_1[3103:3096] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_386[19] = buffer_data_1[3111:3104] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_386[20] = buffer_data_0[3079:3072] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_386[21] = buffer_data_0[3087:3080] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_386[22] = buffer_data_0[3095:3088] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_386[23] = buffer_data_0[3103:3096] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_386[24] = buffer_data_0[3111:3104] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_386 = kernel_img_mul_386[0] + kernel_img_mul_386[1] + kernel_img_mul_386[2] + 
                kernel_img_mul_386[3] + kernel_img_mul_386[4] + kernel_img_mul_386[5] + 
                kernel_img_mul_386[6] + kernel_img_mul_386[7] + kernel_img_mul_386[8] + 
                kernel_img_mul_386[9] + kernel_img_mul_386[10] + kernel_img_mul_386[11] + 
                kernel_img_mul_386[12] + kernel_img_mul_386[13] + kernel_img_mul_386[14] + 
                kernel_img_mul_386[15] + kernel_img_mul_386[16] + kernel_img_mul_386[17] + 
                kernel_img_mul_386[18] + kernel_img_mul_386[19] + kernel_img_mul_386[20] + 
                kernel_img_mul_386[21] + kernel_img_mul_386[22] + kernel_img_mul_386[23] + 
                kernel_img_mul_386[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3095:3088] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3095:3088] <= kernel_img_sum_386[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3095:3088] <= 'd0;
end

wire  [39:0]  kernel_img_mul_387[0:24];
assign kernel_img_mul_387[0] = buffer_data_4[3087:3080] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_387[1] = buffer_data_4[3095:3088] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_387[2] = buffer_data_4[3103:3096] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_387[3] = buffer_data_4[3111:3104] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_387[4] = buffer_data_4[3119:3112] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_387[5] = buffer_data_3[3087:3080] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_387[6] = buffer_data_3[3095:3088] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_387[7] = buffer_data_3[3103:3096] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_387[8] = buffer_data_3[3111:3104] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_387[9] = buffer_data_3[3119:3112] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_387[10] = buffer_data_2[3087:3080] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_387[11] = buffer_data_2[3095:3088] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_387[12] = buffer_data_2[3103:3096] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_387[13] = buffer_data_2[3111:3104] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_387[14] = buffer_data_2[3119:3112] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_387[15] = buffer_data_1[3087:3080] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_387[16] = buffer_data_1[3095:3088] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_387[17] = buffer_data_1[3103:3096] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_387[18] = buffer_data_1[3111:3104] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_387[19] = buffer_data_1[3119:3112] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_387[20] = buffer_data_0[3087:3080] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_387[21] = buffer_data_0[3095:3088] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_387[22] = buffer_data_0[3103:3096] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_387[23] = buffer_data_0[3111:3104] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_387[24] = buffer_data_0[3119:3112] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_387 = kernel_img_mul_387[0] + kernel_img_mul_387[1] + kernel_img_mul_387[2] + 
                kernel_img_mul_387[3] + kernel_img_mul_387[4] + kernel_img_mul_387[5] + 
                kernel_img_mul_387[6] + kernel_img_mul_387[7] + kernel_img_mul_387[8] + 
                kernel_img_mul_387[9] + kernel_img_mul_387[10] + kernel_img_mul_387[11] + 
                kernel_img_mul_387[12] + kernel_img_mul_387[13] + kernel_img_mul_387[14] + 
                kernel_img_mul_387[15] + kernel_img_mul_387[16] + kernel_img_mul_387[17] + 
                kernel_img_mul_387[18] + kernel_img_mul_387[19] + kernel_img_mul_387[20] + 
                kernel_img_mul_387[21] + kernel_img_mul_387[22] + kernel_img_mul_387[23] + 
                kernel_img_mul_387[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3103:3096] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3103:3096] <= kernel_img_sum_387[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3103:3096] <= 'd0;
end

wire  [39:0]  kernel_img_mul_388[0:24];
assign kernel_img_mul_388[0] = buffer_data_4[3095:3088] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_388[1] = buffer_data_4[3103:3096] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_388[2] = buffer_data_4[3111:3104] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_388[3] = buffer_data_4[3119:3112] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_388[4] = buffer_data_4[3127:3120] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_388[5] = buffer_data_3[3095:3088] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_388[6] = buffer_data_3[3103:3096] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_388[7] = buffer_data_3[3111:3104] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_388[8] = buffer_data_3[3119:3112] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_388[9] = buffer_data_3[3127:3120] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_388[10] = buffer_data_2[3095:3088] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_388[11] = buffer_data_2[3103:3096] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_388[12] = buffer_data_2[3111:3104] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_388[13] = buffer_data_2[3119:3112] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_388[14] = buffer_data_2[3127:3120] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_388[15] = buffer_data_1[3095:3088] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_388[16] = buffer_data_1[3103:3096] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_388[17] = buffer_data_1[3111:3104] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_388[18] = buffer_data_1[3119:3112] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_388[19] = buffer_data_1[3127:3120] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_388[20] = buffer_data_0[3095:3088] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_388[21] = buffer_data_0[3103:3096] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_388[22] = buffer_data_0[3111:3104] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_388[23] = buffer_data_0[3119:3112] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_388[24] = buffer_data_0[3127:3120] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_388 = kernel_img_mul_388[0] + kernel_img_mul_388[1] + kernel_img_mul_388[2] + 
                kernel_img_mul_388[3] + kernel_img_mul_388[4] + kernel_img_mul_388[5] + 
                kernel_img_mul_388[6] + kernel_img_mul_388[7] + kernel_img_mul_388[8] + 
                kernel_img_mul_388[9] + kernel_img_mul_388[10] + kernel_img_mul_388[11] + 
                kernel_img_mul_388[12] + kernel_img_mul_388[13] + kernel_img_mul_388[14] + 
                kernel_img_mul_388[15] + kernel_img_mul_388[16] + kernel_img_mul_388[17] + 
                kernel_img_mul_388[18] + kernel_img_mul_388[19] + kernel_img_mul_388[20] + 
                kernel_img_mul_388[21] + kernel_img_mul_388[22] + kernel_img_mul_388[23] + 
                kernel_img_mul_388[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3111:3104] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3111:3104] <= kernel_img_sum_388[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3111:3104] <= 'd0;
end

wire  [39:0]  kernel_img_mul_389[0:24];
assign kernel_img_mul_389[0] = buffer_data_4[3103:3096] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_389[1] = buffer_data_4[3111:3104] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_389[2] = buffer_data_4[3119:3112] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_389[3] = buffer_data_4[3127:3120] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_389[4] = buffer_data_4[3135:3128] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_389[5] = buffer_data_3[3103:3096] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_389[6] = buffer_data_3[3111:3104] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_389[7] = buffer_data_3[3119:3112] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_389[8] = buffer_data_3[3127:3120] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_389[9] = buffer_data_3[3135:3128] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_389[10] = buffer_data_2[3103:3096] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_389[11] = buffer_data_2[3111:3104] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_389[12] = buffer_data_2[3119:3112] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_389[13] = buffer_data_2[3127:3120] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_389[14] = buffer_data_2[3135:3128] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_389[15] = buffer_data_1[3103:3096] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_389[16] = buffer_data_1[3111:3104] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_389[17] = buffer_data_1[3119:3112] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_389[18] = buffer_data_1[3127:3120] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_389[19] = buffer_data_1[3135:3128] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_389[20] = buffer_data_0[3103:3096] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_389[21] = buffer_data_0[3111:3104] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_389[22] = buffer_data_0[3119:3112] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_389[23] = buffer_data_0[3127:3120] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_389[24] = buffer_data_0[3135:3128] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_389 = kernel_img_mul_389[0] + kernel_img_mul_389[1] + kernel_img_mul_389[2] + 
                kernel_img_mul_389[3] + kernel_img_mul_389[4] + kernel_img_mul_389[5] + 
                kernel_img_mul_389[6] + kernel_img_mul_389[7] + kernel_img_mul_389[8] + 
                kernel_img_mul_389[9] + kernel_img_mul_389[10] + kernel_img_mul_389[11] + 
                kernel_img_mul_389[12] + kernel_img_mul_389[13] + kernel_img_mul_389[14] + 
                kernel_img_mul_389[15] + kernel_img_mul_389[16] + kernel_img_mul_389[17] + 
                kernel_img_mul_389[18] + kernel_img_mul_389[19] + kernel_img_mul_389[20] + 
                kernel_img_mul_389[21] + kernel_img_mul_389[22] + kernel_img_mul_389[23] + 
                kernel_img_mul_389[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3119:3112] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3119:3112] <= kernel_img_sum_389[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3119:3112] <= 'd0;
end

wire  [39:0]  kernel_img_mul_390[0:24];
assign kernel_img_mul_390[0] = buffer_data_4[3111:3104] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_390[1] = buffer_data_4[3119:3112] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_390[2] = buffer_data_4[3127:3120] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_390[3] = buffer_data_4[3135:3128] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_390[4] = buffer_data_4[3143:3136] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_390[5] = buffer_data_3[3111:3104] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_390[6] = buffer_data_3[3119:3112] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_390[7] = buffer_data_3[3127:3120] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_390[8] = buffer_data_3[3135:3128] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_390[9] = buffer_data_3[3143:3136] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_390[10] = buffer_data_2[3111:3104] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_390[11] = buffer_data_2[3119:3112] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_390[12] = buffer_data_2[3127:3120] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_390[13] = buffer_data_2[3135:3128] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_390[14] = buffer_data_2[3143:3136] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_390[15] = buffer_data_1[3111:3104] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_390[16] = buffer_data_1[3119:3112] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_390[17] = buffer_data_1[3127:3120] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_390[18] = buffer_data_1[3135:3128] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_390[19] = buffer_data_1[3143:3136] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_390[20] = buffer_data_0[3111:3104] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_390[21] = buffer_data_0[3119:3112] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_390[22] = buffer_data_0[3127:3120] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_390[23] = buffer_data_0[3135:3128] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_390[24] = buffer_data_0[3143:3136] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_390 = kernel_img_mul_390[0] + kernel_img_mul_390[1] + kernel_img_mul_390[2] + 
                kernel_img_mul_390[3] + kernel_img_mul_390[4] + kernel_img_mul_390[5] + 
                kernel_img_mul_390[6] + kernel_img_mul_390[7] + kernel_img_mul_390[8] + 
                kernel_img_mul_390[9] + kernel_img_mul_390[10] + kernel_img_mul_390[11] + 
                kernel_img_mul_390[12] + kernel_img_mul_390[13] + kernel_img_mul_390[14] + 
                kernel_img_mul_390[15] + kernel_img_mul_390[16] + kernel_img_mul_390[17] + 
                kernel_img_mul_390[18] + kernel_img_mul_390[19] + kernel_img_mul_390[20] + 
                kernel_img_mul_390[21] + kernel_img_mul_390[22] + kernel_img_mul_390[23] + 
                kernel_img_mul_390[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3127:3120] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3127:3120] <= kernel_img_sum_390[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3127:3120] <= 'd0;
end

wire  [39:0]  kernel_img_mul_391[0:24];
assign kernel_img_mul_391[0] = buffer_data_4[3119:3112] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_391[1] = buffer_data_4[3127:3120] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_391[2] = buffer_data_4[3135:3128] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_391[3] = buffer_data_4[3143:3136] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_391[4] = buffer_data_4[3151:3144] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_391[5] = buffer_data_3[3119:3112] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_391[6] = buffer_data_3[3127:3120] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_391[7] = buffer_data_3[3135:3128] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_391[8] = buffer_data_3[3143:3136] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_391[9] = buffer_data_3[3151:3144] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_391[10] = buffer_data_2[3119:3112] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_391[11] = buffer_data_2[3127:3120] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_391[12] = buffer_data_2[3135:3128] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_391[13] = buffer_data_2[3143:3136] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_391[14] = buffer_data_2[3151:3144] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_391[15] = buffer_data_1[3119:3112] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_391[16] = buffer_data_1[3127:3120] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_391[17] = buffer_data_1[3135:3128] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_391[18] = buffer_data_1[3143:3136] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_391[19] = buffer_data_1[3151:3144] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_391[20] = buffer_data_0[3119:3112] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_391[21] = buffer_data_0[3127:3120] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_391[22] = buffer_data_0[3135:3128] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_391[23] = buffer_data_0[3143:3136] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_391[24] = buffer_data_0[3151:3144] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_391 = kernel_img_mul_391[0] + kernel_img_mul_391[1] + kernel_img_mul_391[2] + 
                kernel_img_mul_391[3] + kernel_img_mul_391[4] + kernel_img_mul_391[5] + 
                kernel_img_mul_391[6] + kernel_img_mul_391[7] + kernel_img_mul_391[8] + 
                kernel_img_mul_391[9] + kernel_img_mul_391[10] + kernel_img_mul_391[11] + 
                kernel_img_mul_391[12] + kernel_img_mul_391[13] + kernel_img_mul_391[14] + 
                kernel_img_mul_391[15] + kernel_img_mul_391[16] + kernel_img_mul_391[17] + 
                kernel_img_mul_391[18] + kernel_img_mul_391[19] + kernel_img_mul_391[20] + 
                kernel_img_mul_391[21] + kernel_img_mul_391[22] + kernel_img_mul_391[23] + 
                kernel_img_mul_391[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3135:3128] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3135:3128] <= kernel_img_sum_391[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3135:3128] <= 'd0;
end

wire  [39:0]  kernel_img_mul_392[0:24];
assign kernel_img_mul_392[0] = buffer_data_4[3127:3120] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_392[1] = buffer_data_4[3135:3128] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_392[2] = buffer_data_4[3143:3136] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_392[3] = buffer_data_4[3151:3144] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_392[4] = buffer_data_4[3159:3152] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_392[5] = buffer_data_3[3127:3120] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_392[6] = buffer_data_3[3135:3128] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_392[7] = buffer_data_3[3143:3136] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_392[8] = buffer_data_3[3151:3144] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_392[9] = buffer_data_3[3159:3152] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_392[10] = buffer_data_2[3127:3120] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_392[11] = buffer_data_2[3135:3128] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_392[12] = buffer_data_2[3143:3136] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_392[13] = buffer_data_2[3151:3144] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_392[14] = buffer_data_2[3159:3152] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_392[15] = buffer_data_1[3127:3120] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_392[16] = buffer_data_1[3135:3128] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_392[17] = buffer_data_1[3143:3136] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_392[18] = buffer_data_1[3151:3144] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_392[19] = buffer_data_1[3159:3152] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_392[20] = buffer_data_0[3127:3120] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_392[21] = buffer_data_0[3135:3128] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_392[22] = buffer_data_0[3143:3136] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_392[23] = buffer_data_0[3151:3144] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_392[24] = buffer_data_0[3159:3152] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_392 = kernel_img_mul_392[0] + kernel_img_mul_392[1] + kernel_img_mul_392[2] + 
                kernel_img_mul_392[3] + kernel_img_mul_392[4] + kernel_img_mul_392[5] + 
                kernel_img_mul_392[6] + kernel_img_mul_392[7] + kernel_img_mul_392[8] + 
                kernel_img_mul_392[9] + kernel_img_mul_392[10] + kernel_img_mul_392[11] + 
                kernel_img_mul_392[12] + kernel_img_mul_392[13] + kernel_img_mul_392[14] + 
                kernel_img_mul_392[15] + kernel_img_mul_392[16] + kernel_img_mul_392[17] + 
                kernel_img_mul_392[18] + kernel_img_mul_392[19] + kernel_img_mul_392[20] + 
                kernel_img_mul_392[21] + kernel_img_mul_392[22] + kernel_img_mul_392[23] + 
                kernel_img_mul_392[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3143:3136] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3143:3136] <= kernel_img_sum_392[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3143:3136] <= 'd0;
end

wire  [39:0]  kernel_img_mul_393[0:24];
assign kernel_img_mul_393[0] = buffer_data_4[3135:3128] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_393[1] = buffer_data_4[3143:3136] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_393[2] = buffer_data_4[3151:3144] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_393[3] = buffer_data_4[3159:3152] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_393[4] = buffer_data_4[3167:3160] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_393[5] = buffer_data_3[3135:3128] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_393[6] = buffer_data_3[3143:3136] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_393[7] = buffer_data_3[3151:3144] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_393[8] = buffer_data_3[3159:3152] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_393[9] = buffer_data_3[3167:3160] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_393[10] = buffer_data_2[3135:3128] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_393[11] = buffer_data_2[3143:3136] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_393[12] = buffer_data_2[3151:3144] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_393[13] = buffer_data_2[3159:3152] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_393[14] = buffer_data_2[3167:3160] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_393[15] = buffer_data_1[3135:3128] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_393[16] = buffer_data_1[3143:3136] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_393[17] = buffer_data_1[3151:3144] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_393[18] = buffer_data_1[3159:3152] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_393[19] = buffer_data_1[3167:3160] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_393[20] = buffer_data_0[3135:3128] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_393[21] = buffer_data_0[3143:3136] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_393[22] = buffer_data_0[3151:3144] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_393[23] = buffer_data_0[3159:3152] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_393[24] = buffer_data_0[3167:3160] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_393 = kernel_img_mul_393[0] + kernel_img_mul_393[1] + kernel_img_mul_393[2] + 
                kernel_img_mul_393[3] + kernel_img_mul_393[4] + kernel_img_mul_393[5] + 
                kernel_img_mul_393[6] + kernel_img_mul_393[7] + kernel_img_mul_393[8] + 
                kernel_img_mul_393[9] + kernel_img_mul_393[10] + kernel_img_mul_393[11] + 
                kernel_img_mul_393[12] + kernel_img_mul_393[13] + kernel_img_mul_393[14] + 
                kernel_img_mul_393[15] + kernel_img_mul_393[16] + kernel_img_mul_393[17] + 
                kernel_img_mul_393[18] + kernel_img_mul_393[19] + kernel_img_mul_393[20] + 
                kernel_img_mul_393[21] + kernel_img_mul_393[22] + kernel_img_mul_393[23] + 
                kernel_img_mul_393[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3151:3144] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3151:3144] <= kernel_img_sum_393[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3151:3144] <= 'd0;
end

wire  [39:0]  kernel_img_mul_394[0:24];
assign kernel_img_mul_394[0] = buffer_data_4[3143:3136] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_394[1] = buffer_data_4[3151:3144] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_394[2] = buffer_data_4[3159:3152] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_394[3] = buffer_data_4[3167:3160] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_394[4] = buffer_data_4[3175:3168] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_394[5] = buffer_data_3[3143:3136] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_394[6] = buffer_data_3[3151:3144] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_394[7] = buffer_data_3[3159:3152] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_394[8] = buffer_data_3[3167:3160] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_394[9] = buffer_data_3[3175:3168] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_394[10] = buffer_data_2[3143:3136] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_394[11] = buffer_data_2[3151:3144] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_394[12] = buffer_data_2[3159:3152] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_394[13] = buffer_data_2[3167:3160] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_394[14] = buffer_data_2[3175:3168] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_394[15] = buffer_data_1[3143:3136] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_394[16] = buffer_data_1[3151:3144] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_394[17] = buffer_data_1[3159:3152] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_394[18] = buffer_data_1[3167:3160] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_394[19] = buffer_data_1[3175:3168] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_394[20] = buffer_data_0[3143:3136] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_394[21] = buffer_data_0[3151:3144] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_394[22] = buffer_data_0[3159:3152] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_394[23] = buffer_data_0[3167:3160] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_394[24] = buffer_data_0[3175:3168] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_394 = kernel_img_mul_394[0] + kernel_img_mul_394[1] + kernel_img_mul_394[2] + 
                kernel_img_mul_394[3] + kernel_img_mul_394[4] + kernel_img_mul_394[5] + 
                kernel_img_mul_394[6] + kernel_img_mul_394[7] + kernel_img_mul_394[8] + 
                kernel_img_mul_394[9] + kernel_img_mul_394[10] + kernel_img_mul_394[11] + 
                kernel_img_mul_394[12] + kernel_img_mul_394[13] + kernel_img_mul_394[14] + 
                kernel_img_mul_394[15] + kernel_img_mul_394[16] + kernel_img_mul_394[17] + 
                kernel_img_mul_394[18] + kernel_img_mul_394[19] + kernel_img_mul_394[20] + 
                kernel_img_mul_394[21] + kernel_img_mul_394[22] + kernel_img_mul_394[23] + 
                kernel_img_mul_394[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3159:3152] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3159:3152] <= kernel_img_sum_394[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3159:3152] <= 'd0;
end

wire  [39:0]  kernel_img_mul_395[0:24];
assign kernel_img_mul_395[0] = buffer_data_4[3151:3144] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_395[1] = buffer_data_4[3159:3152] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_395[2] = buffer_data_4[3167:3160] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_395[3] = buffer_data_4[3175:3168] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_395[4] = buffer_data_4[3183:3176] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_395[5] = buffer_data_3[3151:3144] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_395[6] = buffer_data_3[3159:3152] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_395[7] = buffer_data_3[3167:3160] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_395[8] = buffer_data_3[3175:3168] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_395[9] = buffer_data_3[3183:3176] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_395[10] = buffer_data_2[3151:3144] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_395[11] = buffer_data_2[3159:3152] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_395[12] = buffer_data_2[3167:3160] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_395[13] = buffer_data_2[3175:3168] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_395[14] = buffer_data_2[3183:3176] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_395[15] = buffer_data_1[3151:3144] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_395[16] = buffer_data_1[3159:3152] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_395[17] = buffer_data_1[3167:3160] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_395[18] = buffer_data_1[3175:3168] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_395[19] = buffer_data_1[3183:3176] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_395[20] = buffer_data_0[3151:3144] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_395[21] = buffer_data_0[3159:3152] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_395[22] = buffer_data_0[3167:3160] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_395[23] = buffer_data_0[3175:3168] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_395[24] = buffer_data_0[3183:3176] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_395 = kernel_img_mul_395[0] + kernel_img_mul_395[1] + kernel_img_mul_395[2] + 
                kernel_img_mul_395[3] + kernel_img_mul_395[4] + kernel_img_mul_395[5] + 
                kernel_img_mul_395[6] + kernel_img_mul_395[7] + kernel_img_mul_395[8] + 
                kernel_img_mul_395[9] + kernel_img_mul_395[10] + kernel_img_mul_395[11] + 
                kernel_img_mul_395[12] + kernel_img_mul_395[13] + kernel_img_mul_395[14] + 
                kernel_img_mul_395[15] + kernel_img_mul_395[16] + kernel_img_mul_395[17] + 
                kernel_img_mul_395[18] + kernel_img_mul_395[19] + kernel_img_mul_395[20] + 
                kernel_img_mul_395[21] + kernel_img_mul_395[22] + kernel_img_mul_395[23] + 
                kernel_img_mul_395[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3167:3160] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3167:3160] <= kernel_img_sum_395[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3167:3160] <= 'd0;
end

wire  [39:0]  kernel_img_mul_396[0:24];
assign kernel_img_mul_396[0] = buffer_data_4[3159:3152] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_396[1] = buffer_data_4[3167:3160] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_396[2] = buffer_data_4[3175:3168] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_396[3] = buffer_data_4[3183:3176] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_396[4] = buffer_data_4[3191:3184] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_396[5] = buffer_data_3[3159:3152] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_396[6] = buffer_data_3[3167:3160] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_396[7] = buffer_data_3[3175:3168] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_396[8] = buffer_data_3[3183:3176] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_396[9] = buffer_data_3[3191:3184] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_396[10] = buffer_data_2[3159:3152] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_396[11] = buffer_data_2[3167:3160] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_396[12] = buffer_data_2[3175:3168] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_396[13] = buffer_data_2[3183:3176] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_396[14] = buffer_data_2[3191:3184] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_396[15] = buffer_data_1[3159:3152] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_396[16] = buffer_data_1[3167:3160] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_396[17] = buffer_data_1[3175:3168] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_396[18] = buffer_data_1[3183:3176] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_396[19] = buffer_data_1[3191:3184] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_396[20] = buffer_data_0[3159:3152] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_396[21] = buffer_data_0[3167:3160] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_396[22] = buffer_data_0[3175:3168] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_396[23] = buffer_data_0[3183:3176] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_396[24] = buffer_data_0[3191:3184] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_396 = kernel_img_mul_396[0] + kernel_img_mul_396[1] + kernel_img_mul_396[2] + 
                kernel_img_mul_396[3] + kernel_img_mul_396[4] + kernel_img_mul_396[5] + 
                kernel_img_mul_396[6] + kernel_img_mul_396[7] + kernel_img_mul_396[8] + 
                kernel_img_mul_396[9] + kernel_img_mul_396[10] + kernel_img_mul_396[11] + 
                kernel_img_mul_396[12] + kernel_img_mul_396[13] + kernel_img_mul_396[14] + 
                kernel_img_mul_396[15] + kernel_img_mul_396[16] + kernel_img_mul_396[17] + 
                kernel_img_mul_396[18] + kernel_img_mul_396[19] + kernel_img_mul_396[20] + 
                kernel_img_mul_396[21] + kernel_img_mul_396[22] + kernel_img_mul_396[23] + 
                kernel_img_mul_396[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3175:3168] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3175:3168] <= kernel_img_sum_396[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3175:3168] <= 'd0;
end

wire  [39:0]  kernel_img_mul_397[0:24];
assign kernel_img_mul_397[0] = buffer_data_4[3167:3160] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_397[1] = buffer_data_4[3175:3168] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_397[2] = buffer_data_4[3183:3176] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_397[3] = buffer_data_4[3191:3184] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_397[4] = buffer_data_4[3199:3192] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_397[5] = buffer_data_3[3167:3160] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_397[6] = buffer_data_3[3175:3168] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_397[7] = buffer_data_3[3183:3176] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_397[8] = buffer_data_3[3191:3184] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_397[9] = buffer_data_3[3199:3192] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_397[10] = buffer_data_2[3167:3160] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_397[11] = buffer_data_2[3175:3168] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_397[12] = buffer_data_2[3183:3176] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_397[13] = buffer_data_2[3191:3184] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_397[14] = buffer_data_2[3199:3192] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_397[15] = buffer_data_1[3167:3160] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_397[16] = buffer_data_1[3175:3168] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_397[17] = buffer_data_1[3183:3176] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_397[18] = buffer_data_1[3191:3184] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_397[19] = buffer_data_1[3199:3192] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_397[20] = buffer_data_0[3167:3160] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_397[21] = buffer_data_0[3175:3168] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_397[22] = buffer_data_0[3183:3176] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_397[23] = buffer_data_0[3191:3184] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_397[24] = buffer_data_0[3199:3192] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_397 = kernel_img_mul_397[0] + kernel_img_mul_397[1] + kernel_img_mul_397[2] + 
                kernel_img_mul_397[3] + kernel_img_mul_397[4] + kernel_img_mul_397[5] + 
                kernel_img_mul_397[6] + kernel_img_mul_397[7] + kernel_img_mul_397[8] + 
                kernel_img_mul_397[9] + kernel_img_mul_397[10] + kernel_img_mul_397[11] + 
                kernel_img_mul_397[12] + kernel_img_mul_397[13] + kernel_img_mul_397[14] + 
                kernel_img_mul_397[15] + kernel_img_mul_397[16] + kernel_img_mul_397[17] + 
                kernel_img_mul_397[18] + kernel_img_mul_397[19] + kernel_img_mul_397[20] + 
                kernel_img_mul_397[21] + kernel_img_mul_397[22] + kernel_img_mul_397[23] + 
                kernel_img_mul_397[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3183:3176] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3183:3176] <= kernel_img_sum_397[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3183:3176] <= 'd0;
end

wire  [39:0]  kernel_img_mul_398[0:24];
assign kernel_img_mul_398[0] = buffer_data_4[3175:3168] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_398[1] = buffer_data_4[3183:3176] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_398[2] = buffer_data_4[3191:3184] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_398[3] = buffer_data_4[3199:3192] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_398[4] = buffer_data_4[3207:3200] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_398[5] = buffer_data_3[3175:3168] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_398[6] = buffer_data_3[3183:3176] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_398[7] = buffer_data_3[3191:3184] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_398[8] = buffer_data_3[3199:3192] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_398[9] = buffer_data_3[3207:3200] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_398[10] = buffer_data_2[3175:3168] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_398[11] = buffer_data_2[3183:3176] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_398[12] = buffer_data_2[3191:3184] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_398[13] = buffer_data_2[3199:3192] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_398[14] = buffer_data_2[3207:3200] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_398[15] = buffer_data_1[3175:3168] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_398[16] = buffer_data_1[3183:3176] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_398[17] = buffer_data_1[3191:3184] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_398[18] = buffer_data_1[3199:3192] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_398[19] = buffer_data_1[3207:3200] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_398[20] = buffer_data_0[3175:3168] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_398[21] = buffer_data_0[3183:3176] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_398[22] = buffer_data_0[3191:3184] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_398[23] = buffer_data_0[3199:3192] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_398[24] = buffer_data_0[3207:3200] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_398 = kernel_img_mul_398[0] + kernel_img_mul_398[1] + kernel_img_mul_398[2] + 
                kernel_img_mul_398[3] + kernel_img_mul_398[4] + kernel_img_mul_398[5] + 
                kernel_img_mul_398[6] + kernel_img_mul_398[7] + kernel_img_mul_398[8] + 
                kernel_img_mul_398[9] + kernel_img_mul_398[10] + kernel_img_mul_398[11] + 
                kernel_img_mul_398[12] + kernel_img_mul_398[13] + kernel_img_mul_398[14] + 
                kernel_img_mul_398[15] + kernel_img_mul_398[16] + kernel_img_mul_398[17] + 
                kernel_img_mul_398[18] + kernel_img_mul_398[19] + kernel_img_mul_398[20] + 
                kernel_img_mul_398[21] + kernel_img_mul_398[22] + kernel_img_mul_398[23] + 
                kernel_img_mul_398[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3191:3184] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3191:3184] <= kernel_img_sum_398[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3191:3184] <= 'd0;
end

wire  [39:0]  kernel_img_mul_399[0:24];
assign kernel_img_mul_399[0] = buffer_data_4[3183:3176] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_399[1] = buffer_data_4[3191:3184] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_399[2] = buffer_data_4[3199:3192] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_399[3] = buffer_data_4[3207:3200] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_399[4] = buffer_data_4[3215:3208] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_399[5] = buffer_data_3[3183:3176] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_399[6] = buffer_data_3[3191:3184] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_399[7] = buffer_data_3[3199:3192] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_399[8] = buffer_data_3[3207:3200] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_399[9] = buffer_data_3[3215:3208] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_399[10] = buffer_data_2[3183:3176] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_399[11] = buffer_data_2[3191:3184] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_399[12] = buffer_data_2[3199:3192] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_399[13] = buffer_data_2[3207:3200] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_399[14] = buffer_data_2[3215:3208] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_399[15] = buffer_data_1[3183:3176] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_399[16] = buffer_data_1[3191:3184] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_399[17] = buffer_data_1[3199:3192] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_399[18] = buffer_data_1[3207:3200] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_399[19] = buffer_data_1[3215:3208] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_399[20] = buffer_data_0[3183:3176] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_399[21] = buffer_data_0[3191:3184] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_399[22] = buffer_data_0[3199:3192] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_399[23] = buffer_data_0[3207:3200] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_399[24] = buffer_data_0[3215:3208] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_399 = kernel_img_mul_399[0] + kernel_img_mul_399[1] + kernel_img_mul_399[2] + 
                kernel_img_mul_399[3] + kernel_img_mul_399[4] + kernel_img_mul_399[5] + 
                kernel_img_mul_399[6] + kernel_img_mul_399[7] + kernel_img_mul_399[8] + 
                kernel_img_mul_399[9] + kernel_img_mul_399[10] + kernel_img_mul_399[11] + 
                kernel_img_mul_399[12] + kernel_img_mul_399[13] + kernel_img_mul_399[14] + 
                kernel_img_mul_399[15] + kernel_img_mul_399[16] + kernel_img_mul_399[17] + 
                kernel_img_mul_399[18] + kernel_img_mul_399[19] + kernel_img_mul_399[20] + 
                kernel_img_mul_399[21] + kernel_img_mul_399[22] + kernel_img_mul_399[23] + 
                kernel_img_mul_399[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3199:3192] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3199:3192] <= kernel_img_sum_399[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3199:3192] <= 'd0;
end

wire  [39:0]  kernel_img_mul_400[0:24];
assign kernel_img_mul_400[0] = buffer_data_4[3191:3184] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_400[1] = buffer_data_4[3199:3192] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_400[2] = buffer_data_4[3207:3200] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_400[3] = buffer_data_4[3215:3208] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_400[4] = buffer_data_4[3223:3216] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_400[5] = buffer_data_3[3191:3184] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_400[6] = buffer_data_3[3199:3192] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_400[7] = buffer_data_3[3207:3200] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_400[8] = buffer_data_3[3215:3208] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_400[9] = buffer_data_3[3223:3216] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_400[10] = buffer_data_2[3191:3184] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_400[11] = buffer_data_2[3199:3192] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_400[12] = buffer_data_2[3207:3200] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_400[13] = buffer_data_2[3215:3208] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_400[14] = buffer_data_2[3223:3216] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_400[15] = buffer_data_1[3191:3184] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_400[16] = buffer_data_1[3199:3192] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_400[17] = buffer_data_1[3207:3200] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_400[18] = buffer_data_1[3215:3208] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_400[19] = buffer_data_1[3223:3216] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_400[20] = buffer_data_0[3191:3184] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_400[21] = buffer_data_0[3199:3192] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_400[22] = buffer_data_0[3207:3200] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_400[23] = buffer_data_0[3215:3208] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_400[24] = buffer_data_0[3223:3216] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_400 = kernel_img_mul_400[0] + kernel_img_mul_400[1] + kernel_img_mul_400[2] + 
                kernel_img_mul_400[3] + kernel_img_mul_400[4] + kernel_img_mul_400[5] + 
                kernel_img_mul_400[6] + kernel_img_mul_400[7] + kernel_img_mul_400[8] + 
                kernel_img_mul_400[9] + kernel_img_mul_400[10] + kernel_img_mul_400[11] + 
                kernel_img_mul_400[12] + kernel_img_mul_400[13] + kernel_img_mul_400[14] + 
                kernel_img_mul_400[15] + kernel_img_mul_400[16] + kernel_img_mul_400[17] + 
                kernel_img_mul_400[18] + kernel_img_mul_400[19] + kernel_img_mul_400[20] + 
                kernel_img_mul_400[21] + kernel_img_mul_400[22] + kernel_img_mul_400[23] + 
                kernel_img_mul_400[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3207:3200] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3207:3200] <= kernel_img_sum_400[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3207:3200] <= 'd0;
end

wire  [39:0]  kernel_img_mul_401[0:24];
assign kernel_img_mul_401[0] = buffer_data_4[3199:3192] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_401[1] = buffer_data_4[3207:3200] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_401[2] = buffer_data_4[3215:3208] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_401[3] = buffer_data_4[3223:3216] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_401[4] = buffer_data_4[3231:3224] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_401[5] = buffer_data_3[3199:3192] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_401[6] = buffer_data_3[3207:3200] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_401[7] = buffer_data_3[3215:3208] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_401[8] = buffer_data_3[3223:3216] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_401[9] = buffer_data_3[3231:3224] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_401[10] = buffer_data_2[3199:3192] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_401[11] = buffer_data_2[3207:3200] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_401[12] = buffer_data_2[3215:3208] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_401[13] = buffer_data_2[3223:3216] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_401[14] = buffer_data_2[3231:3224] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_401[15] = buffer_data_1[3199:3192] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_401[16] = buffer_data_1[3207:3200] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_401[17] = buffer_data_1[3215:3208] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_401[18] = buffer_data_1[3223:3216] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_401[19] = buffer_data_1[3231:3224] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_401[20] = buffer_data_0[3199:3192] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_401[21] = buffer_data_0[3207:3200] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_401[22] = buffer_data_0[3215:3208] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_401[23] = buffer_data_0[3223:3216] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_401[24] = buffer_data_0[3231:3224] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_401 = kernel_img_mul_401[0] + kernel_img_mul_401[1] + kernel_img_mul_401[2] + 
                kernel_img_mul_401[3] + kernel_img_mul_401[4] + kernel_img_mul_401[5] + 
                kernel_img_mul_401[6] + kernel_img_mul_401[7] + kernel_img_mul_401[8] + 
                kernel_img_mul_401[9] + kernel_img_mul_401[10] + kernel_img_mul_401[11] + 
                kernel_img_mul_401[12] + kernel_img_mul_401[13] + kernel_img_mul_401[14] + 
                kernel_img_mul_401[15] + kernel_img_mul_401[16] + kernel_img_mul_401[17] + 
                kernel_img_mul_401[18] + kernel_img_mul_401[19] + kernel_img_mul_401[20] + 
                kernel_img_mul_401[21] + kernel_img_mul_401[22] + kernel_img_mul_401[23] + 
                kernel_img_mul_401[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3215:3208] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3215:3208] <= kernel_img_sum_401[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3215:3208] <= 'd0;
end

wire  [39:0]  kernel_img_mul_402[0:24];
assign kernel_img_mul_402[0] = buffer_data_4[3207:3200] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_402[1] = buffer_data_4[3215:3208] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_402[2] = buffer_data_4[3223:3216] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_402[3] = buffer_data_4[3231:3224] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_402[4] = buffer_data_4[3239:3232] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_402[5] = buffer_data_3[3207:3200] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_402[6] = buffer_data_3[3215:3208] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_402[7] = buffer_data_3[3223:3216] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_402[8] = buffer_data_3[3231:3224] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_402[9] = buffer_data_3[3239:3232] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_402[10] = buffer_data_2[3207:3200] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_402[11] = buffer_data_2[3215:3208] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_402[12] = buffer_data_2[3223:3216] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_402[13] = buffer_data_2[3231:3224] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_402[14] = buffer_data_2[3239:3232] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_402[15] = buffer_data_1[3207:3200] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_402[16] = buffer_data_1[3215:3208] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_402[17] = buffer_data_1[3223:3216] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_402[18] = buffer_data_1[3231:3224] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_402[19] = buffer_data_1[3239:3232] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_402[20] = buffer_data_0[3207:3200] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_402[21] = buffer_data_0[3215:3208] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_402[22] = buffer_data_0[3223:3216] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_402[23] = buffer_data_0[3231:3224] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_402[24] = buffer_data_0[3239:3232] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_402 = kernel_img_mul_402[0] + kernel_img_mul_402[1] + kernel_img_mul_402[2] + 
                kernel_img_mul_402[3] + kernel_img_mul_402[4] + kernel_img_mul_402[5] + 
                kernel_img_mul_402[6] + kernel_img_mul_402[7] + kernel_img_mul_402[8] + 
                kernel_img_mul_402[9] + kernel_img_mul_402[10] + kernel_img_mul_402[11] + 
                kernel_img_mul_402[12] + kernel_img_mul_402[13] + kernel_img_mul_402[14] + 
                kernel_img_mul_402[15] + kernel_img_mul_402[16] + kernel_img_mul_402[17] + 
                kernel_img_mul_402[18] + kernel_img_mul_402[19] + kernel_img_mul_402[20] + 
                kernel_img_mul_402[21] + kernel_img_mul_402[22] + kernel_img_mul_402[23] + 
                kernel_img_mul_402[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3223:3216] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3223:3216] <= kernel_img_sum_402[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3223:3216] <= 'd0;
end

wire  [39:0]  kernel_img_mul_403[0:24];
assign kernel_img_mul_403[0] = buffer_data_4[3215:3208] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_403[1] = buffer_data_4[3223:3216] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_403[2] = buffer_data_4[3231:3224] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_403[3] = buffer_data_4[3239:3232] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_403[4] = buffer_data_4[3247:3240] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_403[5] = buffer_data_3[3215:3208] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_403[6] = buffer_data_3[3223:3216] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_403[7] = buffer_data_3[3231:3224] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_403[8] = buffer_data_3[3239:3232] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_403[9] = buffer_data_3[3247:3240] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_403[10] = buffer_data_2[3215:3208] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_403[11] = buffer_data_2[3223:3216] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_403[12] = buffer_data_2[3231:3224] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_403[13] = buffer_data_2[3239:3232] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_403[14] = buffer_data_2[3247:3240] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_403[15] = buffer_data_1[3215:3208] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_403[16] = buffer_data_1[3223:3216] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_403[17] = buffer_data_1[3231:3224] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_403[18] = buffer_data_1[3239:3232] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_403[19] = buffer_data_1[3247:3240] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_403[20] = buffer_data_0[3215:3208] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_403[21] = buffer_data_0[3223:3216] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_403[22] = buffer_data_0[3231:3224] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_403[23] = buffer_data_0[3239:3232] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_403[24] = buffer_data_0[3247:3240] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_403 = kernel_img_mul_403[0] + kernel_img_mul_403[1] + kernel_img_mul_403[2] + 
                kernel_img_mul_403[3] + kernel_img_mul_403[4] + kernel_img_mul_403[5] + 
                kernel_img_mul_403[6] + kernel_img_mul_403[7] + kernel_img_mul_403[8] + 
                kernel_img_mul_403[9] + kernel_img_mul_403[10] + kernel_img_mul_403[11] + 
                kernel_img_mul_403[12] + kernel_img_mul_403[13] + kernel_img_mul_403[14] + 
                kernel_img_mul_403[15] + kernel_img_mul_403[16] + kernel_img_mul_403[17] + 
                kernel_img_mul_403[18] + kernel_img_mul_403[19] + kernel_img_mul_403[20] + 
                kernel_img_mul_403[21] + kernel_img_mul_403[22] + kernel_img_mul_403[23] + 
                kernel_img_mul_403[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3231:3224] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3231:3224] <= kernel_img_sum_403[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3231:3224] <= 'd0;
end

wire  [39:0]  kernel_img_mul_404[0:24];
assign kernel_img_mul_404[0] = buffer_data_4[3223:3216] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_404[1] = buffer_data_4[3231:3224] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_404[2] = buffer_data_4[3239:3232] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_404[3] = buffer_data_4[3247:3240] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_404[4] = buffer_data_4[3255:3248] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_404[5] = buffer_data_3[3223:3216] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_404[6] = buffer_data_3[3231:3224] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_404[7] = buffer_data_3[3239:3232] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_404[8] = buffer_data_3[3247:3240] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_404[9] = buffer_data_3[3255:3248] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_404[10] = buffer_data_2[3223:3216] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_404[11] = buffer_data_2[3231:3224] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_404[12] = buffer_data_2[3239:3232] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_404[13] = buffer_data_2[3247:3240] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_404[14] = buffer_data_2[3255:3248] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_404[15] = buffer_data_1[3223:3216] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_404[16] = buffer_data_1[3231:3224] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_404[17] = buffer_data_1[3239:3232] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_404[18] = buffer_data_1[3247:3240] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_404[19] = buffer_data_1[3255:3248] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_404[20] = buffer_data_0[3223:3216] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_404[21] = buffer_data_0[3231:3224] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_404[22] = buffer_data_0[3239:3232] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_404[23] = buffer_data_0[3247:3240] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_404[24] = buffer_data_0[3255:3248] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_404 = kernel_img_mul_404[0] + kernel_img_mul_404[1] + kernel_img_mul_404[2] + 
                kernel_img_mul_404[3] + kernel_img_mul_404[4] + kernel_img_mul_404[5] + 
                kernel_img_mul_404[6] + kernel_img_mul_404[7] + kernel_img_mul_404[8] + 
                kernel_img_mul_404[9] + kernel_img_mul_404[10] + kernel_img_mul_404[11] + 
                kernel_img_mul_404[12] + kernel_img_mul_404[13] + kernel_img_mul_404[14] + 
                kernel_img_mul_404[15] + kernel_img_mul_404[16] + kernel_img_mul_404[17] + 
                kernel_img_mul_404[18] + kernel_img_mul_404[19] + kernel_img_mul_404[20] + 
                kernel_img_mul_404[21] + kernel_img_mul_404[22] + kernel_img_mul_404[23] + 
                kernel_img_mul_404[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3239:3232] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3239:3232] <= kernel_img_sum_404[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3239:3232] <= 'd0;
end

wire  [39:0]  kernel_img_mul_405[0:24];
assign kernel_img_mul_405[0] = buffer_data_4[3231:3224] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_405[1] = buffer_data_4[3239:3232] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_405[2] = buffer_data_4[3247:3240] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_405[3] = buffer_data_4[3255:3248] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_405[4] = buffer_data_4[3263:3256] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_405[5] = buffer_data_3[3231:3224] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_405[6] = buffer_data_3[3239:3232] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_405[7] = buffer_data_3[3247:3240] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_405[8] = buffer_data_3[3255:3248] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_405[9] = buffer_data_3[3263:3256] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_405[10] = buffer_data_2[3231:3224] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_405[11] = buffer_data_2[3239:3232] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_405[12] = buffer_data_2[3247:3240] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_405[13] = buffer_data_2[3255:3248] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_405[14] = buffer_data_2[3263:3256] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_405[15] = buffer_data_1[3231:3224] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_405[16] = buffer_data_1[3239:3232] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_405[17] = buffer_data_1[3247:3240] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_405[18] = buffer_data_1[3255:3248] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_405[19] = buffer_data_1[3263:3256] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_405[20] = buffer_data_0[3231:3224] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_405[21] = buffer_data_0[3239:3232] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_405[22] = buffer_data_0[3247:3240] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_405[23] = buffer_data_0[3255:3248] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_405[24] = buffer_data_0[3263:3256] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_405 = kernel_img_mul_405[0] + kernel_img_mul_405[1] + kernel_img_mul_405[2] + 
                kernel_img_mul_405[3] + kernel_img_mul_405[4] + kernel_img_mul_405[5] + 
                kernel_img_mul_405[6] + kernel_img_mul_405[7] + kernel_img_mul_405[8] + 
                kernel_img_mul_405[9] + kernel_img_mul_405[10] + kernel_img_mul_405[11] + 
                kernel_img_mul_405[12] + kernel_img_mul_405[13] + kernel_img_mul_405[14] + 
                kernel_img_mul_405[15] + kernel_img_mul_405[16] + kernel_img_mul_405[17] + 
                kernel_img_mul_405[18] + kernel_img_mul_405[19] + kernel_img_mul_405[20] + 
                kernel_img_mul_405[21] + kernel_img_mul_405[22] + kernel_img_mul_405[23] + 
                kernel_img_mul_405[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3247:3240] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3247:3240] <= kernel_img_sum_405[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3247:3240] <= 'd0;
end

wire  [39:0]  kernel_img_mul_406[0:24];
assign kernel_img_mul_406[0] = buffer_data_4[3239:3232] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_406[1] = buffer_data_4[3247:3240] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_406[2] = buffer_data_4[3255:3248] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_406[3] = buffer_data_4[3263:3256] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_406[4] = buffer_data_4[3271:3264] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_406[5] = buffer_data_3[3239:3232] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_406[6] = buffer_data_3[3247:3240] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_406[7] = buffer_data_3[3255:3248] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_406[8] = buffer_data_3[3263:3256] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_406[9] = buffer_data_3[3271:3264] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_406[10] = buffer_data_2[3239:3232] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_406[11] = buffer_data_2[3247:3240] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_406[12] = buffer_data_2[3255:3248] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_406[13] = buffer_data_2[3263:3256] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_406[14] = buffer_data_2[3271:3264] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_406[15] = buffer_data_1[3239:3232] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_406[16] = buffer_data_1[3247:3240] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_406[17] = buffer_data_1[3255:3248] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_406[18] = buffer_data_1[3263:3256] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_406[19] = buffer_data_1[3271:3264] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_406[20] = buffer_data_0[3239:3232] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_406[21] = buffer_data_0[3247:3240] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_406[22] = buffer_data_0[3255:3248] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_406[23] = buffer_data_0[3263:3256] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_406[24] = buffer_data_0[3271:3264] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_406 = kernel_img_mul_406[0] + kernel_img_mul_406[1] + kernel_img_mul_406[2] + 
                kernel_img_mul_406[3] + kernel_img_mul_406[4] + kernel_img_mul_406[5] + 
                kernel_img_mul_406[6] + kernel_img_mul_406[7] + kernel_img_mul_406[8] + 
                kernel_img_mul_406[9] + kernel_img_mul_406[10] + kernel_img_mul_406[11] + 
                kernel_img_mul_406[12] + kernel_img_mul_406[13] + kernel_img_mul_406[14] + 
                kernel_img_mul_406[15] + kernel_img_mul_406[16] + kernel_img_mul_406[17] + 
                kernel_img_mul_406[18] + kernel_img_mul_406[19] + kernel_img_mul_406[20] + 
                kernel_img_mul_406[21] + kernel_img_mul_406[22] + kernel_img_mul_406[23] + 
                kernel_img_mul_406[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3255:3248] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3255:3248] <= kernel_img_sum_406[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3255:3248] <= 'd0;
end

wire  [39:0]  kernel_img_mul_407[0:24];
assign kernel_img_mul_407[0] = buffer_data_4[3247:3240] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_407[1] = buffer_data_4[3255:3248] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_407[2] = buffer_data_4[3263:3256] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_407[3] = buffer_data_4[3271:3264] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_407[4] = buffer_data_4[3279:3272] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_407[5] = buffer_data_3[3247:3240] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_407[6] = buffer_data_3[3255:3248] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_407[7] = buffer_data_3[3263:3256] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_407[8] = buffer_data_3[3271:3264] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_407[9] = buffer_data_3[3279:3272] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_407[10] = buffer_data_2[3247:3240] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_407[11] = buffer_data_2[3255:3248] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_407[12] = buffer_data_2[3263:3256] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_407[13] = buffer_data_2[3271:3264] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_407[14] = buffer_data_2[3279:3272] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_407[15] = buffer_data_1[3247:3240] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_407[16] = buffer_data_1[3255:3248] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_407[17] = buffer_data_1[3263:3256] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_407[18] = buffer_data_1[3271:3264] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_407[19] = buffer_data_1[3279:3272] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_407[20] = buffer_data_0[3247:3240] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_407[21] = buffer_data_0[3255:3248] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_407[22] = buffer_data_0[3263:3256] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_407[23] = buffer_data_0[3271:3264] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_407[24] = buffer_data_0[3279:3272] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_407 = kernel_img_mul_407[0] + kernel_img_mul_407[1] + kernel_img_mul_407[2] + 
                kernel_img_mul_407[3] + kernel_img_mul_407[4] + kernel_img_mul_407[5] + 
                kernel_img_mul_407[6] + kernel_img_mul_407[7] + kernel_img_mul_407[8] + 
                kernel_img_mul_407[9] + kernel_img_mul_407[10] + kernel_img_mul_407[11] + 
                kernel_img_mul_407[12] + kernel_img_mul_407[13] + kernel_img_mul_407[14] + 
                kernel_img_mul_407[15] + kernel_img_mul_407[16] + kernel_img_mul_407[17] + 
                kernel_img_mul_407[18] + kernel_img_mul_407[19] + kernel_img_mul_407[20] + 
                kernel_img_mul_407[21] + kernel_img_mul_407[22] + kernel_img_mul_407[23] + 
                kernel_img_mul_407[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3263:3256] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3263:3256] <= kernel_img_sum_407[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3263:3256] <= 'd0;
end

wire  [39:0]  kernel_img_mul_408[0:24];
assign kernel_img_mul_408[0] = buffer_data_4[3255:3248] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_408[1] = buffer_data_4[3263:3256] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_408[2] = buffer_data_4[3271:3264] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_408[3] = buffer_data_4[3279:3272] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_408[4] = buffer_data_4[3287:3280] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_408[5] = buffer_data_3[3255:3248] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_408[6] = buffer_data_3[3263:3256] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_408[7] = buffer_data_3[3271:3264] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_408[8] = buffer_data_3[3279:3272] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_408[9] = buffer_data_3[3287:3280] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_408[10] = buffer_data_2[3255:3248] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_408[11] = buffer_data_2[3263:3256] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_408[12] = buffer_data_2[3271:3264] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_408[13] = buffer_data_2[3279:3272] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_408[14] = buffer_data_2[3287:3280] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_408[15] = buffer_data_1[3255:3248] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_408[16] = buffer_data_1[3263:3256] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_408[17] = buffer_data_1[3271:3264] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_408[18] = buffer_data_1[3279:3272] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_408[19] = buffer_data_1[3287:3280] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_408[20] = buffer_data_0[3255:3248] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_408[21] = buffer_data_0[3263:3256] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_408[22] = buffer_data_0[3271:3264] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_408[23] = buffer_data_0[3279:3272] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_408[24] = buffer_data_0[3287:3280] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_408 = kernel_img_mul_408[0] + kernel_img_mul_408[1] + kernel_img_mul_408[2] + 
                kernel_img_mul_408[3] + kernel_img_mul_408[4] + kernel_img_mul_408[5] + 
                kernel_img_mul_408[6] + kernel_img_mul_408[7] + kernel_img_mul_408[8] + 
                kernel_img_mul_408[9] + kernel_img_mul_408[10] + kernel_img_mul_408[11] + 
                kernel_img_mul_408[12] + kernel_img_mul_408[13] + kernel_img_mul_408[14] + 
                kernel_img_mul_408[15] + kernel_img_mul_408[16] + kernel_img_mul_408[17] + 
                kernel_img_mul_408[18] + kernel_img_mul_408[19] + kernel_img_mul_408[20] + 
                kernel_img_mul_408[21] + kernel_img_mul_408[22] + kernel_img_mul_408[23] + 
                kernel_img_mul_408[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3271:3264] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3271:3264] <= kernel_img_sum_408[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3271:3264] <= 'd0;
end

wire  [39:0]  kernel_img_mul_409[0:24];
assign kernel_img_mul_409[0] = buffer_data_4[3263:3256] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_409[1] = buffer_data_4[3271:3264] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_409[2] = buffer_data_4[3279:3272] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_409[3] = buffer_data_4[3287:3280] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_409[4] = buffer_data_4[3295:3288] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_409[5] = buffer_data_3[3263:3256] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_409[6] = buffer_data_3[3271:3264] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_409[7] = buffer_data_3[3279:3272] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_409[8] = buffer_data_3[3287:3280] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_409[9] = buffer_data_3[3295:3288] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_409[10] = buffer_data_2[3263:3256] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_409[11] = buffer_data_2[3271:3264] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_409[12] = buffer_data_2[3279:3272] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_409[13] = buffer_data_2[3287:3280] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_409[14] = buffer_data_2[3295:3288] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_409[15] = buffer_data_1[3263:3256] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_409[16] = buffer_data_1[3271:3264] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_409[17] = buffer_data_1[3279:3272] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_409[18] = buffer_data_1[3287:3280] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_409[19] = buffer_data_1[3295:3288] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_409[20] = buffer_data_0[3263:3256] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_409[21] = buffer_data_0[3271:3264] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_409[22] = buffer_data_0[3279:3272] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_409[23] = buffer_data_0[3287:3280] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_409[24] = buffer_data_0[3295:3288] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_409 = kernel_img_mul_409[0] + kernel_img_mul_409[1] + kernel_img_mul_409[2] + 
                kernel_img_mul_409[3] + kernel_img_mul_409[4] + kernel_img_mul_409[5] + 
                kernel_img_mul_409[6] + kernel_img_mul_409[7] + kernel_img_mul_409[8] + 
                kernel_img_mul_409[9] + kernel_img_mul_409[10] + kernel_img_mul_409[11] + 
                kernel_img_mul_409[12] + kernel_img_mul_409[13] + kernel_img_mul_409[14] + 
                kernel_img_mul_409[15] + kernel_img_mul_409[16] + kernel_img_mul_409[17] + 
                kernel_img_mul_409[18] + kernel_img_mul_409[19] + kernel_img_mul_409[20] + 
                kernel_img_mul_409[21] + kernel_img_mul_409[22] + kernel_img_mul_409[23] + 
                kernel_img_mul_409[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3279:3272] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3279:3272] <= kernel_img_sum_409[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3279:3272] <= 'd0;
end

wire  [39:0]  kernel_img_mul_410[0:24];
assign kernel_img_mul_410[0] = buffer_data_4[3271:3264] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_410[1] = buffer_data_4[3279:3272] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_410[2] = buffer_data_4[3287:3280] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_410[3] = buffer_data_4[3295:3288] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_410[4] = buffer_data_4[3303:3296] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_410[5] = buffer_data_3[3271:3264] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_410[6] = buffer_data_3[3279:3272] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_410[7] = buffer_data_3[3287:3280] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_410[8] = buffer_data_3[3295:3288] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_410[9] = buffer_data_3[3303:3296] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_410[10] = buffer_data_2[3271:3264] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_410[11] = buffer_data_2[3279:3272] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_410[12] = buffer_data_2[3287:3280] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_410[13] = buffer_data_2[3295:3288] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_410[14] = buffer_data_2[3303:3296] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_410[15] = buffer_data_1[3271:3264] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_410[16] = buffer_data_1[3279:3272] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_410[17] = buffer_data_1[3287:3280] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_410[18] = buffer_data_1[3295:3288] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_410[19] = buffer_data_1[3303:3296] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_410[20] = buffer_data_0[3271:3264] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_410[21] = buffer_data_0[3279:3272] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_410[22] = buffer_data_0[3287:3280] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_410[23] = buffer_data_0[3295:3288] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_410[24] = buffer_data_0[3303:3296] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_410 = kernel_img_mul_410[0] + kernel_img_mul_410[1] + kernel_img_mul_410[2] + 
                kernel_img_mul_410[3] + kernel_img_mul_410[4] + kernel_img_mul_410[5] + 
                kernel_img_mul_410[6] + kernel_img_mul_410[7] + kernel_img_mul_410[8] + 
                kernel_img_mul_410[9] + kernel_img_mul_410[10] + kernel_img_mul_410[11] + 
                kernel_img_mul_410[12] + kernel_img_mul_410[13] + kernel_img_mul_410[14] + 
                kernel_img_mul_410[15] + kernel_img_mul_410[16] + kernel_img_mul_410[17] + 
                kernel_img_mul_410[18] + kernel_img_mul_410[19] + kernel_img_mul_410[20] + 
                kernel_img_mul_410[21] + kernel_img_mul_410[22] + kernel_img_mul_410[23] + 
                kernel_img_mul_410[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3287:3280] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3287:3280] <= kernel_img_sum_410[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3287:3280] <= 'd0;
end

wire  [39:0]  kernel_img_mul_411[0:24];
assign kernel_img_mul_411[0] = buffer_data_4[3279:3272] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_411[1] = buffer_data_4[3287:3280] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_411[2] = buffer_data_4[3295:3288] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_411[3] = buffer_data_4[3303:3296] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_411[4] = buffer_data_4[3311:3304] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_411[5] = buffer_data_3[3279:3272] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_411[6] = buffer_data_3[3287:3280] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_411[7] = buffer_data_3[3295:3288] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_411[8] = buffer_data_3[3303:3296] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_411[9] = buffer_data_3[3311:3304] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_411[10] = buffer_data_2[3279:3272] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_411[11] = buffer_data_2[3287:3280] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_411[12] = buffer_data_2[3295:3288] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_411[13] = buffer_data_2[3303:3296] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_411[14] = buffer_data_2[3311:3304] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_411[15] = buffer_data_1[3279:3272] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_411[16] = buffer_data_1[3287:3280] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_411[17] = buffer_data_1[3295:3288] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_411[18] = buffer_data_1[3303:3296] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_411[19] = buffer_data_1[3311:3304] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_411[20] = buffer_data_0[3279:3272] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_411[21] = buffer_data_0[3287:3280] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_411[22] = buffer_data_0[3295:3288] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_411[23] = buffer_data_0[3303:3296] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_411[24] = buffer_data_0[3311:3304] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_411 = kernel_img_mul_411[0] + kernel_img_mul_411[1] + kernel_img_mul_411[2] + 
                kernel_img_mul_411[3] + kernel_img_mul_411[4] + kernel_img_mul_411[5] + 
                kernel_img_mul_411[6] + kernel_img_mul_411[7] + kernel_img_mul_411[8] + 
                kernel_img_mul_411[9] + kernel_img_mul_411[10] + kernel_img_mul_411[11] + 
                kernel_img_mul_411[12] + kernel_img_mul_411[13] + kernel_img_mul_411[14] + 
                kernel_img_mul_411[15] + kernel_img_mul_411[16] + kernel_img_mul_411[17] + 
                kernel_img_mul_411[18] + kernel_img_mul_411[19] + kernel_img_mul_411[20] + 
                kernel_img_mul_411[21] + kernel_img_mul_411[22] + kernel_img_mul_411[23] + 
                kernel_img_mul_411[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3295:3288] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3295:3288] <= kernel_img_sum_411[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3295:3288] <= 'd0;
end

wire  [39:0]  kernel_img_mul_412[0:24];
assign kernel_img_mul_412[0] = buffer_data_4[3287:3280] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_412[1] = buffer_data_4[3295:3288] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_412[2] = buffer_data_4[3303:3296] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_412[3] = buffer_data_4[3311:3304] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_412[4] = buffer_data_4[3319:3312] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_412[5] = buffer_data_3[3287:3280] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_412[6] = buffer_data_3[3295:3288] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_412[7] = buffer_data_3[3303:3296] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_412[8] = buffer_data_3[3311:3304] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_412[9] = buffer_data_3[3319:3312] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_412[10] = buffer_data_2[3287:3280] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_412[11] = buffer_data_2[3295:3288] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_412[12] = buffer_data_2[3303:3296] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_412[13] = buffer_data_2[3311:3304] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_412[14] = buffer_data_2[3319:3312] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_412[15] = buffer_data_1[3287:3280] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_412[16] = buffer_data_1[3295:3288] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_412[17] = buffer_data_1[3303:3296] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_412[18] = buffer_data_1[3311:3304] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_412[19] = buffer_data_1[3319:3312] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_412[20] = buffer_data_0[3287:3280] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_412[21] = buffer_data_0[3295:3288] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_412[22] = buffer_data_0[3303:3296] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_412[23] = buffer_data_0[3311:3304] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_412[24] = buffer_data_0[3319:3312] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_412 = kernel_img_mul_412[0] + kernel_img_mul_412[1] + kernel_img_mul_412[2] + 
                kernel_img_mul_412[3] + kernel_img_mul_412[4] + kernel_img_mul_412[5] + 
                kernel_img_mul_412[6] + kernel_img_mul_412[7] + kernel_img_mul_412[8] + 
                kernel_img_mul_412[9] + kernel_img_mul_412[10] + kernel_img_mul_412[11] + 
                kernel_img_mul_412[12] + kernel_img_mul_412[13] + kernel_img_mul_412[14] + 
                kernel_img_mul_412[15] + kernel_img_mul_412[16] + kernel_img_mul_412[17] + 
                kernel_img_mul_412[18] + kernel_img_mul_412[19] + kernel_img_mul_412[20] + 
                kernel_img_mul_412[21] + kernel_img_mul_412[22] + kernel_img_mul_412[23] + 
                kernel_img_mul_412[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3303:3296] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3303:3296] <= kernel_img_sum_412[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3303:3296] <= 'd0;
end

wire  [39:0]  kernel_img_mul_413[0:24];
assign kernel_img_mul_413[0] = buffer_data_4[3295:3288] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_413[1] = buffer_data_4[3303:3296] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_413[2] = buffer_data_4[3311:3304] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_413[3] = buffer_data_4[3319:3312] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_413[4] = buffer_data_4[3327:3320] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_413[5] = buffer_data_3[3295:3288] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_413[6] = buffer_data_3[3303:3296] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_413[7] = buffer_data_3[3311:3304] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_413[8] = buffer_data_3[3319:3312] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_413[9] = buffer_data_3[3327:3320] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_413[10] = buffer_data_2[3295:3288] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_413[11] = buffer_data_2[3303:3296] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_413[12] = buffer_data_2[3311:3304] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_413[13] = buffer_data_2[3319:3312] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_413[14] = buffer_data_2[3327:3320] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_413[15] = buffer_data_1[3295:3288] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_413[16] = buffer_data_1[3303:3296] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_413[17] = buffer_data_1[3311:3304] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_413[18] = buffer_data_1[3319:3312] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_413[19] = buffer_data_1[3327:3320] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_413[20] = buffer_data_0[3295:3288] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_413[21] = buffer_data_0[3303:3296] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_413[22] = buffer_data_0[3311:3304] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_413[23] = buffer_data_0[3319:3312] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_413[24] = buffer_data_0[3327:3320] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_413 = kernel_img_mul_413[0] + kernel_img_mul_413[1] + kernel_img_mul_413[2] + 
                kernel_img_mul_413[3] + kernel_img_mul_413[4] + kernel_img_mul_413[5] + 
                kernel_img_mul_413[6] + kernel_img_mul_413[7] + kernel_img_mul_413[8] + 
                kernel_img_mul_413[9] + kernel_img_mul_413[10] + kernel_img_mul_413[11] + 
                kernel_img_mul_413[12] + kernel_img_mul_413[13] + kernel_img_mul_413[14] + 
                kernel_img_mul_413[15] + kernel_img_mul_413[16] + kernel_img_mul_413[17] + 
                kernel_img_mul_413[18] + kernel_img_mul_413[19] + kernel_img_mul_413[20] + 
                kernel_img_mul_413[21] + kernel_img_mul_413[22] + kernel_img_mul_413[23] + 
                kernel_img_mul_413[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3311:3304] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3311:3304] <= kernel_img_sum_413[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3311:3304] <= 'd0;
end

wire  [39:0]  kernel_img_mul_414[0:24];
assign kernel_img_mul_414[0] = buffer_data_4[3303:3296] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_414[1] = buffer_data_4[3311:3304] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_414[2] = buffer_data_4[3319:3312] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_414[3] = buffer_data_4[3327:3320] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_414[4] = buffer_data_4[3335:3328] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_414[5] = buffer_data_3[3303:3296] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_414[6] = buffer_data_3[3311:3304] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_414[7] = buffer_data_3[3319:3312] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_414[8] = buffer_data_3[3327:3320] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_414[9] = buffer_data_3[3335:3328] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_414[10] = buffer_data_2[3303:3296] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_414[11] = buffer_data_2[3311:3304] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_414[12] = buffer_data_2[3319:3312] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_414[13] = buffer_data_2[3327:3320] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_414[14] = buffer_data_2[3335:3328] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_414[15] = buffer_data_1[3303:3296] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_414[16] = buffer_data_1[3311:3304] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_414[17] = buffer_data_1[3319:3312] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_414[18] = buffer_data_1[3327:3320] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_414[19] = buffer_data_1[3335:3328] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_414[20] = buffer_data_0[3303:3296] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_414[21] = buffer_data_0[3311:3304] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_414[22] = buffer_data_0[3319:3312] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_414[23] = buffer_data_0[3327:3320] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_414[24] = buffer_data_0[3335:3328] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_414 = kernel_img_mul_414[0] + kernel_img_mul_414[1] + kernel_img_mul_414[2] + 
                kernel_img_mul_414[3] + kernel_img_mul_414[4] + kernel_img_mul_414[5] + 
                kernel_img_mul_414[6] + kernel_img_mul_414[7] + kernel_img_mul_414[8] + 
                kernel_img_mul_414[9] + kernel_img_mul_414[10] + kernel_img_mul_414[11] + 
                kernel_img_mul_414[12] + kernel_img_mul_414[13] + kernel_img_mul_414[14] + 
                kernel_img_mul_414[15] + kernel_img_mul_414[16] + kernel_img_mul_414[17] + 
                kernel_img_mul_414[18] + kernel_img_mul_414[19] + kernel_img_mul_414[20] + 
                kernel_img_mul_414[21] + kernel_img_mul_414[22] + kernel_img_mul_414[23] + 
                kernel_img_mul_414[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3319:3312] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3319:3312] <= kernel_img_sum_414[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3319:3312] <= 'd0;
end

wire  [39:0]  kernel_img_mul_415[0:24];
assign kernel_img_mul_415[0] = buffer_data_4[3311:3304] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_415[1] = buffer_data_4[3319:3312] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_415[2] = buffer_data_4[3327:3320] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_415[3] = buffer_data_4[3335:3328] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_415[4] = buffer_data_4[3343:3336] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_415[5] = buffer_data_3[3311:3304] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_415[6] = buffer_data_3[3319:3312] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_415[7] = buffer_data_3[3327:3320] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_415[8] = buffer_data_3[3335:3328] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_415[9] = buffer_data_3[3343:3336] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_415[10] = buffer_data_2[3311:3304] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_415[11] = buffer_data_2[3319:3312] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_415[12] = buffer_data_2[3327:3320] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_415[13] = buffer_data_2[3335:3328] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_415[14] = buffer_data_2[3343:3336] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_415[15] = buffer_data_1[3311:3304] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_415[16] = buffer_data_1[3319:3312] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_415[17] = buffer_data_1[3327:3320] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_415[18] = buffer_data_1[3335:3328] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_415[19] = buffer_data_1[3343:3336] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_415[20] = buffer_data_0[3311:3304] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_415[21] = buffer_data_0[3319:3312] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_415[22] = buffer_data_0[3327:3320] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_415[23] = buffer_data_0[3335:3328] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_415[24] = buffer_data_0[3343:3336] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_415 = kernel_img_mul_415[0] + kernel_img_mul_415[1] + kernel_img_mul_415[2] + 
                kernel_img_mul_415[3] + kernel_img_mul_415[4] + kernel_img_mul_415[5] + 
                kernel_img_mul_415[6] + kernel_img_mul_415[7] + kernel_img_mul_415[8] + 
                kernel_img_mul_415[9] + kernel_img_mul_415[10] + kernel_img_mul_415[11] + 
                kernel_img_mul_415[12] + kernel_img_mul_415[13] + kernel_img_mul_415[14] + 
                kernel_img_mul_415[15] + kernel_img_mul_415[16] + kernel_img_mul_415[17] + 
                kernel_img_mul_415[18] + kernel_img_mul_415[19] + kernel_img_mul_415[20] + 
                kernel_img_mul_415[21] + kernel_img_mul_415[22] + kernel_img_mul_415[23] + 
                kernel_img_mul_415[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3327:3320] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3327:3320] <= kernel_img_sum_415[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3327:3320] <= 'd0;
end

wire  [39:0]  kernel_img_mul_416[0:24];
assign kernel_img_mul_416[0] = buffer_data_4[3319:3312] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_416[1] = buffer_data_4[3327:3320] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_416[2] = buffer_data_4[3335:3328] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_416[3] = buffer_data_4[3343:3336] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_416[4] = buffer_data_4[3351:3344] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_416[5] = buffer_data_3[3319:3312] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_416[6] = buffer_data_3[3327:3320] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_416[7] = buffer_data_3[3335:3328] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_416[8] = buffer_data_3[3343:3336] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_416[9] = buffer_data_3[3351:3344] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_416[10] = buffer_data_2[3319:3312] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_416[11] = buffer_data_2[3327:3320] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_416[12] = buffer_data_2[3335:3328] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_416[13] = buffer_data_2[3343:3336] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_416[14] = buffer_data_2[3351:3344] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_416[15] = buffer_data_1[3319:3312] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_416[16] = buffer_data_1[3327:3320] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_416[17] = buffer_data_1[3335:3328] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_416[18] = buffer_data_1[3343:3336] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_416[19] = buffer_data_1[3351:3344] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_416[20] = buffer_data_0[3319:3312] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_416[21] = buffer_data_0[3327:3320] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_416[22] = buffer_data_0[3335:3328] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_416[23] = buffer_data_0[3343:3336] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_416[24] = buffer_data_0[3351:3344] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_416 = kernel_img_mul_416[0] + kernel_img_mul_416[1] + kernel_img_mul_416[2] + 
                kernel_img_mul_416[3] + kernel_img_mul_416[4] + kernel_img_mul_416[5] + 
                kernel_img_mul_416[6] + kernel_img_mul_416[7] + kernel_img_mul_416[8] + 
                kernel_img_mul_416[9] + kernel_img_mul_416[10] + kernel_img_mul_416[11] + 
                kernel_img_mul_416[12] + kernel_img_mul_416[13] + kernel_img_mul_416[14] + 
                kernel_img_mul_416[15] + kernel_img_mul_416[16] + kernel_img_mul_416[17] + 
                kernel_img_mul_416[18] + kernel_img_mul_416[19] + kernel_img_mul_416[20] + 
                kernel_img_mul_416[21] + kernel_img_mul_416[22] + kernel_img_mul_416[23] + 
                kernel_img_mul_416[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3335:3328] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3335:3328] <= kernel_img_sum_416[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3335:3328] <= 'd0;
end

wire  [39:0]  kernel_img_mul_417[0:24];
assign kernel_img_mul_417[0] = buffer_data_4[3327:3320] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_417[1] = buffer_data_4[3335:3328] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_417[2] = buffer_data_4[3343:3336] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_417[3] = buffer_data_4[3351:3344] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_417[4] = buffer_data_4[3359:3352] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_417[5] = buffer_data_3[3327:3320] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_417[6] = buffer_data_3[3335:3328] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_417[7] = buffer_data_3[3343:3336] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_417[8] = buffer_data_3[3351:3344] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_417[9] = buffer_data_3[3359:3352] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_417[10] = buffer_data_2[3327:3320] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_417[11] = buffer_data_2[3335:3328] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_417[12] = buffer_data_2[3343:3336] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_417[13] = buffer_data_2[3351:3344] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_417[14] = buffer_data_2[3359:3352] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_417[15] = buffer_data_1[3327:3320] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_417[16] = buffer_data_1[3335:3328] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_417[17] = buffer_data_1[3343:3336] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_417[18] = buffer_data_1[3351:3344] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_417[19] = buffer_data_1[3359:3352] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_417[20] = buffer_data_0[3327:3320] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_417[21] = buffer_data_0[3335:3328] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_417[22] = buffer_data_0[3343:3336] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_417[23] = buffer_data_0[3351:3344] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_417[24] = buffer_data_0[3359:3352] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_417 = kernel_img_mul_417[0] + kernel_img_mul_417[1] + kernel_img_mul_417[2] + 
                kernel_img_mul_417[3] + kernel_img_mul_417[4] + kernel_img_mul_417[5] + 
                kernel_img_mul_417[6] + kernel_img_mul_417[7] + kernel_img_mul_417[8] + 
                kernel_img_mul_417[9] + kernel_img_mul_417[10] + kernel_img_mul_417[11] + 
                kernel_img_mul_417[12] + kernel_img_mul_417[13] + kernel_img_mul_417[14] + 
                kernel_img_mul_417[15] + kernel_img_mul_417[16] + kernel_img_mul_417[17] + 
                kernel_img_mul_417[18] + kernel_img_mul_417[19] + kernel_img_mul_417[20] + 
                kernel_img_mul_417[21] + kernel_img_mul_417[22] + kernel_img_mul_417[23] + 
                kernel_img_mul_417[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3343:3336] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3343:3336] <= kernel_img_sum_417[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3343:3336] <= 'd0;
end

wire  [39:0]  kernel_img_mul_418[0:24];
assign kernel_img_mul_418[0] = buffer_data_4[3335:3328] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_418[1] = buffer_data_4[3343:3336] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_418[2] = buffer_data_4[3351:3344] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_418[3] = buffer_data_4[3359:3352] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_418[4] = buffer_data_4[3367:3360] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_418[5] = buffer_data_3[3335:3328] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_418[6] = buffer_data_3[3343:3336] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_418[7] = buffer_data_3[3351:3344] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_418[8] = buffer_data_3[3359:3352] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_418[9] = buffer_data_3[3367:3360] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_418[10] = buffer_data_2[3335:3328] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_418[11] = buffer_data_2[3343:3336] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_418[12] = buffer_data_2[3351:3344] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_418[13] = buffer_data_2[3359:3352] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_418[14] = buffer_data_2[3367:3360] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_418[15] = buffer_data_1[3335:3328] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_418[16] = buffer_data_1[3343:3336] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_418[17] = buffer_data_1[3351:3344] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_418[18] = buffer_data_1[3359:3352] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_418[19] = buffer_data_1[3367:3360] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_418[20] = buffer_data_0[3335:3328] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_418[21] = buffer_data_0[3343:3336] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_418[22] = buffer_data_0[3351:3344] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_418[23] = buffer_data_0[3359:3352] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_418[24] = buffer_data_0[3367:3360] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_418 = kernel_img_mul_418[0] + kernel_img_mul_418[1] + kernel_img_mul_418[2] + 
                kernel_img_mul_418[3] + kernel_img_mul_418[4] + kernel_img_mul_418[5] + 
                kernel_img_mul_418[6] + kernel_img_mul_418[7] + kernel_img_mul_418[8] + 
                kernel_img_mul_418[9] + kernel_img_mul_418[10] + kernel_img_mul_418[11] + 
                kernel_img_mul_418[12] + kernel_img_mul_418[13] + kernel_img_mul_418[14] + 
                kernel_img_mul_418[15] + kernel_img_mul_418[16] + kernel_img_mul_418[17] + 
                kernel_img_mul_418[18] + kernel_img_mul_418[19] + kernel_img_mul_418[20] + 
                kernel_img_mul_418[21] + kernel_img_mul_418[22] + kernel_img_mul_418[23] + 
                kernel_img_mul_418[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3351:3344] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3351:3344] <= kernel_img_sum_418[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3351:3344] <= 'd0;
end

wire  [39:0]  kernel_img_mul_419[0:24];
assign kernel_img_mul_419[0] = buffer_data_4[3343:3336] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_419[1] = buffer_data_4[3351:3344] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_419[2] = buffer_data_4[3359:3352] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_419[3] = buffer_data_4[3367:3360] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_419[4] = buffer_data_4[3375:3368] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_419[5] = buffer_data_3[3343:3336] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_419[6] = buffer_data_3[3351:3344] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_419[7] = buffer_data_3[3359:3352] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_419[8] = buffer_data_3[3367:3360] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_419[9] = buffer_data_3[3375:3368] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_419[10] = buffer_data_2[3343:3336] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_419[11] = buffer_data_2[3351:3344] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_419[12] = buffer_data_2[3359:3352] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_419[13] = buffer_data_2[3367:3360] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_419[14] = buffer_data_2[3375:3368] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_419[15] = buffer_data_1[3343:3336] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_419[16] = buffer_data_1[3351:3344] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_419[17] = buffer_data_1[3359:3352] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_419[18] = buffer_data_1[3367:3360] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_419[19] = buffer_data_1[3375:3368] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_419[20] = buffer_data_0[3343:3336] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_419[21] = buffer_data_0[3351:3344] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_419[22] = buffer_data_0[3359:3352] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_419[23] = buffer_data_0[3367:3360] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_419[24] = buffer_data_0[3375:3368] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_419 = kernel_img_mul_419[0] + kernel_img_mul_419[1] + kernel_img_mul_419[2] + 
                kernel_img_mul_419[3] + kernel_img_mul_419[4] + kernel_img_mul_419[5] + 
                kernel_img_mul_419[6] + kernel_img_mul_419[7] + kernel_img_mul_419[8] + 
                kernel_img_mul_419[9] + kernel_img_mul_419[10] + kernel_img_mul_419[11] + 
                kernel_img_mul_419[12] + kernel_img_mul_419[13] + kernel_img_mul_419[14] + 
                kernel_img_mul_419[15] + kernel_img_mul_419[16] + kernel_img_mul_419[17] + 
                kernel_img_mul_419[18] + kernel_img_mul_419[19] + kernel_img_mul_419[20] + 
                kernel_img_mul_419[21] + kernel_img_mul_419[22] + kernel_img_mul_419[23] + 
                kernel_img_mul_419[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3359:3352] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3359:3352] <= kernel_img_sum_419[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3359:3352] <= 'd0;
end

wire  [39:0]  kernel_img_mul_420[0:24];
assign kernel_img_mul_420[0] = buffer_data_4[3351:3344] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_420[1] = buffer_data_4[3359:3352] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_420[2] = buffer_data_4[3367:3360] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_420[3] = buffer_data_4[3375:3368] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_420[4] = buffer_data_4[3383:3376] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_420[5] = buffer_data_3[3351:3344] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_420[6] = buffer_data_3[3359:3352] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_420[7] = buffer_data_3[3367:3360] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_420[8] = buffer_data_3[3375:3368] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_420[9] = buffer_data_3[3383:3376] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_420[10] = buffer_data_2[3351:3344] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_420[11] = buffer_data_2[3359:3352] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_420[12] = buffer_data_2[3367:3360] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_420[13] = buffer_data_2[3375:3368] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_420[14] = buffer_data_2[3383:3376] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_420[15] = buffer_data_1[3351:3344] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_420[16] = buffer_data_1[3359:3352] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_420[17] = buffer_data_1[3367:3360] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_420[18] = buffer_data_1[3375:3368] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_420[19] = buffer_data_1[3383:3376] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_420[20] = buffer_data_0[3351:3344] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_420[21] = buffer_data_0[3359:3352] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_420[22] = buffer_data_0[3367:3360] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_420[23] = buffer_data_0[3375:3368] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_420[24] = buffer_data_0[3383:3376] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_420 = kernel_img_mul_420[0] + kernel_img_mul_420[1] + kernel_img_mul_420[2] + 
                kernel_img_mul_420[3] + kernel_img_mul_420[4] + kernel_img_mul_420[5] + 
                kernel_img_mul_420[6] + kernel_img_mul_420[7] + kernel_img_mul_420[8] + 
                kernel_img_mul_420[9] + kernel_img_mul_420[10] + kernel_img_mul_420[11] + 
                kernel_img_mul_420[12] + kernel_img_mul_420[13] + kernel_img_mul_420[14] + 
                kernel_img_mul_420[15] + kernel_img_mul_420[16] + kernel_img_mul_420[17] + 
                kernel_img_mul_420[18] + kernel_img_mul_420[19] + kernel_img_mul_420[20] + 
                kernel_img_mul_420[21] + kernel_img_mul_420[22] + kernel_img_mul_420[23] + 
                kernel_img_mul_420[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3367:3360] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3367:3360] <= kernel_img_sum_420[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3367:3360] <= 'd0;
end

wire  [39:0]  kernel_img_mul_421[0:24];
assign kernel_img_mul_421[0] = buffer_data_4[3359:3352] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_421[1] = buffer_data_4[3367:3360] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_421[2] = buffer_data_4[3375:3368] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_421[3] = buffer_data_4[3383:3376] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_421[4] = buffer_data_4[3391:3384] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_421[5] = buffer_data_3[3359:3352] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_421[6] = buffer_data_3[3367:3360] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_421[7] = buffer_data_3[3375:3368] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_421[8] = buffer_data_3[3383:3376] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_421[9] = buffer_data_3[3391:3384] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_421[10] = buffer_data_2[3359:3352] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_421[11] = buffer_data_2[3367:3360] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_421[12] = buffer_data_2[3375:3368] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_421[13] = buffer_data_2[3383:3376] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_421[14] = buffer_data_2[3391:3384] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_421[15] = buffer_data_1[3359:3352] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_421[16] = buffer_data_1[3367:3360] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_421[17] = buffer_data_1[3375:3368] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_421[18] = buffer_data_1[3383:3376] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_421[19] = buffer_data_1[3391:3384] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_421[20] = buffer_data_0[3359:3352] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_421[21] = buffer_data_0[3367:3360] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_421[22] = buffer_data_0[3375:3368] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_421[23] = buffer_data_0[3383:3376] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_421[24] = buffer_data_0[3391:3384] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_421 = kernel_img_mul_421[0] + kernel_img_mul_421[1] + kernel_img_mul_421[2] + 
                kernel_img_mul_421[3] + kernel_img_mul_421[4] + kernel_img_mul_421[5] + 
                kernel_img_mul_421[6] + kernel_img_mul_421[7] + kernel_img_mul_421[8] + 
                kernel_img_mul_421[9] + kernel_img_mul_421[10] + kernel_img_mul_421[11] + 
                kernel_img_mul_421[12] + kernel_img_mul_421[13] + kernel_img_mul_421[14] + 
                kernel_img_mul_421[15] + kernel_img_mul_421[16] + kernel_img_mul_421[17] + 
                kernel_img_mul_421[18] + kernel_img_mul_421[19] + kernel_img_mul_421[20] + 
                kernel_img_mul_421[21] + kernel_img_mul_421[22] + kernel_img_mul_421[23] + 
                kernel_img_mul_421[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3375:3368] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3375:3368] <= kernel_img_sum_421[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3375:3368] <= 'd0;
end

wire  [39:0]  kernel_img_mul_422[0:24];
assign kernel_img_mul_422[0] = buffer_data_4[3367:3360] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_422[1] = buffer_data_4[3375:3368] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_422[2] = buffer_data_4[3383:3376] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_422[3] = buffer_data_4[3391:3384] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_422[4] = buffer_data_4[3399:3392] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_422[5] = buffer_data_3[3367:3360] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_422[6] = buffer_data_3[3375:3368] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_422[7] = buffer_data_3[3383:3376] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_422[8] = buffer_data_3[3391:3384] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_422[9] = buffer_data_3[3399:3392] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_422[10] = buffer_data_2[3367:3360] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_422[11] = buffer_data_2[3375:3368] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_422[12] = buffer_data_2[3383:3376] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_422[13] = buffer_data_2[3391:3384] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_422[14] = buffer_data_2[3399:3392] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_422[15] = buffer_data_1[3367:3360] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_422[16] = buffer_data_1[3375:3368] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_422[17] = buffer_data_1[3383:3376] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_422[18] = buffer_data_1[3391:3384] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_422[19] = buffer_data_1[3399:3392] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_422[20] = buffer_data_0[3367:3360] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_422[21] = buffer_data_0[3375:3368] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_422[22] = buffer_data_0[3383:3376] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_422[23] = buffer_data_0[3391:3384] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_422[24] = buffer_data_0[3399:3392] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_422 = kernel_img_mul_422[0] + kernel_img_mul_422[1] + kernel_img_mul_422[2] + 
                kernel_img_mul_422[3] + kernel_img_mul_422[4] + kernel_img_mul_422[5] + 
                kernel_img_mul_422[6] + kernel_img_mul_422[7] + kernel_img_mul_422[8] + 
                kernel_img_mul_422[9] + kernel_img_mul_422[10] + kernel_img_mul_422[11] + 
                kernel_img_mul_422[12] + kernel_img_mul_422[13] + kernel_img_mul_422[14] + 
                kernel_img_mul_422[15] + kernel_img_mul_422[16] + kernel_img_mul_422[17] + 
                kernel_img_mul_422[18] + kernel_img_mul_422[19] + kernel_img_mul_422[20] + 
                kernel_img_mul_422[21] + kernel_img_mul_422[22] + kernel_img_mul_422[23] + 
                kernel_img_mul_422[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3383:3376] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3383:3376] <= kernel_img_sum_422[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3383:3376] <= 'd0;
end

wire  [39:0]  kernel_img_mul_423[0:24];
assign kernel_img_mul_423[0] = buffer_data_4[3375:3368] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_423[1] = buffer_data_4[3383:3376] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_423[2] = buffer_data_4[3391:3384] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_423[3] = buffer_data_4[3399:3392] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_423[4] = buffer_data_4[3407:3400] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_423[5] = buffer_data_3[3375:3368] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_423[6] = buffer_data_3[3383:3376] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_423[7] = buffer_data_3[3391:3384] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_423[8] = buffer_data_3[3399:3392] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_423[9] = buffer_data_3[3407:3400] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_423[10] = buffer_data_2[3375:3368] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_423[11] = buffer_data_2[3383:3376] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_423[12] = buffer_data_2[3391:3384] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_423[13] = buffer_data_2[3399:3392] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_423[14] = buffer_data_2[3407:3400] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_423[15] = buffer_data_1[3375:3368] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_423[16] = buffer_data_1[3383:3376] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_423[17] = buffer_data_1[3391:3384] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_423[18] = buffer_data_1[3399:3392] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_423[19] = buffer_data_1[3407:3400] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_423[20] = buffer_data_0[3375:3368] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_423[21] = buffer_data_0[3383:3376] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_423[22] = buffer_data_0[3391:3384] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_423[23] = buffer_data_0[3399:3392] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_423[24] = buffer_data_0[3407:3400] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_423 = kernel_img_mul_423[0] + kernel_img_mul_423[1] + kernel_img_mul_423[2] + 
                kernel_img_mul_423[3] + kernel_img_mul_423[4] + kernel_img_mul_423[5] + 
                kernel_img_mul_423[6] + kernel_img_mul_423[7] + kernel_img_mul_423[8] + 
                kernel_img_mul_423[9] + kernel_img_mul_423[10] + kernel_img_mul_423[11] + 
                kernel_img_mul_423[12] + kernel_img_mul_423[13] + kernel_img_mul_423[14] + 
                kernel_img_mul_423[15] + kernel_img_mul_423[16] + kernel_img_mul_423[17] + 
                kernel_img_mul_423[18] + kernel_img_mul_423[19] + kernel_img_mul_423[20] + 
                kernel_img_mul_423[21] + kernel_img_mul_423[22] + kernel_img_mul_423[23] + 
                kernel_img_mul_423[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3391:3384] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3391:3384] <= kernel_img_sum_423[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3391:3384] <= 'd0;
end

wire  [39:0]  kernel_img_mul_424[0:24];
assign kernel_img_mul_424[0] = buffer_data_4[3383:3376] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_424[1] = buffer_data_4[3391:3384] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_424[2] = buffer_data_4[3399:3392] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_424[3] = buffer_data_4[3407:3400] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_424[4] = buffer_data_4[3415:3408] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_424[5] = buffer_data_3[3383:3376] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_424[6] = buffer_data_3[3391:3384] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_424[7] = buffer_data_3[3399:3392] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_424[8] = buffer_data_3[3407:3400] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_424[9] = buffer_data_3[3415:3408] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_424[10] = buffer_data_2[3383:3376] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_424[11] = buffer_data_2[3391:3384] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_424[12] = buffer_data_2[3399:3392] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_424[13] = buffer_data_2[3407:3400] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_424[14] = buffer_data_2[3415:3408] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_424[15] = buffer_data_1[3383:3376] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_424[16] = buffer_data_1[3391:3384] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_424[17] = buffer_data_1[3399:3392] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_424[18] = buffer_data_1[3407:3400] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_424[19] = buffer_data_1[3415:3408] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_424[20] = buffer_data_0[3383:3376] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_424[21] = buffer_data_0[3391:3384] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_424[22] = buffer_data_0[3399:3392] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_424[23] = buffer_data_0[3407:3400] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_424[24] = buffer_data_0[3415:3408] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_424 = kernel_img_mul_424[0] + kernel_img_mul_424[1] + kernel_img_mul_424[2] + 
                kernel_img_mul_424[3] + kernel_img_mul_424[4] + kernel_img_mul_424[5] + 
                kernel_img_mul_424[6] + kernel_img_mul_424[7] + kernel_img_mul_424[8] + 
                kernel_img_mul_424[9] + kernel_img_mul_424[10] + kernel_img_mul_424[11] + 
                kernel_img_mul_424[12] + kernel_img_mul_424[13] + kernel_img_mul_424[14] + 
                kernel_img_mul_424[15] + kernel_img_mul_424[16] + kernel_img_mul_424[17] + 
                kernel_img_mul_424[18] + kernel_img_mul_424[19] + kernel_img_mul_424[20] + 
                kernel_img_mul_424[21] + kernel_img_mul_424[22] + kernel_img_mul_424[23] + 
                kernel_img_mul_424[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3399:3392] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3399:3392] <= kernel_img_sum_424[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3399:3392] <= 'd0;
end

wire  [39:0]  kernel_img_mul_425[0:24];
assign kernel_img_mul_425[0] = buffer_data_4[3391:3384] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_425[1] = buffer_data_4[3399:3392] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_425[2] = buffer_data_4[3407:3400] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_425[3] = buffer_data_4[3415:3408] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_425[4] = buffer_data_4[3423:3416] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_425[5] = buffer_data_3[3391:3384] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_425[6] = buffer_data_3[3399:3392] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_425[7] = buffer_data_3[3407:3400] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_425[8] = buffer_data_3[3415:3408] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_425[9] = buffer_data_3[3423:3416] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_425[10] = buffer_data_2[3391:3384] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_425[11] = buffer_data_2[3399:3392] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_425[12] = buffer_data_2[3407:3400] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_425[13] = buffer_data_2[3415:3408] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_425[14] = buffer_data_2[3423:3416] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_425[15] = buffer_data_1[3391:3384] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_425[16] = buffer_data_1[3399:3392] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_425[17] = buffer_data_1[3407:3400] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_425[18] = buffer_data_1[3415:3408] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_425[19] = buffer_data_1[3423:3416] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_425[20] = buffer_data_0[3391:3384] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_425[21] = buffer_data_0[3399:3392] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_425[22] = buffer_data_0[3407:3400] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_425[23] = buffer_data_0[3415:3408] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_425[24] = buffer_data_0[3423:3416] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_425 = kernel_img_mul_425[0] + kernel_img_mul_425[1] + kernel_img_mul_425[2] + 
                kernel_img_mul_425[3] + kernel_img_mul_425[4] + kernel_img_mul_425[5] + 
                kernel_img_mul_425[6] + kernel_img_mul_425[7] + kernel_img_mul_425[8] + 
                kernel_img_mul_425[9] + kernel_img_mul_425[10] + kernel_img_mul_425[11] + 
                kernel_img_mul_425[12] + kernel_img_mul_425[13] + kernel_img_mul_425[14] + 
                kernel_img_mul_425[15] + kernel_img_mul_425[16] + kernel_img_mul_425[17] + 
                kernel_img_mul_425[18] + kernel_img_mul_425[19] + kernel_img_mul_425[20] + 
                kernel_img_mul_425[21] + kernel_img_mul_425[22] + kernel_img_mul_425[23] + 
                kernel_img_mul_425[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3407:3400] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3407:3400] <= kernel_img_sum_425[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3407:3400] <= 'd0;
end

wire  [39:0]  kernel_img_mul_426[0:24];
assign kernel_img_mul_426[0] = buffer_data_4[3399:3392] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_426[1] = buffer_data_4[3407:3400] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_426[2] = buffer_data_4[3415:3408] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_426[3] = buffer_data_4[3423:3416] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_426[4] = buffer_data_4[3431:3424] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_426[5] = buffer_data_3[3399:3392] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_426[6] = buffer_data_3[3407:3400] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_426[7] = buffer_data_3[3415:3408] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_426[8] = buffer_data_3[3423:3416] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_426[9] = buffer_data_3[3431:3424] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_426[10] = buffer_data_2[3399:3392] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_426[11] = buffer_data_2[3407:3400] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_426[12] = buffer_data_2[3415:3408] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_426[13] = buffer_data_2[3423:3416] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_426[14] = buffer_data_2[3431:3424] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_426[15] = buffer_data_1[3399:3392] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_426[16] = buffer_data_1[3407:3400] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_426[17] = buffer_data_1[3415:3408] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_426[18] = buffer_data_1[3423:3416] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_426[19] = buffer_data_1[3431:3424] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_426[20] = buffer_data_0[3399:3392] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_426[21] = buffer_data_0[3407:3400] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_426[22] = buffer_data_0[3415:3408] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_426[23] = buffer_data_0[3423:3416] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_426[24] = buffer_data_0[3431:3424] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_426 = kernel_img_mul_426[0] + kernel_img_mul_426[1] + kernel_img_mul_426[2] + 
                kernel_img_mul_426[3] + kernel_img_mul_426[4] + kernel_img_mul_426[5] + 
                kernel_img_mul_426[6] + kernel_img_mul_426[7] + kernel_img_mul_426[8] + 
                kernel_img_mul_426[9] + kernel_img_mul_426[10] + kernel_img_mul_426[11] + 
                kernel_img_mul_426[12] + kernel_img_mul_426[13] + kernel_img_mul_426[14] + 
                kernel_img_mul_426[15] + kernel_img_mul_426[16] + kernel_img_mul_426[17] + 
                kernel_img_mul_426[18] + kernel_img_mul_426[19] + kernel_img_mul_426[20] + 
                kernel_img_mul_426[21] + kernel_img_mul_426[22] + kernel_img_mul_426[23] + 
                kernel_img_mul_426[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3415:3408] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3415:3408] <= kernel_img_sum_426[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3415:3408] <= 'd0;
end

wire  [39:0]  kernel_img_mul_427[0:24];
assign kernel_img_mul_427[0] = buffer_data_4[3407:3400] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_427[1] = buffer_data_4[3415:3408] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_427[2] = buffer_data_4[3423:3416] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_427[3] = buffer_data_4[3431:3424] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_427[4] = buffer_data_4[3439:3432] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_427[5] = buffer_data_3[3407:3400] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_427[6] = buffer_data_3[3415:3408] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_427[7] = buffer_data_3[3423:3416] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_427[8] = buffer_data_3[3431:3424] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_427[9] = buffer_data_3[3439:3432] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_427[10] = buffer_data_2[3407:3400] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_427[11] = buffer_data_2[3415:3408] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_427[12] = buffer_data_2[3423:3416] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_427[13] = buffer_data_2[3431:3424] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_427[14] = buffer_data_2[3439:3432] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_427[15] = buffer_data_1[3407:3400] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_427[16] = buffer_data_1[3415:3408] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_427[17] = buffer_data_1[3423:3416] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_427[18] = buffer_data_1[3431:3424] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_427[19] = buffer_data_1[3439:3432] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_427[20] = buffer_data_0[3407:3400] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_427[21] = buffer_data_0[3415:3408] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_427[22] = buffer_data_0[3423:3416] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_427[23] = buffer_data_0[3431:3424] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_427[24] = buffer_data_0[3439:3432] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_427 = kernel_img_mul_427[0] + kernel_img_mul_427[1] + kernel_img_mul_427[2] + 
                kernel_img_mul_427[3] + kernel_img_mul_427[4] + kernel_img_mul_427[5] + 
                kernel_img_mul_427[6] + kernel_img_mul_427[7] + kernel_img_mul_427[8] + 
                kernel_img_mul_427[9] + kernel_img_mul_427[10] + kernel_img_mul_427[11] + 
                kernel_img_mul_427[12] + kernel_img_mul_427[13] + kernel_img_mul_427[14] + 
                kernel_img_mul_427[15] + kernel_img_mul_427[16] + kernel_img_mul_427[17] + 
                kernel_img_mul_427[18] + kernel_img_mul_427[19] + kernel_img_mul_427[20] + 
                kernel_img_mul_427[21] + kernel_img_mul_427[22] + kernel_img_mul_427[23] + 
                kernel_img_mul_427[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3423:3416] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3423:3416] <= kernel_img_sum_427[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3423:3416] <= 'd0;
end

wire  [39:0]  kernel_img_mul_428[0:24];
assign kernel_img_mul_428[0] = buffer_data_4[3415:3408] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_428[1] = buffer_data_4[3423:3416] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_428[2] = buffer_data_4[3431:3424] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_428[3] = buffer_data_4[3439:3432] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_428[4] = buffer_data_4[3447:3440] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_428[5] = buffer_data_3[3415:3408] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_428[6] = buffer_data_3[3423:3416] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_428[7] = buffer_data_3[3431:3424] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_428[8] = buffer_data_3[3439:3432] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_428[9] = buffer_data_3[3447:3440] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_428[10] = buffer_data_2[3415:3408] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_428[11] = buffer_data_2[3423:3416] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_428[12] = buffer_data_2[3431:3424] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_428[13] = buffer_data_2[3439:3432] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_428[14] = buffer_data_2[3447:3440] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_428[15] = buffer_data_1[3415:3408] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_428[16] = buffer_data_1[3423:3416] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_428[17] = buffer_data_1[3431:3424] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_428[18] = buffer_data_1[3439:3432] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_428[19] = buffer_data_1[3447:3440] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_428[20] = buffer_data_0[3415:3408] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_428[21] = buffer_data_0[3423:3416] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_428[22] = buffer_data_0[3431:3424] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_428[23] = buffer_data_0[3439:3432] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_428[24] = buffer_data_0[3447:3440] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_428 = kernel_img_mul_428[0] + kernel_img_mul_428[1] + kernel_img_mul_428[2] + 
                kernel_img_mul_428[3] + kernel_img_mul_428[4] + kernel_img_mul_428[5] + 
                kernel_img_mul_428[6] + kernel_img_mul_428[7] + kernel_img_mul_428[8] + 
                kernel_img_mul_428[9] + kernel_img_mul_428[10] + kernel_img_mul_428[11] + 
                kernel_img_mul_428[12] + kernel_img_mul_428[13] + kernel_img_mul_428[14] + 
                kernel_img_mul_428[15] + kernel_img_mul_428[16] + kernel_img_mul_428[17] + 
                kernel_img_mul_428[18] + kernel_img_mul_428[19] + kernel_img_mul_428[20] + 
                kernel_img_mul_428[21] + kernel_img_mul_428[22] + kernel_img_mul_428[23] + 
                kernel_img_mul_428[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3431:3424] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3431:3424] <= kernel_img_sum_428[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3431:3424] <= 'd0;
end

wire  [39:0]  kernel_img_mul_429[0:24];
assign kernel_img_mul_429[0] = buffer_data_4[3423:3416] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_429[1] = buffer_data_4[3431:3424] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_429[2] = buffer_data_4[3439:3432] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_429[3] = buffer_data_4[3447:3440] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_429[4] = buffer_data_4[3455:3448] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_429[5] = buffer_data_3[3423:3416] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_429[6] = buffer_data_3[3431:3424] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_429[7] = buffer_data_3[3439:3432] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_429[8] = buffer_data_3[3447:3440] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_429[9] = buffer_data_3[3455:3448] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_429[10] = buffer_data_2[3423:3416] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_429[11] = buffer_data_2[3431:3424] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_429[12] = buffer_data_2[3439:3432] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_429[13] = buffer_data_2[3447:3440] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_429[14] = buffer_data_2[3455:3448] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_429[15] = buffer_data_1[3423:3416] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_429[16] = buffer_data_1[3431:3424] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_429[17] = buffer_data_1[3439:3432] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_429[18] = buffer_data_1[3447:3440] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_429[19] = buffer_data_1[3455:3448] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_429[20] = buffer_data_0[3423:3416] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_429[21] = buffer_data_0[3431:3424] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_429[22] = buffer_data_0[3439:3432] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_429[23] = buffer_data_0[3447:3440] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_429[24] = buffer_data_0[3455:3448] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_429 = kernel_img_mul_429[0] + kernel_img_mul_429[1] + kernel_img_mul_429[2] + 
                kernel_img_mul_429[3] + kernel_img_mul_429[4] + kernel_img_mul_429[5] + 
                kernel_img_mul_429[6] + kernel_img_mul_429[7] + kernel_img_mul_429[8] + 
                kernel_img_mul_429[9] + kernel_img_mul_429[10] + kernel_img_mul_429[11] + 
                kernel_img_mul_429[12] + kernel_img_mul_429[13] + kernel_img_mul_429[14] + 
                kernel_img_mul_429[15] + kernel_img_mul_429[16] + kernel_img_mul_429[17] + 
                kernel_img_mul_429[18] + kernel_img_mul_429[19] + kernel_img_mul_429[20] + 
                kernel_img_mul_429[21] + kernel_img_mul_429[22] + kernel_img_mul_429[23] + 
                kernel_img_mul_429[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3439:3432] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3439:3432] <= kernel_img_sum_429[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3439:3432] <= 'd0;
end

wire  [39:0]  kernel_img_mul_430[0:24];
assign kernel_img_mul_430[0] = buffer_data_4[3431:3424] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_430[1] = buffer_data_4[3439:3432] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_430[2] = buffer_data_4[3447:3440] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_430[3] = buffer_data_4[3455:3448] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_430[4] = buffer_data_4[3463:3456] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_430[5] = buffer_data_3[3431:3424] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_430[6] = buffer_data_3[3439:3432] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_430[7] = buffer_data_3[3447:3440] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_430[8] = buffer_data_3[3455:3448] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_430[9] = buffer_data_3[3463:3456] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_430[10] = buffer_data_2[3431:3424] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_430[11] = buffer_data_2[3439:3432] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_430[12] = buffer_data_2[3447:3440] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_430[13] = buffer_data_2[3455:3448] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_430[14] = buffer_data_2[3463:3456] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_430[15] = buffer_data_1[3431:3424] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_430[16] = buffer_data_1[3439:3432] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_430[17] = buffer_data_1[3447:3440] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_430[18] = buffer_data_1[3455:3448] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_430[19] = buffer_data_1[3463:3456] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_430[20] = buffer_data_0[3431:3424] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_430[21] = buffer_data_0[3439:3432] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_430[22] = buffer_data_0[3447:3440] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_430[23] = buffer_data_0[3455:3448] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_430[24] = buffer_data_0[3463:3456] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_430 = kernel_img_mul_430[0] + kernel_img_mul_430[1] + kernel_img_mul_430[2] + 
                kernel_img_mul_430[3] + kernel_img_mul_430[4] + kernel_img_mul_430[5] + 
                kernel_img_mul_430[6] + kernel_img_mul_430[7] + kernel_img_mul_430[8] + 
                kernel_img_mul_430[9] + kernel_img_mul_430[10] + kernel_img_mul_430[11] + 
                kernel_img_mul_430[12] + kernel_img_mul_430[13] + kernel_img_mul_430[14] + 
                kernel_img_mul_430[15] + kernel_img_mul_430[16] + kernel_img_mul_430[17] + 
                kernel_img_mul_430[18] + kernel_img_mul_430[19] + kernel_img_mul_430[20] + 
                kernel_img_mul_430[21] + kernel_img_mul_430[22] + kernel_img_mul_430[23] + 
                kernel_img_mul_430[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3447:3440] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3447:3440] <= kernel_img_sum_430[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3447:3440] <= 'd0;
end

wire  [39:0]  kernel_img_mul_431[0:24];
assign kernel_img_mul_431[0] = buffer_data_4[3439:3432] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_431[1] = buffer_data_4[3447:3440] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_431[2] = buffer_data_4[3455:3448] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_431[3] = buffer_data_4[3463:3456] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_431[4] = buffer_data_4[3471:3464] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_431[5] = buffer_data_3[3439:3432] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_431[6] = buffer_data_3[3447:3440] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_431[7] = buffer_data_3[3455:3448] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_431[8] = buffer_data_3[3463:3456] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_431[9] = buffer_data_3[3471:3464] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_431[10] = buffer_data_2[3439:3432] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_431[11] = buffer_data_2[3447:3440] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_431[12] = buffer_data_2[3455:3448] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_431[13] = buffer_data_2[3463:3456] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_431[14] = buffer_data_2[3471:3464] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_431[15] = buffer_data_1[3439:3432] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_431[16] = buffer_data_1[3447:3440] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_431[17] = buffer_data_1[3455:3448] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_431[18] = buffer_data_1[3463:3456] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_431[19] = buffer_data_1[3471:3464] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_431[20] = buffer_data_0[3439:3432] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_431[21] = buffer_data_0[3447:3440] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_431[22] = buffer_data_0[3455:3448] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_431[23] = buffer_data_0[3463:3456] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_431[24] = buffer_data_0[3471:3464] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_431 = kernel_img_mul_431[0] + kernel_img_mul_431[1] + kernel_img_mul_431[2] + 
                kernel_img_mul_431[3] + kernel_img_mul_431[4] + kernel_img_mul_431[5] + 
                kernel_img_mul_431[6] + kernel_img_mul_431[7] + kernel_img_mul_431[8] + 
                kernel_img_mul_431[9] + kernel_img_mul_431[10] + kernel_img_mul_431[11] + 
                kernel_img_mul_431[12] + kernel_img_mul_431[13] + kernel_img_mul_431[14] + 
                kernel_img_mul_431[15] + kernel_img_mul_431[16] + kernel_img_mul_431[17] + 
                kernel_img_mul_431[18] + kernel_img_mul_431[19] + kernel_img_mul_431[20] + 
                kernel_img_mul_431[21] + kernel_img_mul_431[22] + kernel_img_mul_431[23] + 
                kernel_img_mul_431[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3455:3448] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3455:3448] <= kernel_img_sum_431[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3455:3448] <= 'd0;
end

wire  [39:0]  kernel_img_mul_432[0:24];
assign kernel_img_mul_432[0] = buffer_data_4[3447:3440] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_432[1] = buffer_data_4[3455:3448] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_432[2] = buffer_data_4[3463:3456] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_432[3] = buffer_data_4[3471:3464] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_432[4] = buffer_data_4[3479:3472] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_432[5] = buffer_data_3[3447:3440] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_432[6] = buffer_data_3[3455:3448] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_432[7] = buffer_data_3[3463:3456] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_432[8] = buffer_data_3[3471:3464] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_432[9] = buffer_data_3[3479:3472] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_432[10] = buffer_data_2[3447:3440] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_432[11] = buffer_data_2[3455:3448] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_432[12] = buffer_data_2[3463:3456] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_432[13] = buffer_data_2[3471:3464] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_432[14] = buffer_data_2[3479:3472] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_432[15] = buffer_data_1[3447:3440] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_432[16] = buffer_data_1[3455:3448] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_432[17] = buffer_data_1[3463:3456] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_432[18] = buffer_data_1[3471:3464] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_432[19] = buffer_data_1[3479:3472] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_432[20] = buffer_data_0[3447:3440] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_432[21] = buffer_data_0[3455:3448] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_432[22] = buffer_data_0[3463:3456] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_432[23] = buffer_data_0[3471:3464] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_432[24] = buffer_data_0[3479:3472] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_432 = kernel_img_mul_432[0] + kernel_img_mul_432[1] + kernel_img_mul_432[2] + 
                kernel_img_mul_432[3] + kernel_img_mul_432[4] + kernel_img_mul_432[5] + 
                kernel_img_mul_432[6] + kernel_img_mul_432[7] + kernel_img_mul_432[8] + 
                kernel_img_mul_432[9] + kernel_img_mul_432[10] + kernel_img_mul_432[11] + 
                kernel_img_mul_432[12] + kernel_img_mul_432[13] + kernel_img_mul_432[14] + 
                kernel_img_mul_432[15] + kernel_img_mul_432[16] + kernel_img_mul_432[17] + 
                kernel_img_mul_432[18] + kernel_img_mul_432[19] + kernel_img_mul_432[20] + 
                kernel_img_mul_432[21] + kernel_img_mul_432[22] + kernel_img_mul_432[23] + 
                kernel_img_mul_432[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3463:3456] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3463:3456] <= kernel_img_sum_432[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3463:3456] <= 'd0;
end

wire  [39:0]  kernel_img_mul_433[0:24];
assign kernel_img_mul_433[0] = buffer_data_4[3455:3448] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_433[1] = buffer_data_4[3463:3456] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_433[2] = buffer_data_4[3471:3464] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_433[3] = buffer_data_4[3479:3472] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_433[4] = buffer_data_4[3487:3480] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_433[5] = buffer_data_3[3455:3448] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_433[6] = buffer_data_3[3463:3456] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_433[7] = buffer_data_3[3471:3464] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_433[8] = buffer_data_3[3479:3472] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_433[9] = buffer_data_3[3487:3480] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_433[10] = buffer_data_2[3455:3448] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_433[11] = buffer_data_2[3463:3456] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_433[12] = buffer_data_2[3471:3464] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_433[13] = buffer_data_2[3479:3472] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_433[14] = buffer_data_2[3487:3480] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_433[15] = buffer_data_1[3455:3448] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_433[16] = buffer_data_1[3463:3456] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_433[17] = buffer_data_1[3471:3464] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_433[18] = buffer_data_1[3479:3472] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_433[19] = buffer_data_1[3487:3480] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_433[20] = buffer_data_0[3455:3448] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_433[21] = buffer_data_0[3463:3456] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_433[22] = buffer_data_0[3471:3464] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_433[23] = buffer_data_0[3479:3472] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_433[24] = buffer_data_0[3487:3480] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_433 = kernel_img_mul_433[0] + kernel_img_mul_433[1] + kernel_img_mul_433[2] + 
                kernel_img_mul_433[3] + kernel_img_mul_433[4] + kernel_img_mul_433[5] + 
                kernel_img_mul_433[6] + kernel_img_mul_433[7] + kernel_img_mul_433[8] + 
                kernel_img_mul_433[9] + kernel_img_mul_433[10] + kernel_img_mul_433[11] + 
                kernel_img_mul_433[12] + kernel_img_mul_433[13] + kernel_img_mul_433[14] + 
                kernel_img_mul_433[15] + kernel_img_mul_433[16] + kernel_img_mul_433[17] + 
                kernel_img_mul_433[18] + kernel_img_mul_433[19] + kernel_img_mul_433[20] + 
                kernel_img_mul_433[21] + kernel_img_mul_433[22] + kernel_img_mul_433[23] + 
                kernel_img_mul_433[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3471:3464] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3471:3464] <= kernel_img_sum_433[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3471:3464] <= 'd0;
end

wire  [39:0]  kernel_img_mul_434[0:24];
assign kernel_img_mul_434[0] = buffer_data_4[3463:3456] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_434[1] = buffer_data_4[3471:3464] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_434[2] = buffer_data_4[3479:3472] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_434[3] = buffer_data_4[3487:3480] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_434[4] = buffer_data_4[3495:3488] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_434[5] = buffer_data_3[3463:3456] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_434[6] = buffer_data_3[3471:3464] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_434[7] = buffer_data_3[3479:3472] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_434[8] = buffer_data_3[3487:3480] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_434[9] = buffer_data_3[3495:3488] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_434[10] = buffer_data_2[3463:3456] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_434[11] = buffer_data_2[3471:3464] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_434[12] = buffer_data_2[3479:3472] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_434[13] = buffer_data_2[3487:3480] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_434[14] = buffer_data_2[3495:3488] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_434[15] = buffer_data_1[3463:3456] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_434[16] = buffer_data_1[3471:3464] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_434[17] = buffer_data_1[3479:3472] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_434[18] = buffer_data_1[3487:3480] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_434[19] = buffer_data_1[3495:3488] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_434[20] = buffer_data_0[3463:3456] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_434[21] = buffer_data_0[3471:3464] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_434[22] = buffer_data_0[3479:3472] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_434[23] = buffer_data_0[3487:3480] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_434[24] = buffer_data_0[3495:3488] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_434 = kernel_img_mul_434[0] + kernel_img_mul_434[1] + kernel_img_mul_434[2] + 
                kernel_img_mul_434[3] + kernel_img_mul_434[4] + kernel_img_mul_434[5] + 
                kernel_img_mul_434[6] + kernel_img_mul_434[7] + kernel_img_mul_434[8] + 
                kernel_img_mul_434[9] + kernel_img_mul_434[10] + kernel_img_mul_434[11] + 
                kernel_img_mul_434[12] + kernel_img_mul_434[13] + kernel_img_mul_434[14] + 
                kernel_img_mul_434[15] + kernel_img_mul_434[16] + kernel_img_mul_434[17] + 
                kernel_img_mul_434[18] + kernel_img_mul_434[19] + kernel_img_mul_434[20] + 
                kernel_img_mul_434[21] + kernel_img_mul_434[22] + kernel_img_mul_434[23] + 
                kernel_img_mul_434[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3479:3472] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3479:3472] <= kernel_img_sum_434[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3479:3472] <= 'd0;
end

wire  [39:0]  kernel_img_mul_435[0:24];
assign kernel_img_mul_435[0] = buffer_data_4[3471:3464] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_435[1] = buffer_data_4[3479:3472] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_435[2] = buffer_data_4[3487:3480] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_435[3] = buffer_data_4[3495:3488] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_435[4] = buffer_data_4[3503:3496] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_435[5] = buffer_data_3[3471:3464] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_435[6] = buffer_data_3[3479:3472] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_435[7] = buffer_data_3[3487:3480] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_435[8] = buffer_data_3[3495:3488] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_435[9] = buffer_data_3[3503:3496] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_435[10] = buffer_data_2[3471:3464] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_435[11] = buffer_data_2[3479:3472] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_435[12] = buffer_data_2[3487:3480] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_435[13] = buffer_data_2[3495:3488] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_435[14] = buffer_data_2[3503:3496] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_435[15] = buffer_data_1[3471:3464] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_435[16] = buffer_data_1[3479:3472] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_435[17] = buffer_data_1[3487:3480] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_435[18] = buffer_data_1[3495:3488] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_435[19] = buffer_data_1[3503:3496] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_435[20] = buffer_data_0[3471:3464] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_435[21] = buffer_data_0[3479:3472] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_435[22] = buffer_data_0[3487:3480] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_435[23] = buffer_data_0[3495:3488] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_435[24] = buffer_data_0[3503:3496] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_435 = kernel_img_mul_435[0] + kernel_img_mul_435[1] + kernel_img_mul_435[2] + 
                kernel_img_mul_435[3] + kernel_img_mul_435[4] + kernel_img_mul_435[5] + 
                kernel_img_mul_435[6] + kernel_img_mul_435[7] + kernel_img_mul_435[8] + 
                kernel_img_mul_435[9] + kernel_img_mul_435[10] + kernel_img_mul_435[11] + 
                kernel_img_mul_435[12] + kernel_img_mul_435[13] + kernel_img_mul_435[14] + 
                kernel_img_mul_435[15] + kernel_img_mul_435[16] + kernel_img_mul_435[17] + 
                kernel_img_mul_435[18] + kernel_img_mul_435[19] + kernel_img_mul_435[20] + 
                kernel_img_mul_435[21] + kernel_img_mul_435[22] + kernel_img_mul_435[23] + 
                kernel_img_mul_435[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3487:3480] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3487:3480] <= kernel_img_sum_435[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3487:3480] <= 'd0;
end

wire  [39:0]  kernel_img_mul_436[0:24];
assign kernel_img_mul_436[0] = buffer_data_4[3479:3472] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_436[1] = buffer_data_4[3487:3480] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_436[2] = buffer_data_4[3495:3488] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_436[3] = buffer_data_4[3503:3496] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_436[4] = buffer_data_4[3511:3504] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_436[5] = buffer_data_3[3479:3472] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_436[6] = buffer_data_3[3487:3480] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_436[7] = buffer_data_3[3495:3488] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_436[8] = buffer_data_3[3503:3496] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_436[9] = buffer_data_3[3511:3504] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_436[10] = buffer_data_2[3479:3472] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_436[11] = buffer_data_2[3487:3480] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_436[12] = buffer_data_2[3495:3488] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_436[13] = buffer_data_2[3503:3496] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_436[14] = buffer_data_2[3511:3504] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_436[15] = buffer_data_1[3479:3472] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_436[16] = buffer_data_1[3487:3480] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_436[17] = buffer_data_1[3495:3488] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_436[18] = buffer_data_1[3503:3496] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_436[19] = buffer_data_1[3511:3504] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_436[20] = buffer_data_0[3479:3472] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_436[21] = buffer_data_0[3487:3480] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_436[22] = buffer_data_0[3495:3488] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_436[23] = buffer_data_0[3503:3496] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_436[24] = buffer_data_0[3511:3504] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_436 = kernel_img_mul_436[0] + kernel_img_mul_436[1] + kernel_img_mul_436[2] + 
                kernel_img_mul_436[3] + kernel_img_mul_436[4] + kernel_img_mul_436[5] + 
                kernel_img_mul_436[6] + kernel_img_mul_436[7] + kernel_img_mul_436[8] + 
                kernel_img_mul_436[9] + kernel_img_mul_436[10] + kernel_img_mul_436[11] + 
                kernel_img_mul_436[12] + kernel_img_mul_436[13] + kernel_img_mul_436[14] + 
                kernel_img_mul_436[15] + kernel_img_mul_436[16] + kernel_img_mul_436[17] + 
                kernel_img_mul_436[18] + kernel_img_mul_436[19] + kernel_img_mul_436[20] + 
                kernel_img_mul_436[21] + kernel_img_mul_436[22] + kernel_img_mul_436[23] + 
                kernel_img_mul_436[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3495:3488] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3495:3488] <= kernel_img_sum_436[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3495:3488] <= 'd0;
end

wire  [39:0]  kernel_img_mul_437[0:24];
assign kernel_img_mul_437[0] = buffer_data_4[3487:3480] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_437[1] = buffer_data_4[3495:3488] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_437[2] = buffer_data_4[3503:3496] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_437[3] = buffer_data_4[3511:3504] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_437[4] = buffer_data_4[3519:3512] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_437[5] = buffer_data_3[3487:3480] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_437[6] = buffer_data_3[3495:3488] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_437[7] = buffer_data_3[3503:3496] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_437[8] = buffer_data_3[3511:3504] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_437[9] = buffer_data_3[3519:3512] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_437[10] = buffer_data_2[3487:3480] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_437[11] = buffer_data_2[3495:3488] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_437[12] = buffer_data_2[3503:3496] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_437[13] = buffer_data_2[3511:3504] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_437[14] = buffer_data_2[3519:3512] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_437[15] = buffer_data_1[3487:3480] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_437[16] = buffer_data_1[3495:3488] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_437[17] = buffer_data_1[3503:3496] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_437[18] = buffer_data_1[3511:3504] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_437[19] = buffer_data_1[3519:3512] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_437[20] = buffer_data_0[3487:3480] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_437[21] = buffer_data_0[3495:3488] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_437[22] = buffer_data_0[3503:3496] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_437[23] = buffer_data_0[3511:3504] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_437[24] = buffer_data_0[3519:3512] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_437 = kernel_img_mul_437[0] + kernel_img_mul_437[1] + kernel_img_mul_437[2] + 
                kernel_img_mul_437[3] + kernel_img_mul_437[4] + kernel_img_mul_437[5] + 
                kernel_img_mul_437[6] + kernel_img_mul_437[7] + kernel_img_mul_437[8] + 
                kernel_img_mul_437[9] + kernel_img_mul_437[10] + kernel_img_mul_437[11] + 
                kernel_img_mul_437[12] + kernel_img_mul_437[13] + kernel_img_mul_437[14] + 
                kernel_img_mul_437[15] + kernel_img_mul_437[16] + kernel_img_mul_437[17] + 
                kernel_img_mul_437[18] + kernel_img_mul_437[19] + kernel_img_mul_437[20] + 
                kernel_img_mul_437[21] + kernel_img_mul_437[22] + kernel_img_mul_437[23] + 
                kernel_img_mul_437[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3503:3496] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3503:3496] <= kernel_img_sum_437[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3503:3496] <= 'd0;
end

wire  [39:0]  kernel_img_mul_438[0:24];
assign kernel_img_mul_438[0] = buffer_data_4[3495:3488] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_438[1] = buffer_data_4[3503:3496] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_438[2] = buffer_data_4[3511:3504] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_438[3] = buffer_data_4[3519:3512] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_438[4] = buffer_data_4[3527:3520] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_438[5] = buffer_data_3[3495:3488] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_438[6] = buffer_data_3[3503:3496] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_438[7] = buffer_data_3[3511:3504] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_438[8] = buffer_data_3[3519:3512] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_438[9] = buffer_data_3[3527:3520] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_438[10] = buffer_data_2[3495:3488] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_438[11] = buffer_data_2[3503:3496] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_438[12] = buffer_data_2[3511:3504] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_438[13] = buffer_data_2[3519:3512] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_438[14] = buffer_data_2[3527:3520] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_438[15] = buffer_data_1[3495:3488] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_438[16] = buffer_data_1[3503:3496] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_438[17] = buffer_data_1[3511:3504] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_438[18] = buffer_data_1[3519:3512] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_438[19] = buffer_data_1[3527:3520] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_438[20] = buffer_data_0[3495:3488] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_438[21] = buffer_data_0[3503:3496] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_438[22] = buffer_data_0[3511:3504] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_438[23] = buffer_data_0[3519:3512] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_438[24] = buffer_data_0[3527:3520] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_438 = kernel_img_mul_438[0] + kernel_img_mul_438[1] + kernel_img_mul_438[2] + 
                kernel_img_mul_438[3] + kernel_img_mul_438[4] + kernel_img_mul_438[5] + 
                kernel_img_mul_438[6] + kernel_img_mul_438[7] + kernel_img_mul_438[8] + 
                kernel_img_mul_438[9] + kernel_img_mul_438[10] + kernel_img_mul_438[11] + 
                kernel_img_mul_438[12] + kernel_img_mul_438[13] + kernel_img_mul_438[14] + 
                kernel_img_mul_438[15] + kernel_img_mul_438[16] + kernel_img_mul_438[17] + 
                kernel_img_mul_438[18] + kernel_img_mul_438[19] + kernel_img_mul_438[20] + 
                kernel_img_mul_438[21] + kernel_img_mul_438[22] + kernel_img_mul_438[23] + 
                kernel_img_mul_438[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3511:3504] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3511:3504] <= kernel_img_sum_438[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3511:3504] <= 'd0;
end

wire  [39:0]  kernel_img_mul_439[0:24];
assign kernel_img_mul_439[0] = buffer_data_4[3503:3496] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_439[1] = buffer_data_4[3511:3504] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_439[2] = buffer_data_4[3519:3512] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_439[3] = buffer_data_4[3527:3520] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_439[4] = buffer_data_4[3535:3528] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_439[5] = buffer_data_3[3503:3496] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_439[6] = buffer_data_3[3511:3504] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_439[7] = buffer_data_3[3519:3512] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_439[8] = buffer_data_3[3527:3520] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_439[9] = buffer_data_3[3535:3528] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_439[10] = buffer_data_2[3503:3496] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_439[11] = buffer_data_2[3511:3504] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_439[12] = buffer_data_2[3519:3512] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_439[13] = buffer_data_2[3527:3520] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_439[14] = buffer_data_2[3535:3528] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_439[15] = buffer_data_1[3503:3496] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_439[16] = buffer_data_1[3511:3504] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_439[17] = buffer_data_1[3519:3512] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_439[18] = buffer_data_1[3527:3520] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_439[19] = buffer_data_1[3535:3528] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_439[20] = buffer_data_0[3503:3496] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_439[21] = buffer_data_0[3511:3504] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_439[22] = buffer_data_0[3519:3512] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_439[23] = buffer_data_0[3527:3520] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_439[24] = buffer_data_0[3535:3528] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_439 = kernel_img_mul_439[0] + kernel_img_mul_439[1] + kernel_img_mul_439[2] + 
                kernel_img_mul_439[3] + kernel_img_mul_439[4] + kernel_img_mul_439[5] + 
                kernel_img_mul_439[6] + kernel_img_mul_439[7] + kernel_img_mul_439[8] + 
                kernel_img_mul_439[9] + kernel_img_mul_439[10] + kernel_img_mul_439[11] + 
                kernel_img_mul_439[12] + kernel_img_mul_439[13] + kernel_img_mul_439[14] + 
                kernel_img_mul_439[15] + kernel_img_mul_439[16] + kernel_img_mul_439[17] + 
                kernel_img_mul_439[18] + kernel_img_mul_439[19] + kernel_img_mul_439[20] + 
                kernel_img_mul_439[21] + kernel_img_mul_439[22] + kernel_img_mul_439[23] + 
                kernel_img_mul_439[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3519:3512] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3519:3512] <= kernel_img_sum_439[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3519:3512] <= 'd0;
end

wire  [39:0]  kernel_img_mul_440[0:24];
assign kernel_img_mul_440[0] = buffer_data_4[3511:3504] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_440[1] = buffer_data_4[3519:3512] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_440[2] = buffer_data_4[3527:3520] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_440[3] = buffer_data_4[3535:3528] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_440[4] = buffer_data_4[3543:3536] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_440[5] = buffer_data_3[3511:3504] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_440[6] = buffer_data_3[3519:3512] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_440[7] = buffer_data_3[3527:3520] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_440[8] = buffer_data_3[3535:3528] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_440[9] = buffer_data_3[3543:3536] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_440[10] = buffer_data_2[3511:3504] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_440[11] = buffer_data_2[3519:3512] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_440[12] = buffer_data_2[3527:3520] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_440[13] = buffer_data_2[3535:3528] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_440[14] = buffer_data_2[3543:3536] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_440[15] = buffer_data_1[3511:3504] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_440[16] = buffer_data_1[3519:3512] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_440[17] = buffer_data_1[3527:3520] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_440[18] = buffer_data_1[3535:3528] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_440[19] = buffer_data_1[3543:3536] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_440[20] = buffer_data_0[3511:3504] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_440[21] = buffer_data_0[3519:3512] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_440[22] = buffer_data_0[3527:3520] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_440[23] = buffer_data_0[3535:3528] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_440[24] = buffer_data_0[3543:3536] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_440 = kernel_img_mul_440[0] + kernel_img_mul_440[1] + kernel_img_mul_440[2] + 
                kernel_img_mul_440[3] + kernel_img_mul_440[4] + kernel_img_mul_440[5] + 
                kernel_img_mul_440[6] + kernel_img_mul_440[7] + kernel_img_mul_440[8] + 
                kernel_img_mul_440[9] + kernel_img_mul_440[10] + kernel_img_mul_440[11] + 
                kernel_img_mul_440[12] + kernel_img_mul_440[13] + kernel_img_mul_440[14] + 
                kernel_img_mul_440[15] + kernel_img_mul_440[16] + kernel_img_mul_440[17] + 
                kernel_img_mul_440[18] + kernel_img_mul_440[19] + kernel_img_mul_440[20] + 
                kernel_img_mul_440[21] + kernel_img_mul_440[22] + kernel_img_mul_440[23] + 
                kernel_img_mul_440[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3527:3520] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3527:3520] <= kernel_img_sum_440[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3527:3520] <= 'd0;
end

wire  [39:0]  kernel_img_mul_441[0:24];
assign kernel_img_mul_441[0] = buffer_data_4[3519:3512] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_441[1] = buffer_data_4[3527:3520] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_441[2] = buffer_data_4[3535:3528] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_441[3] = buffer_data_4[3543:3536] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_441[4] = buffer_data_4[3551:3544] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_441[5] = buffer_data_3[3519:3512] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_441[6] = buffer_data_3[3527:3520] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_441[7] = buffer_data_3[3535:3528] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_441[8] = buffer_data_3[3543:3536] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_441[9] = buffer_data_3[3551:3544] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_441[10] = buffer_data_2[3519:3512] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_441[11] = buffer_data_2[3527:3520] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_441[12] = buffer_data_2[3535:3528] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_441[13] = buffer_data_2[3543:3536] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_441[14] = buffer_data_2[3551:3544] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_441[15] = buffer_data_1[3519:3512] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_441[16] = buffer_data_1[3527:3520] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_441[17] = buffer_data_1[3535:3528] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_441[18] = buffer_data_1[3543:3536] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_441[19] = buffer_data_1[3551:3544] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_441[20] = buffer_data_0[3519:3512] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_441[21] = buffer_data_0[3527:3520] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_441[22] = buffer_data_0[3535:3528] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_441[23] = buffer_data_0[3543:3536] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_441[24] = buffer_data_0[3551:3544] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_441 = kernel_img_mul_441[0] + kernel_img_mul_441[1] + kernel_img_mul_441[2] + 
                kernel_img_mul_441[3] + kernel_img_mul_441[4] + kernel_img_mul_441[5] + 
                kernel_img_mul_441[6] + kernel_img_mul_441[7] + kernel_img_mul_441[8] + 
                kernel_img_mul_441[9] + kernel_img_mul_441[10] + kernel_img_mul_441[11] + 
                kernel_img_mul_441[12] + kernel_img_mul_441[13] + kernel_img_mul_441[14] + 
                kernel_img_mul_441[15] + kernel_img_mul_441[16] + kernel_img_mul_441[17] + 
                kernel_img_mul_441[18] + kernel_img_mul_441[19] + kernel_img_mul_441[20] + 
                kernel_img_mul_441[21] + kernel_img_mul_441[22] + kernel_img_mul_441[23] + 
                kernel_img_mul_441[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3535:3528] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3535:3528] <= kernel_img_sum_441[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3535:3528] <= 'd0;
end

wire  [39:0]  kernel_img_mul_442[0:24];
assign kernel_img_mul_442[0] = buffer_data_4[3527:3520] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_442[1] = buffer_data_4[3535:3528] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_442[2] = buffer_data_4[3543:3536] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_442[3] = buffer_data_4[3551:3544] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_442[4] = buffer_data_4[3559:3552] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_442[5] = buffer_data_3[3527:3520] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_442[6] = buffer_data_3[3535:3528] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_442[7] = buffer_data_3[3543:3536] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_442[8] = buffer_data_3[3551:3544] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_442[9] = buffer_data_3[3559:3552] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_442[10] = buffer_data_2[3527:3520] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_442[11] = buffer_data_2[3535:3528] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_442[12] = buffer_data_2[3543:3536] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_442[13] = buffer_data_2[3551:3544] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_442[14] = buffer_data_2[3559:3552] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_442[15] = buffer_data_1[3527:3520] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_442[16] = buffer_data_1[3535:3528] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_442[17] = buffer_data_1[3543:3536] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_442[18] = buffer_data_1[3551:3544] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_442[19] = buffer_data_1[3559:3552] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_442[20] = buffer_data_0[3527:3520] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_442[21] = buffer_data_0[3535:3528] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_442[22] = buffer_data_0[3543:3536] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_442[23] = buffer_data_0[3551:3544] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_442[24] = buffer_data_0[3559:3552] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_442 = kernel_img_mul_442[0] + kernel_img_mul_442[1] + kernel_img_mul_442[2] + 
                kernel_img_mul_442[3] + kernel_img_mul_442[4] + kernel_img_mul_442[5] + 
                kernel_img_mul_442[6] + kernel_img_mul_442[7] + kernel_img_mul_442[8] + 
                kernel_img_mul_442[9] + kernel_img_mul_442[10] + kernel_img_mul_442[11] + 
                kernel_img_mul_442[12] + kernel_img_mul_442[13] + kernel_img_mul_442[14] + 
                kernel_img_mul_442[15] + kernel_img_mul_442[16] + kernel_img_mul_442[17] + 
                kernel_img_mul_442[18] + kernel_img_mul_442[19] + kernel_img_mul_442[20] + 
                kernel_img_mul_442[21] + kernel_img_mul_442[22] + kernel_img_mul_442[23] + 
                kernel_img_mul_442[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3543:3536] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3543:3536] <= kernel_img_sum_442[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3543:3536] <= 'd0;
end

wire  [39:0]  kernel_img_mul_443[0:24];
assign kernel_img_mul_443[0] = buffer_data_4[3535:3528] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_443[1] = buffer_data_4[3543:3536] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_443[2] = buffer_data_4[3551:3544] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_443[3] = buffer_data_4[3559:3552] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_443[4] = buffer_data_4[3567:3560] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_443[5] = buffer_data_3[3535:3528] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_443[6] = buffer_data_3[3543:3536] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_443[7] = buffer_data_3[3551:3544] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_443[8] = buffer_data_3[3559:3552] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_443[9] = buffer_data_3[3567:3560] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_443[10] = buffer_data_2[3535:3528] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_443[11] = buffer_data_2[3543:3536] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_443[12] = buffer_data_2[3551:3544] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_443[13] = buffer_data_2[3559:3552] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_443[14] = buffer_data_2[3567:3560] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_443[15] = buffer_data_1[3535:3528] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_443[16] = buffer_data_1[3543:3536] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_443[17] = buffer_data_1[3551:3544] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_443[18] = buffer_data_1[3559:3552] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_443[19] = buffer_data_1[3567:3560] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_443[20] = buffer_data_0[3535:3528] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_443[21] = buffer_data_0[3543:3536] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_443[22] = buffer_data_0[3551:3544] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_443[23] = buffer_data_0[3559:3552] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_443[24] = buffer_data_0[3567:3560] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_443 = kernel_img_mul_443[0] + kernel_img_mul_443[1] + kernel_img_mul_443[2] + 
                kernel_img_mul_443[3] + kernel_img_mul_443[4] + kernel_img_mul_443[5] + 
                kernel_img_mul_443[6] + kernel_img_mul_443[7] + kernel_img_mul_443[8] + 
                kernel_img_mul_443[9] + kernel_img_mul_443[10] + kernel_img_mul_443[11] + 
                kernel_img_mul_443[12] + kernel_img_mul_443[13] + kernel_img_mul_443[14] + 
                kernel_img_mul_443[15] + kernel_img_mul_443[16] + kernel_img_mul_443[17] + 
                kernel_img_mul_443[18] + kernel_img_mul_443[19] + kernel_img_mul_443[20] + 
                kernel_img_mul_443[21] + kernel_img_mul_443[22] + kernel_img_mul_443[23] + 
                kernel_img_mul_443[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3551:3544] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3551:3544] <= kernel_img_sum_443[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3551:3544] <= 'd0;
end

wire  [39:0]  kernel_img_mul_444[0:24];
assign kernel_img_mul_444[0] = buffer_data_4[3543:3536] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_444[1] = buffer_data_4[3551:3544] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_444[2] = buffer_data_4[3559:3552] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_444[3] = buffer_data_4[3567:3560] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_444[4] = buffer_data_4[3575:3568] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_444[5] = buffer_data_3[3543:3536] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_444[6] = buffer_data_3[3551:3544] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_444[7] = buffer_data_3[3559:3552] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_444[8] = buffer_data_3[3567:3560] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_444[9] = buffer_data_3[3575:3568] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_444[10] = buffer_data_2[3543:3536] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_444[11] = buffer_data_2[3551:3544] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_444[12] = buffer_data_2[3559:3552] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_444[13] = buffer_data_2[3567:3560] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_444[14] = buffer_data_2[3575:3568] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_444[15] = buffer_data_1[3543:3536] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_444[16] = buffer_data_1[3551:3544] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_444[17] = buffer_data_1[3559:3552] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_444[18] = buffer_data_1[3567:3560] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_444[19] = buffer_data_1[3575:3568] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_444[20] = buffer_data_0[3543:3536] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_444[21] = buffer_data_0[3551:3544] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_444[22] = buffer_data_0[3559:3552] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_444[23] = buffer_data_0[3567:3560] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_444[24] = buffer_data_0[3575:3568] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_444 = kernel_img_mul_444[0] + kernel_img_mul_444[1] + kernel_img_mul_444[2] + 
                kernel_img_mul_444[3] + kernel_img_mul_444[4] + kernel_img_mul_444[5] + 
                kernel_img_mul_444[6] + kernel_img_mul_444[7] + kernel_img_mul_444[8] + 
                kernel_img_mul_444[9] + kernel_img_mul_444[10] + kernel_img_mul_444[11] + 
                kernel_img_mul_444[12] + kernel_img_mul_444[13] + kernel_img_mul_444[14] + 
                kernel_img_mul_444[15] + kernel_img_mul_444[16] + kernel_img_mul_444[17] + 
                kernel_img_mul_444[18] + kernel_img_mul_444[19] + kernel_img_mul_444[20] + 
                kernel_img_mul_444[21] + kernel_img_mul_444[22] + kernel_img_mul_444[23] + 
                kernel_img_mul_444[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3559:3552] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3559:3552] <= kernel_img_sum_444[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3559:3552] <= 'd0;
end

wire  [39:0]  kernel_img_mul_445[0:24];
assign kernel_img_mul_445[0] = buffer_data_4[3551:3544] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_445[1] = buffer_data_4[3559:3552] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_445[2] = buffer_data_4[3567:3560] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_445[3] = buffer_data_4[3575:3568] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_445[4] = buffer_data_4[3583:3576] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_445[5] = buffer_data_3[3551:3544] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_445[6] = buffer_data_3[3559:3552] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_445[7] = buffer_data_3[3567:3560] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_445[8] = buffer_data_3[3575:3568] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_445[9] = buffer_data_3[3583:3576] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_445[10] = buffer_data_2[3551:3544] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_445[11] = buffer_data_2[3559:3552] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_445[12] = buffer_data_2[3567:3560] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_445[13] = buffer_data_2[3575:3568] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_445[14] = buffer_data_2[3583:3576] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_445[15] = buffer_data_1[3551:3544] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_445[16] = buffer_data_1[3559:3552] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_445[17] = buffer_data_1[3567:3560] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_445[18] = buffer_data_1[3575:3568] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_445[19] = buffer_data_1[3583:3576] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_445[20] = buffer_data_0[3551:3544] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_445[21] = buffer_data_0[3559:3552] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_445[22] = buffer_data_0[3567:3560] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_445[23] = buffer_data_0[3575:3568] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_445[24] = buffer_data_0[3583:3576] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_445 = kernel_img_mul_445[0] + kernel_img_mul_445[1] + kernel_img_mul_445[2] + 
                kernel_img_mul_445[3] + kernel_img_mul_445[4] + kernel_img_mul_445[5] + 
                kernel_img_mul_445[6] + kernel_img_mul_445[7] + kernel_img_mul_445[8] + 
                kernel_img_mul_445[9] + kernel_img_mul_445[10] + kernel_img_mul_445[11] + 
                kernel_img_mul_445[12] + kernel_img_mul_445[13] + kernel_img_mul_445[14] + 
                kernel_img_mul_445[15] + kernel_img_mul_445[16] + kernel_img_mul_445[17] + 
                kernel_img_mul_445[18] + kernel_img_mul_445[19] + kernel_img_mul_445[20] + 
                kernel_img_mul_445[21] + kernel_img_mul_445[22] + kernel_img_mul_445[23] + 
                kernel_img_mul_445[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3567:3560] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3567:3560] <= kernel_img_sum_445[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3567:3560] <= 'd0;
end

wire  [39:0]  kernel_img_mul_446[0:24];
assign kernel_img_mul_446[0] = buffer_data_4[3559:3552] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_446[1] = buffer_data_4[3567:3560] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_446[2] = buffer_data_4[3575:3568] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_446[3] = buffer_data_4[3583:3576] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_446[4] = buffer_data_4[3591:3584] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_446[5] = buffer_data_3[3559:3552] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_446[6] = buffer_data_3[3567:3560] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_446[7] = buffer_data_3[3575:3568] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_446[8] = buffer_data_3[3583:3576] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_446[9] = buffer_data_3[3591:3584] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_446[10] = buffer_data_2[3559:3552] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_446[11] = buffer_data_2[3567:3560] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_446[12] = buffer_data_2[3575:3568] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_446[13] = buffer_data_2[3583:3576] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_446[14] = buffer_data_2[3591:3584] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_446[15] = buffer_data_1[3559:3552] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_446[16] = buffer_data_1[3567:3560] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_446[17] = buffer_data_1[3575:3568] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_446[18] = buffer_data_1[3583:3576] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_446[19] = buffer_data_1[3591:3584] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_446[20] = buffer_data_0[3559:3552] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_446[21] = buffer_data_0[3567:3560] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_446[22] = buffer_data_0[3575:3568] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_446[23] = buffer_data_0[3583:3576] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_446[24] = buffer_data_0[3591:3584] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_446 = kernel_img_mul_446[0] + kernel_img_mul_446[1] + kernel_img_mul_446[2] + 
                kernel_img_mul_446[3] + kernel_img_mul_446[4] + kernel_img_mul_446[5] + 
                kernel_img_mul_446[6] + kernel_img_mul_446[7] + kernel_img_mul_446[8] + 
                kernel_img_mul_446[9] + kernel_img_mul_446[10] + kernel_img_mul_446[11] + 
                kernel_img_mul_446[12] + kernel_img_mul_446[13] + kernel_img_mul_446[14] + 
                kernel_img_mul_446[15] + kernel_img_mul_446[16] + kernel_img_mul_446[17] + 
                kernel_img_mul_446[18] + kernel_img_mul_446[19] + kernel_img_mul_446[20] + 
                kernel_img_mul_446[21] + kernel_img_mul_446[22] + kernel_img_mul_446[23] + 
                kernel_img_mul_446[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3575:3568] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3575:3568] <= kernel_img_sum_446[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3575:3568] <= 'd0;
end

wire  [39:0]  kernel_img_mul_447[0:24];
assign kernel_img_mul_447[0] = buffer_data_4[3567:3560] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_447[1] = buffer_data_4[3575:3568] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_447[2] = buffer_data_4[3583:3576] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_447[3] = buffer_data_4[3591:3584] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_447[4] = buffer_data_4[3599:3592] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_447[5] = buffer_data_3[3567:3560] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_447[6] = buffer_data_3[3575:3568] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_447[7] = buffer_data_3[3583:3576] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_447[8] = buffer_data_3[3591:3584] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_447[9] = buffer_data_3[3599:3592] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_447[10] = buffer_data_2[3567:3560] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_447[11] = buffer_data_2[3575:3568] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_447[12] = buffer_data_2[3583:3576] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_447[13] = buffer_data_2[3591:3584] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_447[14] = buffer_data_2[3599:3592] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_447[15] = buffer_data_1[3567:3560] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_447[16] = buffer_data_1[3575:3568] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_447[17] = buffer_data_1[3583:3576] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_447[18] = buffer_data_1[3591:3584] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_447[19] = buffer_data_1[3599:3592] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_447[20] = buffer_data_0[3567:3560] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_447[21] = buffer_data_0[3575:3568] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_447[22] = buffer_data_0[3583:3576] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_447[23] = buffer_data_0[3591:3584] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_447[24] = buffer_data_0[3599:3592] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_447 = kernel_img_mul_447[0] + kernel_img_mul_447[1] + kernel_img_mul_447[2] + 
                kernel_img_mul_447[3] + kernel_img_mul_447[4] + kernel_img_mul_447[5] + 
                kernel_img_mul_447[6] + kernel_img_mul_447[7] + kernel_img_mul_447[8] + 
                kernel_img_mul_447[9] + kernel_img_mul_447[10] + kernel_img_mul_447[11] + 
                kernel_img_mul_447[12] + kernel_img_mul_447[13] + kernel_img_mul_447[14] + 
                kernel_img_mul_447[15] + kernel_img_mul_447[16] + kernel_img_mul_447[17] + 
                kernel_img_mul_447[18] + kernel_img_mul_447[19] + kernel_img_mul_447[20] + 
                kernel_img_mul_447[21] + kernel_img_mul_447[22] + kernel_img_mul_447[23] + 
                kernel_img_mul_447[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3583:3576] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3583:3576] <= kernel_img_sum_447[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3583:3576] <= 'd0;
end

wire  [39:0]  kernel_img_mul_448[0:24];
assign kernel_img_mul_448[0] = buffer_data_4[3575:3568] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_448[1] = buffer_data_4[3583:3576] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_448[2] = buffer_data_4[3591:3584] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_448[3] = buffer_data_4[3599:3592] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_448[4] = buffer_data_4[3607:3600] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_448[5] = buffer_data_3[3575:3568] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_448[6] = buffer_data_3[3583:3576] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_448[7] = buffer_data_3[3591:3584] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_448[8] = buffer_data_3[3599:3592] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_448[9] = buffer_data_3[3607:3600] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_448[10] = buffer_data_2[3575:3568] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_448[11] = buffer_data_2[3583:3576] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_448[12] = buffer_data_2[3591:3584] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_448[13] = buffer_data_2[3599:3592] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_448[14] = buffer_data_2[3607:3600] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_448[15] = buffer_data_1[3575:3568] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_448[16] = buffer_data_1[3583:3576] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_448[17] = buffer_data_1[3591:3584] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_448[18] = buffer_data_1[3599:3592] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_448[19] = buffer_data_1[3607:3600] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_448[20] = buffer_data_0[3575:3568] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_448[21] = buffer_data_0[3583:3576] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_448[22] = buffer_data_0[3591:3584] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_448[23] = buffer_data_0[3599:3592] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_448[24] = buffer_data_0[3607:3600] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_448 = kernel_img_mul_448[0] + kernel_img_mul_448[1] + kernel_img_mul_448[2] + 
                kernel_img_mul_448[3] + kernel_img_mul_448[4] + kernel_img_mul_448[5] + 
                kernel_img_mul_448[6] + kernel_img_mul_448[7] + kernel_img_mul_448[8] + 
                kernel_img_mul_448[9] + kernel_img_mul_448[10] + kernel_img_mul_448[11] + 
                kernel_img_mul_448[12] + kernel_img_mul_448[13] + kernel_img_mul_448[14] + 
                kernel_img_mul_448[15] + kernel_img_mul_448[16] + kernel_img_mul_448[17] + 
                kernel_img_mul_448[18] + kernel_img_mul_448[19] + kernel_img_mul_448[20] + 
                kernel_img_mul_448[21] + kernel_img_mul_448[22] + kernel_img_mul_448[23] + 
                kernel_img_mul_448[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3591:3584] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3591:3584] <= kernel_img_sum_448[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3591:3584] <= 'd0;
end

wire  [39:0]  kernel_img_mul_449[0:24];
assign kernel_img_mul_449[0] = buffer_data_4[3583:3576] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_449[1] = buffer_data_4[3591:3584] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_449[2] = buffer_data_4[3599:3592] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_449[3] = buffer_data_4[3607:3600] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_449[4] = buffer_data_4[3615:3608] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_449[5] = buffer_data_3[3583:3576] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_449[6] = buffer_data_3[3591:3584] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_449[7] = buffer_data_3[3599:3592] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_449[8] = buffer_data_3[3607:3600] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_449[9] = buffer_data_3[3615:3608] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_449[10] = buffer_data_2[3583:3576] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_449[11] = buffer_data_2[3591:3584] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_449[12] = buffer_data_2[3599:3592] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_449[13] = buffer_data_2[3607:3600] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_449[14] = buffer_data_2[3615:3608] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_449[15] = buffer_data_1[3583:3576] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_449[16] = buffer_data_1[3591:3584] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_449[17] = buffer_data_1[3599:3592] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_449[18] = buffer_data_1[3607:3600] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_449[19] = buffer_data_1[3615:3608] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_449[20] = buffer_data_0[3583:3576] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_449[21] = buffer_data_0[3591:3584] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_449[22] = buffer_data_0[3599:3592] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_449[23] = buffer_data_0[3607:3600] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_449[24] = buffer_data_0[3615:3608] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_449 = kernel_img_mul_449[0] + kernel_img_mul_449[1] + kernel_img_mul_449[2] + 
                kernel_img_mul_449[3] + kernel_img_mul_449[4] + kernel_img_mul_449[5] + 
                kernel_img_mul_449[6] + kernel_img_mul_449[7] + kernel_img_mul_449[8] + 
                kernel_img_mul_449[9] + kernel_img_mul_449[10] + kernel_img_mul_449[11] + 
                kernel_img_mul_449[12] + kernel_img_mul_449[13] + kernel_img_mul_449[14] + 
                kernel_img_mul_449[15] + kernel_img_mul_449[16] + kernel_img_mul_449[17] + 
                kernel_img_mul_449[18] + kernel_img_mul_449[19] + kernel_img_mul_449[20] + 
                kernel_img_mul_449[21] + kernel_img_mul_449[22] + kernel_img_mul_449[23] + 
                kernel_img_mul_449[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3599:3592] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3599:3592] <= kernel_img_sum_449[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3599:3592] <= 'd0;
end

wire  [39:0]  kernel_img_mul_450[0:24];
assign kernel_img_mul_450[0] = buffer_data_4[3591:3584] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_450[1] = buffer_data_4[3599:3592] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_450[2] = buffer_data_4[3607:3600] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_450[3] = buffer_data_4[3615:3608] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_450[4] = buffer_data_4[3623:3616] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_450[5] = buffer_data_3[3591:3584] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_450[6] = buffer_data_3[3599:3592] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_450[7] = buffer_data_3[3607:3600] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_450[8] = buffer_data_3[3615:3608] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_450[9] = buffer_data_3[3623:3616] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_450[10] = buffer_data_2[3591:3584] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_450[11] = buffer_data_2[3599:3592] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_450[12] = buffer_data_2[3607:3600] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_450[13] = buffer_data_2[3615:3608] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_450[14] = buffer_data_2[3623:3616] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_450[15] = buffer_data_1[3591:3584] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_450[16] = buffer_data_1[3599:3592] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_450[17] = buffer_data_1[3607:3600] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_450[18] = buffer_data_1[3615:3608] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_450[19] = buffer_data_1[3623:3616] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_450[20] = buffer_data_0[3591:3584] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_450[21] = buffer_data_0[3599:3592] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_450[22] = buffer_data_0[3607:3600] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_450[23] = buffer_data_0[3615:3608] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_450[24] = buffer_data_0[3623:3616] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_450 = kernel_img_mul_450[0] + kernel_img_mul_450[1] + kernel_img_mul_450[2] + 
                kernel_img_mul_450[3] + kernel_img_mul_450[4] + kernel_img_mul_450[5] + 
                kernel_img_mul_450[6] + kernel_img_mul_450[7] + kernel_img_mul_450[8] + 
                kernel_img_mul_450[9] + kernel_img_mul_450[10] + kernel_img_mul_450[11] + 
                kernel_img_mul_450[12] + kernel_img_mul_450[13] + kernel_img_mul_450[14] + 
                kernel_img_mul_450[15] + kernel_img_mul_450[16] + kernel_img_mul_450[17] + 
                kernel_img_mul_450[18] + kernel_img_mul_450[19] + kernel_img_mul_450[20] + 
                kernel_img_mul_450[21] + kernel_img_mul_450[22] + kernel_img_mul_450[23] + 
                kernel_img_mul_450[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3607:3600] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3607:3600] <= kernel_img_sum_450[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3607:3600] <= 'd0;
end

wire  [39:0]  kernel_img_mul_451[0:24];
assign kernel_img_mul_451[0] = buffer_data_4[3599:3592] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_451[1] = buffer_data_4[3607:3600] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_451[2] = buffer_data_4[3615:3608] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_451[3] = buffer_data_4[3623:3616] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_451[4] = buffer_data_4[3631:3624] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_451[5] = buffer_data_3[3599:3592] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_451[6] = buffer_data_3[3607:3600] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_451[7] = buffer_data_3[3615:3608] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_451[8] = buffer_data_3[3623:3616] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_451[9] = buffer_data_3[3631:3624] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_451[10] = buffer_data_2[3599:3592] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_451[11] = buffer_data_2[3607:3600] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_451[12] = buffer_data_2[3615:3608] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_451[13] = buffer_data_2[3623:3616] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_451[14] = buffer_data_2[3631:3624] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_451[15] = buffer_data_1[3599:3592] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_451[16] = buffer_data_1[3607:3600] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_451[17] = buffer_data_1[3615:3608] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_451[18] = buffer_data_1[3623:3616] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_451[19] = buffer_data_1[3631:3624] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_451[20] = buffer_data_0[3599:3592] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_451[21] = buffer_data_0[3607:3600] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_451[22] = buffer_data_0[3615:3608] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_451[23] = buffer_data_0[3623:3616] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_451[24] = buffer_data_0[3631:3624] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_451 = kernel_img_mul_451[0] + kernel_img_mul_451[1] + kernel_img_mul_451[2] + 
                kernel_img_mul_451[3] + kernel_img_mul_451[4] + kernel_img_mul_451[5] + 
                kernel_img_mul_451[6] + kernel_img_mul_451[7] + kernel_img_mul_451[8] + 
                kernel_img_mul_451[9] + kernel_img_mul_451[10] + kernel_img_mul_451[11] + 
                kernel_img_mul_451[12] + kernel_img_mul_451[13] + kernel_img_mul_451[14] + 
                kernel_img_mul_451[15] + kernel_img_mul_451[16] + kernel_img_mul_451[17] + 
                kernel_img_mul_451[18] + kernel_img_mul_451[19] + kernel_img_mul_451[20] + 
                kernel_img_mul_451[21] + kernel_img_mul_451[22] + kernel_img_mul_451[23] + 
                kernel_img_mul_451[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3615:3608] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3615:3608] <= kernel_img_sum_451[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3615:3608] <= 'd0;
end

wire  [39:0]  kernel_img_mul_452[0:24];
assign kernel_img_mul_452[0] = buffer_data_4[3607:3600] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_452[1] = buffer_data_4[3615:3608] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_452[2] = buffer_data_4[3623:3616] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_452[3] = buffer_data_4[3631:3624] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_452[4] = buffer_data_4[3639:3632] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_452[5] = buffer_data_3[3607:3600] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_452[6] = buffer_data_3[3615:3608] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_452[7] = buffer_data_3[3623:3616] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_452[8] = buffer_data_3[3631:3624] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_452[9] = buffer_data_3[3639:3632] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_452[10] = buffer_data_2[3607:3600] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_452[11] = buffer_data_2[3615:3608] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_452[12] = buffer_data_2[3623:3616] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_452[13] = buffer_data_2[3631:3624] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_452[14] = buffer_data_2[3639:3632] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_452[15] = buffer_data_1[3607:3600] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_452[16] = buffer_data_1[3615:3608] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_452[17] = buffer_data_1[3623:3616] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_452[18] = buffer_data_1[3631:3624] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_452[19] = buffer_data_1[3639:3632] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_452[20] = buffer_data_0[3607:3600] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_452[21] = buffer_data_0[3615:3608] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_452[22] = buffer_data_0[3623:3616] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_452[23] = buffer_data_0[3631:3624] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_452[24] = buffer_data_0[3639:3632] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_452 = kernel_img_mul_452[0] + kernel_img_mul_452[1] + kernel_img_mul_452[2] + 
                kernel_img_mul_452[3] + kernel_img_mul_452[4] + kernel_img_mul_452[5] + 
                kernel_img_mul_452[6] + kernel_img_mul_452[7] + kernel_img_mul_452[8] + 
                kernel_img_mul_452[9] + kernel_img_mul_452[10] + kernel_img_mul_452[11] + 
                kernel_img_mul_452[12] + kernel_img_mul_452[13] + kernel_img_mul_452[14] + 
                kernel_img_mul_452[15] + kernel_img_mul_452[16] + kernel_img_mul_452[17] + 
                kernel_img_mul_452[18] + kernel_img_mul_452[19] + kernel_img_mul_452[20] + 
                kernel_img_mul_452[21] + kernel_img_mul_452[22] + kernel_img_mul_452[23] + 
                kernel_img_mul_452[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3623:3616] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3623:3616] <= kernel_img_sum_452[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3623:3616] <= 'd0;
end

wire  [39:0]  kernel_img_mul_453[0:24];
assign kernel_img_mul_453[0] = buffer_data_4[3615:3608] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_453[1] = buffer_data_4[3623:3616] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_453[2] = buffer_data_4[3631:3624] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_453[3] = buffer_data_4[3639:3632] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_453[4] = buffer_data_4[3647:3640] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_453[5] = buffer_data_3[3615:3608] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_453[6] = buffer_data_3[3623:3616] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_453[7] = buffer_data_3[3631:3624] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_453[8] = buffer_data_3[3639:3632] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_453[9] = buffer_data_3[3647:3640] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_453[10] = buffer_data_2[3615:3608] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_453[11] = buffer_data_2[3623:3616] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_453[12] = buffer_data_2[3631:3624] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_453[13] = buffer_data_2[3639:3632] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_453[14] = buffer_data_2[3647:3640] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_453[15] = buffer_data_1[3615:3608] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_453[16] = buffer_data_1[3623:3616] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_453[17] = buffer_data_1[3631:3624] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_453[18] = buffer_data_1[3639:3632] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_453[19] = buffer_data_1[3647:3640] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_453[20] = buffer_data_0[3615:3608] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_453[21] = buffer_data_0[3623:3616] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_453[22] = buffer_data_0[3631:3624] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_453[23] = buffer_data_0[3639:3632] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_453[24] = buffer_data_0[3647:3640] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_453 = kernel_img_mul_453[0] + kernel_img_mul_453[1] + kernel_img_mul_453[2] + 
                kernel_img_mul_453[3] + kernel_img_mul_453[4] + kernel_img_mul_453[5] + 
                kernel_img_mul_453[6] + kernel_img_mul_453[7] + kernel_img_mul_453[8] + 
                kernel_img_mul_453[9] + kernel_img_mul_453[10] + kernel_img_mul_453[11] + 
                kernel_img_mul_453[12] + kernel_img_mul_453[13] + kernel_img_mul_453[14] + 
                kernel_img_mul_453[15] + kernel_img_mul_453[16] + kernel_img_mul_453[17] + 
                kernel_img_mul_453[18] + kernel_img_mul_453[19] + kernel_img_mul_453[20] + 
                kernel_img_mul_453[21] + kernel_img_mul_453[22] + kernel_img_mul_453[23] + 
                kernel_img_mul_453[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3631:3624] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3631:3624] <= kernel_img_sum_453[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3631:3624] <= 'd0;
end

wire  [39:0]  kernel_img_mul_454[0:24];
assign kernel_img_mul_454[0] = buffer_data_4[3623:3616] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_454[1] = buffer_data_4[3631:3624] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_454[2] = buffer_data_4[3639:3632] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_454[3] = buffer_data_4[3647:3640] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_454[4] = buffer_data_4[3655:3648] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_454[5] = buffer_data_3[3623:3616] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_454[6] = buffer_data_3[3631:3624] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_454[7] = buffer_data_3[3639:3632] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_454[8] = buffer_data_3[3647:3640] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_454[9] = buffer_data_3[3655:3648] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_454[10] = buffer_data_2[3623:3616] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_454[11] = buffer_data_2[3631:3624] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_454[12] = buffer_data_2[3639:3632] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_454[13] = buffer_data_2[3647:3640] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_454[14] = buffer_data_2[3655:3648] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_454[15] = buffer_data_1[3623:3616] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_454[16] = buffer_data_1[3631:3624] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_454[17] = buffer_data_1[3639:3632] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_454[18] = buffer_data_1[3647:3640] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_454[19] = buffer_data_1[3655:3648] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_454[20] = buffer_data_0[3623:3616] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_454[21] = buffer_data_0[3631:3624] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_454[22] = buffer_data_0[3639:3632] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_454[23] = buffer_data_0[3647:3640] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_454[24] = buffer_data_0[3655:3648] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_454 = kernel_img_mul_454[0] + kernel_img_mul_454[1] + kernel_img_mul_454[2] + 
                kernel_img_mul_454[3] + kernel_img_mul_454[4] + kernel_img_mul_454[5] + 
                kernel_img_mul_454[6] + kernel_img_mul_454[7] + kernel_img_mul_454[8] + 
                kernel_img_mul_454[9] + kernel_img_mul_454[10] + kernel_img_mul_454[11] + 
                kernel_img_mul_454[12] + kernel_img_mul_454[13] + kernel_img_mul_454[14] + 
                kernel_img_mul_454[15] + kernel_img_mul_454[16] + kernel_img_mul_454[17] + 
                kernel_img_mul_454[18] + kernel_img_mul_454[19] + kernel_img_mul_454[20] + 
                kernel_img_mul_454[21] + kernel_img_mul_454[22] + kernel_img_mul_454[23] + 
                kernel_img_mul_454[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3639:3632] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3639:3632] <= kernel_img_sum_454[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3639:3632] <= 'd0;
end

wire  [39:0]  kernel_img_mul_455[0:24];
assign kernel_img_mul_455[0] = buffer_data_4[3631:3624] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_455[1] = buffer_data_4[3639:3632] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_455[2] = buffer_data_4[3647:3640] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_455[3] = buffer_data_4[3655:3648] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_455[4] = buffer_data_4[3663:3656] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_455[5] = buffer_data_3[3631:3624] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_455[6] = buffer_data_3[3639:3632] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_455[7] = buffer_data_3[3647:3640] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_455[8] = buffer_data_3[3655:3648] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_455[9] = buffer_data_3[3663:3656] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_455[10] = buffer_data_2[3631:3624] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_455[11] = buffer_data_2[3639:3632] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_455[12] = buffer_data_2[3647:3640] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_455[13] = buffer_data_2[3655:3648] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_455[14] = buffer_data_2[3663:3656] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_455[15] = buffer_data_1[3631:3624] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_455[16] = buffer_data_1[3639:3632] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_455[17] = buffer_data_1[3647:3640] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_455[18] = buffer_data_1[3655:3648] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_455[19] = buffer_data_1[3663:3656] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_455[20] = buffer_data_0[3631:3624] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_455[21] = buffer_data_0[3639:3632] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_455[22] = buffer_data_0[3647:3640] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_455[23] = buffer_data_0[3655:3648] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_455[24] = buffer_data_0[3663:3656] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_455 = kernel_img_mul_455[0] + kernel_img_mul_455[1] + kernel_img_mul_455[2] + 
                kernel_img_mul_455[3] + kernel_img_mul_455[4] + kernel_img_mul_455[5] + 
                kernel_img_mul_455[6] + kernel_img_mul_455[7] + kernel_img_mul_455[8] + 
                kernel_img_mul_455[9] + kernel_img_mul_455[10] + kernel_img_mul_455[11] + 
                kernel_img_mul_455[12] + kernel_img_mul_455[13] + kernel_img_mul_455[14] + 
                kernel_img_mul_455[15] + kernel_img_mul_455[16] + kernel_img_mul_455[17] + 
                kernel_img_mul_455[18] + kernel_img_mul_455[19] + kernel_img_mul_455[20] + 
                kernel_img_mul_455[21] + kernel_img_mul_455[22] + kernel_img_mul_455[23] + 
                kernel_img_mul_455[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3647:3640] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3647:3640] <= kernel_img_sum_455[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3647:3640] <= 'd0;
end

wire  [39:0]  kernel_img_mul_456[0:24];
assign kernel_img_mul_456[0] = buffer_data_4[3639:3632] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_456[1] = buffer_data_4[3647:3640] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_456[2] = buffer_data_4[3655:3648] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_456[3] = buffer_data_4[3663:3656] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_456[4] = buffer_data_4[3671:3664] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_456[5] = buffer_data_3[3639:3632] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_456[6] = buffer_data_3[3647:3640] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_456[7] = buffer_data_3[3655:3648] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_456[8] = buffer_data_3[3663:3656] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_456[9] = buffer_data_3[3671:3664] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_456[10] = buffer_data_2[3639:3632] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_456[11] = buffer_data_2[3647:3640] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_456[12] = buffer_data_2[3655:3648] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_456[13] = buffer_data_2[3663:3656] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_456[14] = buffer_data_2[3671:3664] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_456[15] = buffer_data_1[3639:3632] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_456[16] = buffer_data_1[3647:3640] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_456[17] = buffer_data_1[3655:3648] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_456[18] = buffer_data_1[3663:3656] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_456[19] = buffer_data_1[3671:3664] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_456[20] = buffer_data_0[3639:3632] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_456[21] = buffer_data_0[3647:3640] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_456[22] = buffer_data_0[3655:3648] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_456[23] = buffer_data_0[3663:3656] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_456[24] = buffer_data_0[3671:3664] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_456 = kernel_img_mul_456[0] + kernel_img_mul_456[1] + kernel_img_mul_456[2] + 
                kernel_img_mul_456[3] + kernel_img_mul_456[4] + kernel_img_mul_456[5] + 
                kernel_img_mul_456[6] + kernel_img_mul_456[7] + kernel_img_mul_456[8] + 
                kernel_img_mul_456[9] + kernel_img_mul_456[10] + kernel_img_mul_456[11] + 
                kernel_img_mul_456[12] + kernel_img_mul_456[13] + kernel_img_mul_456[14] + 
                kernel_img_mul_456[15] + kernel_img_mul_456[16] + kernel_img_mul_456[17] + 
                kernel_img_mul_456[18] + kernel_img_mul_456[19] + kernel_img_mul_456[20] + 
                kernel_img_mul_456[21] + kernel_img_mul_456[22] + kernel_img_mul_456[23] + 
                kernel_img_mul_456[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3655:3648] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3655:3648] <= kernel_img_sum_456[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3655:3648] <= 'd0;
end

wire  [39:0]  kernel_img_mul_457[0:24];
assign kernel_img_mul_457[0] = buffer_data_4[3647:3640] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_457[1] = buffer_data_4[3655:3648] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_457[2] = buffer_data_4[3663:3656] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_457[3] = buffer_data_4[3671:3664] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_457[4] = buffer_data_4[3679:3672] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_457[5] = buffer_data_3[3647:3640] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_457[6] = buffer_data_3[3655:3648] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_457[7] = buffer_data_3[3663:3656] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_457[8] = buffer_data_3[3671:3664] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_457[9] = buffer_data_3[3679:3672] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_457[10] = buffer_data_2[3647:3640] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_457[11] = buffer_data_2[3655:3648] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_457[12] = buffer_data_2[3663:3656] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_457[13] = buffer_data_2[3671:3664] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_457[14] = buffer_data_2[3679:3672] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_457[15] = buffer_data_1[3647:3640] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_457[16] = buffer_data_1[3655:3648] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_457[17] = buffer_data_1[3663:3656] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_457[18] = buffer_data_1[3671:3664] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_457[19] = buffer_data_1[3679:3672] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_457[20] = buffer_data_0[3647:3640] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_457[21] = buffer_data_0[3655:3648] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_457[22] = buffer_data_0[3663:3656] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_457[23] = buffer_data_0[3671:3664] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_457[24] = buffer_data_0[3679:3672] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_457 = kernel_img_mul_457[0] + kernel_img_mul_457[1] + kernel_img_mul_457[2] + 
                kernel_img_mul_457[3] + kernel_img_mul_457[4] + kernel_img_mul_457[5] + 
                kernel_img_mul_457[6] + kernel_img_mul_457[7] + kernel_img_mul_457[8] + 
                kernel_img_mul_457[9] + kernel_img_mul_457[10] + kernel_img_mul_457[11] + 
                kernel_img_mul_457[12] + kernel_img_mul_457[13] + kernel_img_mul_457[14] + 
                kernel_img_mul_457[15] + kernel_img_mul_457[16] + kernel_img_mul_457[17] + 
                kernel_img_mul_457[18] + kernel_img_mul_457[19] + kernel_img_mul_457[20] + 
                kernel_img_mul_457[21] + kernel_img_mul_457[22] + kernel_img_mul_457[23] + 
                kernel_img_mul_457[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3663:3656] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3663:3656] <= kernel_img_sum_457[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3663:3656] <= 'd0;
end

wire  [39:0]  kernel_img_mul_458[0:24];
assign kernel_img_mul_458[0] = buffer_data_4[3655:3648] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_458[1] = buffer_data_4[3663:3656] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_458[2] = buffer_data_4[3671:3664] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_458[3] = buffer_data_4[3679:3672] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_458[4] = buffer_data_4[3687:3680] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_458[5] = buffer_data_3[3655:3648] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_458[6] = buffer_data_3[3663:3656] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_458[7] = buffer_data_3[3671:3664] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_458[8] = buffer_data_3[3679:3672] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_458[9] = buffer_data_3[3687:3680] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_458[10] = buffer_data_2[3655:3648] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_458[11] = buffer_data_2[3663:3656] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_458[12] = buffer_data_2[3671:3664] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_458[13] = buffer_data_2[3679:3672] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_458[14] = buffer_data_2[3687:3680] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_458[15] = buffer_data_1[3655:3648] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_458[16] = buffer_data_1[3663:3656] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_458[17] = buffer_data_1[3671:3664] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_458[18] = buffer_data_1[3679:3672] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_458[19] = buffer_data_1[3687:3680] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_458[20] = buffer_data_0[3655:3648] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_458[21] = buffer_data_0[3663:3656] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_458[22] = buffer_data_0[3671:3664] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_458[23] = buffer_data_0[3679:3672] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_458[24] = buffer_data_0[3687:3680] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_458 = kernel_img_mul_458[0] + kernel_img_mul_458[1] + kernel_img_mul_458[2] + 
                kernel_img_mul_458[3] + kernel_img_mul_458[4] + kernel_img_mul_458[5] + 
                kernel_img_mul_458[6] + kernel_img_mul_458[7] + kernel_img_mul_458[8] + 
                kernel_img_mul_458[9] + kernel_img_mul_458[10] + kernel_img_mul_458[11] + 
                kernel_img_mul_458[12] + kernel_img_mul_458[13] + kernel_img_mul_458[14] + 
                kernel_img_mul_458[15] + kernel_img_mul_458[16] + kernel_img_mul_458[17] + 
                kernel_img_mul_458[18] + kernel_img_mul_458[19] + kernel_img_mul_458[20] + 
                kernel_img_mul_458[21] + kernel_img_mul_458[22] + kernel_img_mul_458[23] + 
                kernel_img_mul_458[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3671:3664] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3671:3664] <= kernel_img_sum_458[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3671:3664] <= 'd0;
end

wire  [39:0]  kernel_img_mul_459[0:24];
assign kernel_img_mul_459[0] = buffer_data_4[3663:3656] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_459[1] = buffer_data_4[3671:3664] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_459[2] = buffer_data_4[3679:3672] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_459[3] = buffer_data_4[3687:3680] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_459[4] = buffer_data_4[3695:3688] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_459[5] = buffer_data_3[3663:3656] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_459[6] = buffer_data_3[3671:3664] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_459[7] = buffer_data_3[3679:3672] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_459[8] = buffer_data_3[3687:3680] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_459[9] = buffer_data_3[3695:3688] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_459[10] = buffer_data_2[3663:3656] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_459[11] = buffer_data_2[3671:3664] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_459[12] = buffer_data_2[3679:3672] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_459[13] = buffer_data_2[3687:3680] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_459[14] = buffer_data_2[3695:3688] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_459[15] = buffer_data_1[3663:3656] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_459[16] = buffer_data_1[3671:3664] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_459[17] = buffer_data_1[3679:3672] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_459[18] = buffer_data_1[3687:3680] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_459[19] = buffer_data_1[3695:3688] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_459[20] = buffer_data_0[3663:3656] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_459[21] = buffer_data_0[3671:3664] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_459[22] = buffer_data_0[3679:3672] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_459[23] = buffer_data_0[3687:3680] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_459[24] = buffer_data_0[3695:3688] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_459 = kernel_img_mul_459[0] + kernel_img_mul_459[1] + kernel_img_mul_459[2] + 
                kernel_img_mul_459[3] + kernel_img_mul_459[4] + kernel_img_mul_459[5] + 
                kernel_img_mul_459[6] + kernel_img_mul_459[7] + kernel_img_mul_459[8] + 
                kernel_img_mul_459[9] + kernel_img_mul_459[10] + kernel_img_mul_459[11] + 
                kernel_img_mul_459[12] + kernel_img_mul_459[13] + kernel_img_mul_459[14] + 
                kernel_img_mul_459[15] + kernel_img_mul_459[16] + kernel_img_mul_459[17] + 
                kernel_img_mul_459[18] + kernel_img_mul_459[19] + kernel_img_mul_459[20] + 
                kernel_img_mul_459[21] + kernel_img_mul_459[22] + kernel_img_mul_459[23] + 
                kernel_img_mul_459[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3679:3672] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3679:3672] <= kernel_img_sum_459[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3679:3672] <= 'd0;
end

wire  [39:0]  kernel_img_mul_460[0:24];
assign kernel_img_mul_460[0] = buffer_data_4[3671:3664] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_460[1] = buffer_data_4[3679:3672] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_460[2] = buffer_data_4[3687:3680] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_460[3] = buffer_data_4[3695:3688] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_460[4] = buffer_data_4[3703:3696] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_460[5] = buffer_data_3[3671:3664] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_460[6] = buffer_data_3[3679:3672] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_460[7] = buffer_data_3[3687:3680] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_460[8] = buffer_data_3[3695:3688] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_460[9] = buffer_data_3[3703:3696] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_460[10] = buffer_data_2[3671:3664] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_460[11] = buffer_data_2[3679:3672] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_460[12] = buffer_data_2[3687:3680] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_460[13] = buffer_data_2[3695:3688] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_460[14] = buffer_data_2[3703:3696] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_460[15] = buffer_data_1[3671:3664] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_460[16] = buffer_data_1[3679:3672] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_460[17] = buffer_data_1[3687:3680] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_460[18] = buffer_data_1[3695:3688] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_460[19] = buffer_data_1[3703:3696] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_460[20] = buffer_data_0[3671:3664] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_460[21] = buffer_data_0[3679:3672] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_460[22] = buffer_data_0[3687:3680] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_460[23] = buffer_data_0[3695:3688] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_460[24] = buffer_data_0[3703:3696] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_460 = kernel_img_mul_460[0] + kernel_img_mul_460[1] + kernel_img_mul_460[2] + 
                kernel_img_mul_460[3] + kernel_img_mul_460[4] + kernel_img_mul_460[5] + 
                kernel_img_mul_460[6] + kernel_img_mul_460[7] + kernel_img_mul_460[8] + 
                kernel_img_mul_460[9] + kernel_img_mul_460[10] + kernel_img_mul_460[11] + 
                kernel_img_mul_460[12] + kernel_img_mul_460[13] + kernel_img_mul_460[14] + 
                kernel_img_mul_460[15] + kernel_img_mul_460[16] + kernel_img_mul_460[17] + 
                kernel_img_mul_460[18] + kernel_img_mul_460[19] + kernel_img_mul_460[20] + 
                kernel_img_mul_460[21] + kernel_img_mul_460[22] + kernel_img_mul_460[23] + 
                kernel_img_mul_460[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3687:3680] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3687:3680] <= kernel_img_sum_460[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3687:3680] <= 'd0;
end

wire  [39:0]  kernel_img_mul_461[0:24];
assign kernel_img_mul_461[0] = buffer_data_4[3679:3672] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_461[1] = buffer_data_4[3687:3680] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_461[2] = buffer_data_4[3695:3688] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_461[3] = buffer_data_4[3703:3696] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_461[4] = buffer_data_4[3711:3704] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_461[5] = buffer_data_3[3679:3672] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_461[6] = buffer_data_3[3687:3680] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_461[7] = buffer_data_3[3695:3688] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_461[8] = buffer_data_3[3703:3696] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_461[9] = buffer_data_3[3711:3704] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_461[10] = buffer_data_2[3679:3672] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_461[11] = buffer_data_2[3687:3680] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_461[12] = buffer_data_2[3695:3688] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_461[13] = buffer_data_2[3703:3696] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_461[14] = buffer_data_2[3711:3704] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_461[15] = buffer_data_1[3679:3672] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_461[16] = buffer_data_1[3687:3680] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_461[17] = buffer_data_1[3695:3688] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_461[18] = buffer_data_1[3703:3696] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_461[19] = buffer_data_1[3711:3704] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_461[20] = buffer_data_0[3679:3672] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_461[21] = buffer_data_0[3687:3680] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_461[22] = buffer_data_0[3695:3688] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_461[23] = buffer_data_0[3703:3696] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_461[24] = buffer_data_0[3711:3704] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_461 = kernel_img_mul_461[0] + kernel_img_mul_461[1] + kernel_img_mul_461[2] + 
                kernel_img_mul_461[3] + kernel_img_mul_461[4] + kernel_img_mul_461[5] + 
                kernel_img_mul_461[6] + kernel_img_mul_461[7] + kernel_img_mul_461[8] + 
                kernel_img_mul_461[9] + kernel_img_mul_461[10] + kernel_img_mul_461[11] + 
                kernel_img_mul_461[12] + kernel_img_mul_461[13] + kernel_img_mul_461[14] + 
                kernel_img_mul_461[15] + kernel_img_mul_461[16] + kernel_img_mul_461[17] + 
                kernel_img_mul_461[18] + kernel_img_mul_461[19] + kernel_img_mul_461[20] + 
                kernel_img_mul_461[21] + kernel_img_mul_461[22] + kernel_img_mul_461[23] + 
                kernel_img_mul_461[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3695:3688] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3695:3688] <= kernel_img_sum_461[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3695:3688] <= 'd0;
end

wire  [39:0]  kernel_img_mul_462[0:24];
assign kernel_img_mul_462[0] = buffer_data_4[3687:3680] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_462[1] = buffer_data_4[3695:3688] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_462[2] = buffer_data_4[3703:3696] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_462[3] = buffer_data_4[3711:3704] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_462[4] = buffer_data_4[3719:3712] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_462[5] = buffer_data_3[3687:3680] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_462[6] = buffer_data_3[3695:3688] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_462[7] = buffer_data_3[3703:3696] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_462[8] = buffer_data_3[3711:3704] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_462[9] = buffer_data_3[3719:3712] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_462[10] = buffer_data_2[3687:3680] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_462[11] = buffer_data_2[3695:3688] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_462[12] = buffer_data_2[3703:3696] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_462[13] = buffer_data_2[3711:3704] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_462[14] = buffer_data_2[3719:3712] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_462[15] = buffer_data_1[3687:3680] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_462[16] = buffer_data_1[3695:3688] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_462[17] = buffer_data_1[3703:3696] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_462[18] = buffer_data_1[3711:3704] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_462[19] = buffer_data_1[3719:3712] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_462[20] = buffer_data_0[3687:3680] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_462[21] = buffer_data_0[3695:3688] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_462[22] = buffer_data_0[3703:3696] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_462[23] = buffer_data_0[3711:3704] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_462[24] = buffer_data_0[3719:3712] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_462 = kernel_img_mul_462[0] + kernel_img_mul_462[1] + kernel_img_mul_462[2] + 
                kernel_img_mul_462[3] + kernel_img_mul_462[4] + kernel_img_mul_462[5] + 
                kernel_img_mul_462[6] + kernel_img_mul_462[7] + kernel_img_mul_462[8] + 
                kernel_img_mul_462[9] + kernel_img_mul_462[10] + kernel_img_mul_462[11] + 
                kernel_img_mul_462[12] + kernel_img_mul_462[13] + kernel_img_mul_462[14] + 
                kernel_img_mul_462[15] + kernel_img_mul_462[16] + kernel_img_mul_462[17] + 
                kernel_img_mul_462[18] + kernel_img_mul_462[19] + kernel_img_mul_462[20] + 
                kernel_img_mul_462[21] + kernel_img_mul_462[22] + kernel_img_mul_462[23] + 
                kernel_img_mul_462[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3703:3696] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3703:3696] <= kernel_img_sum_462[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3703:3696] <= 'd0;
end

wire  [39:0]  kernel_img_mul_463[0:24];
assign kernel_img_mul_463[0] = buffer_data_4[3695:3688] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_463[1] = buffer_data_4[3703:3696] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_463[2] = buffer_data_4[3711:3704] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_463[3] = buffer_data_4[3719:3712] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_463[4] = buffer_data_4[3727:3720] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_463[5] = buffer_data_3[3695:3688] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_463[6] = buffer_data_3[3703:3696] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_463[7] = buffer_data_3[3711:3704] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_463[8] = buffer_data_3[3719:3712] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_463[9] = buffer_data_3[3727:3720] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_463[10] = buffer_data_2[3695:3688] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_463[11] = buffer_data_2[3703:3696] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_463[12] = buffer_data_2[3711:3704] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_463[13] = buffer_data_2[3719:3712] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_463[14] = buffer_data_2[3727:3720] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_463[15] = buffer_data_1[3695:3688] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_463[16] = buffer_data_1[3703:3696] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_463[17] = buffer_data_1[3711:3704] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_463[18] = buffer_data_1[3719:3712] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_463[19] = buffer_data_1[3727:3720] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_463[20] = buffer_data_0[3695:3688] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_463[21] = buffer_data_0[3703:3696] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_463[22] = buffer_data_0[3711:3704] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_463[23] = buffer_data_0[3719:3712] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_463[24] = buffer_data_0[3727:3720] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_463 = kernel_img_mul_463[0] + kernel_img_mul_463[1] + kernel_img_mul_463[2] + 
                kernel_img_mul_463[3] + kernel_img_mul_463[4] + kernel_img_mul_463[5] + 
                kernel_img_mul_463[6] + kernel_img_mul_463[7] + kernel_img_mul_463[8] + 
                kernel_img_mul_463[9] + kernel_img_mul_463[10] + kernel_img_mul_463[11] + 
                kernel_img_mul_463[12] + kernel_img_mul_463[13] + kernel_img_mul_463[14] + 
                kernel_img_mul_463[15] + kernel_img_mul_463[16] + kernel_img_mul_463[17] + 
                kernel_img_mul_463[18] + kernel_img_mul_463[19] + kernel_img_mul_463[20] + 
                kernel_img_mul_463[21] + kernel_img_mul_463[22] + kernel_img_mul_463[23] + 
                kernel_img_mul_463[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3711:3704] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3711:3704] <= kernel_img_sum_463[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3711:3704] <= 'd0;
end

wire  [39:0]  kernel_img_mul_464[0:24];
assign kernel_img_mul_464[0] = buffer_data_4[3703:3696] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_464[1] = buffer_data_4[3711:3704] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_464[2] = buffer_data_4[3719:3712] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_464[3] = buffer_data_4[3727:3720] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_464[4] = buffer_data_4[3735:3728] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_464[5] = buffer_data_3[3703:3696] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_464[6] = buffer_data_3[3711:3704] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_464[7] = buffer_data_3[3719:3712] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_464[8] = buffer_data_3[3727:3720] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_464[9] = buffer_data_3[3735:3728] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_464[10] = buffer_data_2[3703:3696] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_464[11] = buffer_data_2[3711:3704] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_464[12] = buffer_data_2[3719:3712] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_464[13] = buffer_data_2[3727:3720] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_464[14] = buffer_data_2[3735:3728] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_464[15] = buffer_data_1[3703:3696] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_464[16] = buffer_data_1[3711:3704] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_464[17] = buffer_data_1[3719:3712] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_464[18] = buffer_data_1[3727:3720] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_464[19] = buffer_data_1[3735:3728] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_464[20] = buffer_data_0[3703:3696] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_464[21] = buffer_data_0[3711:3704] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_464[22] = buffer_data_0[3719:3712] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_464[23] = buffer_data_0[3727:3720] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_464[24] = buffer_data_0[3735:3728] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_464 = kernel_img_mul_464[0] + kernel_img_mul_464[1] + kernel_img_mul_464[2] + 
                kernel_img_mul_464[3] + kernel_img_mul_464[4] + kernel_img_mul_464[5] + 
                kernel_img_mul_464[6] + kernel_img_mul_464[7] + kernel_img_mul_464[8] + 
                kernel_img_mul_464[9] + kernel_img_mul_464[10] + kernel_img_mul_464[11] + 
                kernel_img_mul_464[12] + kernel_img_mul_464[13] + kernel_img_mul_464[14] + 
                kernel_img_mul_464[15] + kernel_img_mul_464[16] + kernel_img_mul_464[17] + 
                kernel_img_mul_464[18] + kernel_img_mul_464[19] + kernel_img_mul_464[20] + 
                kernel_img_mul_464[21] + kernel_img_mul_464[22] + kernel_img_mul_464[23] + 
                kernel_img_mul_464[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3719:3712] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3719:3712] <= kernel_img_sum_464[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3719:3712] <= 'd0;
end

wire  [39:0]  kernel_img_mul_465[0:24];
assign kernel_img_mul_465[0] = buffer_data_4[3711:3704] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_465[1] = buffer_data_4[3719:3712] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_465[2] = buffer_data_4[3727:3720] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_465[3] = buffer_data_4[3735:3728] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_465[4] = buffer_data_4[3743:3736] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_465[5] = buffer_data_3[3711:3704] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_465[6] = buffer_data_3[3719:3712] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_465[7] = buffer_data_3[3727:3720] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_465[8] = buffer_data_3[3735:3728] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_465[9] = buffer_data_3[3743:3736] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_465[10] = buffer_data_2[3711:3704] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_465[11] = buffer_data_2[3719:3712] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_465[12] = buffer_data_2[3727:3720] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_465[13] = buffer_data_2[3735:3728] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_465[14] = buffer_data_2[3743:3736] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_465[15] = buffer_data_1[3711:3704] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_465[16] = buffer_data_1[3719:3712] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_465[17] = buffer_data_1[3727:3720] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_465[18] = buffer_data_1[3735:3728] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_465[19] = buffer_data_1[3743:3736] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_465[20] = buffer_data_0[3711:3704] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_465[21] = buffer_data_0[3719:3712] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_465[22] = buffer_data_0[3727:3720] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_465[23] = buffer_data_0[3735:3728] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_465[24] = buffer_data_0[3743:3736] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_465 = kernel_img_mul_465[0] + kernel_img_mul_465[1] + kernel_img_mul_465[2] + 
                kernel_img_mul_465[3] + kernel_img_mul_465[4] + kernel_img_mul_465[5] + 
                kernel_img_mul_465[6] + kernel_img_mul_465[7] + kernel_img_mul_465[8] + 
                kernel_img_mul_465[9] + kernel_img_mul_465[10] + kernel_img_mul_465[11] + 
                kernel_img_mul_465[12] + kernel_img_mul_465[13] + kernel_img_mul_465[14] + 
                kernel_img_mul_465[15] + kernel_img_mul_465[16] + kernel_img_mul_465[17] + 
                kernel_img_mul_465[18] + kernel_img_mul_465[19] + kernel_img_mul_465[20] + 
                kernel_img_mul_465[21] + kernel_img_mul_465[22] + kernel_img_mul_465[23] + 
                kernel_img_mul_465[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3727:3720] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3727:3720] <= kernel_img_sum_465[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3727:3720] <= 'd0;
end

wire  [39:0]  kernel_img_mul_466[0:24];
assign kernel_img_mul_466[0] = buffer_data_4[3719:3712] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_466[1] = buffer_data_4[3727:3720] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_466[2] = buffer_data_4[3735:3728] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_466[3] = buffer_data_4[3743:3736] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_466[4] = buffer_data_4[3751:3744] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_466[5] = buffer_data_3[3719:3712] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_466[6] = buffer_data_3[3727:3720] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_466[7] = buffer_data_3[3735:3728] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_466[8] = buffer_data_3[3743:3736] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_466[9] = buffer_data_3[3751:3744] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_466[10] = buffer_data_2[3719:3712] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_466[11] = buffer_data_2[3727:3720] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_466[12] = buffer_data_2[3735:3728] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_466[13] = buffer_data_2[3743:3736] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_466[14] = buffer_data_2[3751:3744] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_466[15] = buffer_data_1[3719:3712] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_466[16] = buffer_data_1[3727:3720] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_466[17] = buffer_data_1[3735:3728] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_466[18] = buffer_data_1[3743:3736] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_466[19] = buffer_data_1[3751:3744] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_466[20] = buffer_data_0[3719:3712] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_466[21] = buffer_data_0[3727:3720] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_466[22] = buffer_data_0[3735:3728] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_466[23] = buffer_data_0[3743:3736] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_466[24] = buffer_data_0[3751:3744] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_466 = kernel_img_mul_466[0] + kernel_img_mul_466[1] + kernel_img_mul_466[2] + 
                kernel_img_mul_466[3] + kernel_img_mul_466[4] + kernel_img_mul_466[5] + 
                kernel_img_mul_466[6] + kernel_img_mul_466[7] + kernel_img_mul_466[8] + 
                kernel_img_mul_466[9] + kernel_img_mul_466[10] + kernel_img_mul_466[11] + 
                kernel_img_mul_466[12] + kernel_img_mul_466[13] + kernel_img_mul_466[14] + 
                kernel_img_mul_466[15] + kernel_img_mul_466[16] + kernel_img_mul_466[17] + 
                kernel_img_mul_466[18] + kernel_img_mul_466[19] + kernel_img_mul_466[20] + 
                kernel_img_mul_466[21] + kernel_img_mul_466[22] + kernel_img_mul_466[23] + 
                kernel_img_mul_466[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3735:3728] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3735:3728] <= kernel_img_sum_466[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3735:3728] <= 'd0;
end

wire  [39:0]  kernel_img_mul_467[0:24];
assign kernel_img_mul_467[0] = buffer_data_4[3727:3720] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_467[1] = buffer_data_4[3735:3728] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_467[2] = buffer_data_4[3743:3736] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_467[3] = buffer_data_4[3751:3744] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_467[4] = buffer_data_4[3759:3752] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_467[5] = buffer_data_3[3727:3720] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_467[6] = buffer_data_3[3735:3728] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_467[7] = buffer_data_3[3743:3736] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_467[8] = buffer_data_3[3751:3744] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_467[9] = buffer_data_3[3759:3752] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_467[10] = buffer_data_2[3727:3720] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_467[11] = buffer_data_2[3735:3728] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_467[12] = buffer_data_2[3743:3736] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_467[13] = buffer_data_2[3751:3744] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_467[14] = buffer_data_2[3759:3752] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_467[15] = buffer_data_1[3727:3720] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_467[16] = buffer_data_1[3735:3728] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_467[17] = buffer_data_1[3743:3736] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_467[18] = buffer_data_1[3751:3744] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_467[19] = buffer_data_1[3759:3752] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_467[20] = buffer_data_0[3727:3720] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_467[21] = buffer_data_0[3735:3728] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_467[22] = buffer_data_0[3743:3736] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_467[23] = buffer_data_0[3751:3744] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_467[24] = buffer_data_0[3759:3752] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_467 = kernel_img_mul_467[0] + kernel_img_mul_467[1] + kernel_img_mul_467[2] + 
                kernel_img_mul_467[3] + kernel_img_mul_467[4] + kernel_img_mul_467[5] + 
                kernel_img_mul_467[6] + kernel_img_mul_467[7] + kernel_img_mul_467[8] + 
                kernel_img_mul_467[9] + kernel_img_mul_467[10] + kernel_img_mul_467[11] + 
                kernel_img_mul_467[12] + kernel_img_mul_467[13] + kernel_img_mul_467[14] + 
                kernel_img_mul_467[15] + kernel_img_mul_467[16] + kernel_img_mul_467[17] + 
                kernel_img_mul_467[18] + kernel_img_mul_467[19] + kernel_img_mul_467[20] + 
                kernel_img_mul_467[21] + kernel_img_mul_467[22] + kernel_img_mul_467[23] + 
                kernel_img_mul_467[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3743:3736] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3743:3736] <= kernel_img_sum_467[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3743:3736] <= 'd0;
end

wire  [39:0]  kernel_img_mul_468[0:24];
assign kernel_img_mul_468[0] = buffer_data_4[3735:3728] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_468[1] = buffer_data_4[3743:3736] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_468[2] = buffer_data_4[3751:3744] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_468[3] = buffer_data_4[3759:3752] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_468[4] = buffer_data_4[3767:3760] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_468[5] = buffer_data_3[3735:3728] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_468[6] = buffer_data_3[3743:3736] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_468[7] = buffer_data_3[3751:3744] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_468[8] = buffer_data_3[3759:3752] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_468[9] = buffer_data_3[3767:3760] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_468[10] = buffer_data_2[3735:3728] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_468[11] = buffer_data_2[3743:3736] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_468[12] = buffer_data_2[3751:3744] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_468[13] = buffer_data_2[3759:3752] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_468[14] = buffer_data_2[3767:3760] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_468[15] = buffer_data_1[3735:3728] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_468[16] = buffer_data_1[3743:3736] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_468[17] = buffer_data_1[3751:3744] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_468[18] = buffer_data_1[3759:3752] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_468[19] = buffer_data_1[3767:3760] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_468[20] = buffer_data_0[3735:3728] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_468[21] = buffer_data_0[3743:3736] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_468[22] = buffer_data_0[3751:3744] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_468[23] = buffer_data_0[3759:3752] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_468[24] = buffer_data_0[3767:3760] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_468 = kernel_img_mul_468[0] + kernel_img_mul_468[1] + kernel_img_mul_468[2] + 
                kernel_img_mul_468[3] + kernel_img_mul_468[4] + kernel_img_mul_468[5] + 
                kernel_img_mul_468[6] + kernel_img_mul_468[7] + kernel_img_mul_468[8] + 
                kernel_img_mul_468[9] + kernel_img_mul_468[10] + kernel_img_mul_468[11] + 
                kernel_img_mul_468[12] + kernel_img_mul_468[13] + kernel_img_mul_468[14] + 
                kernel_img_mul_468[15] + kernel_img_mul_468[16] + kernel_img_mul_468[17] + 
                kernel_img_mul_468[18] + kernel_img_mul_468[19] + kernel_img_mul_468[20] + 
                kernel_img_mul_468[21] + kernel_img_mul_468[22] + kernel_img_mul_468[23] + 
                kernel_img_mul_468[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3751:3744] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3751:3744] <= kernel_img_sum_468[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3751:3744] <= 'd0;
end

wire  [39:0]  kernel_img_mul_469[0:24];
assign kernel_img_mul_469[0] = buffer_data_4[3743:3736] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_469[1] = buffer_data_4[3751:3744] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_469[2] = buffer_data_4[3759:3752] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_469[3] = buffer_data_4[3767:3760] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_469[4] = buffer_data_4[3775:3768] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_469[5] = buffer_data_3[3743:3736] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_469[6] = buffer_data_3[3751:3744] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_469[7] = buffer_data_3[3759:3752] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_469[8] = buffer_data_3[3767:3760] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_469[9] = buffer_data_3[3775:3768] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_469[10] = buffer_data_2[3743:3736] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_469[11] = buffer_data_2[3751:3744] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_469[12] = buffer_data_2[3759:3752] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_469[13] = buffer_data_2[3767:3760] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_469[14] = buffer_data_2[3775:3768] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_469[15] = buffer_data_1[3743:3736] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_469[16] = buffer_data_1[3751:3744] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_469[17] = buffer_data_1[3759:3752] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_469[18] = buffer_data_1[3767:3760] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_469[19] = buffer_data_1[3775:3768] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_469[20] = buffer_data_0[3743:3736] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_469[21] = buffer_data_0[3751:3744] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_469[22] = buffer_data_0[3759:3752] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_469[23] = buffer_data_0[3767:3760] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_469[24] = buffer_data_0[3775:3768] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_469 = kernel_img_mul_469[0] + kernel_img_mul_469[1] + kernel_img_mul_469[2] + 
                kernel_img_mul_469[3] + kernel_img_mul_469[4] + kernel_img_mul_469[5] + 
                kernel_img_mul_469[6] + kernel_img_mul_469[7] + kernel_img_mul_469[8] + 
                kernel_img_mul_469[9] + kernel_img_mul_469[10] + kernel_img_mul_469[11] + 
                kernel_img_mul_469[12] + kernel_img_mul_469[13] + kernel_img_mul_469[14] + 
                kernel_img_mul_469[15] + kernel_img_mul_469[16] + kernel_img_mul_469[17] + 
                kernel_img_mul_469[18] + kernel_img_mul_469[19] + kernel_img_mul_469[20] + 
                kernel_img_mul_469[21] + kernel_img_mul_469[22] + kernel_img_mul_469[23] + 
                kernel_img_mul_469[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3759:3752] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3759:3752] <= kernel_img_sum_469[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3759:3752] <= 'd0;
end

wire  [39:0]  kernel_img_mul_470[0:24];
assign kernel_img_mul_470[0] = buffer_data_4[3751:3744] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_470[1] = buffer_data_4[3759:3752] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_470[2] = buffer_data_4[3767:3760] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_470[3] = buffer_data_4[3775:3768] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_470[4] = buffer_data_4[3783:3776] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_470[5] = buffer_data_3[3751:3744] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_470[6] = buffer_data_3[3759:3752] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_470[7] = buffer_data_3[3767:3760] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_470[8] = buffer_data_3[3775:3768] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_470[9] = buffer_data_3[3783:3776] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_470[10] = buffer_data_2[3751:3744] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_470[11] = buffer_data_2[3759:3752] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_470[12] = buffer_data_2[3767:3760] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_470[13] = buffer_data_2[3775:3768] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_470[14] = buffer_data_2[3783:3776] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_470[15] = buffer_data_1[3751:3744] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_470[16] = buffer_data_1[3759:3752] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_470[17] = buffer_data_1[3767:3760] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_470[18] = buffer_data_1[3775:3768] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_470[19] = buffer_data_1[3783:3776] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_470[20] = buffer_data_0[3751:3744] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_470[21] = buffer_data_0[3759:3752] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_470[22] = buffer_data_0[3767:3760] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_470[23] = buffer_data_0[3775:3768] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_470[24] = buffer_data_0[3783:3776] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_470 = kernel_img_mul_470[0] + kernel_img_mul_470[1] + kernel_img_mul_470[2] + 
                kernel_img_mul_470[3] + kernel_img_mul_470[4] + kernel_img_mul_470[5] + 
                kernel_img_mul_470[6] + kernel_img_mul_470[7] + kernel_img_mul_470[8] + 
                kernel_img_mul_470[9] + kernel_img_mul_470[10] + kernel_img_mul_470[11] + 
                kernel_img_mul_470[12] + kernel_img_mul_470[13] + kernel_img_mul_470[14] + 
                kernel_img_mul_470[15] + kernel_img_mul_470[16] + kernel_img_mul_470[17] + 
                kernel_img_mul_470[18] + kernel_img_mul_470[19] + kernel_img_mul_470[20] + 
                kernel_img_mul_470[21] + kernel_img_mul_470[22] + kernel_img_mul_470[23] + 
                kernel_img_mul_470[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3767:3760] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3767:3760] <= kernel_img_sum_470[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3767:3760] <= 'd0;
end

wire  [39:0]  kernel_img_mul_471[0:24];
assign kernel_img_mul_471[0] = buffer_data_4[3759:3752] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_471[1] = buffer_data_4[3767:3760] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_471[2] = buffer_data_4[3775:3768] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_471[3] = buffer_data_4[3783:3776] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_471[4] = buffer_data_4[3791:3784] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_471[5] = buffer_data_3[3759:3752] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_471[6] = buffer_data_3[3767:3760] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_471[7] = buffer_data_3[3775:3768] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_471[8] = buffer_data_3[3783:3776] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_471[9] = buffer_data_3[3791:3784] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_471[10] = buffer_data_2[3759:3752] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_471[11] = buffer_data_2[3767:3760] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_471[12] = buffer_data_2[3775:3768] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_471[13] = buffer_data_2[3783:3776] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_471[14] = buffer_data_2[3791:3784] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_471[15] = buffer_data_1[3759:3752] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_471[16] = buffer_data_1[3767:3760] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_471[17] = buffer_data_1[3775:3768] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_471[18] = buffer_data_1[3783:3776] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_471[19] = buffer_data_1[3791:3784] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_471[20] = buffer_data_0[3759:3752] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_471[21] = buffer_data_0[3767:3760] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_471[22] = buffer_data_0[3775:3768] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_471[23] = buffer_data_0[3783:3776] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_471[24] = buffer_data_0[3791:3784] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_471 = kernel_img_mul_471[0] + kernel_img_mul_471[1] + kernel_img_mul_471[2] + 
                kernel_img_mul_471[3] + kernel_img_mul_471[4] + kernel_img_mul_471[5] + 
                kernel_img_mul_471[6] + kernel_img_mul_471[7] + kernel_img_mul_471[8] + 
                kernel_img_mul_471[9] + kernel_img_mul_471[10] + kernel_img_mul_471[11] + 
                kernel_img_mul_471[12] + kernel_img_mul_471[13] + kernel_img_mul_471[14] + 
                kernel_img_mul_471[15] + kernel_img_mul_471[16] + kernel_img_mul_471[17] + 
                kernel_img_mul_471[18] + kernel_img_mul_471[19] + kernel_img_mul_471[20] + 
                kernel_img_mul_471[21] + kernel_img_mul_471[22] + kernel_img_mul_471[23] + 
                kernel_img_mul_471[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3775:3768] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3775:3768] <= kernel_img_sum_471[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3775:3768] <= 'd0;
end

wire  [39:0]  kernel_img_mul_472[0:24];
assign kernel_img_mul_472[0] = buffer_data_4[3767:3760] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_472[1] = buffer_data_4[3775:3768] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_472[2] = buffer_data_4[3783:3776] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_472[3] = buffer_data_4[3791:3784] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_472[4] = buffer_data_4[3799:3792] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_472[5] = buffer_data_3[3767:3760] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_472[6] = buffer_data_3[3775:3768] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_472[7] = buffer_data_3[3783:3776] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_472[8] = buffer_data_3[3791:3784] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_472[9] = buffer_data_3[3799:3792] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_472[10] = buffer_data_2[3767:3760] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_472[11] = buffer_data_2[3775:3768] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_472[12] = buffer_data_2[3783:3776] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_472[13] = buffer_data_2[3791:3784] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_472[14] = buffer_data_2[3799:3792] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_472[15] = buffer_data_1[3767:3760] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_472[16] = buffer_data_1[3775:3768] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_472[17] = buffer_data_1[3783:3776] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_472[18] = buffer_data_1[3791:3784] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_472[19] = buffer_data_1[3799:3792] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_472[20] = buffer_data_0[3767:3760] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_472[21] = buffer_data_0[3775:3768] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_472[22] = buffer_data_0[3783:3776] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_472[23] = buffer_data_0[3791:3784] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_472[24] = buffer_data_0[3799:3792] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_472 = kernel_img_mul_472[0] + kernel_img_mul_472[1] + kernel_img_mul_472[2] + 
                kernel_img_mul_472[3] + kernel_img_mul_472[4] + kernel_img_mul_472[5] + 
                kernel_img_mul_472[6] + kernel_img_mul_472[7] + kernel_img_mul_472[8] + 
                kernel_img_mul_472[9] + kernel_img_mul_472[10] + kernel_img_mul_472[11] + 
                kernel_img_mul_472[12] + kernel_img_mul_472[13] + kernel_img_mul_472[14] + 
                kernel_img_mul_472[15] + kernel_img_mul_472[16] + kernel_img_mul_472[17] + 
                kernel_img_mul_472[18] + kernel_img_mul_472[19] + kernel_img_mul_472[20] + 
                kernel_img_mul_472[21] + kernel_img_mul_472[22] + kernel_img_mul_472[23] + 
                kernel_img_mul_472[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3783:3776] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3783:3776] <= kernel_img_sum_472[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3783:3776] <= 'd0;
end

wire  [39:0]  kernel_img_mul_473[0:24];
assign kernel_img_mul_473[0] = buffer_data_4[3775:3768] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_473[1] = buffer_data_4[3783:3776] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_473[2] = buffer_data_4[3791:3784] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_473[3] = buffer_data_4[3799:3792] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_473[4] = buffer_data_4[3807:3800] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_473[5] = buffer_data_3[3775:3768] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_473[6] = buffer_data_3[3783:3776] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_473[7] = buffer_data_3[3791:3784] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_473[8] = buffer_data_3[3799:3792] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_473[9] = buffer_data_3[3807:3800] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_473[10] = buffer_data_2[3775:3768] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_473[11] = buffer_data_2[3783:3776] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_473[12] = buffer_data_2[3791:3784] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_473[13] = buffer_data_2[3799:3792] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_473[14] = buffer_data_2[3807:3800] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_473[15] = buffer_data_1[3775:3768] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_473[16] = buffer_data_1[3783:3776] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_473[17] = buffer_data_1[3791:3784] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_473[18] = buffer_data_1[3799:3792] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_473[19] = buffer_data_1[3807:3800] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_473[20] = buffer_data_0[3775:3768] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_473[21] = buffer_data_0[3783:3776] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_473[22] = buffer_data_0[3791:3784] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_473[23] = buffer_data_0[3799:3792] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_473[24] = buffer_data_0[3807:3800] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_473 = kernel_img_mul_473[0] + kernel_img_mul_473[1] + kernel_img_mul_473[2] + 
                kernel_img_mul_473[3] + kernel_img_mul_473[4] + kernel_img_mul_473[5] + 
                kernel_img_mul_473[6] + kernel_img_mul_473[7] + kernel_img_mul_473[8] + 
                kernel_img_mul_473[9] + kernel_img_mul_473[10] + kernel_img_mul_473[11] + 
                kernel_img_mul_473[12] + kernel_img_mul_473[13] + kernel_img_mul_473[14] + 
                kernel_img_mul_473[15] + kernel_img_mul_473[16] + kernel_img_mul_473[17] + 
                kernel_img_mul_473[18] + kernel_img_mul_473[19] + kernel_img_mul_473[20] + 
                kernel_img_mul_473[21] + kernel_img_mul_473[22] + kernel_img_mul_473[23] + 
                kernel_img_mul_473[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3791:3784] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3791:3784] <= kernel_img_sum_473[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3791:3784] <= 'd0;
end

wire  [39:0]  kernel_img_mul_474[0:24];
assign kernel_img_mul_474[0] = buffer_data_4[3783:3776] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_474[1] = buffer_data_4[3791:3784] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_474[2] = buffer_data_4[3799:3792] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_474[3] = buffer_data_4[3807:3800] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_474[4] = buffer_data_4[3815:3808] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_474[5] = buffer_data_3[3783:3776] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_474[6] = buffer_data_3[3791:3784] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_474[7] = buffer_data_3[3799:3792] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_474[8] = buffer_data_3[3807:3800] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_474[9] = buffer_data_3[3815:3808] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_474[10] = buffer_data_2[3783:3776] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_474[11] = buffer_data_2[3791:3784] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_474[12] = buffer_data_2[3799:3792] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_474[13] = buffer_data_2[3807:3800] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_474[14] = buffer_data_2[3815:3808] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_474[15] = buffer_data_1[3783:3776] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_474[16] = buffer_data_1[3791:3784] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_474[17] = buffer_data_1[3799:3792] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_474[18] = buffer_data_1[3807:3800] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_474[19] = buffer_data_1[3815:3808] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_474[20] = buffer_data_0[3783:3776] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_474[21] = buffer_data_0[3791:3784] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_474[22] = buffer_data_0[3799:3792] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_474[23] = buffer_data_0[3807:3800] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_474[24] = buffer_data_0[3815:3808] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_474 = kernel_img_mul_474[0] + kernel_img_mul_474[1] + kernel_img_mul_474[2] + 
                kernel_img_mul_474[3] + kernel_img_mul_474[4] + kernel_img_mul_474[5] + 
                kernel_img_mul_474[6] + kernel_img_mul_474[7] + kernel_img_mul_474[8] + 
                kernel_img_mul_474[9] + kernel_img_mul_474[10] + kernel_img_mul_474[11] + 
                kernel_img_mul_474[12] + kernel_img_mul_474[13] + kernel_img_mul_474[14] + 
                kernel_img_mul_474[15] + kernel_img_mul_474[16] + kernel_img_mul_474[17] + 
                kernel_img_mul_474[18] + kernel_img_mul_474[19] + kernel_img_mul_474[20] + 
                kernel_img_mul_474[21] + kernel_img_mul_474[22] + kernel_img_mul_474[23] + 
                kernel_img_mul_474[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3799:3792] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3799:3792] <= kernel_img_sum_474[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3799:3792] <= 'd0;
end

wire  [39:0]  kernel_img_mul_475[0:24];
assign kernel_img_mul_475[0] = buffer_data_4[3791:3784] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_475[1] = buffer_data_4[3799:3792] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_475[2] = buffer_data_4[3807:3800] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_475[3] = buffer_data_4[3815:3808] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_475[4] = buffer_data_4[3823:3816] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_475[5] = buffer_data_3[3791:3784] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_475[6] = buffer_data_3[3799:3792] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_475[7] = buffer_data_3[3807:3800] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_475[8] = buffer_data_3[3815:3808] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_475[9] = buffer_data_3[3823:3816] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_475[10] = buffer_data_2[3791:3784] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_475[11] = buffer_data_2[3799:3792] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_475[12] = buffer_data_2[3807:3800] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_475[13] = buffer_data_2[3815:3808] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_475[14] = buffer_data_2[3823:3816] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_475[15] = buffer_data_1[3791:3784] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_475[16] = buffer_data_1[3799:3792] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_475[17] = buffer_data_1[3807:3800] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_475[18] = buffer_data_1[3815:3808] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_475[19] = buffer_data_1[3823:3816] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_475[20] = buffer_data_0[3791:3784] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_475[21] = buffer_data_0[3799:3792] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_475[22] = buffer_data_0[3807:3800] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_475[23] = buffer_data_0[3815:3808] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_475[24] = buffer_data_0[3823:3816] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_475 = kernel_img_mul_475[0] + kernel_img_mul_475[1] + kernel_img_mul_475[2] + 
                kernel_img_mul_475[3] + kernel_img_mul_475[4] + kernel_img_mul_475[5] + 
                kernel_img_mul_475[6] + kernel_img_mul_475[7] + kernel_img_mul_475[8] + 
                kernel_img_mul_475[9] + kernel_img_mul_475[10] + kernel_img_mul_475[11] + 
                kernel_img_mul_475[12] + kernel_img_mul_475[13] + kernel_img_mul_475[14] + 
                kernel_img_mul_475[15] + kernel_img_mul_475[16] + kernel_img_mul_475[17] + 
                kernel_img_mul_475[18] + kernel_img_mul_475[19] + kernel_img_mul_475[20] + 
                kernel_img_mul_475[21] + kernel_img_mul_475[22] + kernel_img_mul_475[23] + 
                kernel_img_mul_475[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3807:3800] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3807:3800] <= kernel_img_sum_475[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3807:3800] <= 'd0;
end

wire  [39:0]  kernel_img_mul_476[0:24];
assign kernel_img_mul_476[0] = buffer_data_4[3799:3792] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_476[1] = buffer_data_4[3807:3800] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_476[2] = buffer_data_4[3815:3808] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_476[3] = buffer_data_4[3823:3816] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_476[4] = buffer_data_4[3831:3824] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_476[5] = buffer_data_3[3799:3792] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_476[6] = buffer_data_3[3807:3800] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_476[7] = buffer_data_3[3815:3808] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_476[8] = buffer_data_3[3823:3816] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_476[9] = buffer_data_3[3831:3824] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_476[10] = buffer_data_2[3799:3792] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_476[11] = buffer_data_2[3807:3800] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_476[12] = buffer_data_2[3815:3808] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_476[13] = buffer_data_2[3823:3816] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_476[14] = buffer_data_2[3831:3824] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_476[15] = buffer_data_1[3799:3792] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_476[16] = buffer_data_1[3807:3800] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_476[17] = buffer_data_1[3815:3808] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_476[18] = buffer_data_1[3823:3816] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_476[19] = buffer_data_1[3831:3824] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_476[20] = buffer_data_0[3799:3792] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_476[21] = buffer_data_0[3807:3800] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_476[22] = buffer_data_0[3815:3808] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_476[23] = buffer_data_0[3823:3816] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_476[24] = buffer_data_0[3831:3824] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_476 = kernel_img_mul_476[0] + kernel_img_mul_476[1] + kernel_img_mul_476[2] + 
                kernel_img_mul_476[3] + kernel_img_mul_476[4] + kernel_img_mul_476[5] + 
                kernel_img_mul_476[6] + kernel_img_mul_476[7] + kernel_img_mul_476[8] + 
                kernel_img_mul_476[9] + kernel_img_mul_476[10] + kernel_img_mul_476[11] + 
                kernel_img_mul_476[12] + kernel_img_mul_476[13] + kernel_img_mul_476[14] + 
                kernel_img_mul_476[15] + kernel_img_mul_476[16] + kernel_img_mul_476[17] + 
                kernel_img_mul_476[18] + kernel_img_mul_476[19] + kernel_img_mul_476[20] + 
                kernel_img_mul_476[21] + kernel_img_mul_476[22] + kernel_img_mul_476[23] + 
                kernel_img_mul_476[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3815:3808] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3815:3808] <= kernel_img_sum_476[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3815:3808] <= 'd0;
end

wire  [39:0]  kernel_img_mul_477[0:24];
assign kernel_img_mul_477[0] = buffer_data_4[3807:3800] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_477[1] = buffer_data_4[3815:3808] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_477[2] = buffer_data_4[3823:3816] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_477[3] = buffer_data_4[3831:3824] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_477[4] = buffer_data_4[3839:3832] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_477[5] = buffer_data_3[3807:3800] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_477[6] = buffer_data_3[3815:3808] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_477[7] = buffer_data_3[3823:3816] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_477[8] = buffer_data_3[3831:3824] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_477[9] = buffer_data_3[3839:3832] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_477[10] = buffer_data_2[3807:3800] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_477[11] = buffer_data_2[3815:3808] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_477[12] = buffer_data_2[3823:3816] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_477[13] = buffer_data_2[3831:3824] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_477[14] = buffer_data_2[3839:3832] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_477[15] = buffer_data_1[3807:3800] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_477[16] = buffer_data_1[3815:3808] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_477[17] = buffer_data_1[3823:3816] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_477[18] = buffer_data_1[3831:3824] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_477[19] = buffer_data_1[3839:3832] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_477[20] = buffer_data_0[3807:3800] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_477[21] = buffer_data_0[3815:3808] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_477[22] = buffer_data_0[3823:3816] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_477[23] = buffer_data_0[3831:3824] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_477[24] = buffer_data_0[3839:3832] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_477 = kernel_img_mul_477[0] + kernel_img_mul_477[1] + kernel_img_mul_477[2] + 
                kernel_img_mul_477[3] + kernel_img_mul_477[4] + kernel_img_mul_477[5] + 
                kernel_img_mul_477[6] + kernel_img_mul_477[7] + kernel_img_mul_477[8] + 
                kernel_img_mul_477[9] + kernel_img_mul_477[10] + kernel_img_mul_477[11] + 
                kernel_img_mul_477[12] + kernel_img_mul_477[13] + kernel_img_mul_477[14] + 
                kernel_img_mul_477[15] + kernel_img_mul_477[16] + kernel_img_mul_477[17] + 
                kernel_img_mul_477[18] + kernel_img_mul_477[19] + kernel_img_mul_477[20] + 
                kernel_img_mul_477[21] + kernel_img_mul_477[22] + kernel_img_mul_477[23] + 
                kernel_img_mul_477[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3823:3816] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3823:3816] <= kernel_img_sum_477[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3823:3816] <= 'd0;
end

wire  [39:0]  kernel_img_mul_478[0:24];
assign kernel_img_mul_478[0] = buffer_data_4[3815:3808] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_478[1] = buffer_data_4[3823:3816] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_478[2] = buffer_data_4[3831:3824] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_478[3] = buffer_data_4[3839:3832] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_478[4] = buffer_data_4[3847:3840] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_478[5] = buffer_data_3[3815:3808] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_478[6] = buffer_data_3[3823:3816] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_478[7] = buffer_data_3[3831:3824] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_478[8] = buffer_data_3[3839:3832] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_478[9] = buffer_data_3[3847:3840] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_478[10] = buffer_data_2[3815:3808] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_478[11] = buffer_data_2[3823:3816] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_478[12] = buffer_data_2[3831:3824] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_478[13] = buffer_data_2[3839:3832] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_478[14] = buffer_data_2[3847:3840] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_478[15] = buffer_data_1[3815:3808] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_478[16] = buffer_data_1[3823:3816] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_478[17] = buffer_data_1[3831:3824] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_478[18] = buffer_data_1[3839:3832] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_478[19] = buffer_data_1[3847:3840] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_478[20] = buffer_data_0[3815:3808] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_478[21] = buffer_data_0[3823:3816] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_478[22] = buffer_data_0[3831:3824] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_478[23] = buffer_data_0[3839:3832] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_478[24] = buffer_data_0[3847:3840] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_478 = kernel_img_mul_478[0] + kernel_img_mul_478[1] + kernel_img_mul_478[2] + 
                kernel_img_mul_478[3] + kernel_img_mul_478[4] + kernel_img_mul_478[5] + 
                kernel_img_mul_478[6] + kernel_img_mul_478[7] + kernel_img_mul_478[8] + 
                kernel_img_mul_478[9] + kernel_img_mul_478[10] + kernel_img_mul_478[11] + 
                kernel_img_mul_478[12] + kernel_img_mul_478[13] + kernel_img_mul_478[14] + 
                kernel_img_mul_478[15] + kernel_img_mul_478[16] + kernel_img_mul_478[17] + 
                kernel_img_mul_478[18] + kernel_img_mul_478[19] + kernel_img_mul_478[20] + 
                kernel_img_mul_478[21] + kernel_img_mul_478[22] + kernel_img_mul_478[23] + 
                kernel_img_mul_478[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3831:3824] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3831:3824] <= kernel_img_sum_478[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3831:3824] <= 'd0;
end

wire  [39:0]  kernel_img_mul_479[0:24];
assign kernel_img_mul_479[0] = buffer_data_4[3823:3816] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_479[1] = buffer_data_4[3831:3824] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_479[2] = buffer_data_4[3839:3832] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_479[3] = buffer_data_4[3847:3840] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_479[4] = buffer_data_4[3855:3848] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_479[5] = buffer_data_3[3823:3816] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_479[6] = buffer_data_3[3831:3824] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_479[7] = buffer_data_3[3839:3832] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_479[8] = buffer_data_3[3847:3840] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_479[9] = buffer_data_3[3855:3848] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_479[10] = buffer_data_2[3823:3816] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_479[11] = buffer_data_2[3831:3824] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_479[12] = buffer_data_2[3839:3832] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_479[13] = buffer_data_2[3847:3840] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_479[14] = buffer_data_2[3855:3848] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_479[15] = buffer_data_1[3823:3816] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_479[16] = buffer_data_1[3831:3824] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_479[17] = buffer_data_1[3839:3832] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_479[18] = buffer_data_1[3847:3840] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_479[19] = buffer_data_1[3855:3848] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_479[20] = buffer_data_0[3823:3816] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_479[21] = buffer_data_0[3831:3824] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_479[22] = buffer_data_0[3839:3832] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_479[23] = buffer_data_0[3847:3840] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_479[24] = buffer_data_0[3855:3848] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_479 = kernel_img_mul_479[0] + kernel_img_mul_479[1] + kernel_img_mul_479[2] + 
                kernel_img_mul_479[3] + kernel_img_mul_479[4] + kernel_img_mul_479[5] + 
                kernel_img_mul_479[6] + kernel_img_mul_479[7] + kernel_img_mul_479[8] + 
                kernel_img_mul_479[9] + kernel_img_mul_479[10] + kernel_img_mul_479[11] + 
                kernel_img_mul_479[12] + kernel_img_mul_479[13] + kernel_img_mul_479[14] + 
                kernel_img_mul_479[15] + kernel_img_mul_479[16] + kernel_img_mul_479[17] + 
                kernel_img_mul_479[18] + kernel_img_mul_479[19] + kernel_img_mul_479[20] + 
                kernel_img_mul_479[21] + kernel_img_mul_479[22] + kernel_img_mul_479[23] + 
                kernel_img_mul_479[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3839:3832] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3839:3832] <= kernel_img_sum_479[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3839:3832] <= 'd0;
end

wire  [39:0]  kernel_img_mul_480[0:24];
assign kernel_img_mul_480[0] = buffer_data_4[3831:3824] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_480[1] = buffer_data_4[3839:3832] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_480[2] = buffer_data_4[3847:3840] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_480[3] = buffer_data_4[3855:3848] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_480[4] = buffer_data_4[3863:3856] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_480[5] = buffer_data_3[3831:3824] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_480[6] = buffer_data_3[3839:3832] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_480[7] = buffer_data_3[3847:3840] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_480[8] = buffer_data_3[3855:3848] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_480[9] = buffer_data_3[3863:3856] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_480[10] = buffer_data_2[3831:3824] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_480[11] = buffer_data_2[3839:3832] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_480[12] = buffer_data_2[3847:3840] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_480[13] = buffer_data_2[3855:3848] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_480[14] = buffer_data_2[3863:3856] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_480[15] = buffer_data_1[3831:3824] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_480[16] = buffer_data_1[3839:3832] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_480[17] = buffer_data_1[3847:3840] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_480[18] = buffer_data_1[3855:3848] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_480[19] = buffer_data_1[3863:3856] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_480[20] = buffer_data_0[3831:3824] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_480[21] = buffer_data_0[3839:3832] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_480[22] = buffer_data_0[3847:3840] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_480[23] = buffer_data_0[3855:3848] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_480[24] = buffer_data_0[3863:3856] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_480 = kernel_img_mul_480[0] + kernel_img_mul_480[1] + kernel_img_mul_480[2] + 
                kernel_img_mul_480[3] + kernel_img_mul_480[4] + kernel_img_mul_480[5] + 
                kernel_img_mul_480[6] + kernel_img_mul_480[7] + kernel_img_mul_480[8] + 
                kernel_img_mul_480[9] + kernel_img_mul_480[10] + kernel_img_mul_480[11] + 
                kernel_img_mul_480[12] + kernel_img_mul_480[13] + kernel_img_mul_480[14] + 
                kernel_img_mul_480[15] + kernel_img_mul_480[16] + kernel_img_mul_480[17] + 
                kernel_img_mul_480[18] + kernel_img_mul_480[19] + kernel_img_mul_480[20] + 
                kernel_img_mul_480[21] + kernel_img_mul_480[22] + kernel_img_mul_480[23] + 
                kernel_img_mul_480[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3847:3840] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3847:3840] <= kernel_img_sum_480[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3847:3840] <= 'd0;
end

wire  [39:0]  kernel_img_mul_481[0:24];
assign kernel_img_mul_481[0] = buffer_data_4[3839:3832] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_481[1] = buffer_data_4[3847:3840] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_481[2] = buffer_data_4[3855:3848] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_481[3] = buffer_data_4[3863:3856] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_481[4] = buffer_data_4[3871:3864] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_481[5] = buffer_data_3[3839:3832] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_481[6] = buffer_data_3[3847:3840] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_481[7] = buffer_data_3[3855:3848] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_481[8] = buffer_data_3[3863:3856] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_481[9] = buffer_data_3[3871:3864] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_481[10] = buffer_data_2[3839:3832] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_481[11] = buffer_data_2[3847:3840] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_481[12] = buffer_data_2[3855:3848] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_481[13] = buffer_data_2[3863:3856] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_481[14] = buffer_data_2[3871:3864] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_481[15] = buffer_data_1[3839:3832] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_481[16] = buffer_data_1[3847:3840] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_481[17] = buffer_data_1[3855:3848] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_481[18] = buffer_data_1[3863:3856] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_481[19] = buffer_data_1[3871:3864] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_481[20] = buffer_data_0[3839:3832] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_481[21] = buffer_data_0[3847:3840] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_481[22] = buffer_data_0[3855:3848] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_481[23] = buffer_data_0[3863:3856] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_481[24] = buffer_data_0[3871:3864] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_481 = kernel_img_mul_481[0] + kernel_img_mul_481[1] + kernel_img_mul_481[2] + 
                kernel_img_mul_481[3] + kernel_img_mul_481[4] + kernel_img_mul_481[5] + 
                kernel_img_mul_481[6] + kernel_img_mul_481[7] + kernel_img_mul_481[8] + 
                kernel_img_mul_481[9] + kernel_img_mul_481[10] + kernel_img_mul_481[11] + 
                kernel_img_mul_481[12] + kernel_img_mul_481[13] + kernel_img_mul_481[14] + 
                kernel_img_mul_481[15] + kernel_img_mul_481[16] + kernel_img_mul_481[17] + 
                kernel_img_mul_481[18] + kernel_img_mul_481[19] + kernel_img_mul_481[20] + 
                kernel_img_mul_481[21] + kernel_img_mul_481[22] + kernel_img_mul_481[23] + 
                kernel_img_mul_481[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3855:3848] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3855:3848] <= kernel_img_sum_481[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3855:3848] <= 'd0;
end

wire  [39:0]  kernel_img_mul_482[0:24];
assign kernel_img_mul_482[0] = buffer_data_4[3847:3840] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_482[1] = buffer_data_4[3855:3848] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_482[2] = buffer_data_4[3863:3856] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_482[3] = buffer_data_4[3871:3864] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_482[4] = buffer_data_4[3879:3872] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_482[5] = buffer_data_3[3847:3840] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_482[6] = buffer_data_3[3855:3848] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_482[7] = buffer_data_3[3863:3856] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_482[8] = buffer_data_3[3871:3864] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_482[9] = buffer_data_3[3879:3872] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_482[10] = buffer_data_2[3847:3840] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_482[11] = buffer_data_2[3855:3848] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_482[12] = buffer_data_2[3863:3856] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_482[13] = buffer_data_2[3871:3864] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_482[14] = buffer_data_2[3879:3872] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_482[15] = buffer_data_1[3847:3840] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_482[16] = buffer_data_1[3855:3848] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_482[17] = buffer_data_1[3863:3856] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_482[18] = buffer_data_1[3871:3864] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_482[19] = buffer_data_1[3879:3872] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_482[20] = buffer_data_0[3847:3840] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_482[21] = buffer_data_0[3855:3848] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_482[22] = buffer_data_0[3863:3856] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_482[23] = buffer_data_0[3871:3864] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_482[24] = buffer_data_0[3879:3872] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_482 = kernel_img_mul_482[0] + kernel_img_mul_482[1] + kernel_img_mul_482[2] + 
                kernel_img_mul_482[3] + kernel_img_mul_482[4] + kernel_img_mul_482[5] + 
                kernel_img_mul_482[6] + kernel_img_mul_482[7] + kernel_img_mul_482[8] + 
                kernel_img_mul_482[9] + kernel_img_mul_482[10] + kernel_img_mul_482[11] + 
                kernel_img_mul_482[12] + kernel_img_mul_482[13] + kernel_img_mul_482[14] + 
                kernel_img_mul_482[15] + kernel_img_mul_482[16] + kernel_img_mul_482[17] + 
                kernel_img_mul_482[18] + kernel_img_mul_482[19] + kernel_img_mul_482[20] + 
                kernel_img_mul_482[21] + kernel_img_mul_482[22] + kernel_img_mul_482[23] + 
                kernel_img_mul_482[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3863:3856] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3863:3856] <= kernel_img_sum_482[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3863:3856] <= 'd0;
end

wire  [39:0]  kernel_img_mul_483[0:24];
assign kernel_img_mul_483[0] = buffer_data_4[3855:3848] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_483[1] = buffer_data_4[3863:3856] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_483[2] = buffer_data_4[3871:3864] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_483[3] = buffer_data_4[3879:3872] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_483[4] = buffer_data_4[3887:3880] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_483[5] = buffer_data_3[3855:3848] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_483[6] = buffer_data_3[3863:3856] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_483[7] = buffer_data_3[3871:3864] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_483[8] = buffer_data_3[3879:3872] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_483[9] = buffer_data_3[3887:3880] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_483[10] = buffer_data_2[3855:3848] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_483[11] = buffer_data_2[3863:3856] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_483[12] = buffer_data_2[3871:3864] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_483[13] = buffer_data_2[3879:3872] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_483[14] = buffer_data_2[3887:3880] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_483[15] = buffer_data_1[3855:3848] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_483[16] = buffer_data_1[3863:3856] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_483[17] = buffer_data_1[3871:3864] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_483[18] = buffer_data_1[3879:3872] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_483[19] = buffer_data_1[3887:3880] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_483[20] = buffer_data_0[3855:3848] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_483[21] = buffer_data_0[3863:3856] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_483[22] = buffer_data_0[3871:3864] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_483[23] = buffer_data_0[3879:3872] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_483[24] = buffer_data_0[3887:3880] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_483 = kernel_img_mul_483[0] + kernel_img_mul_483[1] + kernel_img_mul_483[2] + 
                kernel_img_mul_483[3] + kernel_img_mul_483[4] + kernel_img_mul_483[5] + 
                kernel_img_mul_483[6] + kernel_img_mul_483[7] + kernel_img_mul_483[8] + 
                kernel_img_mul_483[9] + kernel_img_mul_483[10] + kernel_img_mul_483[11] + 
                kernel_img_mul_483[12] + kernel_img_mul_483[13] + kernel_img_mul_483[14] + 
                kernel_img_mul_483[15] + kernel_img_mul_483[16] + kernel_img_mul_483[17] + 
                kernel_img_mul_483[18] + kernel_img_mul_483[19] + kernel_img_mul_483[20] + 
                kernel_img_mul_483[21] + kernel_img_mul_483[22] + kernel_img_mul_483[23] + 
                kernel_img_mul_483[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3871:3864] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3871:3864] <= kernel_img_sum_483[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3871:3864] <= 'd0;
end

wire  [39:0]  kernel_img_mul_484[0:24];
assign kernel_img_mul_484[0] = buffer_data_4[3863:3856] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_484[1] = buffer_data_4[3871:3864] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_484[2] = buffer_data_4[3879:3872] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_484[3] = buffer_data_4[3887:3880] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_484[4] = buffer_data_4[3895:3888] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_484[5] = buffer_data_3[3863:3856] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_484[6] = buffer_data_3[3871:3864] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_484[7] = buffer_data_3[3879:3872] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_484[8] = buffer_data_3[3887:3880] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_484[9] = buffer_data_3[3895:3888] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_484[10] = buffer_data_2[3863:3856] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_484[11] = buffer_data_2[3871:3864] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_484[12] = buffer_data_2[3879:3872] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_484[13] = buffer_data_2[3887:3880] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_484[14] = buffer_data_2[3895:3888] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_484[15] = buffer_data_1[3863:3856] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_484[16] = buffer_data_1[3871:3864] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_484[17] = buffer_data_1[3879:3872] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_484[18] = buffer_data_1[3887:3880] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_484[19] = buffer_data_1[3895:3888] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_484[20] = buffer_data_0[3863:3856] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_484[21] = buffer_data_0[3871:3864] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_484[22] = buffer_data_0[3879:3872] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_484[23] = buffer_data_0[3887:3880] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_484[24] = buffer_data_0[3895:3888] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_484 = kernel_img_mul_484[0] + kernel_img_mul_484[1] + kernel_img_mul_484[2] + 
                kernel_img_mul_484[3] + kernel_img_mul_484[4] + kernel_img_mul_484[5] + 
                kernel_img_mul_484[6] + kernel_img_mul_484[7] + kernel_img_mul_484[8] + 
                kernel_img_mul_484[9] + kernel_img_mul_484[10] + kernel_img_mul_484[11] + 
                kernel_img_mul_484[12] + kernel_img_mul_484[13] + kernel_img_mul_484[14] + 
                kernel_img_mul_484[15] + kernel_img_mul_484[16] + kernel_img_mul_484[17] + 
                kernel_img_mul_484[18] + kernel_img_mul_484[19] + kernel_img_mul_484[20] + 
                kernel_img_mul_484[21] + kernel_img_mul_484[22] + kernel_img_mul_484[23] + 
                kernel_img_mul_484[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3879:3872] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3879:3872] <= kernel_img_sum_484[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3879:3872] <= 'd0;
end

wire  [39:0]  kernel_img_mul_485[0:24];
assign kernel_img_mul_485[0] = buffer_data_4[3871:3864] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_485[1] = buffer_data_4[3879:3872] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_485[2] = buffer_data_4[3887:3880] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_485[3] = buffer_data_4[3895:3888] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_485[4] = buffer_data_4[3903:3896] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_485[5] = buffer_data_3[3871:3864] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_485[6] = buffer_data_3[3879:3872] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_485[7] = buffer_data_3[3887:3880] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_485[8] = buffer_data_3[3895:3888] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_485[9] = buffer_data_3[3903:3896] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_485[10] = buffer_data_2[3871:3864] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_485[11] = buffer_data_2[3879:3872] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_485[12] = buffer_data_2[3887:3880] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_485[13] = buffer_data_2[3895:3888] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_485[14] = buffer_data_2[3903:3896] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_485[15] = buffer_data_1[3871:3864] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_485[16] = buffer_data_1[3879:3872] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_485[17] = buffer_data_1[3887:3880] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_485[18] = buffer_data_1[3895:3888] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_485[19] = buffer_data_1[3903:3896] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_485[20] = buffer_data_0[3871:3864] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_485[21] = buffer_data_0[3879:3872] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_485[22] = buffer_data_0[3887:3880] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_485[23] = buffer_data_0[3895:3888] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_485[24] = buffer_data_0[3903:3896] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_485 = kernel_img_mul_485[0] + kernel_img_mul_485[1] + kernel_img_mul_485[2] + 
                kernel_img_mul_485[3] + kernel_img_mul_485[4] + kernel_img_mul_485[5] + 
                kernel_img_mul_485[6] + kernel_img_mul_485[7] + kernel_img_mul_485[8] + 
                kernel_img_mul_485[9] + kernel_img_mul_485[10] + kernel_img_mul_485[11] + 
                kernel_img_mul_485[12] + kernel_img_mul_485[13] + kernel_img_mul_485[14] + 
                kernel_img_mul_485[15] + kernel_img_mul_485[16] + kernel_img_mul_485[17] + 
                kernel_img_mul_485[18] + kernel_img_mul_485[19] + kernel_img_mul_485[20] + 
                kernel_img_mul_485[21] + kernel_img_mul_485[22] + kernel_img_mul_485[23] + 
                kernel_img_mul_485[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3887:3880] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3887:3880] <= kernel_img_sum_485[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3887:3880] <= 'd0;
end

wire  [39:0]  kernel_img_mul_486[0:24];
assign kernel_img_mul_486[0] = buffer_data_4[3879:3872] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_486[1] = buffer_data_4[3887:3880] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_486[2] = buffer_data_4[3895:3888] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_486[3] = buffer_data_4[3903:3896] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_486[4] = buffer_data_4[3911:3904] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_486[5] = buffer_data_3[3879:3872] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_486[6] = buffer_data_3[3887:3880] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_486[7] = buffer_data_3[3895:3888] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_486[8] = buffer_data_3[3903:3896] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_486[9] = buffer_data_3[3911:3904] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_486[10] = buffer_data_2[3879:3872] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_486[11] = buffer_data_2[3887:3880] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_486[12] = buffer_data_2[3895:3888] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_486[13] = buffer_data_2[3903:3896] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_486[14] = buffer_data_2[3911:3904] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_486[15] = buffer_data_1[3879:3872] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_486[16] = buffer_data_1[3887:3880] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_486[17] = buffer_data_1[3895:3888] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_486[18] = buffer_data_1[3903:3896] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_486[19] = buffer_data_1[3911:3904] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_486[20] = buffer_data_0[3879:3872] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_486[21] = buffer_data_0[3887:3880] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_486[22] = buffer_data_0[3895:3888] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_486[23] = buffer_data_0[3903:3896] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_486[24] = buffer_data_0[3911:3904] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_486 = kernel_img_mul_486[0] + kernel_img_mul_486[1] + kernel_img_mul_486[2] + 
                kernel_img_mul_486[3] + kernel_img_mul_486[4] + kernel_img_mul_486[5] + 
                kernel_img_mul_486[6] + kernel_img_mul_486[7] + kernel_img_mul_486[8] + 
                kernel_img_mul_486[9] + kernel_img_mul_486[10] + kernel_img_mul_486[11] + 
                kernel_img_mul_486[12] + kernel_img_mul_486[13] + kernel_img_mul_486[14] + 
                kernel_img_mul_486[15] + kernel_img_mul_486[16] + kernel_img_mul_486[17] + 
                kernel_img_mul_486[18] + kernel_img_mul_486[19] + kernel_img_mul_486[20] + 
                kernel_img_mul_486[21] + kernel_img_mul_486[22] + kernel_img_mul_486[23] + 
                kernel_img_mul_486[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3895:3888] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3895:3888] <= kernel_img_sum_486[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3895:3888] <= 'd0;
end

wire  [39:0]  kernel_img_mul_487[0:24];
assign kernel_img_mul_487[0] = buffer_data_4[3887:3880] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_487[1] = buffer_data_4[3895:3888] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_487[2] = buffer_data_4[3903:3896] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_487[3] = buffer_data_4[3911:3904] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_487[4] = buffer_data_4[3919:3912] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_487[5] = buffer_data_3[3887:3880] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_487[6] = buffer_data_3[3895:3888] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_487[7] = buffer_data_3[3903:3896] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_487[8] = buffer_data_3[3911:3904] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_487[9] = buffer_data_3[3919:3912] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_487[10] = buffer_data_2[3887:3880] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_487[11] = buffer_data_2[3895:3888] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_487[12] = buffer_data_2[3903:3896] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_487[13] = buffer_data_2[3911:3904] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_487[14] = buffer_data_2[3919:3912] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_487[15] = buffer_data_1[3887:3880] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_487[16] = buffer_data_1[3895:3888] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_487[17] = buffer_data_1[3903:3896] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_487[18] = buffer_data_1[3911:3904] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_487[19] = buffer_data_1[3919:3912] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_487[20] = buffer_data_0[3887:3880] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_487[21] = buffer_data_0[3895:3888] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_487[22] = buffer_data_0[3903:3896] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_487[23] = buffer_data_0[3911:3904] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_487[24] = buffer_data_0[3919:3912] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_487 = kernel_img_mul_487[0] + kernel_img_mul_487[1] + kernel_img_mul_487[2] + 
                kernel_img_mul_487[3] + kernel_img_mul_487[4] + kernel_img_mul_487[5] + 
                kernel_img_mul_487[6] + kernel_img_mul_487[7] + kernel_img_mul_487[8] + 
                kernel_img_mul_487[9] + kernel_img_mul_487[10] + kernel_img_mul_487[11] + 
                kernel_img_mul_487[12] + kernel_img_mul_487[13] + kernel_img_mul_487[14] + 
                kernel_img_mul_487[15] + kernel_img_mul_487[16] + kernel_img_mul_487[17] + 
                kernel_img_mul_487[18] + kernel_img_mul_487[19] + kernel_img_mul_487[20] + 
                kernel_img_mul_487[21] + kernel_img_mul_487[22] + kernel_img_mul_487[23] + 
                kernel_img_mul_487[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3903:3896] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3903:3896] <= kernel_img_sum_487[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3903:3896] <= 'd0;
end

wire  [39:0]  kernel_img_mul_488[0:24];
assign kernel_img_mul_488[0] = buffer_data_4[3895:3888] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_488[1] = buffer_data_4[3903:3896] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_488[2] = buffer_data_4[3911:3904] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_488[3] = buffer_data_4[3919:3912] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_488[4] = buffer_data_4[3927:3920] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_488[5] = buffer_data_3[3895:3888] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_488[6] = buffer_data_3[3903:3896] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_488[7] = buffer_data_3[3911:3904] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_488[8] = buffer_data_3[3919:3912] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_488[9] = buffer_data_3[3927:3920] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_488[10] = buffer_data_2[3895:3888] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_488[11] = buffer_data_2[3903:3896] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_488[12] = buffer_data_2[3911:3904] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_488[13] = buffer_data_2[3919:3912] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_488[14] = buffer_data_2[3927:3920] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_488[15] = buffer_data_1[3895:3888] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_488[16] = buffer_data_1[3903:3896] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_488[17] = buffer_data_1[3911:3904] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_488[18] = buffer_data_1[3919:3912] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_488[19] = buffer_data_1[3927:3920] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_488[20] = buffer_data_0[3895:3888] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_488[21] = buffer_data_0[3903:3896] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_488[22] = buffer_data_0[3911:3904] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_488[23] = buffer_data_0[3919:3912] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_488[24] = buffer_data_0[3927:3920] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_488 = kernel_img_mul_488[0] + kernel_img_mul_488[1] + kernel_img_mul_488[2] + 
                kernel_img_mul_488[3] + kernel_img_mul_488[4] + kernel_img_mul_488[5] + 
                kernel_img_mul_488[6] + kernel_img_mul_488[7] + kernel_img_mul_488[8] + 
                kernel_img_mul_488[9] + kernel_img_mul_488[10] + kernel_img_mul_488[11] + 
                kernel_img_mul_488[12] + kernel_img_mul_488[13] + kernel_img_mul_488[14] + 
                kernel_img_mul_488[15] + kernel_img_mul_488[16] + kernel_img_mul_488[17] + 
                kernel_img_mul_488[18] + kernel_img_mul_488[19] + kernel_img_mul_488[20] + 
                kernel_img_mul_488[21] + kernel_img_mul_488[22] + kernel_img_mul_488[23] + 
                kernel_img_mul_488[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3911:3904] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3911:3904] <= kernel_img_sum_488[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3911:3904] <= 'd0;
end

wire  [39:0]  kernel_img_mul_489[0:24];
assign kernel_img_mul_489[0] = buffer_data_4[3903:3896] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_489[1] = buffer_data_4[3911:3904] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_489[2] = buffer_data_4[3919:3912] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_489[3] = buffer_data_4[3927:3920] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_489[4] = buffer_data_4[3935:3928] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_489[5] = buffer_data_3[3903:3896] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_489[6] = buffer_data_3[3911:3904] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_489[7] = buffer_data_3[3919:3912] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_489[8] = buffer_data_3[3927:3920] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_489[9] = buffer_data_3[3935:3928] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_489[10] = buffer_data_2[3903:3896] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_489[11] = buffer_data_2[3911:3904] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_489[12] = buffer_data_2[3919:3912] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_489[13] = buffer_data_2[3927:3920] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_489[14] = buffer_data_2[3935:3928] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_489[15] = buffer_data_1[3903:3896] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_489[16] = buffer_data_1[3911:3904] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_489[17] = buffer_data_1[3919:3912] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_489[18] = buffer_data_1[3927:3920] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_489[19] = buffer_data_1[3935:3928] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_489[20] = buffer_data_0[3903:3896] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_489[21] = buffer_data_0[3911:3904] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_489[22] = buffer_data_0[3919:3912] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_489[23] = buffer_data_0[3927:3920] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_489[24] = buffer_data_0[3935:3928] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_489 = kernel_img_mul_489[0] + kernel_img_mul_489[1] + kernel_img_mul_489[2] + 
                kernel_img_mul_489[3] + kernel_img_mul_489[4] + kernel_img_mul_489[5] + 
                kernel_img_mul_489[6] + kernel_img_mul_489[7] + kernel_img_mul_489[8] + 
                kernel_img_mul_489[9] + kernel_img_mul_489[10] + kernel_img_mul_489[11] + 
                kernel_img_mul_489[12] + kernel_img_mul_489[13] + kernel_img_mul_489[14] + 
                kernel_img_mul_489[15] + kernel_img_mul_489[16] + kernel_img_mul_489[17] + 
                kernel_img_mul_489[18] + kernel_img_mul_489[19] + kernel_img_mul_489[20] + 
                kernel_img_mul_489[21] + kernel_img_mul_489[22] + kernel_img_mul_489[23] + 
                kernel_img_mul_489[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3919:3912] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3919:3912] <= kernel_img_sum_489[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3919:3912] <= 'd0;
end

wire  [39:0]  kernel_img_mul_490[0:24];
assign kernel_img_mul_490[0] = buffer_data_4[3911:3904] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_490[1] = buffer_data_4[3919:3912] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_490[2] = buffer_data_4[3927:3920] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_490[3] = buffer_data_4[3935:3928] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_490[4] = buffer_data_4[3943:3936] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_490[5] = buffer_data_3[3911:3904] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_490[6] = buffer_data_3[3919:3912] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_490[7] = buffer_data_3[3927:3920] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_490[8] = buffer_data_3[3935:3928] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_490[9] = buffer_data_3[3943:3936] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_490[10] = buffer_data_2[3911:3904] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_490[11] = buffer_data_2[3919:3912] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_490[12] = buffer_data_2[3927:3920] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_490[13] = buffer_data_2[3935:3928] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_490[14] = buffer_data_2[3943:3936] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_490[15] = buffer_data_1[3911:3904] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_490[16] = buffer_data_1[3919:3912] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_490[17] = buffer_data_1[3927:3920] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_490[18] = buffer_data_1[3935:3928] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_490[19] = buffer_data_1[3943:3936] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_490[20] = buffer_data_0[3911:3904] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_490[21] = buffer_data_0[3919:3912] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_490[22] = buffer_data_0[3927:3920] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_490[23] = buffer_data_0[3935:3928] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_490[24] = buffer_data_0[3943:3936] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_490 = kernel_img_mul_490[0] + kernel_img_mul_490[1] + kernel_img_mul_490[2] + 
                kernel_img_mul_490[3] + kernel_img_mul_490[4] + kernel_img_mul_490[5] + 
                kernel_img_mul_490[6] + kernel_img_mul_490[7] + kernel_img_mul_490[8] + 
                kernel_img_mul_490[9] + kernel_img_mul_490[10] + kernel_img_mul_490[11] + 
                kernel_img_mul_490[12] + kernel_img_mul_490[13] + kernel_img_mul_490[14] + 
                kernel_img_mul_490[15] + kernel_img_mul_490[16] + kernel_img_mul_490[17] + 
                kernel_img_mul_490[18] + kernel_img_mul_490[19] + kernel_img_mul_490[20] + 
                kernel_img_mul_490[21] + kernel_img_mul_490[22] + kernel_img_mul_490[23] + 
                kernel_img_mul_490[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3927:3920] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3927:3920] <= kernel_img_sum_490[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3927:3920] <= 'd0;
end

wire  [39:0]  kernel_img_mul_491[0:24];
assign kernel_img_mul_491[0] = buffer_data_4[3919:3912] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_491[1] = buffer_data_4[3927:3920] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_491[2] = buffer_data_4[3935:3928] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_491[3] = buffer_data_4[3943:3936] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_491[4] = buffer_data_4[3951:3944] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_491[5] = buffer_data_3[3919:3912] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_491[6] = buffer_data_3[3927:3920] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_491[7] = buffer_data_3[3935:3928] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_491[8] = buffer_data_3[3943:3936] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_491[9] = buffer_data_3[3951:3944] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_491[10] = buffer_data_2[3919:3912] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_491[11] = buffer_data_2[3927:3920] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_491[12] = buffer_data_2[3935:3928] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_491[13] = buffer_data_2[3943:3936] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_491[14] = buffer_data_2[3951:3944] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_491[15] = buffer_data_1[3919:3912] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_491[16] = buffer_data_1[3927:3920] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_491[17] = buffer_data_1[3935:3928] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_491[18] = buffer_data_1[3943:3936] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_491[19] = buffer_data_1[3951:3944] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_491[20] = buffer_data_0[3919:3912] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_491[21] = buffer_data_0[3927:3920] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_491[22] = buffer_data_0[3935:3928] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_491[23] = buffer_data_0[3943:3936] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_491[24] = buffer_data_0[3951:3944] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_491 = kernel_img_mul_491[0] + kernel_img_mul_491[1] + kernel_img_mul_491[2] + 
                kernel_img_mul_491[3] + kernel_img_mul_491[4] + kernel_img_mul_491[5] + 
                kernel_img_mul_491[6] + kernel_img_mul_491[7] + kernel_img_mul_491[8] + 
                kernel_img_mul_491[9] + kernel_img_mul_491[10] + kernel_img_mul_491[11] + 
                kernel_img_mul_491[12] + kernel_img_mul_491[13] + kernel_img_mul_491[14] + 
                kernel_img_mul_491[15] + kernel_img_mul_491[16] + kernel_img_mul_491[17] + 
                kernel_img_mul_491[18] + kernel_img_mul_491[19] + kernel_img_mul_491[20] + 
                kernel_img_mul_491[21] + kernel_img_mul_491[22] + kernel_img_mul_491[23] + 
                kernel_img_mul_491[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3935:3928] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3935:3928] <= kernel_img_sum_491[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3935:3928] <= 'd0;
end

wire  [39:0]  kernel_img_mul_492[0:24];
assign kernel_img_mul_492[0] = buffer_data_4[3927:3920] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_492[1] = buffer_data_4[3935:3928] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_492[2] = buffer_data_4[3943:3936] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_492[3] = buffer_data_4[3951:3944] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_492[4] = buffer_data_4[3959:3952] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_492[5] = buffer_data_3[3927:3920] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_492[6] = buffer_data_3[3935:3928] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_492[7] = buffer_data_3[3943:3936] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_492[8] = buffer_data_3[3951:3944] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_492[9] = buffer_data_3[3959:3952] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_492[10] = buffer_data_2[3927:3920] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_492[11] = buffer_data_2[3935:3928] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_492[12] = buffer_data_2[3943:3936] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_492[13] = buffer_data_2[3951:3944] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_492[14] = buffer_data_2[3959:3952] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_492[15] = buffer_data_1[3927:3920] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_492[16] = buffer_data_1[3935:3928] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_492[17] = buffer_data_1[3943:3936] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_492[18] = buffer_data_1[3951:3944] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_492[19] = buffer_data_1[3959:3952] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_492[20] = buffer_data_0[3927:3920] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_492[21] = buffer_data_0[3935:3928] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_492[22] = buffer_data_0[3943:3936] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_492[23] = buffer_data_0[3951:3944] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_492[24] = buffer_data_0[3959:3952] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_492 = kernel_img_mul_492[0] + kernel_img_mul_492[1] + kernel_img_mul_492[2] + 
                kernel_img_mul_492[3] + kernel_img_mul_492[4] + kernel_img_mul_492[5] + 
                kernel_img_mul_492[6] + kernel_img_mul_492[7] + kernel_img_mul_492[8] + 
                kernel_img_mul_492[9] + kernel_img_mul_492[10] + kernel_img_mul_492[11] + 
                kernel_img_mul_492[12] + kernel_img_mul_492[13] + kernel_img_mul_492[14] + 
                kernel_img_mul_492[15] + kernel_img_mul_492[16] + kernel_img_mul_492[17] + 
                kernel_img_mul_492[18] + kernel_img_mul_492[19] + kernel_img_mul_492[20] + 
                kernel_img_mul_492[21] + kernel_img_mul_492[22] + kernel_img_mul_492[23] + 
                kernel_img_mul_492[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3943:3936] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3943:3936] <= kernel_img_sum_492[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3943:3936] <= 'd0;
end

wire  [39:0]  kernel_img_mul_493[0:24];
assign kernel_img_mul_493[0] = buffer_data_4[3935:3928] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_493[1] = buffer_data_4[3943:3936] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_493[2] = buffer_data_4[3951:3944] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_493[3] = buffer_data_4[3959:3952] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_493[4] = buffer_data_4[3967:3960] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_493[5] = buffer_data_3[3935:3928] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_493[6] = buffer_data_3[3943:3936] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_493[7] = buffer_data_3[3951:3944] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_493[8] = buffer_data_3[3959:3952] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_493[9] = buffer_data_3[3967:3960] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_493[10] = buffer_data_2[3935:3928] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_493[11] = buffer_data_2[3943:3936] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_493[12] = buffer_data_2[3951:3944] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_493[13] = buffer_data_2[3959:3952] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_493[14] = buffer_data_2[3967:3960] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_493[15] = buffer_data_1[3935:3928] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_493[16] = buffer_data_1[3943:3936] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_493[17] = buffer_data_1[3951:3944] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_493[18] = buffer_data_1[3959:3952] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_493[19] = buffer_data_1[3967:3960] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_493[20] = buffer_data_0[3935:3928] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_493[21] = buffer_data_0[3943:3936] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_493[22] = buffer_data_0[3951:3944] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_493[23] = buffer_data_0[3959:3952] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_493[24] = buffer_data_0[3967:3960] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_493 = kernel_img_mul_493[0] + kernel_img_mul_493[1] + kernel_img_mul_493[2] + 
                kernel_img_mul_493[3] + kernel_img_mul_493[4] + kernel_img_mul_493[5] + 
                kernel_img_mul_493[6] + kernel_img_mul_493[7] + kernel_img_mul_493[8] + 
                kernel_img_mul_493[9] + kernel_img_mul_493[10] + kernel_img_mul_493[11] + 
                kernel_img_mul_493[12] + kernel_img_mul_493[13] + kernel_img_mul_493[14] + 
                kernel_img_mul_493[15] + kernel_img_mul_493[16] + kernel_img_mul_493[17] + 
                kernel_img_mul_493[18] + kernel_img_mul_493[19] + kernel_img_mul_493[20] + 
                kernel_img_mul_493[21] + kernel_img_mul_493[22] + kernel_img_mul_493[23] + 
                kernel_img_mul_493[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3951:3944] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3951:3944] <= kernel_img_sum_493[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3951:3944] <= 'd0;
end

wire  [39:0]  kernel_img_mul_494[0:24];
assign kernel_img_mul_494[0] = buffer_data_4[3943:3936] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_494[1] = buffer_data_4[3951:3944] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_494[2] = buffer_data_4[3959:3952] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_494[3] = buffer_data_4[3967:3960] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_494[4] = buffer_data_4[3975:3968] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_494[5] = buffer_data_3[3943:3936] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_494[6] = buffer_data_3[3951:3944] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_494[7] = buffer_data_3[3959:3952] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_494[8] = buffer_data_3[3967:3960] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_494[9] = buffer_data_3[3975:3968] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_494[10] = buffer_data_2[3943:3936] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_494[11] = buffer_data_2[3951:3944] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_494[12] = buffer_data_2[3959:3952] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_494[13] = buffer_data_2[3967:3960] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_494[14] = buffer_data_2[3975:3968] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_494[15] = buffer_data_1[3943:3936] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_494[16] = buffer_data_1[3951:3944] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_494[17] = buffer_data_1[3959:3952] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_494[18] = buffer_data_1[3967:3960] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_494[19] = buffer_data_1[3975:3968] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_494[20] = buffer_data_0[3943:3936] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_494[21] = buffer_data_0[3951:3944] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_494[22] = buffer_data_0[3959:3952] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_494[23] = buffer_data_0[3967:3960] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_494[24] = buffer_data_0[3975:3968] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_494 = kernel_img_mul_494[0] + kernel_img_mul_494[1] + kernel_img_mul_494[2] + 
                kernel_img_mul_494[3] + kernel_img_mul_494[4] + kernel_img_mul_494[5] + 
                kernel_img_mul_494[6] + kernel_img_mul_494[7] + kernel_img_mul_494[8] + 
                kernel_img_mul_494[9] + kernel_img_mul_494[10] + kernel_img_mul_494[11] + 
                kernel_img_mul_494[12] + kernel_img_mul_494[13] + kernel_img_mul_494[14] + 
                kernel_img_mul_494[15] + kernel_img_mul_494[16] + kernel_img_mul_494[17] + 
                kernel_img_mul_494[18] + kernel_img_mul_494[19] + kernel_img_mul_494[20] + 
                kernel_img_mul_494[21] + kernel_img_mul_494[22] + kernel_img_mul_494[23] + 
                kernel_img_mul_494[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3959:3952] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3959:3952] <= kernel_img_sum_494[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3959:3952] <= 'd0;
end

wire  [39:0]  kernel_img_mul_495[0:24];
assign kernel_img_mul_495[0] = buffer_data_4[3951:3944] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_495[1] = buffer_data_4[3959:3952] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_495[2] = buffer_data_4[3967:3960] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_495[3] = buffer_data_4[3975:3968] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_495[4] = buffer_data_4[3983:3976] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_495[5] = buffer_data_3[3951:3944] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_495[6] = buffer_data_3[3959:3952] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_495[7] = buffer_data_3[3967:3960] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_495[8] = buffer_data_3[3975:3968] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_495[9] = buffer_data_3[3983:3976] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_495[10] = buffer_data_2[3951:3944] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_495[11] = buffer_data_2[3959:3952] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_495[12] = buffer_data_2[3967:3960] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_495[13] = buffer_data_2[3975:3968] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_495[14] = buffer_data_2[3983:3976] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_495[15] = buffer_data_1[3951:3944] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_495[16] = buffer_data_1[3959:3952] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_495[17] = buffer_data_1[3967:3960] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_495[18] = buffer_data_1[3975:3968] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_495[19] = buffer_data_1[3983:3976] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_495[20] = buffer_data_0[3951:3944] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_495[21] = buffer_data_0[3959:3952] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_495[22] = buffer_data_0[3967:3960] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_495[23] = buffer_data_0[3975:3968] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_495[24] = buffer_data_0[3983:3976] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_495 = kernel_img_mul_495[0] + kernel_img_mul_495[1] + kernel_img_mul_495[2] + 
                kernel_img_mul_495[3] + kernel_img_mul_495[4] + kernel_img_mul_495[5] + 
                kernel_img_mul_495[6] + kernel_img_mul_495[7] + kernel_img_mul_495[8] + 
                kernel_img_mul_495[9] + kernel_img_mul_495[10] + kernel_img_mul_495[11] + 
                kernel_img_mul_495[12] + kernel_img_mul_495[13] + kernel_img_mul_495[14] + 
                kernel_img_mul_495[15] + kernel_img_mul_495[16] + kernel_img_mul_495[17] + 
                kernel_img_mul_495[18] + kernel_img_mul_495[19] + kernel_img_mul_495[20] + 
                kernel_img_mul_495[21] + kernel_img_mul_495[22] + kernel_img_mul_495[23] + 
                kernel_img_mul_495[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3967:3960] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3967:3960] <= kernel_img_sum_495[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3967:3960] <= 'd0;
end

wire  [39:0]  kernel_img_mul_496[0:24];
assign kernel_img_mul_496[0] = buffer_data_4[3959:3952] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_496[1] = buffer_data_4[3967:3960] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_496[2] = buffer_data_4[3975:3968] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_496[3] = buffer_data_4[3983:3976] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_496[4] = buffer_data_4[3991:3984] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_496[5] = buffer_data_3[3959:3952] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_496[6] = buffer_data_3[3967:3960] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_496[7] = buffer_data_3[3975:3968] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_496[8] = buffer_data_3[3983:3976] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_496[9] = buffer_data_3[3991:3984] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_496[10] = buffer_data_2[3959:3952] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_496[11] = buffer_data_2[3967:3960] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_496[12] = buffer_data_2[3975:3968] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_496[13] = buffer_data_2[3983:3976] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_496[14] = buffer_data_2[3991:3984] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_496[15] = buffer_data_1[3959:3952] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_496[16] = buffer_data_1[3967:3960] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_496[17] = buffer_data_1[3975:3968] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_496[18] = buffer_data_1[3983:3976] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_496[19] = buffer_data_1[3991:3984] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_496[20] = buffer_data_0[3959:3952] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_496[21] = buffer_data_0[3967:3960] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_496[22] = buffer_data_0[3975:3968] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_496[23] = buffer_data_0[3983:3976] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_496[24] = buffer_data_0[3991:3984] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_496 = kernel_img_mul_496[0] + kernel_img_mul_496[1] + kernel_img_mul_496[2] + 
                kernel_img_mul_496[3] + kernel_img_mul_496[4] + kernel_img_mul_496[5] + 
                kernel_img_mul_496[6] + kernel_img_mul_496[7] + kernel_img_mul_496[8] + 
                kernel_img_mul_496[9] + kernel_img_mul_496[10] + kernel_img_mul_496[11] + 
                kernel_img_mul_496[12] + kernel_img_mul_496[13] + kernel_img_mul_496[14] + 
                kernel_img_mul_496[15] + kernel_img_mul_496[16] + kernel_img_mul_496[17] + 
                kernel_img_mul_496[18] + kernel_img_mul_496[19] + kernel_img_mul_496[20] + 
                kernel_img_mul_496[21] + kernel_img_mul_496[22] + kernel_img_mul_496[23] + 
                kernel_img_mul_496[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3975:3968] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3975:3968] <= kernel_img_sum_496[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3975:3968] <= 'd0;
end

wire  [39:0]  kernel_img_mul_497[0:24];
assign kernel_img_mul_497[0] = buffer_data_4[3967:3960] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_497[1] = buffer_data_4[3975:3968] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_497[2] = buffer_data_4[3983:3976] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_497[3] = buffer_data_4[3991:3984] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_497[4] = buffer_data_4[3999:3992] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_497[5] = buffer_data_3[3967:3960] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_497[6] = buffer_data_3[3975:3968] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_497[7] = buffer_data_3[3983:3976] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_497[8] = buffer_data_3[3991:3984] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_497[9] = buffer_data_3[3999:3992] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_497[10] = buffer_data_2[3967:3960] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_497[11] = buffer_data_2[3975:3968] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_497[12] = buffer_data_2[3983:3976] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_497[13] = buffer_data_2[3991:3984] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_497[14] = buffer_data_2[3999:3992] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_497[15] = buffer_data_1[3967:3960] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_497[16] = buffer_data_1[3975:3968] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_497[17] = buffer_data_1[3983:3976] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_497[18] = buffer_data_1[3991:3984] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_497[19] = buffer_data_1[3999:3992] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_497[20] = buffer_data_0[3967:3960] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_497[21] = buffer_data_0[3975:3968] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_497[22] = buffer_data_0[3983:3976] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_497[23] = buffer_data_0[3991:3984] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_497[24] = buffer_data_0[3999:3992] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_497 = kernel_img_mul_497[0] + kernel_img_mul_497[1] + kernel_img_mul_497[2] + 
                kernel_img_mul_497[3] + kernel_img_mul_497[4] + kernel_img_mul_497[5] + 
                kernel_img_mul_497[6] + kernel_img_mul_497[7] + kernel_img_mul_497[8] + 
                kernel_img_mul_497[9] + kernel_img_mul_497[10] + kernel_img_mul_497[11] + 
                kernel_img_mul_497[12] + kernel_img_mul_497[13] + kernel_img_mul_497[14] + 
                kernel_img_mul_497[15] + kernel_img_mul_497[16] + kernel_img_mul_497[17] + 
                kernel_img_mul_497[18] + kernel_img_mul_497[19] + kernel_img_mul_497[20] + 
                kernel_img_mul_497[21] + kernel_img_mul_497[22] + kernel_img_mul_497[23] + 
                kernel_img_mul_497[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3983:3976] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3983:3976] <= kernel_img_sum_497[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3983:3976] <= 'd0;
end

wire  [39:0]  kernel_img_mul_498[0:24];
assign kernel_img_mul_498[0] = buffer_data_4[3975:3968] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_498[1] = buffer_data_4[3983:3976] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_498[2] = buffer_data_4[3991:3984] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_498[3] = buffer_data_4[3999:3992] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_498[4] = buffer_data_4[4007:4000] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_498[5] = buffer_data_3[3975:3968] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_498[6] = buffer_data_3[3983:3976] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_498[7] = buffer_data_3[3991:3984] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_498[8] = buffer_data_3[3999:3992] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_498[9] = buffer_data_3[4007:4000] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_498[10] = buffer_data_2[3975:3968] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_498[11] = buffer_data_2[3983:3976] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_498[12] = buffer_data_2[3991:3984] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_498[13] = buffer_data_2[3999:3992] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_498[14] = buffer_data_2[4007:4000] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_498[15] = buffer_data_1[3975:3968] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_498[16] = buffer_data_1[3983:3976] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_498[17] = buffer_data_1[3991:3984] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_498[18] = buffer_data_1[3999:3992] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_498[19] = buffer_data_1[4007:4000] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_498[20] = buffer_data_0[3975:3968] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_498[21] = buffer_data_0[3983:3976] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_498[22] = buffer_data_0[3991:3984] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_498[23] = buffer_data_0[3999:3992] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_498[24] = buffer_data_0[4007:4000] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_498 = kernel_img_mul_498[0] + kernel_img_mul_498[1] + kernel_img_mul_498[2] + 
                kernel_img_mul_498[3] + kernel_img_mul_498[4] + kernel_img_mul_498[5] + 
                kernel_img_mul_498[6] + kernel_img_mul_498[7] + kernel_img_mul_498[8] + 
                kernel_img_mul_498[9] + kernel_img_mul_498[10] + kernel_img_mul_498[11] + 
                kernel_img_mul_498[12] + kernel_img_mul_498[13] + kernel_img_mul_498[14] + 
                kernel_img_mul_498[15] + kernel_img_mul_498[16] + kernel_img_mul_498[17] + 
                kernel_img_mul_498[18] + kernel_img_mul_498[19] + kernel_img_mul_498[20] + 
                kernel_img_mul_498[21] + kernel_img_mul_498[22] + kernel_img_mul_498[23] + 
                kernel_img_mul_498[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3991:3984] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3991:3984] <= kernel_img_sum_498[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3991:3984] <= 'd0;
end

wire  [39:0]  kernel_img_mul_499[0:24];
assign kernel_img_mul_499[0] = buffer_data_4[3983:3976] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_499[1] = buffer_data_4[3991:3984] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_499[2] = buffer_data_4[3999:3992] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_499[3] = buffer_data_4[4007:4000] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_499[4] = buffer_data_4[4015:4008] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_499[5] = buffer_data_3[3983:3976] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_499[6] = buffer_data_3[3991:3984] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_499[7] = buffer_data_3[3999:3992] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_499[8] = buffer_data_3[4007:4000] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_499[9] = buffer_data_3[4015:4008] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_499[10] = buffer_data_2[3983:3976] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_499[11] = buffer_data_2[3991:3984] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_499[12] = buffer_data_2[3999:3992] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_499[13] = buffer_data_2[4007:4000] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_499[14] = buffer_data_2[4015:4008] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_499[15] = buffer_data_1[3983:3976] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_499[16] = buffer_data_1[3991:3984] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_499[17] = buffer_data_1[3999:3992] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_499[18] = buffer_data_1[4007:4000] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_499[19] = buffer_data_1[4015:4008] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_499[20] = buffer_data_0[3983:3976] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_499[21] = buffer_data_0[3991:3984] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_499[22] = buffer_data_0[3999:3992] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_499[23] = buffer_data_0[4007:4000] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_499[24] = buffer_data_0[4015:4008] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_499 = kernel_img_mul_499[0] + kernel_img_mul_499[1] + kernel_img_mul_499[2] + 
                kernel_img_mul_499[3] + kernel_img_mul_499[4] + kernel_img_mul_499[5] + 
                kernel_img_mul_499[6] + kernel_img_mul_499[7] + kernel_img_mul_499[8] + 
                kernel_img_mul_499[9] + kernel_img_mul_499[10] + kernel_img_mul_499[11] + 
                kernel_img_mul_499[12] + kernel_img_mul_499[13] + kernel_img_mul_499[14] + 
                kernel_img_mul_499[15] + kernel_img_mul_499[16] + kernel_img_mul_499[17] + 
                kernel_img_mul_499[18] + kernel_img_mul_499[19] + kernel_img_mul_499[20] + 
                kernel_img_mul_499[21] + kernel_img_mul_499[22] + kernel_img_mul_499[23] + 
                kernel_img_mul_499[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[3999:3992] <= 'd0;
  else if (current_state==ST_START)
    blur_din[3999:3992] <= kernel_img_sum_499[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3999:3992] <= 'd0;
end

wire  [39:0]  kernel_img_mul_500[0:24];
assign kernel_img_mul_500[0] = buffer_data_4[3991:3984] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_500[1] = buffer_data_4[3999:3992] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_500[2] = buffer_data_4[4007:4000] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_500[3] = buffer_data_4[4015:4008] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_500[4] = buffer_data_4[4023:4016] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_500[5] = buffer_data_3[3991:3984] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_500[6] = buffer_data_3[3999:3992] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_500[7] = buffer_data_3[4007:4000] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_500[8] = buffer_data_3[4015:4008] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_500[9] = buffer_data_3[4023:4016] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_500[10] = buffer_data_2[3991:3984] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_500[11] = buffer_data_2[3999:3992] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_500[12] = buffer_data_2[4007:4000] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_500[13] = buffer_data_2[4015:4008] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_500[14] = buffer_data_2[4023:4016] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_500[15] = buffer_data_1[3991:3984] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_500[16] = buffer_data_1[3999:3992] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_500[17] = buffer_data_1[4007:4000] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_500[18] = buffer_data_1[4015:4008] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_500[19] = buffer_data_1[4023:4016] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_500[20] = buffer_data_0[3991:3984] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_500[21] = buffer_data_0[3999:3992] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_500[22] = buffer_data_0[4007:4000] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_500[23] = buffer_data_0[4015:4008] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_500[24] = buffer_data_0[4023:4016] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_500 = kernel_img_mul_500[0] + kernel_img_mul_500[1] + kernel_img_mul_500[2] + 
                kernel_img_mul_500[3] + kernel_img_mul_500[4] + kernel_img_mul_500[5] + 
                kernel_img_mul_500[6] + kernel_img_mul_500[7] + kernel_img_mul_500[8] + 
                kernel_img_mul_500[9] + kernel_img_mul_500[10] + kernel_img_mul_500[11] + 
                kernel_img_mul_500[12] + kernel_img_mul_500[13] + kernel_img_mul_500[14] + 
                kernel_img_mul_500[15] + kernel_img_mul_500[16] + kernel_img_mul_500[17] + 
                kernel_img_mul_500[18] + kernel_img_mul_500[19] + kernel_img_mul_500[20] + 
                kernel_img_mul_500[21] + kernel_img_mul_500[22] + kernel_img_mul_500[23] + 
                kernel_img_mul_500[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4007:4000] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4007:4000] <= kernel_img_sum_500[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4007:4000] <= 'd0;
end

wire  [39:0]  kernel_img_mul_501[0:24];
assign kernel_img_mul_501[0] = buffer_data_4[3999:3992] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_501[1] = buffer_data_4[4007:4000] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_501[2] = buffer_data_4[4015:4008] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_501[3] = buffer_data_4[4023:4016] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_501[4] = buffer_data_4[4031:4024] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_501[5] = buffer_data_3[3999:3992] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_501[6] = buffer_data_3[4007:4000] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_501[7] = buffer_data_3[4015:4008] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_501[8] = buffer_data_3[4023:4016] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_501[9] = buffer_data_3[4031:4024] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_501[10] = buffer_data_2[3999:3992] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_501[11] = buffer_data_2[4007:4000] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_501[12] = buffer_data_2[4015:4008] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_501[13] = buffer_data_2[4023:4016] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_501[14] = buffer_data_2[4031:4024] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_501[15] = buffer_data_1[3999:3992] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_501[16] = buffer_data_1[4007:4000] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_501[17] = buffer_data_1[4015:4008] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_501[18] = buffer_data_1[4023:4016] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_501[19] = buffer_data_1[4031:4024] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_501[20] = buffer_data_0[3999:3992] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_501[21] = buffer_data_0[4007:4000] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_501[22] = buffer_data_0[4015:4008] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_501[23] = buffer_data_0[4023:4016] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_501[24] = buffer_data_0[4031:4024] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_501 = kernel_img_mul_501[0] + kernel_img_mul_501[1] + kernel_img_mul_501[2] + 
                kernel_img_mul_501[3] + kernel_img_mul_501[4] + kernel_img_mul_501[5] + 
                kernel_img_mul_501[6] + kernel_img_mul_501[7] + kernel_img_mul_501[8] + 
                kernel_img_mul_501[9] + kernel_img_mul_501[10] + kernel_img_mul_501[11] + 
                kernel_img_mul_501[12] + kernel_img_mul_501[13] + kernel_img_mul_501[14] + 
                kernel_img_mul_501[15] + kernel_img_mul_501[16] + kernel_img_mul_501[17] + 
                kernel_img_mul_501[18] + kernel_img_mul_501[19] + kernel_img_mul_501[20] + 
                kernel_img_mul_501[21] + kernel_img_mul_501[22] + kernel_img_mul_501[23] + 
                kernel_img_mul_501[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4015:4008] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4015:4008] <= kernel_img_sum_501[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4015:4008] <= 'd0;
end

wire  [39:0]  kernel_img_mul_502[0:24];
assign kernel_img_mul_502[0] = buffer_data_4[4007:4000] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_502[1] = buffer_data_4[4015:4008] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_502[2] = buffer_data_4[4023:4016] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_502[3] = buffer_data_4[4031:4024] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_502[4] = buffer_data_4[4039:4032] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_502[5] = buffer_data_3[4007:4000] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_502[6] = buffer_data_3[4015:4008] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_502[7] = buffer_data_3[4023:4016] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_502[8] = buffer_data_3[4031:4024] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_502[9] = buffer_data_3[4039:4032] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_502[10] = buffer_data_2[4007:4000] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_502[11] = buffer_data_2[4015:4008] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_502[12] = buffer_data_2[4023:4016] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_502[13] = buffer_data_2[4031:4024] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_502[14] = buffer_data_2[4039:4032] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_502[15] = buffer_data_1[4007:4000] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_502[16] = buffer_data_1[4015:4008] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_502[17] = buffer_data_1[4023:4016] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_502[18] = buffer_data_1[4031:4024] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_502[19] = buffer_data_1[4039:4032] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_502[20] = buffer_data_0[4007:4000] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_502[21] = buffer_data_0[4015:4008] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_502[22] = buffer_data_0[4023:4016] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_502[23] = buffer_data_0[4031:4024] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_502[24] = buffer_data_0[4039:4032] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_502 = kernel_img_mul_502[0] + kernel_img_mul_502[1] + kernel_img_mul_502[2] + 
                kernel_img_mul_502[3] + kernel_img_mul_502[4] + kernel_img_mul_502[5] + 
                kernel_img_mul_502[6] + kernel_img_mul_502[7] + kernel_img_mul_502[8] + 
                kernel_img_mul_502[9] + kernel_img_mul_502[10] + kernel_img_mul_502[11] + 
                kernel_img_mul_502[12] + kernel_img_mul_502[13] + kernel_img_mul_502[14] + 
                kernel_img_mul_502[15] + kernel_img_mul_502[16] + kernel_img_mul_502[17] + 
                kernel_img_mul_502[18] + kernel_img_mul_502[19] + kernel_img_mul_502[20] + 
                kernel_img_mul_502[21] + kernel_img_mul_502[22] + kernel_img_mul_502[23] + 
                kernel_img_mul_502[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4023:4016] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4023:4016] <= kernel_img_sum_502[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4023:4016] <= 'd0;
end

wire  [39:0]  kernel_img_mul_503[0:24];
assign kernel_img_mul_503[0] = buffer_data_4[4015:4008] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_503[1] = buffer_data_4[4023:4016] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_503[2] = buffer_data_4[4031:4024] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_503[3] = buffer_data_4[4039:4032] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_503[4] = buffer_data_4[4047:4040] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_503[5] = buffer_data_3[4015:4008] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_503[6] = buffer_data_3[4023:4016] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_503[7] = buffer_data_3[4031:4024] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_503[8] = buffer_data_3[4039:4032] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_503[9] = buffer_data_3[4047:4040] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_503[10] = buffer_data_2[4015:4008] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_503[11] = buffer_data_2[4023:4016] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_503[12] = buffer_data_2[4031:4024] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_503[13] = buffer_data_2[4039:4032] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_503[14] = buffer_data_2[4047:4040] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_503[15] = buffer_data_1[4015:4008] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_503[16] = buffer_data_1[4023:4016] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_503[17] = buffer_data_1[4031:4024] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_503[18] = buffer_data_1[4039:4032] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_503[19] = buffer_data_1[4047:4040] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_503[20] = buffer_data_0[4015:4008] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_503[21] = buffer_data_0[4023:4016] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_503[22] = buffer_data_0[4031:4024] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_503[23] = buffer_data_0[4039:4032] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_503[24] = buffer_data_0[4047:4040] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_503 = kernel_img_mul_503[0] + kernel_img_mul_503[1] + kernel_img_mul_503[2] + 
                kernel_img_mul_503[3] + kernel_img_mul_503[4] + kernel_img_mul_503[5] + 
                kernel_img_mul_503[6] + kernel_img_mul_503[7] + kernel_img_mul_503[8] + 
                kernel_img_mul_503[9] + kernel_img_mul_503[10] + kernel_img_mul_503[11] + 
                kernel_img_mul_503[12] + kernel_img_mul_503[13] + kernel_img_mul_503[14] + 
                kernel_img_mul_503[15] + kernel_img_mul_503[16] + kernel_img_mul_503[17] + 
                kernel_img_mul_503[18] + kernel_img_mul_503[19] + kernel_img_mul_503[20] + 
                kernel_img_mul_503[21] + kernel_img_mul_503[22] + kernel_img_mul_503[23] + 
                kernel_img_mul_503[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4031:4024] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4031:4024] <= kernel_img_sum_503[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4031:4024] <= 'd0;
end

wire  [39:0]  kernel_img_mul_504[0:24];
assign kernel_img_mul_504[0] = buffer_data_4[4023:4016] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_504[1] = buffer_data_4[4031:4024] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_504[2] = buffer_data_4[4039:4032] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_504[3] = buffer_data_4[4047:4040] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_504[4] = buffer_data_4[4055:4048] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_504[5] = buffer_data_3[4023:4016] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_504[6] = buffer_data_3[4031:4024] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_504[7] = buffer_data_3[4039:4032] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_504[8] = buffer_data_3[4047:4040] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_504[9] = buffer_data_3[4055:4048] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_504[10] = buffer_data_2[4023:4016] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_504[11] = buffer_data_2[4031:4024] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_504[12] = buffer_data_2[4039:4032] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_504[13] = buffer_data_2[4047:4040] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_504[14] = buffer_data_2[4055:4048] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_504[15] = buffer_data_1[4023:4016] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_504[16] = buffer_data_1[4031:4024] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_504[17] = buffer_data_1[4039:4032] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_504[18] = buffer_data_1[4047:4040] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_504[19] = buffer_data_1[4055:4048] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_504[20] = buffer_data_0[4023:4016] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_504[21] = buffer_data_0[4031:4024] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_504[22] = buffer_data_0[4039:4032] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_504[23] = buffer_data_0[4047:4040] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_504[24] = buffer_data_0[4055:4048] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_504 = kernel_img_mul_504[0] + kernel_img_mul_504[1] + kernel_img_mul_504[2] + 
                kernel_img_mul_504[3] + kernel_img_mul_504[4] + kernel_img_mul_504[5] + 
                kernel_img_mul_504[6] + kernel_img_mul_504[7] + kernel_img_mul_504[8] + 
                kernel_img_mul_504[9] + kernel_img_mul_504[10] + kernel_img_mul_504[11] + 
                kernel_img_mul_504[12] + kernel_img_mul_504[13] + kernel_img_mul_504[14] + 
                kernel_img_mul_504[15] + kernel_img_mul_504[16] + kernel_img_mul_504[17] + 
                kernel_img_mul_504[18] + kernel_img_mul_504[19] + kernel_img_mul_504[20] + 
                kernel_img_mul_504[21] + kernel_img_mul_504[22] + kernel_img_mul_504[23] + 
                kernel_img_mul_504[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4039:4032] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4039:4032] <= kernel_img_sum_504[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4039:4032] <= 'd0;
end

wire  [39:0]  kernel_img_mul_505[0:24];
assign kernel_img_mul_505[0] = buffer_data_4[4031:4024] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_505[1] = buffer_data_4[4039:4032] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_505[2] = buffer_data_4[4047:4040] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_505[3] = buffer_data_4[4055:4048] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_505[4] = buffer_data_4[4063:4056] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_505[5] = buffer_data_3[4031:4024] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_505[6] = buffer_data_3[4039:4032] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_505[7] = buffer_data_3[4047:4040] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_505[8] = buffer_data_3[4055:4048] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_505[9] = buffer_data_3[4063:4056] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_505[10] = buffer_data_2[4031:4024] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_505[11] = buffer_data_2[4039:4032] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_505[12] = buffer_data_2[4047:4040] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_505[13] = buffer_data_2[4055:4048] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_505[14] = buffer_data_2[4063:4056] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_505[15] = buffer_data_1[4031:4024] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_505[16] = buffer_data_1[4039:4032] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_505[17] = buffer_data_1[4047:4040] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_505[18] = buffer_data_1[4055:4048] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_505[19] = buffer_data_1[4063:4056] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_505[20] = buffer_data_0[4031:4024] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_505[21] = buffer_data_0[4039:4032] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_505[22] = buffer_data_0[4047:4040] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_505[23] = buffer_data_0[4055:4048] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_505[24] = buffer_data_0[4063:4056] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_505 = kernel_img_mul_505[0] + kernel_img_mul_505[1] + kernel_img_mul_505[2] + 
                kernel_img_mul_505[3] + kernel_img_mul_505[4] + kernel_img_mul_505[5] + 
                kernel_img_mul_505[6] + kernel_img_mul_505[7] + kernel_img_mul_505[8] + 
                kernel_img_mul_505[9] + kernel_img_mul_505[10] + kernel_img_mul_505[11] + 
                kernel_img_mul_505[12] + kernel_img_mul_505[13] + kernel_img_mul_505[14] + 
                kernel_img_mul_505[15] + kernel_img_mul_505[16] + kernel_img_mul_505[17] + 
                kernel_img_mul_505[18] + kernel_img_mul_505[19] + kernel_img_mul_505[20] + 
                kernel_img_mul_505[21] + kernel_img_mul_505[22] + kernel_img_mul_505[23] + 
                kernel_img_mul_505[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4047:4040] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4047:4040] <= kernel_img_sum_505[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4047:4040] <= 'd0;
end

wire  [39:0]  kernel_img_mul_506[0:24];
assign kernel_img_mul_506[0] = buffer_data_4[4039:4032] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_506[1] = buffer_data_4[4047:4040] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_506[2] = buffer_data_4[4055:4048] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_506[3] = buffer_data_4[4063:4056] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_506[4] = buffer_data_4[4071:4064] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_506[5] = buffer_data_3[4039:4032] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_506[6] = buffer_data_3[4047:4040] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_506[7] = buffer_data_3[4055:4048] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_506[8] = buffer_data_3[4063:4056] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_506[9] = buffer_data_3[4071:4064] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_506[10] = buffer_data_2[4039:4032] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_506[11] = buffer_data_2[4047:4040] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_506[12] = buffer_data_2[4055:4048] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_506[13] = buffer_data_2[4063:4056] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_506[14] = buffer_data_2[4071:4064] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_506[15] = buffer_data_1[4039:4032] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_506[16] = buffer_data_1[4047:4040] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_506[17] = buffer_data_1[4055:4048] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_506[18] = buffer_data_1[4063:4056] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_506[19] = buffer_data_1[4071:4064] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_506[20] = buffer_data_0[4039:4032] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_506[21] = buffer_data_0[4047:4040] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_506[22] = buffer_data_0[4055:4048] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_506[23] = buffer_data_0[4063:4056] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_506[24] = buffer_data_0[4071:4064] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_506 = kernel_img_mul_506[0] + kernel_img_mul_506[1] + kernel_img_mul_506[2] + 
                kernel_img_mul_506[3] + kernel_img_mul_506[4] + kernel_img_mul_506[5] + 
                kernel_img_mul_506[6] + kernel_img_mul_506[7] + kernel_img_mul_506[8] + 
                kernel_img_mul_506[9] + kernel_img_mul_506[10] + kernel_img_mul_506[11] + 
                kernel_img_mul_506[12] + kernel_img_mul_506[13] + kernel_img_mul_506[14] + 
                kernel_img_mul_506[15] + kernel_img_mul_506[16] + kernel_img_mul_506[17] + 
                kernel_img_mul_506[18] + kernel_img_mul_506[19] + kernel_img_mul_506[20] + 
                kernel_img_mul_506[21] + kernel_img_mul_506[22] + kernel_img_mul_506[23] + 
                kernel_img_mul_506[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4055:4048] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4055:4048] <= kernel_img_sum_506[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4055:4048] <= 'd0;
end

wire  [39:0]  kernel_img_mul_507[0:24];
assign kernel_img_mul_507[0] = buffer_data_4[4047:4040] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_507[1] = buffer_data_4[4055:4048] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_507[2] = buffer_data_4[4063:4056] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_507[3] = buffer_data_4[4071:4064] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_507[4] = buffer_data_4[4079:4072] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_507[5] = buffer_data_3[4047:4040] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_507[6] = buffer_data_3[4055:4048] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_507[7] = buffer_data_3[4063:4056] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_507[8] = buffer_data_3[4071:4064] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_507[9] = buffer_data_3[4079:4072] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_507[10] = buffer_data_2[4047:4040] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_507[11] = buffer_data_2[4055:4048] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_507[12] = buffer_data_2[4063:4056] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_507[13] = buffer_data_2[4071:4064] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_507[14] = buffer_data_2[4079:4072] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_507[15] = buffer_data_1[4047:4040] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_507[16] = buffer_data_1[4055:4048] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_507[17] = buffer_data_1[4063:4056] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_507[18] = buffer_data_1[4071:4064] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_507[19] = buffer_data_1[4079:4072] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_507[20] = buffer_data_0[4047:4040] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_507[21] = buffer_data_0[4055:4048] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_507[22] = buffer_data_0[4063:4056] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_507[23] = buffer_data_0[4071:4064] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_507[24] = buffer_data_0[4079:4072] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_507 = kernel_img_mul_507[0] + kernel_img_mul_507[1] + kernel_img_mul_507[2] + 
                kernel_img_mul_507[3] + kernel_img_mul_507[4] + kernel_img_mul_507[5] + 
                kernel_img_mul_507[6] + kernel_img_mul_507[7] + kernel_img_mul_507[8] + 
                kernel_img_mul_507[9] + kernel_img_mul_507[10] + kernel_img_mul_507[11] + 
                kernel_img_mul_507[12] + kernel_img_mul_507[13] + kernel_img_mul_507[14] + 
                kernel_img_mul_507[15] + kernel_img_mul_507[16] + kernel_img_mul_507[17] + 
                kernel_img_mul_507[18] + kernel_img_mul_507[19] + kernel_img_mul_507[20] + 
                kernel_img_mul_507[21] + kernel_img_mul_507[22] + kernel_img_mul_507[23] + 
                kernel_img_mul_507[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4063:4056] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4063:4056] <= kernel_img_sum_507[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4063:4056] <= 'd0;
end

wire  [39:0]  kernel_img_mul_508[0:24];
assign kernel_img_mul_508[0] = buffer_data_4[4055:4048] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_508[1] = buffer_data_4[4063:4056] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_508[2] = buffer_data_4[4071:4064] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_508[3] = buffer_data_4[4079:4072] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_508[4] = buffer_data_4[4087:4080] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_508[5] = buffer_data_3[4055:4048] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_508[6] = buffer_data_3[4063:4056] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_508[7] = buffer_data_3[4071:4064] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_508[8] = buffer_data_3[4079:4072] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_508[9] = buffer_data_3[4087:4080] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_508[10] = buffer_data_2[4055:4048] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_508[11] = buffer_data_2[4063:4056] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_508[12] = buffer_data_2[4071:4064] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_508[13] = buffer_data_2[4079:4072] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_508[14] = buffer_data_2[4087:4080] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_508[15] = buffer_data_1[4055:4048] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_508[16] = buffer_data_1[4063:4056] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_508[17] = buffer_data_1[4071:4064] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_508[18] = buffer_data_1[4079:4072] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_508[19] = buffer_data_1[4087:4080] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_508[20] = buffer_data_0[4055:4048] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_508[21] = buffer_data_0[4063:4056] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_508[22] = buffer_data_0[4071:4064] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_508[23] = buffer_data_0[4079:4072] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_508[24] = buffer_data_0[4087:4080] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_508 = kernel_img_mul_508[0] + kernel_img_mul_508[1] + kernel_img_mul_508[2] + 
                kernel_img_mul_508[3] + kernel_img_mul_508[4] + kernel_img_mul_508[5] + 
                kernel_img_mul_508[6] + kernel_img_mul_508[7] + kernel_img_mul_508[8] + 
                kernel_img_mul_508[9] + kernel_img_mul_508[10] + kernel_img_mul_508[11] + 
                kernel_img_mul_508[12] + kernel_img_mul_508[13] + kernel_img_mul_508[14] + 
                kernel_img_mul_508[15] + kernel_img_mul_508[16] + kernel_img_mul_508[17] + 
                kernel_img_mul_508[18] + kernel_img_mul_508[19] + kernel_img_mul_508[20] + 
                kernel_img_mul_508[21] + kernel_img_mul_508[22] + kernel_img_mul_508[23] + 
                kernel_img_mul_508[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4071:4064] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4071:4064] <= kernel_img_sum_508[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4071:4064] <= 'd0;
end

wire  [39:0]  kernel_img_mul_509[0:24];
assign kernel_img_mul_509[0] = buffer_data_4[4063:4056] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_509[1] = buffer_data_4[4071:4064] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_509[2] = buffer_data_4[4079:4072] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_509[3] = buffer_data_4[4087:4080] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_509[4] = buffer_data_4[4095:4088] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_509[5] = buffer_data_3[4063:4056] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_509[6] = buffer_data_3[4071:4064] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_509[7] = buffer_data_3[4079:4072] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_509[8] = buffer_data_3[4087:4080] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_509[9] = buffer_data_3[4095:4088] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_509[10] = buffer_data_2[4063:4056] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_509[11] = buffer_data_2[4071:4064] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_509[12] = buffer_data_2[4079:4072] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_509[13] = buffer_data_2[4087:4080] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_509[14] = buffer_data_2[4095:4088] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_509[15] = buffer_data_1[4063:4056] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_509[16] = buffer_data_1[4071:4064] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_509[17] = buffer_data_1[4079:4072] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_509[18] = buffer_data_1[4087:4080] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_509[19] = buffer_data_1[4095:4088] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_509[20] = buffer_data_0[4063:4056] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_509[21] = buffer_data_0[4071:4064] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_509[22] = buffer_data_0[4079:4072] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_509[23] = buffer_data_0[4087:4080] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_509[24] = buffer_data_0[4095:4088] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_509 = kernel_img_mul_509[0] + kernel_img_mul_509[1] + kernel_img_mul_509[2] + 
                kernel_img_mul_509[3] + kernel_img_mul_509[4] + kernel_img_mul_509[5] + 
                kernel_img_mul_509[6] + kernel_img_mul_509[7] + kernel_img_mul_509[8] + 
                kernel_img_mul_509[9] + kernel_img_mul_509[10] + kernel_img_mul_509[11] + 
                kernel_img_mul_509[12] + kernel_img_mul_509[13] + kernel_img_mul_509[14] + 
                kernel_img_mul_509[15] + kernel_img_mul_509[16] + kernel_img_mul_509[17] + 
                kernel_img_mul_509[18] + kernel_img_mul_509[19] + kernel_img_mul_509[20] + 
                kernel_img_mul_509[21] + kernel_img_mul_509[22] + kernel_img_mul_509[23] + 
                kernel_img_mul_509[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4079:4072] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4079:4072] <= kernel_img_sum_509[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4079:4072] <= 'd0;
end

wire  [39:0]  kernel_img_mul_510[0:24];
assign kernel_img_mul_510[0] = buffer_data_4[4071:4064] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_510[1] = buffer_data_4[4079:4072] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_510[2] = buffer_data_4[4087:4080] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_510[3] = buffer_data_4[4095:4088] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_510[4] = buffer_data_4[4103:4096] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_510[5] = buffer_data_3[4071:4064] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_510[6] = buffer_data_3[4079:4072] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_510[7] = buffer_data_3[4087:4080] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_510[8] = buffer_data_3[4095:4088] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_510[9] = buffer_data_3[4103:4096] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_510[10] = buffer_data_2[4071:4064] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_510[11] = buffer_data_2[4079:4072] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_510[12] = buffer_data_2[4087:4080] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_510[13] = buffer_data_2[4095:4088] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_510[14] = buffer_data_2[4103:4096] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_510[15] = buffer_data_1[4071:4064] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_510[16] = buffer_data_1[4079:4072] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_510[17] = buffer_data_1[4087:4080] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_510[18] = buffer_data_1[4095:4088] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_510[19] = buffer_data_1[4103:4096] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_510[20] = buffer_data_0[4071:4064] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_510[21] = buffer_data_0[4079:4072] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_510[22] = buffer_data_0[4087:4080] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_510[23] = buffer_data_0[4095:4088] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_510[24] = buffer_data_0[4103:4096] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_510 = kernel_img_mul_510[0] + kernel_img_mul_510[1] + kernel_img_mul_510[2] + 
                kernel_img_mul_510[3] + kernel_img_mul_510[4] + kernel_img_mul_510[5] + 
                kernel_img_mul_510[6] + kernel_img_mul_510[7] + kernel_img_mul_510[8] + 
                kernel_img_mul_510[9] + kernel_img_mul_510[10] + kernel_img_mul_510[11] + 
                kernel_img_mul_510[12] + kernel_img_mul_510[13] + kernel_img_mul_510[14] + 
                kernel_img_mul_510[15] + kernel_img_mul_510[16] + kernel_img_mul_510[17] + 
                kernel_img_mul_510[18] + kernel_img_mul_510[19] + kernel_img_mul_510[20] + 
                kernel_img_mul_510[21] + kernel_img_mul_510[22] + kernel_img_mul_510[23] + 
                kernel_img_mul_510[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4087:4080] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4087:4080] <= kernel_img_sum_510[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4087:4080] <= 'd0;
end

wire  [39:0]  kernel_img_mul_511[0:24];
assign kernel_img_mul_511[0] = buffer_data_4[4079:4072] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_511[1] = buffer_data_4[4087:4080] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_511[2] = buffer_data_4[4095:4088] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_511[3] = buffer_data_4[4103:4096] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_511[4] = buffer_data_4[4111:4104] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_511[5] = buffer_data_3[4079:4072] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_511[6] = buffer_data_3[4087:4080] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_511[7] = buffer_data_3[4095:4088] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_511[8] = buffer_data_3[4103:4096] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_511[9] = buffer_data_3[4111:4104] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_511[10] = buffer_data_2[4079:4072] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_511[11] = buffer_data_2[4087:4080] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_511[12] = buffer_data_2[4095:4088] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_511[13] = buffer_data_2[4103:4096] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_511[14] = buffer_data_2[4111:4104] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_511[15] = buffer_data_1[4079:4072] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_511[16] = buffer_data_1[4087:4080] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_511[17] = buffer_data_1[4095:4088] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_511[18] = buffer_data_1[4103:4096] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_511[19] = buffer_data_1[4111:4104] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_511[20] = buffer_data_0[4079:4072] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_511[21] = buffer_data_0[4087:4080] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_511[22] = buffer_data_0[4095:4088] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_511[23] = buffer_data_0[4103:4096] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_511[24] = buffer_data_0[4111:4104] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_511 = kernel_img_mul_511[0] + kernel_img_mul_511[1] + kernel_img_mul_511[2] + 
                kernel_img_mul_511[3] + kernel_img_mul_511[4] + kernel_img_mul_511[5] + 
                kernel_img_mul_511[6] + kernel_img_mul_511[7] + kernel_img_mul_511[8] + 
                kernel_img_mul_511[9] + kernel_img_mul_511[10] + kernel_img_mul_511[11] + 
                kernel_img_mul_511[12] + kernel_img_mul_511[13] + kernel_img_mul_511[14] + 
                kernel_img_mul_511[15] + kernel_img_mul_511[16] + kernel_img_mul_511[17] + 
                kernel_img_mul_511[18] + kernel_img_mul_511[19] + kernel_img_mul_511[20] + 
                kernel_img_mul_511[21] + kernel_img_mul_511[22] + kernel_img_mul_511[23] + 
                kernel_img_mul_511[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4095:4088] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4095:4088] <= kernel_img_sum_511[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4095:4088] <= 'd0;
end

wire  [39:0]  kernel_img_mul_512[0:24];
assign kernel_img_mul_512[0] = buffer_data_4[4087:4080] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_512[1] = buffer_data_4[4095:4088] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_512[2] = buffer_data_4[4103:4096] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_512[3] = buffer_data_4[4111:4104] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_512[4] = buffer_data_4[4119:4112] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_512[5] = buffer_data_3[4087:4080] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_512[6] = buffer_data_3[4095:4088] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_512[7] = buffer_data_3[4103:4096] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_512[8] = buffer_data_3[4111:4104] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_512[9] = buffer_data_3[4119:4112] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_512[10] = buffer_data_2[4087:4080] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_512[11] = buffer_data_2[4095:4088] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_512[12] = buffer_data_2[4103:4096] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_512[13] = buffer_data_2[4111:4104] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_512[14] = buffer_data_2[4119:4112] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_512[15] = buffer_data_1[4087:4080] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_512[16] = buffer_data_1[4095:4088] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_512[17] = buffer_data_1[4103:4096] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_512[18] = buffer_data_1[4111:4104] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_512[19] = buffer_data_1[4119:4112] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_512[20] = buffer_data_0[4087:4080] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_512[21] = buffer_data_0[4095:4088] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_512[22] = buffer_data_0[4103:4096] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_512[23] = buffer_data_0[4111:4104] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_512[24] = buffer_data_0[4119:4112] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_512 = kernel_img_mul_512[0] + kernel_img_mul_512[1] + kernel_img_mul_512[2] + 
                kernel_img_mul_512[3] + kernel_img_mul_512[4] + kernel_img_mul_512[5] + 
                kernel_img_mul_512[6] + kernel_img_mul_512[7] + kernel_img_mul_512[8] + 
                kernel_img_mul_512[9] + kernel_img_mul_512[10] + kernel_img_mul_512[11] + 
                kernel_img_mul_512[12] + kernel_img_mul_512[13] + kernel_img_mul_512[14] + 
                kernel_img_mul_512[15] + kernel_img_mul_512[16] + kernel_img_mul_512[17] + 
                kernel_img_mul_512[18] + kernel_img_mul_512[19] + kernel_img_mul_512[20] + 
                kernel_img_mul_512[21] + kernel_img_mul_512[22] + kernel_img_mul_512[23] + 
                kernel_img_mul_512[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4103:4096] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4103:4096] <= kernel_img_sum_512[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4103:4096] <= 'd0;
end

wire  [39:0]  kernel_img_mul_513[0:24];
assign kernel_img_mul_513[0] = buffer_data_4[4095:4088] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_513[1] = buffer_data_4[4103:4096] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_513[2] = buffer_data_4[4111:4104] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_513[3] = buffer_data_4[4119:4112] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_513[4] = buffer_data_4[4127:4120] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_513[5] = buffer_data_3[4095:4088] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_513[6] = buffer_data_3[4103:4096] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_513[7] = buffer_data_3[4111:4104] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_513[8] = buffer_data_3[4119:4112] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_513[9] = buffer_data_3[4127:4120] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_513[10] = buffer_data_2[4095:4088] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_513[11] = buffer_data_2[4103:4096] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_513[12] = buffer_data_2[4111:4104] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_513[13] = buffer_data_2[4119:4112] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_513[14] = buffer_data_2[4127:4120] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_513[15] = buffer_data_1[4095:4088] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_513[16] = buffer_data_1[4103:4096] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_513[17] = buffer_data_1[4111:4104] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_513[18] = buffer_data_1[4119:4112] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_513[19] = buffer_data_1[4127:4120] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_513[20] = buffer_data_0[4095:4088] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_513[21] = buffer_data_0[4103:4096] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_513[22] = buffer_data_0[4111:4104] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_513[23] = buffer_data_0[4119:4112] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_513[24] = buffer_data_0[4127:4120] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_513 = kernel_img_mul_513[0] + kernel_img_mul_513[1] + kernel_img_mul_513[2] + 
                kernel_img_mul_513[3] + kernel_img_mul_513[4] + kernel_img_mul_513[5] + 
                kernel_img_mul_513[6] + kernel_img_mul_513[7] + kernel_img_mul_513[8] + 
                kernel_img_mul_513[9] + kernel_img_mul_513[10] + kernel_img_mul_513[11] + 
                kernel_img_mul_513[12] + kernel_img_mul_513[13] + kernel_img_mul_513[14] + 
                kernel_img_mul_513[15] + kernel_img_mul_513[16] + kernel_img_mul_513[17] + 
                kernel_img_mul_513[18] + kernel_img_mul_513[19] + kernel_img_mul_513[20] + 
                kernel_img_mul_513[21] + kernel_img_mul_513[22] + kernel_img_mul_513[23] + 
                kernel_img_mul_513[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4111:4104] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4111:4104] <= kernel_img_sum_513[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4111:4104] <= 'd0;
end

wire  [39:0]  kernel_img_mul_514[0:24];
assign kernel_img_mul_514[0] = buffer_data_4[4103:4096] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_514[1] = buffer_data_4[4111:4104] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_514[2] = buffer_data_4[4119:4112] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_514[3] = buffer_data_4[4127:4120] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_514[4] = buffer_data_4[4135:4128] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_514[5] = buffer_data_3[4103:4096] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_514[6] = buffer_data_3[4111:4104] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_514[7] = buffer_data_3[4119:4112] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_514[8] = buffer_data_3[4127:4120] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_514[9] = buffer_data_3[4135:4128] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_514[10] = buffer_data_2[4103:4096] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_514[11] = buffer_data_2[4111:4104] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_514[12] = buffer_data_2[4119:4112] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_514[13] = buffer_data_2[4127:4120] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_514[14] = buffer_data_2[4135:4128] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_514[15] = buffer_data_1[4103:4096] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_514[16] = buffer_data_1[4111:4104] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_514[17] = buffer_data_1[4119:4112] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_514[18] = buffer_data_1[4127:4120] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_514[19] = buffer_data_1[4135:4128] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_514[20] = buffer_data_0[4103:4096] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_514[21] = buffer_data_0[4111:4104] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_514[22] = buffer_data_0[4119:4112] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_514[23] = buffer_data_0[4127:4120] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_514[24] = buffer_data_0[4135:4128] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_514 = kernel_img_mul_514[0] + kernel_img_mul_514[1] + kernel_img_mul_514[2] + 
                kernel_img_mul_514[3] + kernel_img_mul_514[4] + kernel_img_mul_514[5] + 
                kernel_img_mul_514[6] + kernel_img_mul_514[7] + kernel_img_mul_514[8] + 
                kernel_img_mul_514[9] + kernel_img_mul_514[10] + kernel_img_mul_514[11] + 
                kernel_img_mul_514[12] + kernel_img_mul_514[13] + kernel_img_mul_514[14] + 
                kernel_img_mul_514[15] + kernel_img_mul_514[16] + kernel_img_mul_514[17] + 
                kernel_img_mul_514[18] + kernel_img_mul_514[19] + kernel_img_mul_514[20] + 
                kernel_img_mul_514[21] + kernel_img_mul_514[22] + kernel_img_mul_514[23] + 
                kernel_img_mul_514[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4119:4112] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4119:4112] <= kernel_img_sum_514[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4119:4112] <= 'd0;
end

wire  [39:0]  kernel_img_mul_515[0:24];
assign kernel_img_mul_515[0] = buffer_data_4[4111:4104] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_515[1] = buffer_data_4[4119:4112] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_515[2] = buffer_data_4[4127:4120] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_515[3] = buffer_data_4[4135:4128] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_515[4] = buffer_data_4[4143:4136] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_515[5] = buffer_data_3[4111:4104] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_515[6] = buffer_data_3[4119:4112] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_515[7] = buffer_data_3[4127:4120] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_515[8] = buffer_data_3[4135:4128] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_515[9] = buffer_data_3[4143:4136] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_515[10] = buffer_data_2[4111:4104] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_515[11] = buffer_data_2[4119:4112] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_515[12] = buffer_data_2[4127:4120] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_515[13] = buffer_data_2[4135:4128] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_515[14] = buffer_data_2[4143:4136] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_515[15] = buffer_data_1[4111:4104] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_515[16] = buffer_data_1[4119:4112] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_515[17] = buffer_data_1[4127:4120] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_515[18] = buffer_data_1[4135:4128] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_515[19] = buffer_data_1[4143:4136] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_515[20] = buffer_data_0[4111:4104] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_515[21] = buffer_data_0[4119:4112] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_515[22] = buffer_data_0[4127:4120] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_515[23] = buffer_data_0[4135:4128] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_515[24] = buffer_data_0[4143:4136] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_515 = kernel_img_mul_515[0] + kernel_img_mul_515[1] + kernel_img_mul_515[2] + 
                kernel_img_mul_515[3] + kernel_img_mul_515[4] + kernel_img_mul_515[5] + 
                kernel_img_mul_515[6] + kernel_img_mul_515[7] + kernel_img_mul_515[8] + 
                kernel_img_mul_515[9] + kernel_img_mul_515[10] + kernel_img_mul_515[11] + 
                kernel_img_mul_515[12] + kernel_img_mul_515[13] + kernel_img_mul_515[14] + 
                kernel_img_mul_515[15] + kernel_img_mul_515[16] + kernel_img_mul_515[17] + 
                kernel_img_mul_515[18] + kernel_img_mul_515[19] + kernel_img_mul_515[20] + 
                kernel_img_mul_515[21] + kernel_img_mul_515[22] + kernel_img_mul_515[23] + 
                kernel_img_mul_515[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4127:4120] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4127:4120] <= kernel_img_sum_515[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4127:4120] <= 'd0;
end

wire  [39:0]  kernel_img_mul_516[0:24];
assign kernel_img_mul_516[0] = buffer_data_4[4119:4112] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_516[1] = buffer_data_4[4127:4120] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_516[2] = buffer_data_4[4135:4128] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_516[3] = buffer_data_4[4143:4136] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_516[4] = buffer_data_4[4151:4144] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_516[5] = buffer_data_3[4119:4112] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_516[6] = buffer_data_3[4127:4120] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_516[7] = buffer_data_3[4135:4128] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_516[8] = buffer_data_3[4143:4136] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_516[9] = buffer_data_3[4151:4144] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_516[10] = buffer_data_2[4119:4112] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_516[11] = buffer_data_2[4127:4120] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_516[12] = buffer_data_2[4135:4128] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_516[13] = buffer_data_2[4143:4136] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_516[14] = buffer_data_2[4151:4144] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_516[15] = buffer_data_1[4119:4112] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_516[16] = buffer_data_1[4127:4120] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_516[17] = buffer_data_1[4135:4128] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_516[18] = buffer_data_1[4143:4136] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_516[19] = buffer_data_1[4151:4144] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_516[20] = buffer_data_0[4119:4112] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_516[21] = buffer_data_0[4127:4120] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_516[22] = buffer_data_0[4135:4128] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_516[23] = buffer_data_0[4143:4136] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_516[24] = buffer_data_0[4151:4144] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_516 = kernel_img_mul_516[0] + kernel_img_mul_516[1] + kernel_img_mul_516[2] + 
                kernel_img_mul_516[3] + kernel_img_mul_516[4] + kernel_img_mul_516[5] + 
                kernel_img_mul_516[6] + kernel_img_mul_516[7] + kernel_img_mul_516[8] + 
                kernel_img_mul_516[9] + kernel_img_mul_516[10] + kernel_img_mul_516[11] + 
                kernel_img_mul_516[12] + kernel_img_mul_516[13] + kernel_img_mul_516[14] + 
                kernel_img_mul_516[15] + kernel_img_mul_516[16] + kernel_img_mul_516[17] + 
                kernel_img_mul_516[18] + kernel_img_mul_516[19] + kernel_img_mul_516[20] + 
                kernel_img_mul_516[21] + kernel_img_mul_516[22] + kernel_img_mul_516[23] + 
                kernel_img_mul_516[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4135:4128] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4135:4128] <= kernel_img_sum_516[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4135:4128] <= 'd0;
end

wire  [39:0]  kernel_img_mul_517[0:24];
assign kernel_img_mul_517[0] = buffer_data_4[4127:4120] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_517[1] = buffer_data_4[4135:4128] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_517[2] = buffer_data_4[4143:4136] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_517[3] = buffer_data_4[4151:4144] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_517[4] = buffer_data_4[4159:4152] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_517[5] = buffer_data_3[4127:4120] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_517[6] = buffer_data_3[4135:4128] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_517[7] = buffer_data_3[4143:4136] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_517[8] = buffer_data_3[4151:4144] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_517[9] = buffer_data_3[4159:4152] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_517[10] = buffer_data_2[4127:4120] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_517[11] = buffer_data_2[4135:4128] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_517[12] = buffer_data_2[4143:4136] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_517[13] = buffer_data_2[4151:4144] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_517[14] = buffer_data_2[4159:4152] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_517[15] = buffer_data_1[4127:4120] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_517[16] = buffer_data_1[4135:4128] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_517[17] = buffer_data_1[4143:4136] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_517[18] = buffer_data_1[4151:4144] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_517[19] = buffer_data_1[4159:4152] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_517[20] = buffer_data_0[4127:4120] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_517[21] = buffer_data_0[4135:4128] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_517[22] = buffer_data_0[4143:4136] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_517[23] = buffer_data_0[4151:4144] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_517[24] = buffer_data_0[4159:4152] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_517 = kernel_img_mul_517[0] + kernel_img_mul_517[1] + kernel_img_mul_517[2] + 
                kernel_img_mul_517[3] + kernel_img_mul_517[4] + kernel_img_mul_517[5] + 
                kernel_img_mul_517[6] + kernel_img_mul_517[7] + kernel_img_mul_517[8] + 
                kernel_img_mul_517[9] + kernel_img_mul_517[10] + kernel_img_mul_517[11] + 
                kernel_img_mul_517[12] + kernel_img_mul_517[13] + kernel_img_mul_517[14] + 
                kernel_img_mul_517[15] + kernel_img_mul_517[16] + kernel_img_mul_517[17] + 
                kernel_img_mul_517[18] + kernel_img_mul_517[19] + kernel_img_mul_517[20] + 
                kernel_img_mul_517[21] + kernel_img_mul_517[22] + kernel_img_mul_517[23] + 
                kernel_img_mul_517[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4143:4136] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4143:4136] <= kernel_img_sum_517[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4143:4136] <= 'd0;
end

wire  [39:0]  kernel_img_mul_518[0:24];
assign kernel_img_mul_518[0] = buffer_data_4[4135:4128] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_518[1] = buffer_data_4[4143:4136] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_518[2] = buffer_data_4[4151:4144] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_518[3] = buffer_data_4[4159:4152] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_518[4] = buffer_data_4[4167:4160] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_518[5] = buffer_data_3[4135:4128] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_518[6] = buffer_data_3[4143:4136] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_518[7] = buffer_data_3[4151:4144] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_518[8] = buffer_data_3[4159:4152] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_518[9] = buffer_data_3[4167:4160] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_518[10] = buffer_data_2[4135:4128] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_518[11] = buffer_data_2[4143:4136] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_518[12] = buffer_data_2[4151:4144] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_518[13] = buffer_data_2[4159:4152] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_518[14] = buffer_data_2[4167:4160] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_518[15] = buffer_data_1[4135:4128] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_518[16] = buffer_data_1[4143:4136] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_518[17] = buffer_data_1[4151:4144] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_518[18] = buffer_data_1[4159:4152] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_518[19] = buffer_data_1[4167:4160] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_518[20] = buffer_data_0[4135:4128] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_518[21] = buffer_data_0[4143:4136] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_518[22] = buffer_data_0[4151:4144] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_518[23] = buffer_data_0[4159:4152] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_518[24] = buffer_data_0[4167:4160] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_518 = kernel_img_mul_518[0] + kernel_img_mul_518[1] + kernel_img_mul_518[2] + 
                kernel_img_mul_518[3] + kernel_img_mul_518[4] + kernel_img_mul_518[5] + 
                kernel_img_mul_518[6] + kernel_img_mul_518[7] + kernel_img_mul_518[8] + 
                kernel_img_mul_518[9] + kernel_img_mul_518[10] + kernel_img_mul_518[11] + 
                kernel_img_mul_518[12] + kernel_img_mul_518[13] + kernel_img_mul_518[14] + 
                kernel_img_mul_518[15] + kernel_img_mul_518[16] + kernel_img_mul_518[17] + 
                kernel_img_mul_518[18] + kernel_img_mul_518[19] + kernel_img_mul_518[20] + 
                kernel_img_mul_518[21] + kernel_img_mul_518[22] + kernel_img_mul_518[23] + 
                kernel_img_mul_518[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4151:4144] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4151:4144] <= kernel_img_sum_518[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4151:4144] <= 'd0;
end

wire  [39:0]  kernel_img_mul_519[0:24];
assign kernel_img_mul_519[0] = buffer_data_4[4143:4136] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_519[1] = buffer_data_4[4151:4144] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_519[2] = buffer_data_4[4159:4152] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_519[3] = buffer_data_4[4167:4160] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_519[4] = buffer_data_4[4175:4168] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_519[5] = buffer_data_3[4143:4136] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_519[6] = buffer_data_3[4151:4144] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_519[7] = buffer_data_3[4159:4152] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_519[8] = buffer_data_3[4167:4160] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_519[9] = buffer_data_3[4175:4168] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_519[10] = buffer_data_2[4143:4136] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_519[11] = buffer_data_2[4151:4144] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_519[12] = buffer_data_2[4159:4152] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_519[13] = buffer_data_2[4167:4160] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_519[14] = buffer_data_2[4175:4168] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_519[15] = buffer_data_1[4143:4136] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_519[16] = buffer_data_1[4151:4144] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_519[17] = buffer_data_1[4159:4152] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_519[18] = buffer_data_1[4167:4160] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_519[19] = buffer_data_1[4175:4168] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_519[20] = buffer_data_0[4143:4136] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_519[21] = buffer_data_0[4151:4144] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_519[22] = buffer_data_0[4159:4152] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_519[23] = buffer_data_0[4167:4160] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_519[24] = buffer_data_0[4175:4168] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_519 = kernel_img_mul_519[0] + kernel_img_mul_519[1] + kernel_img_mul_519[2] + 
                kernel_img_mul_519[3] + kernel_img_mul_519[4] + kernel_img_mul_519[5] + 
                kernel_img_mul_519[6] + kernel_img_mul_519[7] + kernel_img_mul_519[8] + 
                kernel_img_mul_519[9] + kernel_img_mul_519[10] + kernel_img_mul_519[11] + 
                kernel_img_mul_519[12] + kernel_img_mul_519[13] + kernel_img_mul_519[14] + 
                kernel_img_mul_519[15] + kernel_img_mul_519[16] + kernel_img_mul_519[17] + 
                kernel_img_mul_519[18] + kernel_img_mul_519[19] + kernel_img_mul_519[20] + 
                kernel_img_mul_519[21] + kernel_img_mul_519[22] + kernel_img_mul_519[23] + 
                kernel_img_mul_519[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4159:4152] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4159:4152] <= kernel_img_sum_519[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4159:4152] <= 'd0;
end

wire  [39:0]  kernel_img_mul_520[0:24];
assign kernel_img_mul_520[0] = buffer_data_4[4151:4144] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_520[1] = buffer_data_4[4159:4152] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_520[2] = buffer_data_4[4167:4160] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_520[3] = buffer_data_4[4175:4168] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_520[4] = buffer_data_4[4183:4176] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_520[5] = buffer_data_3[4151:4144] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_520[6] = buffer_data_3[4159:4152] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_520[7] = buffer_data_3[4167:4160] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_520[8] = buffer_data_3[4175:4168] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_520[9] = buffer_data_3[4183:4176] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_520[10] = buffer_data_2[4151:4144] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_520[11] = buffer_data_2[4159:4152] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_520[12] = buffer_data_2[4167:4160] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_520[13] = buffer_data_2[4175:4168] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_520[14] = buffer_data_2[4183:4176] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_520[15] = buffer_data_1[4151:4144] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_520[16] = buffer_data_1[4159:4152] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_520[17] = buffer_data_1[4167:4160] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_520[18] = buffer_data_1[4175:4168] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_520[19] = buffer_data_1[4183:4176] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_520[20] = buffer_data_0[4151:4144] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_520[21] = buffer_data_0[4159:4152] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_520[22] = buffer_data_0[4167:4160] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_520[23] = buffer_data_0[4175:4168] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_520[24] = buffer_data_0[4183:4176] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_520 = kernel_img_mul_520[0] + kernel_img_mul_520[1] + kernel_img_mul_520[2] + 
                kernel_img_mul_520[3] + kernel_img_mul_520[4] + kernel_img_mul_520[5] + 
                kernel_img_mul_520[6] + kernel_img_mul_520[7] + kernel_img_mul_520[8] + 
                kernel_img_mul_520[9] + kernel_img_mul_520[10] + kernel_img_mul_520[11] + 
                kernel_img_mul_520[12] + kernel_img_mul_520[13] + kernel_img_mul_520[14] + 
                kernel_img_mul_520[15] + kernel_img_mul_520[16] + kernel_img_mul_520[17] + 
                kernel_img_mul_520[18] + kernel_img_mul_520[19] + kernel_img_mul_520[20] + 
                kernel_img_mul_520[21] + kernel_img_mul_520[22] + kernel_img_mul_520[23] + 
                kernel_img_mul_520[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4167:4160] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4167:4160] <= kernel_img_sum_520[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4167:4160] <= 'd0;
end

wire  [39:0]  kernel_img_mul_521[0:24];
assign kernel_img_mul_521[0] = buffer_data_4[4159:4152] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_521[1] = buffer_data_4[4167:4160] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_521[2] = buffer_data_4[4175:4168] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_521[3] = buffer_data_4[4183:4176] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_521[4] = buffer_data_4[4191:4184] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_521[5] = buffer_data_3[4159:4152] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_521[6] = buffer_data_3[4167:4160] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_521[7] = buffer_data_3[4175:4168] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_521[8] = buffer_data_3[4183:4176] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_521[9] = buffer_data_3[4191:4184] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_521[10] = buffer_data_2[4159:4152] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_521[11] = buffer_data_2[4167:4160] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_521[12] = buffer_data_2[4175:4168] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_521[13] = buffer_data_2[4183:4176] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_521[14] = buffer_data_2[4191:4184] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_521[15] = buffer_data_1[4159:4152] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_521[16] = buffer_data_1[4167:4160] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_521[17] = buffer_data_1[4175:4168] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_521[18] = buffer_data_1[4183:4176] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_521[19] = buffer_data_1[4191:4184] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_521[20] = buffer_data_0[4159:4152] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_521[21] = buffer_data_0[4167:4160] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_521[22] = buffer_data_0[4175:4168] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_521[23] = buffer_data_0[4183:4176] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_521[24] = buffer_data_0[4191:4184] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_521 = kernel_img_mul_521[0] + kernel_img_mul_521[1] + kernel_img_mul_521[2] + 
                kernel_img_mul_521[3] + kernel_img_mul_521[4] + kernel_img_mul_521[5] + 
                kernel_img_mul_521[6] + kernel_img_mul_521[7] + kernel_img_mul_521[8] + 
                kernel_img_mul_521[9] + kernel_img_mul_521[10] + kernel_img_mul_521[11] + 
                kernel_img_mul_521[12] + kernel_img_mul_521[13] + kernel_img_mul_521[14] + 
                kernel_img_mul_521[15] + kernel_img_mul_521[16] + kernel_img_mul_521[17] + 
                kernel_img_mul_521[18] + kernel_img_mul_521[19] + kernel_img_mul_521[20] + 
                kernel_img_mul_521[21] + kernel_img_mul_521[22] + kernel_img_mul_521[23] + 
                kernel_img_mul_521[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4175:4168] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4175:4168] <= kernel_img_sum_521[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4175:4168] <= 'd0;
end

wire  [39:0]  kernel_img_mul_522[0:24];
assign kernel_img_mul_522[0] = buffer_data_4[4167:4160] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_522[1] = buffer_data_4[4175:4168] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_522[2] = buffer_data_4[4183:4176] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_522[3] = buffer_data_4[4191:4184] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_522[4] = buffer_data_4[4199:4192] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_522[5] = buffer_data_3[4167:4160] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_522[6] = buffer_data_3[4175:4168] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_522[7] = buffer_data_3[4183:4176] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_522[8] = buffer_data_3[4191:4184] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_522[9] = buffer_data_3[4199:4192] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_522[10] = buffer_data_2[4167:4160] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_522[11] = buffer_data_2[4175:4168] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_522[12] = buffer_data_2[4183:4176] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_522[13] = buffer_data_2[4191:4184] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_522[14] = buffer_data_2[4199:4192] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_522[15] = buffer_data_1[4167:4160] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_522[16] = buffer_data_1[4175:4168] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_522[17] = buffer_data_1[4183:4176] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_522[18] = buffer_data_1[4191:4184] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_522[19] = buffer_data_1[4199:4192] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_522[20] = buffer_data_0[4167:4160] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_522[21] = buffer_data_0[4175:4168] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_522[22] = buffer_data_0[4183:4176] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_522[23] = buffer_data_0[4191:4184] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_522[24] = buffer_data_0[4199:4192] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_522 = kernel_img_mul_522[0] + kernel_img_mul_522[1] + kernel_img_mul_522[2] + 
                kernel_img_mul_522[3] + kernel_img_mul_522[4] + kernel_img_mul_522[5] + 
                kernel_img_mul_522[6] + kernel_img_mul_522[7] + kernel_img_mul_522[8] + 
                kernel_img_mul_522[9] + kernel_img_mul_522[10] + kernel_img_mul_522[11] + 
                kernel_img_mul_522[12] + kernel_img_mul_522[13] + kernel_img_mul_522[14] + 
                kernel_img_mul_522[15] + kernel_img_mul_522[16] + kernel_img_mul_522[17] + 
                kernel_img_mul_522[18] + kernel_img_mul_522[19] + kernel_img_mul_522[20] + 
                kernel_img_mul_522[21] + kernel_img_mul_522[22] + kernel_img_mul_522[23] + 
                kernel_img_mul_522[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4183:4176] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4183:4176] <= kernel_img_sum_522[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4183:4176] <= 'd0;
end

wire  [39:0]  kernel_img_mul_523[0:24];
assign kernel_img_mul_523[0] = buffer_data_4[4175:4168] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_523[1] = buffer_data_4[4183:4176] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_523[2] = buffer_data_4[4191:4184] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_523[3] = buffer_data_4[4199:4192] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_523[4] = buffer_data_4[4207:4200] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_523[5] = buffer_data_3[4175:4168] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_523[6] = buffer_data_3[4183:4176] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_523[7] = buffer_data_3[4191:4184] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_523[8] = buffer_data_3[4199:4192] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_523[9] = buffer_data_3[4207:4200] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_523[10] = buffer_data_2[4175:4168] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_523[11] = buffer_data_2[4183:4176] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_523[12] = buffer_data_2[4191:4184] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_523[13] = buffer_data_2[4199:4192] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_523[14] = buffer_data_2[4207:4200] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_523[15] = buffer_data_1[4175:4168] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_523[16] = buffer_data_1[4183:4176] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_523[17] = buffer_data_1[4191:4184] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_523[18] = buffer_data_1[4199:4192] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_523[19] = buffer_data_1[4207:4200] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_523[20] = buffer_data_0[4175:4168] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_523[21] = buffer_data_0[4183:4176] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_523[22] = buffer_data_0[4191:4184] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_523[23] = buffer_data_0[4199:4192] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_523[24] = buffer_data_0[4207:4200] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_523 = kernel_img_mul_523[0] + kernel_img_mul_523[1] + kernel_img_mul_523[2] + 
                kernel_img_mul_523[3] + kernel_img_mul_523[4] + kernel_img_mul_523[5] + 
                kernel_img_mul_523[6] + kernel_img_mul_523[7] + kernel_img_mul_523[8] + 
                kernel_img_mul_523[9] + kernel_img_mul_523[10] + kernel_img_mul_523[11] + 
                kernel_img_mul_523[12] + kernel_img_mul_523[13] + kernel_img_mul_523[14] + 
                kernel_img_mul_523[15] + kernel_img_mul_523[16] + kernel_img_mul_523[17] + 
                kernel_img_mul_523[18] + kernel_img_mul_523[19] + kernel_img_mul_523[20] + 
                kernel_img_mul_523[21] + kernel_img_mul_523[22] + kernel_img_mul_523[23] + 
                kernel_img_mul_523[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4191:4184] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4191:4184] <= kernel_img_sum_523[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4191:4184] <= 'd0;
end

wire  [39:0]  kernel_img_mul_524[0:24];
assign kernel_img_mul_524[0] = buffer_data_4[4183:4176] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_524[1] = buffer_data_4[4191:4184] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_524[2] = buffer_data_4[4199:4192] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_524[3] = buffer_data_4[4207:4200] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_524[4] = buffer_data_4[4215:4208] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_524[5] = buffer_data_3[4183:4176] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_524[6] = buffer_data_3[4191:4184] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_524[7] = buffer_data_3[4199:4192] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_524[8] = buffer_data_3[4207:4200] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_524[9] = buffer_data_3[4215:4208] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_524[10] = buffer_data_2[4183:4176] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_524[11] = buffer_data_2[4191:4184] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_524[12] = buffer_data_2[4199:4192] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_524[13] = buffer_data_2[4207:4200] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_524[14] = buffer_data_2[4215:4208] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_524[15] = buffer_data_1[4183:4176] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_524[16] = buffer_data_1[4191:4184] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_524[17] = buffer_data_1[4199:4192] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_524[18] = buffer_data_1[4207:4200] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_524[19] = buffer_data_1[4215:4208] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_524[20] = buffer_data_0[4183:4176] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_524[21] = buffer_data_0[4191:4184] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_524[22] = buffer_data_0[4199:4192] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_524[23] = buffer_data_0[4207:4200] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_524[24] = buffer_data_0[4215:4208] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_524 = kernel_img_mul_524[0] + kernel_img_mul_524[1] + kernel_img_mul_524[2] + 
                kernel_img_mul_524[3] + kernel_img_mul_524[4] + kernel_img_mul_524[5] + 
                kernel_img_mul_524[6] + kernel_img_mul_524[7] + kernel_img_mul_524[8] + 
                kernel_img_mul_524[9] + kernel_img_mul_524[10] + kernel_img_mul_524[11] + 
                kernel_img_mul_524[12] + kernel_img_mul_524[13] + kernel_img_mul_524[14] + 
                kernel_img_mul_524[15] + kernel_img_mul_524[16] + kernel_img_mul_524[17] + 
                kernel_img_mul_524[18] + kernel_img_mul_524[19] + kernel_img_mul_524[20] + 
                kernel_img_mul_524[21] + kernel_img_mul_524[22] + kernel_img_mul_524[23] + 
                kernel_img_mul_524[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4199:4192] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4199:4192] <= kernel_img_sum_524[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4199:4192] <= 'd0;
end

wire  [39:0]  kernel_img_mul_525[0:24];
assign kernel_img_mul_525[0] = buffer_data_4[4191:4184] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_525[1] = buffer_data_4[4199:4192] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_525[2] = buffer_data_4[4207:4200] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_525[3] = buffer_data_4[4215:4208] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_525[4] = buffer_data_4[4223:4216] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_525[5] = buffer_data_3[4191:4184] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_525[6] = buffer_data_3[4199:4192] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_525[7] = buffer_data_3[4207:4200] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_525[8] = buffer_data_3[4215:4208] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_525[9] = buffer_data_3[4223:4216] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_525[10] = buffer_data_2[4191:4184] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_525[11] = buffer_data_2[4199:4192] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_525[12] = buffer_data_2[4207:4200] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_525[13] = buffer_data_2[4215:4208] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_525[14] = buffer_data_2[4223:4216] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_525[15] = buffer_data_1[4191:4184] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_525[16] = buffer_data_1[4199:4192] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_525[17] = buffer_data_1[4207:4200] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_525[18] = buffer_data_1[4215:4208] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_525[19] = buffer_data_1[4223:4216] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_525[20] = buffer_data_0[4191:4184] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_525[21] = buffer_data_0[4199:4192] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_525[22] = buffer_data_0[4207:4200] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_525[23] = buffer_data_0[4215:4208] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_525[24] = buffer_data_0[4223:4216] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_525 = kernel_img_mul_525[0] + kernel_img_mul_525[1] + kernel_img_mul_525[2] + 
                kernel_img_mul_525[3] + kernel_img_mul_525[4] + kernel_img_mul_525[5] + 
                kernel_img_mul_525[6] + kernel_img_mul_525[7] + kernel_img_mul_525[8] + 
                kernel_img_mul_525[9] + kernel_img_mul_525[10] + kernel_img_mul_525[11] + 
                kernel_img_mul_525[12] + kernel_img_mul_525[13] + kernel_img_mul_525[14] + 
                kernel_img_mul_525[15] + kernel_img_mul_525[16] + kernel_img_mul_525[17] + 
                kernel_img_mul_525[18] + kernel_img_mul_525[19] + kernel_img_mul_525[20] + 
                kernel_img_mul_525[21] + kernel_img_mul_525[22] + kernel_img_mul_525[23] + 
                kernel_img_mul_525[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4207:4200] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4207:4200] <= kernel_img_sum_525[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4207:4200] <= 'd0;
end

wire  [39:0]  kernel_img_mul_526[0:24];
assign kernel_img_mul_526[0] = buffer_data_4[4199:4192] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_526[1] = buffer_data_4[4207:4200] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_526[2] = buffer_data_4[4215:4208] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_526[3] = buffer_data_4[4223:4216] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_526[4] = buffer_data_4[4231:4224] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_526[5] = buffer_data_3[4199:4192] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_526[6] = buffer_data_3[4207:4200] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_526[7] = buffer_data_3[4215:4208] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_526[8] = buffer_data_3[4223:4216] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_526[9] = buffer_data_3[4231:4224] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_526[10] = buffer_data_2[4199:4192] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_526[11] = buffer_data_2[4207:4200] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_526[12] = buffer_data_2[4215:4208] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_526[13] = buffer_data_2[4223:4216] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_526[14] = buffer_data_2[4231:4224] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_526[15] = buffer_data_1[4199:4192] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_526[16] = buffer_data_1[4207:4200] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_526[17] = buffer_data_1[4215:4208] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_526[18] = buffer_data_1[4223:4216] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_526[19] = buffer_data_1[4231:4224] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_526[20] = buffer_data_0[4199:4192] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_526[21] = buffer_data_0[4207:4200] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_526[22] = buffer_data_0[4215:4208] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_526[23] = buffer_data_0[4223:4216] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_526[24] = buffer_data_0[4231:4224] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_526 = kernel_img_mul_526[0] + kernel_img_mul_526[1] + kernel_img_mul_526[2] + 
                kernel_img_mul_526[3] + kernel_img_mul_526[4] + kernel_img_mul_526[5] + 
                kernel_img_mul_526[6] + kernel_img_mul_526[7] + kernel_img_mul_526[8] + 
                kernel_img_mul_526[9] + kernel_img_mul_526[10] + kernel_img_mul_526[11] + 
                kernel_img_mul_526[12] + kernel_img_mul_526[13] + kernel_img_mul_526[14] + 
                kernel_img_mul_526[15] + kernel_img_mul_526[16] + kernel_img_mul_526[17] + 
                kernel_img_mul_526[18] + kernel_img_mul_526[19] + kernel_img_mul_526[20] + 
                kernel_img_mul_526[21] + kernel_img_mul_526[22] + kernel_img_mul_526[23] + 
                kernel_img_mul_526[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4215:4208] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4215:4208] <= kernel_img_sum_526[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4215:4208] <= 'd0;
end

wire  [39:0]  kernel_img_mul_527[0:24];
assign kernel_img_mul_527[0] = buffer_data_4[4207:4200] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_527[1] = buffer_data_4[4215:4208] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_527[2] = buffer_data_4[4223:4216] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_527[3] = buffer_data_4[4231:4224] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_527[4] = buffer_data_4[4239:4232] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_527[5] = buffer_data_3[4207:4200] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_527[6] = buffer_data_3[4215:4208] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_527[7] = buffer_data_3[4223:4216] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_527[8] = buffer_data_3[4231:4224] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_527[9] = buffer_data_3[4239:4232] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_527[10] = buffer_data_2[4207:4200] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_527[11] = buffer_data_2[4215:4208] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_527[12] = buffer_data_2[4223:4216] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_527[13] = buffer_data_2[4231:4224] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_527[14] = buffer_data_2[4239:4232] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_527[15] = buffer_data_1[4207:4200] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_527[16] = buffer_data_1[4215:4208] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_527[17] = buffer_data_1[4223:4216] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_527[18] = buffer_data_1[4231:4224] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_527[19] = buffer_data_1[4239:4232] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_527[20] = buffer_data_0[4207:4200] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_527[21] = buffer_data_0[4215:4208] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_527[22] = buffer_data_0[4223:4216] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_527[23] = buffer_data_0[4231:4224] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_527[24] = buffer_data_0[4239:4232] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_527 = kernel_img_mul_527[0] + kernel_img_mul_527[1] + kernel_img_mul_527[2] + 
                kernel_img_mul_527[3] + kernel_img_mul_527[4] + kernel_img_mul_527[5] + 
                kernel_img_mul_527[6] + kernel_img_mul_527[7] + kernel_img_mul_527[8] + 
                kernel_img_mul_527[9] + kernel_img_mul_527[10] + kernel_img_mul_527[11] + 
                kernel_img_mul_527[12] + kernel_img_mul_527[13] + kernel_img_mul_527[14] + 
                kernel_img_mul_527[15] + kernel_img_mul_527[16] + kernel_img_mul_527[17] + 
                kernel_img_mul_527[18] + kernel_img_mul_527[19] + kernel_img_mul_527[20] + 
                kernel_img_mul_527[21] + kernel_img_mul_527[22] + kernel_img_mul_527[23] + 
                kernel_img_mul_527[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4223:4216] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4223:4216] <= kernel_img_sum_527[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4223:4216] <= 'd0;
end

wire  [39:0]  kernel_img_mul_528[0:24];
assign kernel_img_mul_528[0] = buffer_data_4[4215:4208] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_528[1] = buffer_data_4[4223:4216] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_528[2] = buffer_data_4[4231:4224] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_528[3] = buffer_data_4[4239:4232] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_528[4] = buffer_data_4[4247:4240] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_528[5] = buffer_data_3[4215:4208] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_528[6] = buffer_data_3[4223:4216] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_528[7] = buffer_data_3[4231:4224] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_528[8] = buffer_data_3[4239:4232] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_528[9] = buffer_data_3[4247:4240] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_528[10] = buffer_data_2[4215:4208] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_528[11] = buffer_data_2[4223:4216] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_528[12] = buffer_data_2[4231:4224] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_528[13] = buffer_data_2[4239:4232] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_528[14] = buffer_data_2[4247:4240] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_528[15] = buffer_data_1[4215:4208] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_528[16] = buffer_data_1[4223:4216] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_528[17] = buffer_data_1[4231:4224] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_528[18] = buffer_data_1[4239:4232] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_528[19] = buffer_data_1[4247:4240] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_528[20] = buffer_data_0[4215:4208] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_528[21] = buffer_data_0[4223:4216] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_528[22] = buffer_data_0[4231:4224] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_528[23] = buffer_data_0[4239:4232] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_528[24] = buffer_data_0[4247:4240] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_528 = kernel_img_mul_528[0] + kernel_img_mul_528[1] + kernel_img_mul_528[2] + 
                kernel_img_mul_528[3] + kernel_img_mul_528[4] + kernel_img_mul_528[5] + 
                kernel_img_mul_528[6] + kernel_img_mul_528[7] + kernel_img_mul_528[8] + 
                kernel_img_mul_528[9] + kernel_img_mul_528[10] + kernel_img_mul_528[11] + 
                kernel_img_mul_528[12] + kernel_img_mul_528[13] + kernel_img_mul_528[14] + 
                kernel_img_mul_528[15] + kernel_img_mul_528[16] + kernel_img_mul_528[17] + 
                kernel_img_mul_528[18] + kernel_img_mul_528[19] + kernel_img_mul_528[20] + 
                kernel_img_mul_528[21] + kernel_img_mul_528[22] + kernel_img_mul_528[23] + 
                kernel_img_mul_528[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4231:4224] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4231:4224] <= kernel_img_sum_528[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4231:4224] <= 'd0;
end

wire  [39:0]  kernel_img_mul_529[0:24];
assign kernel_img_mul_529[0] = buffer_data_4[4223:4216] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_529[1] = buffer_data_4[4231:4224] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_529[2] = buffer_data_4[4239:4232] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_529[3] = buffer_data_4[4247:4240] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_529[4] = buffer_data_4[4255:4248] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_529[5] = buffer_data_3[4223:4216] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_529[6] = buffer_data_3[4231:4224] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_529[7] = buffer_data_3[4239:4232] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_529[8] = buffer_data_3[4247:4240] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_529[9] = buffer_data_3[4255:4248] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_529[10] = buffer_data_2[4223:4216] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_529[11] = buffer_data_2[4231:4224] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_529[12] = buffer_data_2[4239:4232] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_529[13] = buffer_data_2[4247:4240] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_529[14] = buffer_data_2[4255:4248] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_529[15] = buffer_data_1[4223:4216] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_529[16] = buffer_data_1[4231:4224] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_529[17] = buffer_data_1[4239:4232] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_529[18] = buffer_data_1[4247:4240] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_529[19] = buffer_data_1[4255:4248] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_529[20] = buffer_data_0[4223:4216] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_529[21] = buffer_data_0[4231:4224] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_529[22] = buffer_data_0[4239:4232] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_529[23] = buffer_data_0[4247:4240] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_529[24] = buffer_data_0[4255:4248] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_529 = kernel_img_mul_529[0] + kernel_img_mul_529[1] + kernel_img_mul_529[2] + 
                kernel_img_mul_529[3] + kernel_img_mul_529[4] + kernel_img_mul_529[5] + 
                kernel_img_mul_529[6] + kernel_img_mul_529[7] + kernel_img_mul_529[8] + 
                kernel_img_mul_529[9] + kernel_img_mul_529[10] + kernel_img_mul_529[11] + 
                kernel_img_mul_529[12] + kernel_img_mul_529[13] + kernel_img_mul_529[14] + 
                kernel_img_mul_529[15] + kernel_img_mul_529[16] + kernel_img_mul_529[17] + 
                kernel_img_mul_529[18] + kernel_img_mul_529[19] + kernel_img_mul_529[20] + 
                kernel_img_mul_529[21] + kernel_img_mul_529[22] + kernel_img_mul_529[23] + 
                kernel_img_mul_529[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4239:4232] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4239:4232] <= kernel_img_sum_529[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4239:4232] <= 'd0;
end

wire  [39:0]  kernel_img_mul_530[0:24];
assign kernel_img_mul_530[0] = buffer_data_4[4231:4224] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_530[1] = buffer_data_4[4239:4232] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_530[2] = buffer_data_4[4247:4240] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_530[3] = buffer_data_4[4255:4248] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_530[4] = buffer_data_4[4263:4256] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_530[5] = buffer_data_3[4231:4224] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_530[6] = buffer_data_3[4239:4232] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_530[7] = buffer_data_3[4247:4240] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_530[8] = buffer_data_3[4255:4248] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_530[9] = buffer_data_3[4263:4256] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_530[10] = buffer_data_2[4231:4224] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_530[11] = buffer_data_2[4239:4232] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_530[12] = buffer_data_2[4247:4240] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_530[13] = buffer_data_2[4255:4248] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_530[14] = buffer_data_2[4263:4256] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_530[15] = buffer_data_1[4231:4224] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_530[16] = buffer_data_1[4239:4232] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_530[17] = buffer_data_1[4247:4240] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_530[18] = buffer_data_1[4255:4248] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_530[19] = buffer_data_1[4263:4256] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_530[20] = buffer_data_0[4231:4224] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_530[21] = buffer_data_0[4239:4232] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_530[22] = buffer_data_0[4247:4240] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_530[23] = buffer_data_0[4255:4248] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_530[24] = buffer_data_0[4263:4256] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_530 = kernel_img_mul_530[0] + kernel_img_mul_530[1] + kernel_img_mul_530[2] + 
                kernel_img_mul_530[3] + kernel_img_mul_530[4] + kernel_img_mul_530[5] + 
                kernel_img_mul_530[6] + kernel_img_mul_530[7] + kernel_img_mul_530[8] + 
                kernel_img_mul_530[9] + kernel_img_mul_530[10] + kernel_img_mul_530[11] + 
                kernel_img_mul_530[12] + kernel_img_mul_530[13] + kernel_img_mul_530[14] + 
                kernel_img_mul_530[15] + kernel_img_mul_530[16] + kernel_img_mul_530[17] + 
                kernel_img_mul_530[18] + kernel_img_mul_530[19] + kernel_img_mul_530[20] + 
                kernel_img_mul_530[21] + kernel_img_mul_530[22] + kernel_img_mul_530[23] + 
                kernel_img_mul_530[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4247:4240] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4247:4240] <= kernel_img_sum_530[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4247:4240] <= 'd0;
end

wire  [39:0]  kernel_img_mul_531[0:24];
assign kernel_img_mul_531[0] = buffer_data_4[4239:4232] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_531[1] = buffer_data_4[4247:4240] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_531[2] = buffer_data_4[4255:4248] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_531[3] = buffer_data_4[4263:4256] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_531[4] = buffer_data_4[4271:4264] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_531[5] = buffer_data_3[4239:4232] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_531[6] = buffer_data_3[4247:4240] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_531[7] = buffer_data_3[4255:4248] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_531[8] = buffer_data_3[4263:4256] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_531[9] = buffer_data_3[4271:4264] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_531[10] = buffer_data_2[4239:4232] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_531[11] = buffer_data_2[4247:4240] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_531[12] = buffer_data_2[4255:4248] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_531[13] = buffer_data_2[4263:4256] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_531[14] = buffer_data_2[4271:4264] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_531[15] = buffer_data_1[4239:4232] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_531[16] = buffer_data_1[4247:4240] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_531[17] = buffer_data_1[4255:4248] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_531[18] = buffer_data_1[4263:4256] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_531[19] = buffer_data_1[4271:4264] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_531[20] = buffer_data_0[4239:4232] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_531[21] = buffer_data_0[4247:4240] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_531[22] = buffer_data_0[4255:4248] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_531[23] = buffer_data_0[4263:4256] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_531[24] = buffer_data_0[4271:4264] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_531 = kernel_img_mul_531[0] + kernel_img_mul_531[1] + kernel_img_mul_531[2] + 
                kernel_img_mul_531[3] + kernel_img_mul_531[4] + kernel_img_mul_531[5] + 
                kernel_img_mul_531[6] + kernel_img_mul_531[7] + kernel_img_mul_531[8] + 
                kernel_img_mul_531[9] + kernel_img_mul_531[10] + kernel_img_mul_531[11] + 
                kernel_img_mul_531[12] + kernel_img_mul_531[13] + kernel_img_mul_531[14] + 
                kernel_img_mul_531[15] + kernel_img_mul_531[16] + kernel_img_mul_531[17] + 
                kernel_img_mul_531[18] + kernel_img_mul_531[19] + kernel_img_mul_531[20] + 
                kernel_img_mul_531[21] + kernel_img_mul_531[22] + kernel_img_mul_531[23] + 
                kernel_img_mul_531[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4255:4248] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4255:4248] <= kernel_img_sum_531[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4255:4248] <= 'd0;
end

wire  [39:0]  kernel_img_mul_532[0:24];
assign kernel_img_mul_532[0] = buffer_data_4[4247:4240] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_532[1] = buffer_data_4[4255:4248] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_532[2] = buffer_data_4[4263:4256] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_532[3] = buffer_data_4[4271:4264] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_532[4] = buffer_data_4[4279:4272] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_532[5] = buffer_data_3[4247:4240] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_532[6] = buffer_data_3[4255:4248] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_532[7] = buffer_data_3[4263:4256] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_532[8] = buffer_data_3[4271:4264] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_532[9] = buffer_data_3[4279:4272] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_532[10] = buffer_data_2[4247:4240] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_532[11] = buffer_data_2[4255:4248] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_532[12] = buffer_data_2[4263:4256] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_532[13] = buffer_data_2[4271:4264] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_532[14] = buffer_data_2[4279:4272] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_532[15] = buffer_data_1[4247:4240] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_532[16] = buffer_data_1[4255:4248] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_532[17] = buffer_data_1[4263:4256] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_532[18] = buffer_data_1[4271:4264] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_532[19] = buffer_data_1[4279:4272] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_532[20] = buffer_data_0[4247:4240] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_532[21] = buffer_data_0[4255:4248] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_532[22] = buffer_data_0[4263:4256] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_532[23] = buffer_data_0[4271:4264] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_532[24] = buffer_data_0[4279:4272] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_532 = kernel_img_mul_532[0] + kernel_img_mul_532[1] + kernel_img_mul_532[2] + 
                kernel_img_mul_532[3] + kernel_img_mul_532[4] + kernel_img_mul_532[5] + 
                kernel_img_mul_532[6] + kernel_img_mul_532[7] + kernel_img_mul_532[8] + 
                kernel_img_mul_532[9] + kernel_img_mul_532[10] + kernel_img_mul_532[11] + 
                kernel_img_mul_532[12] + kernel_img_mul_532[13] + kernel_img_mul_532[14] + 
                kernel_img_mul_532[15] + kernel_img_mul_532[16] + kernel_img_mul_532[17] + 
                kernel_img_mul_532[18] + kernel_img_mul_532[19] + kernel_img_mul_532[20] + 
                kernel_img_mul_532[21] + kernel_img_mul_532[22] + kernel_img_mul_532[23] + 
                kernel_img_mul_532[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4263:4256] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4263:4256] <= kernel_img_sum_532[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4263:4256] <= 'd0;
end

wire  [39:0]  kernel_img_mul_533[0:24];
assign kernel_img_mul_533[0] = buffer_data_4[4255:4248] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_533[1] = buffer_data_4[4263:4256] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_533[2] = buffer_data_4[4271:4264] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_533[3] = buffer_data_4[4279:4272] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_533[4] = buffer_data_4[4287:4280] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_533[5] = buffer_data_3[4255:4248] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_533[6] = buffer_data_3[4263:4256] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_533[7] = buffer_data_3[4271:4264] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_533[8] = buffer_data_3[4279:4272] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_533[9] = buffer_data_3[4287:4280] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_533[10] = buffer_data_2[4255:4248] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_533[11] = buffer_data_2[4263:4256] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_533[12] = buffer_data_2[4271:4264] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_533[13] = buffer_data_2[4279:4272] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_533[14] = buffer_data_2[4287:4280] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_533[15] = buffer_data_1[4255:4248] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_533[16] = buffer_data_1[4263:4256] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_533[17] = buffer_data_1[4271:4264] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_533[18] = buffer_data_1[4279:4272] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_533[19] = buffer_data_1[4287:4280] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_533[20] = buffer_data_0[4255:4248] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_533[21] = buffer_data_0[4263:4256] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_533[22] = buffer_data_0[4271:4264] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_533[23] = buffer_data_0[4279:4272] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_533[24] = buffer_data_0[4287:4280] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_533 = kernel_img_mul_533[0] + kernel_img_mul_533[1] + kernel_img_mul_533[2] + 
                kernel_img_mul_533[3] + kernel_img_mul_533[4] + kernel_img_mul_533[5] + 
                kernel_img_mul_533[6] + kernel_img_mul_533[7] + kernel_img_mul_533[8] + 
                kernel_img_mul_533[9] + kernel_img_mul_533[10] + kernel_img_mul_533[11] + 
                kernel_img_mul_533[12] + kernel_img_mul_533[13] + kernel_img_mul_533[14] + 
                kernel_img_mul_533[15] + kernel_img_mul_533[16] + kernel_img_mul_533[17] + 
                kernel_img_mul_533[18] + kernel_img_mul_533[19] + kernel_img_mul_533[20] + 
                kernel_img_mul_533[21] + kernel_img_mul_533[22] + kernel_img_mul_533[23] + 
                kernel_img_mul_533[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4271:4264] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4271:4264] <= kernel_img_sum_533[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4271:4264] <= 'd0;
end

wire  [39:0]  kernel_img_mul_534[0:24];
assign kernel_img_mul_534[0] = buffer_data_4[4263:4256] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_534[1] = buffer_data_4[4271:4264] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_534[2] = buffer_data_4[4279:4272] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_534[3] = buffer_data_4[4287:4280] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_534[4] = buffer_data_4[4295:4288] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_534[5] = buffer_data_3[4263:4256] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_534[6] = buffer_data_3[4271:4264] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_534[7] = buffer_data_3[4279:4272] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_534[8] = buffer_data_3[4287:4280] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_534[9] = buffer_data_3[4295:4288] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_534[10] = buffer_data_2[4263:4256] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_534[11] = buffer_data_2[4271:4264] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_534[12] = buffer_data_2[4279:4272] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_534[13] = buffer_data_2[4287:4280] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_534[14] = buffer_data_2[4295:4288] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_534[15] = buffer_data_1[4263:4256] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_534[16] = buffer_data_1[4271:4264] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_534[17] = buffer_data_1[4279:4272] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_534[18] = buffer_data_1[4287:4280] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_534[19] = buffer_data_1[4295:4288] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_534[20] = buffer_data_0[4263:4256] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_534[21] = buffer_data_0[4271:4264] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_534[22] = buffer_data_0[4279:4272] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_534[23] = buffer_data_0[4287:4280] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_534[24] = buffer_data_0[4295:4288] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_534 = kernel_img_mul_534[0] + kernel_img_mul_534[1] + kernel_img_mul_534[2] + 
                kernel_img_mul_534[3] + kernel_img_mul_534[4] + kernel_img_mul_534[5] + 
                kernel_img_mul_534[6] + kernel_img_mul_534[7] + kernel_img_mul_534[8] + 
                kernel_img_mul_534[9] + kernel_img_mul_534[10] + kernel_img_mul_534[11] + 
                kernel_img_mul_534[12] + kernel_img_mul_534[13] + kernel_img_mul_534[14] + 
                kernel_img_mul_534[15] + kernel_img_mul_534[16] + kernel_img_mul_534[17] + 
                kernel_img_mul_534[18] + kernel_img_mul_534[19] + kernel_img_mul_534[20] + 
                kernel_img_mul_534[21] + kernel_img_mul_534[22] + kernel_img_mul_534[23] + 
                kernel_img_mul_534[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4279:4272] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4279:4272] <= kernel_img_sum_534[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4279:4272] <= 'd0;
end

wire  [39:0]  kernel_img_mul_535[0:24];
assign kernel_img_mul_535[0] = buffer_data_4[4271:4264] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_535[1] = buffer_data_4[4279:4272] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_535[2] = buffer_data_4[4287:4280] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_535[3] = buffer_data_4[4295:4288] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_535[4] = buffer_data_4[4303:4296] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_535[5] = buffer_data_3[4271:4264] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_535[6] = buffer_data_3[4279:4272] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_535[7] = buffer_data_3[4287:4280] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_535[8] = buffer_data_3[4295:4288] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_535[9] = buffer_data_3[4303:4296] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_535[10] = buffer_data_2[4271:4264] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_535[11] = buffer_data_2[4279:4272] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_535[12] = buffer_data_2[4287:4280] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_535[13] = buffer_data_2[4295:4288] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_535[14] = buffer_data_2[4303:4296] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_535[15] = buffer_data_1[4271:4264] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_535[16] = buffer_data_1[4279:4272] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_535[17] = buffer_data_1[4287:4280] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_535[18] = buffer_data_1[4295:4288] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_535[19] = buffer_data_1[4303:4296] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_535[20] = buffer_data_0[4271:4264] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_535[21] = buffer_data_0[4279:4272] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_535[22] = buffer_data_0[4287:4280] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_535[23] = buffer_data_0[4295:4288] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_535[24] = buffer_data_0[4303:4296] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_535 = kernel_img_mul_535[0] + kernel_img_mul_535[1] + kernel_img_mul_535[2] + 
                kernel_img_mul_535[3] + kernel_img_mul_535[4] + kernel_img_mul_535[5] + 
                kernel_img_mul_535[6] + kernel_img_mul_535[7] + kernel_img_mul_535[8] + 
                kernel_img_mul_535[9] + kernel_img_mul_535[10] + kernel_img_mul_535[11] + 
                kernel_img_mul_535[12] + kernel_img_mul_535[13] + kernel_img_mul_535[14] + 
                kernel_img_mul_535[15] + kernel_img_mul_535[16] + kernel_img_mul_535[17] + 
                kernel_img_mul_535[18] + kernel_img_mul_535[19] + kernel_img_mul_535[20] + 
                kernel_img_mul_535[21] + kernel_img_mul_535[22] + kernel_img_mul_535[23] + 
                kernel_img_mul_535[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4287:4280] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4287:4280] <= kernel_img_sum_535[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4287:4280] <= 'd0;
end

wire  [39:0]  kernel_img_mul_536[0:24];
assign kernel_img_mul_536[0] = buffer_data_4[4279:4272] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_536[1] = buffer_data_4[4287:4280] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_536[2] = buffer_data_4[4295:4288] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_536[3] = buffer_data_4[4303:4296] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_536[4] = buffer_data_4[4311:4304] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_536[5] = buffer_data_3[4279:4272] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_536[6] = buffer_data_3[4287:4280] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_536[7] = buffer_data_3[4295:4288] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_536[8] = buffer_data_3[4303:4296] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_536[9] = buffer_data_3[4311:4304] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_536[10] = buffer_data_2[4279:4272] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_536[11] = buffer_data_2[4287:4280] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_536[12] = buffer_data_2[4295:4288] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_536[13] = buffer_data_2[4303:4296] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_536[14] = buffer_data_2[4311:4304] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_536[15] = buffer_data_1[4279:4272] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_536[16] = buffer_data_1[4287:4280] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_536[17] = buffer_data_1[4295:4288] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_536[18] = buffer_data_1[4303:4296] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_536[19] = buffer_data_1[4311:4304] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_536[20] = buffer_data_0[4279:4272] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_536[21] = buffer_data_0[4287:4280] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_536[22] = buffer_data_0[4295:4288] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_536[23] = buffer_data_0[4303:4296] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_536[24] = buffer_data_0[4311:4304] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_536 = kernel_img_mul_536[0] + kernel_img_mul_536[1] + kernel_img_mul_536[2] + 
                kernel_img_mul_536[3] + kernel_img_mul_536[4] + kernel_img_mul_536[5] + 
                kernel_img_mul_536[6] + kernel_img_mul_536[7] + kernel_img_mul_536[8] + 
                kernel_img_mul_536[9] + kernel_img_mul_536[10] + kernel_img_mul_536[11] + 
                kernel_img_mul_536[12] + kernel_img_mul_536[13] + kernel_img_mul_536[14] + 
                kernel_img_mul_536[15] + kernel_img_mul_536[16] + kernel_img_mul_536[17] + 
                kernel_img_mul_536[18] + kernel_img_mul_536[19] + kernel_img_mul_536[20] + 
                kernel_img_mul_536[21] + kernel_img_mul_536[22] + kernel_img_mul_536[23] + 
                kernel_img_mul_536[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4295:4288] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4295:4288] <= kernel_img_sum_536[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4295:4288] <= 'd0;
end

wire  [39:0]  kernel_img_mul_537[0:24];
assign kernel_img_mul_537[0] = buffer_data_4[4287:4280] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_537[1] = buffer_data_4[4295:4288] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_537[2] = buffer_data_4[4303:4296] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_537[3] = buffer_data_4[4311:4304] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_537[4] = buffer_data_4[4319:4312] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_537[5] = buffer_data_3[4287:4280] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_537[6] = buffer_data_3[4295:4288] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_537[7] = buffer_data_3[4303:4296] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_537[8] = buffer_data_3[4311:4304] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_537[9] = buffer_data_3[4319:4312] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_537[10] = buffer_data_2[4287:4280] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_537[11] = buffer_data_2[4295:4288] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_537[12] = buffer_data_2[4303:4296] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_537[13] = buffer_data_2[4311:4304] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_537[14] = buffer_data_2[4319:4312] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_537[15] = buffer_data_1[4287:4280] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_537[16] = buffer_data_1[4295:4288] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_537[17] = buffer_data_1[4303:4296] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_537[18] = buffer_data_1[4311:4304] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_537[19] = buffer_data_1[4319:4312] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_537[20] = buffer_data_0[4287:4280] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_537[21] = buffer_data_0[4295:4288] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_537[22] = buffer_data_0[4303:4296] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_537[23] = buffer_data_0[4311:4304] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_537[24] = buffer_data_0[4319:4312] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_537 = kernel_img_mul_537[0] + kernel_img_mul_537[1] + kernel_img_mul_537[2] + 
                kernel_img_mul_537[3] + kernel_img_mul_537[4] + kernel_img_mul_537[5] + 
                kernel_img_mul_537[6] + kernel_img_mul_537[7] + kernel_img_mul_537[8] + 
                kernel_img_mul_537[9] + kernel_img_mul_537[10] + kernel_img_mul_537[11] + 
                kernel_img_mul_537[12] + kernel_img_mul_537[13] + kernel_img_mul_537[14] + 
                kernel_img_mul_537[15] + kernel_img_mul_537[16] + kernel_img_mul_537[17] + 
                kernel_img_mul_537[18] + kernel_img_mul_537[19] + kernel_img_mul_537[20] + 
                kernel_img_mul_537[21] + kernel_img_mul_537[22] + kernel_img_mul_537[23] + 
                kernel_img_mul_537[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4303:4296] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4303:4296] <= kernel_img_sum_537[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4303:4296] <= 'd0;
end

wire  [39:0]  kernel_img_mul_538[0:24];
assign kernel_img_mul_538[0] = buffer_data_4[4295:4288] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_538[1] = buffer_data_4[4303:4296] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_538[2] = buffer_data_4[4311:4304] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_538[3] = buffer_data_4[4319:4312] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_538[4] = buffer_data_4[4327:4320] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_538[5] = buffer_data_3[4295:4288] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_538[6] = buffer_data_3[4303:4296] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_538[7] = buffer_data_3[4311:4304] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_538[8] = buffer_data_3[4319:4312] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_538[9] = buffer_data_3[4327:4320] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_538[10] = buffer_data_2[4295:4288] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_538[11] = buffer_data_2[4303:4296] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_538[12] = buffer_data_2[4311:4304] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_538[13] = buffer_data_2[4319:4312] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_538[14] = buffer_data_2[4327:4320] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_538[15] = buffer_data_1[4295:4288] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_538[16] = buffer_data_1[4303:4296] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_538[17] = buffer_data_1[4311:4304] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_538[18] = buffer_data_1[4319:4312] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_538[19] = buffer_data_1[4327:4320] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_538[20] = buffer_data_0[4295:4288] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_538[21] = buffer_data_0[4303:4296] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_538[22] = buffer_data_0[4311:4304] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_538[23] = buffer_data_0[4319:4312] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_538[24] = buffer_data_0[4327:4320] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_538 = kernel_img_mul_538[0] + kernel_img_mul_538[1] + kernel_img_mul_538[2] + 
                kernel_img_mul_538[3] + kernel_img_mul_538[4] + kernel_img_mul_538[5] + 
                kernel_img_mul_538[6] + kernel_img_mul_538[7] + kernel_img_mul_538[8] + 
                kernel_img_mul_538[9] + kernel_img_mul_538[10] + kernel_img_mul_538[11] + 
                kernel_img_mul_538[12] + kernel_img_mul_538[13] + kernel_img_mul_538[14] + 
                kernel_img_mul_538[15] + kernel_img_mul_538[16] + kernel_img_mul_538[17] + 
                kernel_img_mul_538[18] + kernel_img_mul_538[19] + kernel_img_mul_538[20] + 
                kernel_img_mul_538[21] + kernel_img_mul_538[22] + kernel_img_mul_538[23] + 
                kernel_img_mul_538[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4311:4304] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4311:4304] <= kernel_img_sum_538[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4311:4304] <= 'd0;
end

wire  [39:0]  kernel_img_mul_539[0:24];
assign kernel_img_mul_539[0] = buffer_data_4[4303:4296] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_539[1] = buffer_data_4[4311:4304] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_539[2] = buffer_data_4[4319:4312] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_539[3] = buffer_data_4[4327:4320] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_539[4] = buffer_data_4[4335:4328] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_539[5] = buffer_data_3[4303:4296] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_539[6] = buffer_data_3[4311:4304] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_539[7] = buffer_data_3[4319:4312] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_539[8] = buffer_data_3[4327:4320] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_539[9] = buffer_data_3[4335:4328] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_539[10] = buffer_data_2[4303:4296] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_539[11] = buffer_data_2[4311:4304] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_539[12] = buffer_data_2[4319:4312] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_539[13] = buffer_data_2[4327:4320] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_539[14] = buffer_data_2[4335:4328] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_539[15] = buffer_data_1[4303:4296] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_539[16] = buffer_data_1[4311:4304] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_539[17] = buffer_data_1[4319:4312] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_539[18] = buffer_data_1[4327:4320] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_539[19] = buffer_data_1[4335:4328] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_539[20] = buffer_data_0[4303:4296] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_539[21] = buffer_data_0[4311:4304] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_539[22] = buffer_data_0[4319:4312] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_539[23] = buffer_data_0[4327:4320] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_539[24] = buffer_data_0[4335:4328] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_539 = kernel_img_mul_539[0] + kernel_img_mul_539[1] + kernel_img_mul_539[2] + 
                kernel_img_mul_539[3] + kernel_img_mul_539[4] + kernel_img_mul_539[5] + 
                kernel_img_mul_539[6] + kernel_img_mul_539[7] + kernel_img_mul_539[8] + 
                kernel_img_mul_539[9] + kernel_img_mul_539[10] + kernel_img_mul_539[11] + 
                kernel_img_mul_539[12] + kernel_img_mul_539[13] + kernel_img_mul_539[14] + 
                kernel_img_mul_539[15] + kernel_img_mul_539[16] + kernel_img_mul_539[17] + 
                kernel_img_mul_539[18] + kernel_img_mul_539[19] + kernel_img_mul_539[20] + 
                kernel_img_mul_539[21] + kernel_img_mul_539[22] + kernel_img_mul_539[23] + 
                kernel_img_mul_539[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4319:4312] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4319:4312] <= kernel_img_sum_539[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4319:4312] <= 'd0;
end

wire  [39:0]  kernel_img_mul_540[0:24];
assign kernel_img_mul_540[0] = buffer_data_4[4311:4304] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_540[1] = buffer_data_4[4319:4312] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_540[2] = buffer_data_4[4327:4320] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_540[3] = buffer_data_4[4335:4328] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_540[4] = buffer_data_4[4343:4336] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_540[5] = buffer_data_3[4311:4304] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_540[6] = buffer_data_3[4319:4312] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_540[7] = buffer_data_3[4327:4320] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_540[8] = buffer_data_3[4335:4328] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_540[9] = buffer_data_3[4343:4336] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_540[10] = buffer_data_2[4311:4304] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_540[11] = buffer_data_2[4319:4312] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_540[12] = buffer_data_2[4327:4320] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_540[13] = buffer_data_2[4335:4328] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_540[14] = buffer_data_2[4343:4336] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_540[15] = buffer_data_1[4311:4304] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_540[16] = buffer_data_1[4319:4312] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_540[17] = buffer_data_1[4327:4320] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_540[18] = buffer_data_1[4335:4328] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_540[19] = buffer_data_1[4343:4336] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_540[20] = buffer_data_0[4311:4304] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_540[21] = buffer_data_0[4319:4312] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_540[22] = buffer_data_0[4327:4320] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_540[23] = buffer_data_0[4335:4328] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_540[24] = buffer_data_0[4343:4336] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_540 = kernel_img_mul_540[0] + kernel_img_mul_540[1] + kernel_img_mul_540[2] + 
                kernel_img_mul_540[3] + kernel_img_mul_540[4] + kernel_img_mul_540[5] + 
                kernel_img_mul_540[6] + kernel_img_mul_540[7] + kernel_img_mul_540[8] + 
                kernel_img_mul_540[9] + kernel_img_mul_540[10] + kernel_img_mul_540[11] + 
                kernel_img_mul_540[12] + kernel_img_mul_540[13] + kernel_img_mul_540[14] + 
                kernel_img_mul_540[15] + kernel_img_mul_540[16] + kernel_img_mul_540[17] + 
                kernel_img_mul_540[18] + kernel_img_mul_540[19] + kernel_img_mul_540[20] + 
                kernel_img_mul_540[21] + kernel_img_mul_540[22] + kernel_img_mul_540[23] + 
                kernel_img_mul_540[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4327:4320] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4327:4320] <= kernel_img_sum_540[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4327:4320] <= 'd0;
end

wire  [39:0]  kernel_img_mul_541[0:24];
assign kernel_img_mul_541[0] = buffer_data_4[4319:4312] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_541[1] = buffer_data_4[4327:4320] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_541[2] = buffer_data_4[4335:4328] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_541[3] = buffer_data_4[4343:4336] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_541[4] = buffer_data_4[4351:4344] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_541[5] = buffer_data_3[4319:4312] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_541[6] = buffer_data_3[4327:4320] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_541[7] = buffer_data_3[4335:4328] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_541[8] = buffer_data_3[4343:4336] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_541[9] = buffer_data_3[4351:4344] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_541[10] = buffer_data_2[4319:4312] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_541[11] = buffer_data_2[4327:4320] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_541[12] = buffer_data_2[4335:4328] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_541[13] = buffer_data_2[4343:4336] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_541[14] = buffer_data_2[4351:4344] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_541[15] = buffer_data_1[4319:4312] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_541[16] = buffer_data_1[4327:4320] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_541[17] = buffer_data_1[4335:4328] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_541[18] = buffer_data_1[4343:4336] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_541[19] = buffer_data_1[4351:4344] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_541[20] = buffer_data_0[4319:4312] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_541[21] = buffer_data_0[4327:4320] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_541[22] = buffer_data_0[4335:4328] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_541[23] = buffer_data_0[4343:4336] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_541[24] = buffer_data_0[4351:4344] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_541 = kernel_img_mul_541[0] + kernel_img_mul_541[1] + kernel_img_mul_541[2] + 
                kernel_img_mul_541[3] + kernel_img_mul_541[4] + kernel_img_mul_541[5] + 
                kernel_img_mul_541[6] + kernel_img_mul_541[7] + kernel_img_mul_541[8] + 
                kernel_img_mul_541[9] + kernel_img_mul_541[10] + kernel_img_mul_541[11] + 
                kernel_img_mul_541[12] + kernel_img_mul_541[13] + kernel_img_mul_541[14] + 
                kernel_img_mul_541[15] + kernel_img_mul_541[16] + kernel_img_mul_541[17] + 
                kernel_img_mul_541[18] + kernel_img_mul_541[19] + kernel_img_mul_541[20] + 
                kernel_img_mul_541[21] + kernel_img_mul_541[22] + kernel_img_mul_541[23] + 
                kernel_img_mul_541[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4335:4328] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4335:4328] <= kernel_img_sum_541[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4335:4328] <= 'd0;
end

wire  [39:0]  kernel_img_mul_542[0:24];
assign kernel_img_mul_542[0] = buffer_data_4[4327:4320] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_542[1] = buffer_data_4[4335:4328] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_542[2] = buffer_data_4[4343:4336] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_542[3] = buffer_data_4[4351:4344] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_542[4] = buffer_data_4[4359:4352] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_542[5] = buffer_data_3[4327:4320] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_542[6] = buffer_data_3[4335:4328] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_542[7] = buffer_data_3[4343:4336] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_542[8] = buffer_data_3[4351:4344] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_542[9] = buffer_data_3[4359:4352] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_542[10] = buffer_data_2[4327:4320] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_542[11] = buffer_data_2[4335:4328] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_542[12] = buffer_data_2[4343:4336] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_542[13] = buffer_data_2[4351:4344] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_542[14] = buffer_data_2[4359:4352] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_542[15] = buffer_data_1[4327:4320] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_542[16] = buffer_data_1[4335:4328] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_542[17] = buffer_data_1[4343:4336] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_542[18] = buffer_data_1[4351:4344] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_542[19] = buffer_data_1[4359:4352] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_542[20] = buffer_data_0[4327:4320] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_542[21] = buffer_data_0[4335:4328] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_542[22] = buffer_data_0[4343:4336] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_542[23] = buffer_data_0[4351:4344] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_542[24] = buffer_data_0[4359:4352] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_542 = kernel_img_mul_542[0] + kernel_img_mul_542[1] + kernel_img_mul_542[2] + 
                kernel_img_mul_542[3] + kernel_img_mul_542[4] + kernel_img_mul_542[5] + 
                kernel_img_mul_542[6] + kernel_img_mul_542[7] + kernel_img_mul_542[8] + 
                kernel_img_mul_542[9] + kernel_img_mul_542[10] + kernel_img_mul_542[11] + 
                kernel_img_mul_542[12] + kernel_img_mul_542[13] + kernel_img_mul_542[14] + 
                kernel_img_mul_542[15] + kernel_img_mul_542[16] + kernel_img_mul_542[17] + 
                kernel_img_mul_542[18] + kernel_img_mul_542[19] + kernel_img_mul_542[20] + 
                kernel_img_mul_542[21] + kernel_img_mul_542[22] + kernel_img_mul_542[23] + 
                kernel_img_mul_542[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4343:4336] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4343:4336] <= kernel_img_sum_542[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4343:4336] <= 'd0;
end

wire  [39:0]  kernel_img_mul_543[0:24];
assign kernel_img_mul_543[0] = buffer_data_4[4335:4328] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_543[1] = buffer_data_4[4343:4336] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_543[2] = buffer_data_4[4351:4344] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_543[3] = buffer_data_4[4359:4352] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_543[4] = buffer_data_4[4367:4360] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_543[5] = buffer_data_3[4335:4328] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_543[6] = buffer_data_3[4343:4336] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_543[7] = buffer_data_3[4351:4344] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_543[8] = buffer_data_3[4359:4352] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_543[9] = buffer_data_3[4367:4360] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_543[10] = buffer_data_2[4335:4328] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_543[11] = buffer_data_2[4343:4336] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_543[12] = buffer_data_2[4351:4344] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_543[13] = buffer_data_2[4359:4352] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_543[14] = buffer_data_2[4367:4360] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_543[15] = buffer_data_1[4335:4328] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_543[16] = buffer_data_1[4343:4336] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_543[17] = buffer_data_1[4351:4344] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_543[18] = buffer_data_1[4359:4352] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_543[19] = buffer_data_1[4367:4360] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_543[20] = buffer_data_0[4335:4328] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_543[21] = buffer_data_0[4343:4336] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_543[22] = buffer_data_0[4351:4344] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_543[23] = buffer_data_0[4359:4352] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_543[24] = buffer_data_0[4367:4360] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_543 = kernel_img_mul_543[0] + kernel_img_mul_543[1] + kernel_img_mul_543[2] + 
                kernel_img_mul_543[3] + kernel_img_mul_543[4] + kernel_img_mul_543[5] + 
                kernel_img_mul_543[6] + kernel_img_mul_543[7] + kernel_img_mul_543[8] + 
                kernel_img_mul_543[9] + kernel_img_mul_543[10] + kernel_img_mul_543[11] + 
                kernel_img_mul_543[12] + kernel_img_mul_543[13] + kernel_img_mul_543[14] + 
                kernel_img_mul_543[15] + kernel_img_mul_543[16] + kernel_img_mul_543[17] + 
                kernel_img_mul_543[18] + kernel_img_mul_543[19] + kernel_img_mul_543[20] + 
                kernel_img_mul_543[21] + kernel_img_mul_543[22] + kernel_img_mul_543[23] + 
                kernel_img_mul_543[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4351:4344] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4351:4344] <= kernel_img_sum_543[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4351:4344] <= 'd0;
end

wire  [39:0]  kernel_img_mul_544[0:24];
assign kernel_img_mul_544[0] = buffer_data_4[4343:4336] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_544[1] = buffer_data_4[4351:4344] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_544[2] = buffer_data_4[4359:4352] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_544[3] = buffer_data_4[4367:4360] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_544[4] = buffer_data_4[4375:4368] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_544[5] = buffer_data_3[4343:4336] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_544[6] = buffer_data_3[4351:4344] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_544[7] = buffer_data_3[4359:4352] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_544[8] = buffer_data_3[4367:4360] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_544[9] = buffer_data_3[4375:4368] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_544[10] = buffer_data_2[4343:4336] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_544[11] = buffer_data_2[4351:4344] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_544[12] = buffer_data_2[4359:4352] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_544[13] = buffer_data_2[4367:4360] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_544[14] = buffer_data_2[4375:4368] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_544[15] = buffer_data_1[4343:4336] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_544[16] = buffer_data_1[4351:4344] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_544[17] = buffer_data_1[4359:4352] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_544[18] = buffer_data_1[4367:4360] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_544[19] = buffer_data_1[4375:4368] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_544[20] = buffer_data_0[4343:4336] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_544[21] = buffer_data_0[4351:4344] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_544[22] = buffer_data_0[4359:4352] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_544[23] = buffer_data_0[4367:4360] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_544[24] = buffer_data_0[4375:4368] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_544 = kernel_img_mul_544[0] + kernel_img_mul_544[1] + kernel_img_mul_544[2] + 
                kernel_img_mul_544[3] + kernel_img_mul_544[4] + kernel_img_mul_544[5] + 
                kernel_img_mul_544[6] + kernel_img_mul_544[7] + kernel_img_mul_544[8] + 
                kernel_img_mul_544[9] + kernel_img_mul_544[10] + kernel_img_mul_544[11] + 
                kernel_img_mul_544[12] + kernel_img_mul_544[13] + kernel_img_mul_544[14] + 
                kernel_img_mul_544[15] + kernel_img_mul_544[16] + kernel_img_mul_544[17] + 
                kernel_img_mul_544[18] + kernel_img_mul_544[19] + kernel_img_mul_544[20] + 
                kernel_img_mul_544[21] + kernel_img_mul_544[22] + kernel_img_mul_544[23] + 
                kernel_img_mul_544[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4359:4352] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4359:4352] <= kernel_img_sum_544[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4359:4352] <= 'd0;
end

wire  [39:0]  kernel_img_mul_545[0:24];
assign kernel_img_mul_545[0] = buffer_data_4[4351:4344] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_545[1] = buffer_data_4[4359:4352] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_545[2] = buffer_data_4[4367:4360] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_545[3] = buffer_data_4[4375:4368] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_545[4] = buffer_data_4[4383:4376] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_545[5] = buffer_data_3[4351:4344] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_545[6] = buffer_data_3[4359:4352] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_545[7] = buffer_data_3[4367:4360] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_545[8] = buffer_data_3[4375:4368] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_545[9] = buffer_data_3[4383:4376] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_545[10] = buffer_data_2[4351:4344] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_545[11] = buffer_data_2[4359:4352] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_545[12] = buffer_data_2[4367:4360] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_545[13] = buffer_data_2[4375:4368] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_545[14] = buffer_data_2[4383:4376] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_545[15] = buffer_data_1[4351:4344] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_545[16] = buffer_data_1[4359:4352] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_545[17] = buffer_data_1[4367:4360] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_545[18] = buffer_data_1[4375:4368] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_545[19] = buffer_data_1[4383:4376] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_545[20] = buffer_data_0[4351:4344] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_545[21] = buffer_data_0[4359:4352] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_545[22] = buffer_data_0[4367:4360] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_545[23] = buffer_data_0[4375:4368] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_545[24] = buffer_data_0[4383:4376] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_545 = kernel_img_mul_545[0] + kernel_img_mul_545[1] + kernel_img_mul_545[2] + 
                kernel_img_mul_545[3] + kernel_img_mul_545[4] + kernel_img_mul_545[5] + 
                kernel_img_mul_545[6] + kernel_img_mul_545[7] + kernel_img_mul_545[8] + 
                kernel_img_mul_545[9] + kernel_img_mul_545[10] + kernel_img_mul_545[11] + 
                kernel_img_mul_545[12] + kernel_img_mul_545[13] + kernel_img_mul_545[14] + 
                kernel_img_mul_545[15] + kernel_img_mul_545[16] + kernel_img_mul_545[17] + 
                kernel_img_mul_545[18] + kernel_img_mul_545[19] + kernel_img_mul_545[20] + 
                kernel_img_mul_545[21] + kernel_img_mul_545[22] + kernel_img_mul_545[23] + 
                kernel_img_mul_545[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4367:4360] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4367:4360] <= kernel_img_sum_545[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4367:4360] <= 'd0;
end

wire  [39:0]  kernel_img_mul_546[0:24];
assign kernel_img_mul_546[0] = buffer_data_4[4359:4352] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_546[1] = buffer_data_4[4367:4360] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_546[2] = buffer_data_4[4375:4368] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_546[3] = buffer_data_4[4383:4376] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_546[4] = buffer_data_4[4391:4384] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_546[5] = buffer_data_3[4359:4352] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_546[6] = buffer_data_3[4367:4360] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_546[7] = buffer_data_3[4375:4368] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_546[8] = buffer_data_3[4383:4376] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_546[9] = buffer_data_3[4391:4384] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_546[10] = buffer_data_2[4359:4352] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_546[11] = buffer_data_2[4367:4360] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_546[12] = buffer_data_2[4375:4368] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_546[13] = buffer_data_2[4383:4376] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_546[14] = buffer_data_2[4391:4384] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_546[15] = buffer_data_1[4359:4352] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_546[16] = buffer_data_1[4367:4360] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_546[17] = buffer_data_1[4375:4368] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_546[18] = buffer_data_1[4383:4376] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_546[19] = buffer_data_1[4391:4384] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_546[20] = buffer_data_0[4359:4352] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_546[21] = buffer_data_0[4367:4360] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_546[22] = buffer_data_0[4375:4368] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_546[23] = buffer_data_0[4383:4376] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_546[24] = buffer_data_0[4391:4384] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_546 = kernel_img_mul_546[0] + kernel_img_mul_546[1] + kernel_img_mul_546[2] + 
                kernel_img_mul_546[3] + kernel_img_mul_546[4] + kernel_img_mul_546[5] + 
                kernel_img_mul_546[6] + kernel_img_mul_546[7] + kernel_img_mul_546[8] + 
                kernel_img_mul_546[9] + kernel_img_mul_546[10] + kernel_img_mul_546[11] + 
                kernel_img_mul_546[12] + kernel_img_mul_546[13] + kernel_img_mul_546[14] + 
                kernel_img_mul_546[15] + kernel_img_mul_546[16] + kernel_img_mul_546[17] + 
                kernel_img_mul_546[18] + kernel_img_mul_546[19] + kernel_img_mul_546[20] + 
                kernel_img_mul_546[21] + kernel_img_mul_546[22] + kernel_img_mul_546[23] + 
                kernel_img_mul_546[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4375:4368] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4375:4368] <= kernel_img_sum_546[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4375:4368] <= 'd0;
end

wire  [39:0]  kernel_img_mul_547[0:24];
assign kernel_img_mul_547[0] = buffer_data_4[4367:4360] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_547[1] = buffer_data_4[4375:4368] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_547[2] = buffer_data_4[4383:4376] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_547[3] = buffer_data_4[4391:4384] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_547[4] = buffer_data_4[4399:4392] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_547[5] = buffer_data_3[4367:4360] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_547[6] = buffer_data_3[4375:4368] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_547[7] = buffer_data_3[4383:4376] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_547[8] = buffer_data_3[4391:4384] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_547[9] = buffer_data_3[4399:4392] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_547[10] = buffer_data_2[4367:4360] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_547[11] = buffer_data_2[4375:4368] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_547[12] = buffer_data_2[4383:4376] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_547[13] = buffer_data_2[4391:4384] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_547[14] = buffer_data_2[4399:4392] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_547[15] = buffer_data_1[4367:4360] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_547[16] = buffer_data_1[4375:4368] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_547[17] = buffer_data_1[4383:4376] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_547[18] = buffer_data_1[4391:4384] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_547[19] = buffer_data_1[4399:4392] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_547[20] = buffer_data_0[4367:4360] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_547[21] = buffer_data_0[4375:4368] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_547[22] = buffer_data_0[4383:4376] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_547[23] = buffer_data_0[4391:4384] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_547[24] = buffer_data_0[4399:4392] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_547 = kernel_img_mul_547[0] + kernel_img_mul_547[1] + kernel_img_mul_547[2] + 
                kernel_img_mul_547[3] + kernel_img_mul_547[4] + kernel_img_mul_547[5] + 
                kernel_img_mul_547[6] + kernel_img_mul_547[7] + kernel_img_mul_547[8] + 
                kernel_img_mul_547[9] + kernel_img_mul_547[10] + kernel_img_mul_547[11] + 
                kernel_img_mul_547[12] + kernel_img_mul_547[13] + kernel_img_mul_547[14] + 
                kernel_img_mul_547[15] + kernel_img_mul_547[16] + kernel_img_mul_547[17] + 
                kernel_img_mul_547[18] + kernel_img_mul_547[19] + kernel_img_mul_547[20] + 
                kernel_img_mul_547[21] + kernel_img_mul_547[22] + kernel_img_mul_547[23] + 
                kernel_img_mul_547[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4383:4376] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4383:4376] <= kernel_img_sum_547[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4383:4376] <= 'd0;
end

wire  [39:0]  kernel_img_mul_548[0:24];
assign kernel_img_mul_548[0] = buffer_data_4[4375:4368] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_548[1] = buffer_data_4[4383:4376] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_548[2] = buffer_data_4[4391:4384] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_548[3] = buffer_data_4[4399:4392] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_548[4] = buffer_data_4[4407:4400] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_548[5] = buffer_data_3[4375:4368] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_548[6] = buffer_data_3[4383:4376] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_548[7] = buffer_data_3[4391:4384] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_548[8] = buffer_data_3[4399:4392] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_548[9] = buffer_data_3[4407:4400] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_548[10] = buffer_data_2[4375:4368] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_548[11] = buffer_data_2[4383:4376] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_548[12] = buffer_data_2[4391:4384] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_548[13] = buffer_data_2[4399:4392] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_548[14] = buffer_data_2[4407:4400] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_548[15] = buffer_data_1[4375:4368] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_548[16] = buffer_data_1[4383:4376] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_548[17] = buffer_data_1[4391:4384] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_548[18] = buffer_data_1[4399:4392] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_548[19] = buffer_data_1[4407:4400] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_548[20] = buffer_data_0[4375:4368] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_548[21] = buffer_data_0[4383:4376] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_548[22] = buffer_data_0[4391:4384] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_548[23] = buffer_data_0[4399:4392] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_548[24] = buffer_data_0[4407:4400] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_548 = kernel_img_mul_548[0] + kernel_img_mul_548[1] + kernel_img_mul_548[2] + 
                kernel_img_mul_548[3] + kernel_img_mul_548[4] + kernel_img_mul_548[5] + 
                kernel_img_mul_548[6] + kernel_img_mul_548[7] + kernel_img_mul_548[8] + 
                kernel_img_mul_548[9] + kernel_img_mul_548[10] + kernel_img_mul_548[11] + 
                kernel_img_mul_548[12] + kernel_img_mul_548[13] + kernel_img_mul_548[14] + 
                kernel_img_mul_548[15] + kernel_img_mul_548[16] + kernel_img_mul_548[17] + 
                kernel_img_mul_548[18] + kernel_img_mul_548[19] + kernel_img_mul_548[20] + 
                kernel_img_mul_548[21] + kernel_img_mul_548[22] + kernel_img_mul_548[23] + 
                kernel_img_mul_548[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4391:4384] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4391:4384] <= kernel_img_sum_548[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4391:4384] <= 'd0;
end

wire  [39:0]  kernel_img_mul_549[0:24];
assign kernel_img_mul_549[0] = buffer_data_4[4383:4376] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_549[1] = buffer_data_4[4391:4384] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_549[2] = buffer_data_4[4399:4392] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_549[3] = buffer_data_4[4407:4400] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_549[4] = buffer_data_4[4415:4408] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_549[5] = buffer_data_3[4383:4376] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_549[6] = buffer_data_3[4391:4384] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_549[7] = buffer_data_3[4399:4392] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_549[8] = buffer_data_3[4407:4400] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_549[9] = buffer_data_3[4415:4408] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_549[10] = buffer_data_2[4383:4376] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_549[11] = buffer_data_2[4391:4384] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_549[12] = buffer_data_2[4399:4392] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_549[13] = buffer_data_2[4407:4400] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_549[14] = buffer_data_2[4415:4408] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_549[15] = buffer_data_1[4383:4376] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_549[16] = buffer_data_1[4391:4384] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_549[17] = buffer_data_1[4399:4392] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_549[18] = buffer_data_1[4407:4400] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_549[19] = buffer_data_1[4415:4408] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_549[20] = buffer_data_0[4383:4376] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_549[21] = buffer_data_0[4391:4384] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_549[22] = buffer_data_0[4399:4392] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_549[23] = buffer_data_0[4407:4400] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_549[24] = buffer_data_0[4415:4408] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_549 = kernel_img_mul_549[0] + kernel_img_mul_549[1] + kernel_img_mul_549[2] + 
                kernel_img_mul_549[3] + kernel_img_mul_549[4] + kernel_img_mul_549[5] + 
                kernel_img_mul_549[6] + kernel_img_mul_549[7] + kernel_img_mul_549[8] + 
                kernel_img_mul_549[9] + kernel_img_mul_549[10] + kernel_img_mul_549[11] + 
                kernel_img_mul_549[12] + kernel_img_mul_549[13] + kernel_img_mul_549[14] + 
                kernel_img_mul_549[15] + kernel_img_mul_549[16] + kernel_img_mul_549[17] + 
                kernel_img_mul_549[18] + kernel_img_mul_549[19] + kernel_img_mul_549[20] + 
                kernel_img_mul_549[21] + kernel_img_mul_549[22] + kernel_img_mul_549[23] + 
                kernel_img_mul_549[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4399:4392] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4399:4392] <= kernel_img_sum_549[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4399:4392] <= 'd0;
end

wire  [39:0]  kernel_img_mul_550[0:24];
assign kernel_img_mul_550[0] = buffer_data_4[4391:4384] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_550[1] = buffer_data_4[4399:4392] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_550[2] = buffer_data_4[4407:4400] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_550[3] = buffer_data_4[4415:4408] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_550[4] = buffer_data_4[4423:4416] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_550[5] = buffer_data_3[4391:4384] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_550[6] = buffer_data_3[4399:4392] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_550[7] = buffer_data_3[4407:4400] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_550[8] = buffer_data_3[4415:4408] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_550[9] = buffer_data_3[4423:4416] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_550[10] = buffer_data_2[4391:4384] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_550[11] = buffer_data_2[4399:4392] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_550[12] = buffer_data_2[4407:4400] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_550[13] = buffer_data_2[4415:4408] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_550[14] = buffer_data_2[4423:4416] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_550[15] = buffer_data_1[4391:4384] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_550[16] = buffer_data_1[4399:4392] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_550[17] = buffer_data_1[4407:4400] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_550[18] = buffer_data_1[4415:4408] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_550[19] = buffer_data_1[4423:4416] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_550[20] = buffer_data_0[4391:4384] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_550[21] = buffer_data_0[4399:4392] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_550[22] = buffer_data_0[4407:4400] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_550[23] = buffer_data_0[4415:4408] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_550[24] = buffer_data_0[4423:4416] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_550 = kernel_img_mul_550[0] + kernel_img_mul_550[1] + kernel_img_mul_550[2] + 
                kernel_img_mul_550[3] + kernel_img_mul_550[4] + kernel_img_mul_550[5] + 
                kernel_img_mul_550[6] + kernel_img_mul_550[7] + kernel_img_mul_550[8] + 
                kernel_img_mul_550[9] + kernel_img_mul_550[10] + kernel_img_mul_550[11] + 
                kernel_img_mul_550[12] + kernel_img_mul_550[13] + kernel_img_mul_550[14] + 
                kernel_img_mul_550[15] + kernel_img_mul_550[16] + kernel_img_mul_550[17] + 
                kernel_img_mul_550[18] + kernel_img_mul_550[19] + kernel_img_mul_550[20] + 
                kernel_img_mul_550[21] + kernel_img_mul_550[22] + kernel_img_mul_550[23] + 
                kernel_img_mul_550[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4407:4400] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4407:4400] <= kernel_img_sum_550[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4407:4400] <= 'd0;
end

wire  [39:0]  kernel_img_mul_551[0:24];
assign kernel_img_mul_551[0] = buffer_data_4[4399:4392] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_551[1] = buffer_data_4[4407:4400] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_551[2] = buffer_data_4[4415:4408] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_551[3] = buffer_data_4[4423:4416] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_551[4] = buffer_data_4[4431:4424] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_551[5] = buffer_data_3[4399:4392] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_551[6] = buffer_data_3[4407:4400] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_551[7] = buffer_data_3[4415:4408] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_551[8] = buffer_data_3[4423:4416] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_551[9] = buffer_data_3[4431:4424] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_551[10] = buffer_data_2[4399:4392] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_551[11] = buffer_data_2[4407:4400] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_551[12] = buffer_data_2[4415:4408] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_551[13] = buffer_data_2[4423:4416] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_551[14] = buffer_data_2[4431:4424] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_551[15] = buffer_data_1[4399:4392] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_551[16] = buffer_data_1[4407:4400] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_551[17] = buffer_data_1[4415:4408] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_551[18] = buffer_data_1[4423:4416] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_551[19] = buffer_data_1[4431:4424] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_551[20] = buffer_data_0[4399:4392] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_551[21] = buffer_data_0[4407:4400] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_551[22] = buffer_data_0[4415:4408] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_551[23] = buffer_data_0[4423:4416] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_551[24] = buffer_data_0[4431:4424] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_551 = kernel_img_mul_551[0] + kernel_img_mul_551[1] + kernel_img_mul_551[2] + 
                kernel_img_mul_551[3] + kernel_img_mul_551[4] + kernel_img_mul_551[5] + 
                kernel_img_mul_551[6] + kernel_img_mul_551[7] + kernel_img_mul_551[8] + 
                kernel_img_mul_551[9] + kernel_img_mul_551[10] + kernel_img_mul_551[11] + 
                kernel_img_mul_551[12] + kernel_img_mul_551[13] + kernel_img_mul_551[14] + 
                kernel_img_mul_551[15] + kernel_img_mul_551[16] + kernel_img_mul_551[17] + 
                kernel_img_mul_551[18] + kernel_img_mul_551[19] + kernel_img_mul_551[20] + 
                kernel_img_mul_551[21] + kernel_img_mul_551[22] + kernel_img_mul_551[23] + 
                kernel_img_mul_551[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4415:4408] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4415:4408] <= kernel_img_sum_551[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4415:4408] <= 'd0;
end

wire  [39:0]  kernel_img_mul_552[0:24];
assign kernel_img_mul_552[0] = buffer_data_4[4407:4400] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_552[1] = buffer_data_4[4415:4408] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_552[2] = buffer_data_4[4423:4416] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_552[3] = buffer_data_4[4431:4424] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_552[4] = buffer_data_4[4439:4432] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_552[5] = buffer_data_3[4407:4400] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_552[6] = buffer_data_3[4415:4408] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_552[7] = buffer_data_3[4423:4416] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_552[8] = buffer_data_3[4431:4424] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_552[9] = buffer_data_3[4439:4432] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_552[10] = buffer_data_2[4407:4400] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_552[11] = buffer_data_2[4415:4408] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_552[12] = buffer_data_2[4423:4416] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_552[13] = buffer_data_2[4431:4424] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_552[14] = buffer_data_2[4439:4432] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_552[15] = buffer_data_1[4407:4400] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_552[16] = buffer_data_1[4415:4408] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_552[17] = buffer_data_1[4423:4416] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_552[18] = buffer_data_1[4431:4424] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_552[19] = buffer_data_1[4439:4432] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_552[20] = buffer_data_0[4407:4400] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_552[21] = buffer_data_0[4415:4408] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_552[22] = buffer_data_0[4423:4416] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_552[23] = buffer_data_0[4431:4424] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_552[24] = buffer_data_0[4439:4432] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_552 = kernel_img_mul_552[0] + kernel_img_mul_552[1] + kernel_img_mul_552[2] + 
                kernel_img_mul_552[3] + kernel_img_mul_552[4] + kernel_img_mul_552[5] + 
                kernel_img_mul_552[6] + kernel_img_mul_552[7] + kernel_img_mul_552[8] + 
                kernel_img_mul_552[9] + kernel_img_mul_552[10] + kernel_img_mul_552[11] + 
                kernel_img_mul_552[12] + kernel_img_mul_552[13] + kernel_img_mul_552[14] + 
                kernel_img_mul_552[15] + kernel_img_mul_552[16] + kernel_img_mul_552[17] + 
                kernel_img_mul_552[18] + kernel_img_mul_552[19] + kernel_img_mul_552[20] + 
                kernel_img_mul_552[21] + kernel_img_mul_552[22] + kernel_img_mul_552[23] + 
                kernel_img_mul_552[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4423:4416] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4423:4416] <= kernel_img_sum_552[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4423:4416] <= 'd0;
end

wire  [39:0]  kernel_img_mul_553[0:24];
assign kernel_img_mul_553[0] = buffer_data_4[4415:4408] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_553[1] = buffer_data_4[4423:4416] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_553[2] = buffer_data_4[4431:4424] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_553[3] = buffer_data_4[4439:4432] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_553[4] = buffer_data_4[4447:4440] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_553[5] = buffer_data_3[4415:4408] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_553[6] = buffer_data_3[4423:4416] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_553[7] = buffer_data_3[4431:4424] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_553[8] = buffer_data_3[4439:4432] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_553[9] = buffer_data_3[4447:4440] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_553[10] = buffer_data_2[4415:4408] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_553[11] = buffer_data_2[4423:4416] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_553[12] = buffer_data_2[4431:4424] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_553[13] = buffer_data_2[4439:4432] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_553[14] = buffer_data_2[4447:4440] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_553[15] = buffer_data_1[4415:4408] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_553[16] = buffer_data_1[4423:4416] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_553[17] = buffer_data_1[4431:4424] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_553[18] = buffer_data_1[4439:4432] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_553[19] = buffer_data_1[4447:4440] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_553[20] = buffer_data_0[4415:4408] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_553[21] = buffer_data_0[4423:4416] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_553[22] = buffer_data_0[4431:4424] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_553[23] = buffer_data_0[4439:4432] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_553[24] = buffer_data_0[4447:4440] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_553 = kernel_img_mul_553[0] + kernel_img_mul_553[1] + kernel_img_mul_553[2] + 
                kernel_img_mul_553[3] + kernel_img_mul_553[4] + kernel_img_mul_553[5] + 
                kernel_img_mul_553[6] + kernel_img_mul_553[7] + kernel_img_mul_553[8] + 
                kernel_img_mul_553[9] + kernel_img_mul_553[10] + kernel_img_mul_553[11] + 
                kernel_img_mul_553[12] + kernel_img_mul_553[13] + kernel_img_mul_553[14] + 
                kernel_img_mul_553[15] + kernel_img_mul_553[16] + kernel_img_mul_553[17] + 
                kernel_img_mul_553[18] + kernel_img_mul_553[19] + kernel_img_mul_553[20] + 
                kernel_img_mul_553[21] + kernel_img_mul_553[22] + kernel_img_mul_553[23] + 
                kernel_img_mul_553[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4431:4424] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4431:4424] <= kernel_img_sum_553[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4431:4424] <= 'd0;
end

wire  [39:0]  kernel_img_mul_554[0:24];
assign kernel_img_mul_554[0] = buffer_data_4[4423:4416] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_554[1] = buffer_data_4[4431:4424] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_554[2] = buffer_data_4[4439:4432] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_554[3] = buffer_data_4[4447:4440] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_554[4] = buffer_data_4[4455:4448] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_554[5] = buffer_data_3[4423:4416] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_554[6] = buffer_data_3[4431:4424] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_554[7] = buffer_data_3[4439:4432] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_554[8] = buffer_data_3[4447:4440] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_554[9] = buffer_data_3[4455:4448] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_554[10] = buffer_data_2[4423:4416] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_554[11] = buffer_data_2[4431:4424] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_554[12] = buffer_data_2[4439:4432] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_554[13] = buffer_data_2[4447:4440] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_554[14] = buffer_data_2[4455:4448] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_554[15] = buffer_data_1[4423:4416] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_554[16] = buffer_data_1[4431:4424] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_554[17] = buffer_data_1[4439:4432] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_554[18] = buffer_data_1[4447:4440] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_554[19] = buffer_data_1[4455:4448] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_554[20] = buffer_data_0[4423:4416] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_554[21] = buffer_data_0[4431:4424] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_554[22] = buffer_data_0[4439:4432] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_554[23] = buffer_data_0[4447:4440] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_554[24] = buffer_data_0[4455:4448] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_554 = kernel_img_mul_554[0] + kernel_img_mul_554[1] + kernel_img_mul_554[2] + 
                kernel_img_mul_554[3] + kernel_img_mul_554[4] + kernel_img_mul_554[5] + 
                kernel_img_mul_554[6] + kernel_img_mul_554[7] + kernel_img_mul_554[8] + 
                kernel_img_mul_554[9] + kernel_img_mul_554[10] + kernel_img_mul_554[11] + 
                kernel_img_mul_554[12] + kernel_img_mul_554[13] + kernel_img_mul_554[14] + 
                kernel_img_mul_554[15] + kernel_img_mul_554[16] + kernel_img_mul_554[17] + 
                kernel_img_mul_554[18] + kernel_img_mul_554[19] + kernel_img_mul_554[20] + 
                kernel_img_mul_554[21] + kernel_img_mul_554[22] + kernel_img_mul_554[23] + 
                kernel_img_mul_554[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4439:4432] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4439:4432] <= kernel_img_sum_554[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4439:4432] <= 'd0;
end

wire  [39:0]  kernel_img_mul_555[0:24];
assign kernel_img_mul_555[0] = buffer_data_4[4431:4424] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_555[1] = buffer_data_4[4439:4432] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_555[2] = buffer_data_4[4447:4440] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_555[3] = buffer_data_4[4455:4448] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_555[4] = buffer_data_4[4463:4456] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_555[5] = buffer_data_3[4431:4424] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_555[6] = buffer_data_3[4439:4432] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_555[7] = buffer_data_3[4447:4440] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_555[8] = buffer_data_3[4455:4448] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_555[9] = buffer_data_3[4463:4456] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_555[10] = buffer_data_2[4431:4424] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_555[11] = buffer_data_2[4439:4432] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_555[12] = buffer_data_2[4447:4440] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_555[13] = buffer_data_2[4455:4448] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_555[14] = buffer_data_2[4463:4456] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_555[15] = buffer_data_1[4431:4424] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_555[16] = buffer_data_1[4439:4432] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_555[17] = buffer_data_1[4447:4440] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_555[18] = buffer_data_1[4455:4448] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_555[19] = buffer_data_1[4463:4456] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_555[20] = buffer_data_0[4431:4424] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_555[21] = buffer_data_0[4439:4432] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_555[22] = buffer_data_0[4447:4440] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_555[23] = buffer_data_0[4455:4448] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_555[24] = buffer_data_0[4463:4456] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_555 = kernel_img_mul_555[0] + kernel_img_mul_555[1] + kernel_img_mul_555[2] + 
                kernel_img_mul_555[3] + kernel_img_mul_555[4] + kernel_img_mul_555[5] + 
                kernel_img_mul_555[6] + kernel_img_mul_555[7] + kernel_img_mul_555[8] + 
                kernel_img_mul_555[9] + kernel_img_mul_555[10] + kernel_img_mul_555[11] + 
                kernel_img_mul_555[12] + kernel_img_mul_555[13] + kernel_img_mul_555[14] + 
                kernel_img_mul_555[15] + kernel_img_mul_555[16] + kernel_img_mul_555[17] + 
                kernel_img_mul_555[18] + kernel_img_mul_555[19] + kernel_img_mul_555[20] + 
                kernel_img_mul_555[21] + kernel_img_mul_555[22] + kernel_img_mul_555[23] + 
                kernel_img_mul_555[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4447:4440] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4447:4440] <= kernel_img_sum_555[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4447:4440] <= 'd0;
end

wire  [39:0]  kernel_img_mul_556[0:24];
assign kernel_img_mul_556[0] = buffer_data_4[4439:4432] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_556[1] = buffer_data_4[4447:4440] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_556[2] = buffer_data_4[4455:4448] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_556[3] = buffer_data_4[4463:4456] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_556[4] = buffer_data_4[4471:4464] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_556[5] = buffer_data_3[4439:4432] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_556[6] = buffer_data_3[4447:4440] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_556[7] = buffer_data_3[4455:4448] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_556[8] = buffer_data_3[4463:4456] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_556[9] = buffer_data_3[4471:4464] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_556[10] = buffer_data_2[4439:4432] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_556[11] = buffer_data_2[4447:4440] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_556[12] = buffer_data_2[4455:4448] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_556[13] = buffer_data_2[4463:4456] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_556[14] = buffer_data_2[4471:4464] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_556[15] = buffer_data_1[4439:4432] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_556[16] = buffer_data_1[4447:4440] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_556[17] = buffer_data_1[4455:4448] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_556[18] = buffer_data_1[4463:4456] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_556[19] = buffer_data_1[4471:4464] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_556[20] = buffer_data_0[4439:4432] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_556[21] = buffer_data_0[4447:4440] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_556[22] = buffer_data_0[4455:4448] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_556[23] = buffer_data_0[4463:4456] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_556[24] = buffer_data_0[4471:4464] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_556 = kernel_img_mul_556[0] + kernel_img_mul_556[1] + kernel_img_mul_556[2] + 
                kernel_img_mul_556[3] + kernel_img_mul_556[4] + kernel_img_mul_556[5] + 
                kernel_img_mul_556[6] + kernel_img_mul_556[7] + kernel_img_mul_556[8] + 
                kernel_img_mul_556[9] + kernel_img_mul_556[10] + kernel_img_mul_556[11] + 
                kernel_img_mul_556[12] + kernel_img_mul_556[13] + kernel_img_mul_556[14] + 
                kernel_img_mul_556[15] + kernel_img_mul_556[16] + kernel_img_mul_556[17] + 
                kernel_img_mul_556[18] + kernel_img_mul_556[19] + kernel_img_mul_556[20] + 
                kernel_img_mul_556[21] + kernel_img_mul_556[22] + kernel_img_mul_556[23] + 
                kernel_img_mul_556[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4455:4448] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4455:4448] <= kernel_img_sum_556[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4455:4448] <= 'd0;
end

wire  [39:0]  kernel_img_mul_557[0:24];
assign kernel_img_mul_557[0] = buffer_data_4[4447:4440] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_557[1] = buffer_data_4[4455:4448] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_557[2] = buffer_data_4[4463:4456] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_557[3] = buffer_data_4[4471:4464] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_557[4] = buffer_data_4[4479:4472] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_557[5] = buffer_data_3[4447:4440] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_557[6] = buffer_data_3[4455:4448] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_557[7] = buffer_data_3[4463:4456] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_557[8] = buffer_data_3[4471:4464] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_557[9] = buffer_data_3[4479:4472] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_557[10] = buffer_data_2[4447:4440] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_557[11] = buffer_data_2[4455:4448] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_557[12] = buffer_data_2[4463:4456] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_557[13] = buffer_data_2[4471:4464] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_557[14] = buffer_data_2[4479:4472] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_557[15] = buffer_data_1[4447:4440] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_557[16] = buffer_data_1[4455:4448] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_557[17] = buffer_data_1[4463:4456] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_557[18] = buffer_data_1[4471:4464] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_557[19] = buffer_data_1[4479:4472] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_557[20] = buffer_data_0[4447:4440] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_557[21] = buffer_data_0[4455:4448] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_557[22] = buffer_data_0[4463:4456] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_557[23] = buffer_data_0[4471:4464] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_557[24] = buffer_data_0[4479:4472] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_557 = kernel_img_mul_557[0] + kernel_img_mul_557[1] + kernel_img_mul_557[2] + 
                kernel_img_mul_557[3] + kernel_img_mul_557[4] + kernel_img_mul_557[5] + 
                kernel_img_mul_557[6] + kernel_img_mul_557[7] + kernel_img_mul_557[8] + 
                kernel_img_mul_557[9] + kernel_img_mul_557[10] + kernel_img_mul_557[11] + 
                kernel_img_mul_557[12] + kernel_img_mul_557[13] + kernel_img_mul_557[14] + 
                kernel_img_mul_557[15] + kernel_img_mul_557[16] + kernel_img_mul_557[17] + 
                kernel_img_mul_557[18] + kernel_img_mul_557[19] + kernel_img_mul_557[20] + 
                kernel_img_mul_557[21] + kernel_img_mul_557[22] + kernel_img_mul_557[23] + 
                kernel_img_mul_557[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4463:4456] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4463:4456] <= kernel_img_sum_557[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4463:4456] <= 'd0;
end

wire  [39:0]  kernel_img_mul_558[0:24];
assign kernel_img_mul_558[0] = buffer_data_4[4455:4448] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_558[1] = buffer_data_4[4463:4456] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_558[2] = buffer_data_4[4471:4464] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_558[3] = buffer_data_4[4479:4472] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_558[4] = buffer_data_4[4487:4480] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_558[5] = buffer_data_3[4455:4448] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_558[6] = buffer_data_3[4463:4456] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_558[7] = buffer_data_3[4471:4464] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_558[8] = buffer_data_3[4479:4472] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_558[9] = buffer_data_3[4487:4480] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_558[10] = buffer_data_2[4455:4448] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_558[11] = buffer_data_2[4463:4456] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_558[12] = buffer_data_2[4471:4464] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_558[13] = buffer_data_2[4479:4472] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_558[14] = buffer_data_2[4487:4480] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_558[15] = buffer_data_1[4455:4448] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_558[16] = buffer_data_1[4463:4456] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_558[17] = buffer_data_1[4471:4464] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_558[18] = buffer_data_1[4479:4472] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_558[19] = buffer_data_1[4487:4480] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_558[20] = buffer_data_0[4455:4448] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_558[21] = buffer_data_0[4463:4456] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_558[22] = buffer_data_0[4471:4464] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_558[23] = buffer_data_0[4479:4472] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_558[24] = buffer_data_0[4487:4480] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_558 = kernel_img_mul_558[0] + kernel_img_mul_558[1] + kernel_img_mul_558[2] + 
                kernel_img_mul_558[3] + kernel_img_mul_558[4] + kernel_img_mul_558[5] + 
                kernel_img_mul_558[6] + kernel_img_mul_558[7] + kernel_img_mul_558[8] + 
                kernel_img_mul_558[9] + kernel_img_mul_558[10] + kernel_img_mul_558[11] + 
                kernel_img_mul_558[12] + kernel_img_mul_558[13] + kernel_img_mul_558[14] + 
                kernel_img_mul_558[15] + kernel_img_mul_558[16] + kernel_img_mul_558[17] + 
                kernel_img_mul_558[18] + kernel_img_mul_558[19] + kernel_img_mul_558[20] + 
                kernel_img_mul_558[21] + kernel_img_mul_558[22] + kernel_img_mul_558[23] + 
                kernel_img_mul_558[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4471:4464] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4471:4464] <= kernel_img_sum_558[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4471:4464] <= 'd0;
end

wire  [39:0]  kernel_img_mul_559[0:24];
assign kernel_img_mul_559[0] = buffer_data_4[4463:4456] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_559[1] = buffer_data_4[4471:4464] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_559[2] = buffer_data_4[4479:4472] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_559[3] = buffer_data_4[4487:4480] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_559[4] = buffer_data_4[4495:4488] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_559[5] = buffer_data_3[4463:4456] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_559[6] = buffer_data_3[4471:4464] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_559[7] = buffer_data_3[4479:4472] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_559[8] = buffer_data_3[4487:4480] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_559[9] = buffer_data_3[4495:4488] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_559[10] = buffer_data_2[4463:4456] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_559[11] = buffer_data_2[4471:4464] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_559[12] = buffer_data_2[4479:4472] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_559[13] = buffer_data_2[4487:4480] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_559[14] = buffer_data_2[4495:4488] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_559[15] = buffer_data_1[4463:4456] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_559[16] = buffer_data_1[4471:4464] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_559[17] = buffer_data_1[4479:4472] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_559[18] = buffer_data_1[4487:4480] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_559[19] = buffer_data_1[4495:4488] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_559[20] = buffer_data_0[4463:4456] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_559[21] = buffer_data_0[4471:4464] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_559[22] = buffer_data_0[4479:4472] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_559[23] = buffer_data_0[4487:4480] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_559[24] = buffer_data_0[4495:4488] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_559 = kernel_img_mul_559[0] + kernel_img_mul_559[1] + kernel_img_mul_559[2] + 
                kernel_img_mul_559[3] + kernel_img_mul_559[4] + kernel_img_mul_559[5] + 
                kernel_img_mul_559[6] + kernel_img_mul_559[7] + kernel_img_mul_559[8] + 
                kernel_img_mul_559[9] + kernel_img_mul_559[10] + kernel_img_mul_559[11] + 
                kernel_img_mul_559[12] + kernel_img_mul_559[13] + kernel_img_mul_559[14] + 
                kernel_img_mul_559[15] + kernel_img_mul_559[16] + kernel_img_mul_559[17] + 
                kernel_img_mul_559[18] + kernel_img_mul_559[19] + kernel_img_mul_559[20] + 
                kernel_img_mul_559[21] + kernel_img_mul_559[22] + kernel_img_mul_559[23] + 
                kernel_img_mul_559[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4479:4472] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4479:4472] <= kernel_img_sum_559[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4479:4472] <= 'd0;
end

wire  [39:0]  kernel_img_mul_560[0:24];
assign kernel_img_mul_560[0] = buffer_data_4[4471:4464] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_560[1] = buffer_data_4[4479:4472] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_560[2] = buffer_data_4[4487:4480] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_560[3] = buffer_data_4[4495:4488] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_560[4] = buffer_data_4[4503:4496] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_560[5] = buffer_data_3[4471:4464] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_560[6] = buffer_data_3[4479:4472] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_560[7] = buffer_data_3[4487:4480] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_560[8] = buffer_data_3[4495:4488] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_560[9] = buffer_data_3[4503:4496] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_560[10] = buffer_data_2[4471:4464] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_560[11] = buffer_data_2[4479:4472] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_560[12] = buffer_data_2[4487:4480] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_560[13] = buffer_data_2[4495:4488] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_560[14] = buffer_data_2[4503:4496] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_560[15] = buffer_data_1[4471:4464] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_560[16] = buffer_data_1[4479:4472] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_560[17] = buffer_data_1[4487:4480] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_560[18] = buffer_data_1[4495:4488] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_560[19] = buffer_data_1[4503:4496] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_560[20] = buffer_data_0[4471:4464] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_560[21] = buffer_data_0[4479:4472] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_560[22] = buffer_data_0[4487:4480] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_560[23] = buffer_data_0[4495:4488] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_560[24] = buffer_data_0[4503:4496] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_560 = kernel_img_mul_560[0] + kernel_img_mul_560[1] + kernel_img_mul_560[2] + 
                kernel_img_mul_560[3] + kernel_img_mul_560[4] + kernel_img_mul_560[5] + 
                kernel_img_mul_560[6] + kernel_img_mul_560[7] + kernel_img_mul_560[8] + 
                kernel_img_mul_560[9] + kernel_img_mul_560[10] + kernel_img_mul_560[11] + 
                kernel_img_mul_560[12] + kernel_img_mul_560[13] + kernel_img_mul_560[14] + 
                kernel_img_mul_560[15] + kernel_img_mul_560[16] + kernel_img_mul_560[17] + 
                kernel_img_mul_560[18] + kernel_img_mul_560[19] + kernel_img_mul_560[20] + 
                kernel_img_mul_560[21] + kernel_img_mul_560[22] + kernel_img_mul_560[23] + 
                kernel_img_mul_560[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4487:4480] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4487:4480] <= kernel_img_sum_560[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4487:4480] <= 'd0;
end

wire  [39:0]  kernel_img_mul_561[0:24];
assign kernel_img_mul_561[0] = buffer_data_4[4479:4472] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_561[1] = buffer_data_4[4487:4480] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_561[2] = buffer_data_4[4495:4488] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_561[3] = buffer_data_4[4503:4496] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_561[4] = buffer_data_4[4511:4504] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_561[5] = buffer_data_3[4479:4472] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_561[6] = buffer_data_3[4487:4480] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_561[7] = buffer_data_3[4495:4488] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_561[8] = buffer_data_3[4503:4496] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_561[9] = buffer_data_3[4511:4504] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_561[10] = buffer_data_2[4479:4472] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_561[11] = buffer_data_2[4487:4480] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_561[12] = buffer_data_2[4495:4488] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_561[13] = buffer_data_2[4503:4496] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_561[14] = buffer_data_2[4511:4504] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_561[15] = buffer_data_1[4479:4472] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_561[16] = buffer_data_1[4487:4480] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_561[17] = buffer_data_1[4495:4488] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_561[18] = buffer_data_1[4503:4496] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_561[19] = buffer_data_1[4511:4504] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_561[20] = buffer_data_0[4479:4472] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_561[21] = buffer_data_0[4487:4480] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_561[22] = buffer_data_0[4495:4488] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_561[23] = buffer_data_0[4503:4496] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_561[24] = buffer_data_0[4511:4504] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_561 = kernel_img_mul_561[0] + kernel_img_mul_561[1] + kernel_img_mul_561[2] + 
                kernel_img_mul_561[3] + kernel_img_mul_561[4] + kernel_img_mul_561[5] + 
                kernel_img_mul_561[6] + kernel_img_mul_561[7] + kernel_img_mul_561[8] + 
                kernel_img_mul_561[9] + kernel_img_mul_561[10] + kernel_img_mul_561[11] + 
                kernel_img_mul_561[12] + kernel_img_mul_561[13] + kernel_img_mul_561[14] + 
                kernel_img_mul_561[15] + kernel_img_mul_561[16] + kernel_img_mul_561[17] + 
                kernel_img_mul_561[18] + kernel_img_mul_561[19] + kernel_img_mul_561[20] + 
                kernel_img_mul_561[21] + kernel_img_mul_561[22] + kernel_img_mul_561[23] + 
                kernel_img_mul_561[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4495:4488] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4495:4488] <= kernel_img_sum_561[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4495:4488] <= 'd0;
end

wire  [39:0]  kernel_img_mul_562[0:24];
assign kernel_img_mul_562[0] = buffer_data_4[4487:4480] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_562[1] = buffer_data_4[4495:4488] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_562[2] = buffer_data_4[4503:4496] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_562[3] = buffer_data_4[4511:4504] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_562[4] = buffer_data_4[4519:4512] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_562[5] = buffer_data_3[4487:4480] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_562[6] = buffer_data_3[4495:4488] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_562[7] = buffer_data_3[4503:4496] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_562[8] = buffer_data_3[4511:4504] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_562[9] = buffer_data_3[4519:4512] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_562[10] = buffer_data_2[4487:4480] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_562[11] = buffer_data_2[4495:4488] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_562[12] = buffer_data_2[4503:4496] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_562[13] = buffer_data_2[4511:4504] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_562[14] = buffer_data_2[4519:4512] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_562[15] = buffer_data_1[4487:4480] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_562[16] = buffer_data_1[4495:4488] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_562[17] = buffer_data_1[4503:4496] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_562[18] = buffer_data_1[4511:4504] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_562[19] = buffer_data_1[4519:4512] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_562[20] = buffer_data_0[4487:4480] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_562[21] = buffer_data_0[4495:4488] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_562[22] = buffer_data_0[4503:4496] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_562[23] = buffer_data_0[4511:4504] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_562[24] = buffer_data_0[4519:4512] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_562 = kernel_img_mul_562[0] + kernel_img_mul_562[1] + kernel_img_mul_562[2] + 
                kernel_img_mul_562[3] + kernel_img_mul_562[4] + kernel_img_mul_562[5] + 
                kernel_img_mul_562[6] + kernel_img_mul_562[7] + kernel_img_mul_562[8] + 
                kernel_img_mul_562[9] + kernel_img_mul_562[10] + kernel_img_mul_562[11] + 
                kernel_img_mul_562[12] + kernel_img_mul_562[13] + kernel_img_mul_562[14] + 
                kernel_img_mul_562[15] + kernel_img_mul_562[16] + kernel_img_mul_562[17] + 
                kernel_img_mul_562[18] + kernel_img_mul_562[19] + kernel_img_mul_562[20] + 
                kernel_img_mul_562[21] + kernel_img_mul_562[22] + kernel_img_mul_562[23] + 
                kernel_img_mul_562[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4503:4496] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4503:4496] <= kernel_img_sum_562[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4503:4496] <= 'd0;
end

wire  [39:0]  kernel_img_mul_563[0:24];
assign kernel_img_mul_563[0] = buffer_data_4[4495:4488] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_563[1] = buffer_data_4[4503:4496] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_563[2] = buffer_data_4[4511:4504] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_563[3] = buffer_data_4[4519:4512] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_563[4] = buffer_data_4[4527:4520] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_563[5] = buffer_data_3[4495:4488] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_563[6] = buffer_data_3[4503:4496] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_563[7] = buffer_data_3[4511:4504] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_563[8] = buffer_data_3[4519:4512] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_563[9] = buffer_data_3[4527:4520] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_563[10] = buffer_data_2[4495:4488] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_563[11] = buffer_data_2[4503:4496] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_563[12] = buffer_data_2[4511:4504] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_563[13] = buffer_data_2[4519:4512] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_563[14] = buffer_data_2[4527:4520] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_563[15] = buffer_data_1[4495:4488] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_563[16] = buffer_data_1[4503:4496] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_563[17] = buffer_data_1[4511:4504] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_563[18] = buffer_data_1[4519:4512] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_563[19] = buffer_data_1[4527:4520] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_563[20] = buffer_data_0[4495:4488] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_563[21] = buffer_data_0[4503:4496] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_563[22] = buffer_data_0[4511:4504] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_563[23] = buffer_data_0[4519:4512] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_563[24] = buffer_data_0[4527:4520] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_563 = kernel_img_mul_563[0] + kernel_img_mul_563[1] + kernel_img_mul_563[2] + 
                kernel_img_mul_563[3] + kernel_img_mul_563[4] + kernel_img_mul_563[5] + 
                kernel_img_mul_563[6] + kernel_img_mul_563[7] + kernel_img_mul_563[8] + 
                kernel_img_mul_563[9] + kernel_img_mul_563[10] + kernel_img_mul_563[11] + 
                kernel_img_mul_563[12] + kernel_img_mul_563[13] + kernel_img_mul_563[14] + 
                kernel_img_mul_563[15] + kernel_img_mul_563[16] + kernel_img_mul_563[17] + 
                kernel_img_mul_563[18] + kernel_img_mul_563[19] + kernel_img_mul_563[20] + 
                kernel_img_mul_563[21] + kernel_img_mul_563[22] + kernel_img_mul_563[23] + 
                kernel_img_mul_563[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4511:4504] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4511:4504] <= kernel_img_sum_563[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4511:4504] <= 'd0;
end

wire  [39:0]  kernel_img_mul_564[0:24];
assign kernel_img_mul_564[0] = buffer_data_4[4503:4496] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_564[1] = buffer_data_4[4511:4504] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_564[2] = buffer_data_4[4519:4512] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_564[3] = buffer_data_4[4527:4520] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_564[4] = buffer_data_4[4535:4528] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_564[5] = buffer_data_3[4503:4496] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_564[6] = buffer_data_3[4511:4504] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_564[7] = buffer_data_3[4519:4512] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_564[8] = buffer_data_3[4527:4520] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_564[9] = buffer_data_3[4535:4528] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_564[10] = buffer_data_2[4503:4496] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_564[11] = buffer_data_2[4511:4504] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_564[12] = buffer_data_2[4519:4512] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_564[13] = buffer_data_2[4527:4520] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_564[14] = buffer_data_2[4535:4528] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_564[15] = buffer_data_1[4503:4496] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_564[16] = buffer_data_1[4511:4504] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_564[17] = buffer_data_1[4519:4512] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_564[18] = buffer_data_1[4527:4520] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_564[19] = buffer_data_1[4535:4528] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_564[20] = buffer_data_0[4503:4496] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_564[21] = buffer_data_0[4511:4504] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_564[22] = buffer_data_0[4519:4512] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_564[23] = buffer_data_0[4527:4520] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_564[24] = buffer_data_0[4535:4528] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_564 = kernel_img_mul_564[0] + kernel_img_mul_564[1] + kernel_img_mul_564[2] + 
                kernel_img_mul_564[3] + kernel_img_mul_564[4] + kernel_img_mul_564[5] + 
                kernel_img_mul_564[6] + kernel_img_mul_564[7] + kernel_img_mul_564[8] + 
                kernel_img_mul_564[9] + kernel_img_mul_564[10] + kernel_img_mul_564[11] + 
                kernel_img_mul_564[12] + kernel_img_mul_564[13] + kernel_img_mul_564[14] + 
                kernel_img_mul_564[15] + kernel_img_mul_564[16] + kernel_img_mul_564[17] + 
                kernel_img_mul_564[18] + kernel_img_mul_564[19] + kernel_img_mul_564[20] + 
                kernel_img_mul_564[21] + kernel_img_mul_564[22] + kernel_img_mul_564[23] + 
                kernel_img_mul_564[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4519:4512] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4519:4512] <= kernel_img_sum_564[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4519:4512] <= 'd0;
end

wire  [39:0]  kernel_img_mul_565[0:24];
assign kernel_img_mul_565[0] = buffer_data_4[4511:4504] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_565[1] = buffer_data_4[4519:4512] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_565[2] = buffer_data_4[4527:4520] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_565[3] = buffer_data_4[4535:4528] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_565[4] = buffer_data_4[4543:4536] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_565[5] = buffer_data_3[4511:4504] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_565[6] = buffer_data_3[4519:4512] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_565[7] = buffer_data_3[4527:4520] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_565[8] = buffer_data_3[4535:4528] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_565[9] = buffer_data_3[4543:4536] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_565[10] = buffer_data_2[4511:4504] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_565[11] = buffer_data_2[4519:4512] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_565[12] = buffer_data_2[4527:4520] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_565[13] = buffer_data_2[4535:4528] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_565[14] = buffer_data_2[4543:4536] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_565[15] = buffer_data_1[4511:4504] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_565[16] = buffer_data_1[4519:4512] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_565[17] = buffer_data_1[4527:4520] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_565[18] = buffer_data_1[4535:4528] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_565[19] = buffer_data_1[4543:4536] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_565[20] = buffer_data_0[4511:4504] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_565[21] = buffer_data_0[4519:4512] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_565[22] = buffer_data_0[4527:4520] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_565[23] = buffer_data_0[4535:4528] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_565[24] = buffer_data_0[4543:4536] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_565 = kernel_img_mul_565[0] + kernel_img_mul_565[1] + kernel_img_mul_565[2] + 
                kernel_img_mul_565[3] + kernel_img_mul_565[4] + kernel_img_mul_565[5] + 
                kernel_img_mul_565[6] + kernel_img_mul_565[7] + kernel_img_mul_565[8] + 
                kernel_img_mul_565[9] + kernel_img_mul_565[10] + kernel_img_mul_565[11] + 
                kernel_img_mul_565[12] + kernel_img_mul_565[13] + kernel_img_mul_565[14] + 
                kernel_img_mul_565[15] + kernel_img_mul_565[16] + kernel_img_mul_565[17] + 
                kernel_img_mul_565[18] + kernel_img_mul_565[19] + kernel_img_mul_565[20] + 
                kernel_img_mul_565[21] + kernel_img_mul_565[22] + kernel_img_mul_565[23] + 
                kernel_img_mul_565[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4527:4520] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4527:4520] <= kernel_img_sum_565[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4527:4520] <= 'd0;
end

wire  [39:0]  kernel_img_mul_566[0:24];
assign kernel_img_mul_566[0] = buffer_data_4[4519:4512] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_566[1] = buffer_data_4[4527:4520] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_566[2] = buffer_data_4[4535:4528] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_566[3] = buffer_data_4[4543:4536] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_566[4] = buffer_data_4[4551:4544] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_566[5] = buffer_data_3[4519:4512] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_566[6] = buffer_data_3[4527:4520] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_566[7] = buffer_data_3[4535:4528] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_566[8] = buffer_data_3[4543:4536] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_566[9] = buffer_data_3[4551:4544] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_566[10] = buffer_data_2[4519:4512] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_566[11] = buffer_data_2[4527:4520] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_566[12] = buffer_data_2[4535:4528] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_566[13] = buffer_data_2[4543:4536] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_566[14] = buffer_data_2[4551:4544] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_566[15] = buffer_data_1[4519:4512] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_566[16] = buffer_data_1[4527:4520] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_566[17] = buffer_data_1[4535:4528] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_566[18] = buffer_data_1[4543:4536] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_566[19] = buffer_data_1[4551:4544] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_566[20] = buffer_data_0[4519:4512] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_566[21] = buffer_data_0[4527:4520] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_566[22] = buffer_data_0[4535:4528] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_566[23] = buffer_data_0[4543:4536] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_566[24] = buffer_data_0[4551:4544] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_566 = kernel_img_mul_566[0] + kernel_img_mul_566[1] + kernel_img_mul_566[2] + 
                kernel_img_mul_566[3] + kernel_img_mul_566[4] + kernel_img_mul_566[5] + 
                kernel_img_mul_566[6] + kernel_img_mul_566[7] + kernel_img_mul_566[8] + 
                kernel_img_mul_566[9] + kernel_img_mul_566[10] + kernel_img_mul_566[11] + 
                kernel_img_mul_566[12] + kernel_img_mul_566[13] + kernel_img_mul_566[14] + 
                kernel_img_mul_566[15] + kernel_img_mul_566[16] + kernel_img_mul_566[17] + 
                kernel_img_mul_566[18] + kernel_img_mul_566[19] + kernel_img_mul_566[20] + 
                kernel_img_mul_566[21] + kernel_img_mul_566[22] + kernel_img_mul_566[23] + 
                kernel_img_mul_566[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4535:4528] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4535:4528] <= kernel_img_sum_566[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4535:4528] <= 'd0;
end

wire  [39:0]  kernel_img_mul_567[0:24];
assign kernel_img_mul_567[0] = buffer_data_4[4527:4520] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_567[1] = buffer_data_4[4535:4528] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_567[2] = buffer_data_4[4543:4536] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_567[3] = buffer_data_4[4551:4544] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_567[4] = buffer_data_4[4559:4552] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_567[5] = buffer_data_3[4527:4520] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_567[6] = buffer_data_3[4535:4528] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_567[7] = buffer_data_3[4543:4536] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_567[8] = buffer_data_3[4551:4544] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_567[9] = buffer_data_3[4559:4552] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_567[10] = buffer_data_2[4527:4520] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_567[11] = buffer_data_2[4535:4528] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_567[12] = buffer_data_2[4543:4536] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_567[13] = buffer_data_2[4551:4544] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_567[14] = buffer_data_2[4559:4552] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_567[15] = buffer_data_1[4527:4520] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_567[16] = buffer_data_1[4535:4528] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_567[17] = buffer_data_1[4543:4536] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_567[18] = buffer_data_1[4551:4544] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_567[19] = buffer_data_1[4559:4552] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_567[20] = buffer_data_0[4527:4520] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_567[21] = buffer_data_0[4535:4528] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_567[22] = buffer_data_0[4543:4536] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_567[23] = buffer_data_0[4551:4544] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_567[24] = buffer_data_0[4559:4552] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_567 = kernel_img_mul_567[0] + kernel_img_mul_567[1] + kernel_img_mul_567[2] + 
                kernel_img_mul_567[3] + kernel_img_mul_567[4] + kernel_img_mul_567[5] + 
                kernel_img_mul_567[6] + kernel_img_mul_567[7] + kernel_img_mul_567[8] + 
                kernel_img_mul_567[9] + kernel_img_mul_567[10] + kernel_img_mul_567[11] + 
                kernel_img_mul_567[12] + kernel_img_mul_567[13] + kernel_img_mul_567[14] + 
                kernel_img_mul_567[15] + kernel_img_mul_567[16] + kernel_img_mul_567[17] + 
                kernel_img_mul_567[18] + kernel_img_mul_567[19] + kernel_img_mul_567[20] + 
                kernel_img_mul_567[21] + kernel_img_mul_567[22] + kernel_img_mul_567[23] + 
                kernel_img_mul_567[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4543:4536] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4543:4536] <= kernel_img_sum_567[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4543:4536] <= 'd0;
end

wire  [39:0]  kernel_img_mul_568[0:24];
assign kernel_img_mul_568[0] = buffer_data_4[4535:4528] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_568[1] = buffer_data_4[4543:4536] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_568[2] = buffer_data_4[4551:4544] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_568[3] = buffer_data_4[4559:4552] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_568[4] = buffer_data_4[4567:4560] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_568[5] = buffer_data_3[4535:4528] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_568[6] = buffer_data_3[4543:4536] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_568[7] = buffer_data_3[4551:4544] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_568[8] = buffer_data_3[4559:4552] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_568[9] = buffer_data_3[4567:4560] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_568[10] = buffer_data_2[4535:4528] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_568[11] = buffer_data_2[4543:4536] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_568[12] = buffer_data_2[4551:4544] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_568[13] = buffer_data_2[4559:4552] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_568[14] = buffer_data_2[4567:4560] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_568[15] = buffer_data_1[4535:4528] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_568[16] = buffer_data_1[4543:4536] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_568[17] = buffer_data_1[4551:4544] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_568[18] = buffer_data_1[4559:4552] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_568[19] = buffer_data_1[4567:4560] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_568[20] = buffer_data_0[4535:4528] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_568[21] = buffer_data_0[4543:4536] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_568[22] = buffer_data_0[4551:4544] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_568[23] = buffer_data_0[4559:4552] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_568[24] = buffer_data_0[4567:4560] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_568 = kernel_img_mul_568[0] + kernel_img_mul_568[1] + kernel_img_mul_568[2] + 
                kernel_img_mul_568[3] + kernel_img_mul_568[4] + kernel_img_mul_568[5] + 
                kernel_img_mul_568[6] + kernel_img_mul_568[7] + kernel_img_mul_568[8] + 
                kernel_img_mul_568[9] + kernel_img_mul_568[10] + kernel_img_mul_568[11] + 
                kernel_img_mul_568[12] + kernel_img_mul_568[13] + kernel_img_mul_568[14] + 
                kernel_img_mul_568[15] + kernel_img_mul_568[16] + kernel_img_mul_568[17] + 
                kernel_img_mul_568[18] + kernel_img_mul_568[19] + kernel_img_mul_568[20] + 
                kernel_img_mul_568[21] + kernel_img_mul_568[22] + kernel_img_mul_568[23] + 
                kernel_img_mul_568[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4551:4544] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4551:4544] <= kernel_img_sum_568[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4551:4544] <= 'd0;
end

wire  [39:0]  kernel_img_mul_569[0:24];
assign kernel_img_mul_569[0] = buffer_data_4[4543:4536] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_569[1] = buffer_data_4[4551:4544] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_569[2] = buffer_data_4[4559:4552] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_569[3] = buffer_data_4[4567:4560] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_569[4] = buffer_data_4[4575:4568] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_569[5] = buffer_data_3[4543:4536] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_569[6] = buffer_data_3[4551:4544] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_569[7] = buffer_data_3[4559:4552] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_569[8] = buffer_data_3[4567:4560] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_569[9] = buffer_data_3[4575:4568] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_569[10] = buffer_data_2[4543:4536] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_569[11] = buffer_data_2[4551:4544] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_569[12] = buffer_data_2[4559:4552] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_569[13] = buffer_data_2[4567:4560] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_569[14] = buffer_data_2[4575:4568] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_569[15] = buffer_data_1[4543:4536] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_569[16] = buffer_data_1[4551:4544] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_569[17] = buffer_data_1[4559:4552] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_569[18] = buffer_data_1[4567:4560] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_569[19] = buffer_data_1[4575:4568] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_569[20] = buffer_data_0[4543:4536] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_569[21] = buffer_data_0[4551:4544] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_569[22] = buffer_data_0[4559:4552] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_569[23] = buffer_data_0[4567:4560] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_569[24] = buffer_data_0[4575:4568] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_569 = kernel_img_mul_569[0] + kernel_img_mul_569[1] + kernel_img_mul_569[2] + 
                kernel_img_mul_569[3] + kernel_img_mul_569[4] + kernel_img_mul_569[5] + 
                kernel_img_mul_569[6] + kernel_img_mul_569[7] + kernel_img_mul_569[8] + 
                kernel_img_mul_569[9] + kernel_img_mul_569[10] + kernel_img_mul_569[11] + 
                kernel_img_mul_569[12] + kernel_img_mul_569[13] + kernel_img_mul_569[14] + 
                kernel_img_mul_569[15] + kernel_img_mul_569[16] + kernel_img_mul_569[17] + 
                kernel_img_mul_569[18] + kernel_img_mul_569[19] + kernel_img_mul_569[20] + 
                kernel_img_mul_569[21] + kernel_img_mul_569[22] + kernel_img_mul_569[23] + 
                kernel_img_mul_569[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4559:4552] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4559:4552] <= kernel_img_sum_569[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4559:4552] <= 'd0;
end

wire  [39:0]  kernel_img_mul_570[0:24];
assign kernel_img_mul_570[0] = buffer_data_4[4551:4544] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_570[1] = buffer_data_4[4559:4552] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_570[2] = buffer_data_4[4567:4560] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_570[3] = buffer_data_4[4575:4568] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_570[4] = buffer_data_4[4583:4576] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_570[5] = buffer_data_3[4551:4544] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_570[6] = buffer_data_3[4559:4552] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_570[7] = buffer_data_3[4567:4560] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_570[8] = buffer_data_3[4575:4568] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_570[9] = buffer_data_3[4583:4576] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_570[10] = buffer_data_2[4551:4544] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_570[11] = buffer_data_2[4559:4552] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_570[12] = buffer_data_2[4567:4560] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_570[13] = buffer_data_2[4575:4568] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_570[14] = buffer_data_2[4583:4576] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_570[15] = buffer_data_1[4551:4544] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_570[16] = buffer_data_1[4559:4552] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_570[17] = buffer_data_1[4567:4560] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_570[18] = buffer_data_1[4575:4568] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_570[19] = buffer_data_1[4583:4576] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_570[20] = buffer_data_0[4551:4544] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_570[21] = buffer_data_0[4559:4552] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_570[22] = buffer_data_0[4567:4560] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_570[23] = buffer_data_0[4575:4568] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_570[24] = buffer_data_0[4583:4576] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_570 = kernel_img_mul_570[0] + kernel_img_mul_570[1] + kernel_img_mul_570[2] + 
                kernel_img_mul_570[3] + kernel_img_mul_570[4] + kernel_img_mul_570[5] + 
                kernel_img_mul_570[6] + kernel_img_mul_570[7] + kernel_img_mul_570[8] + 
                kernel_img_mul_570[9] + kernel_img_mul_570[10] + kernel_img_mul_570[11] + 
                kernel_img_mul_570[12] + kernel_img_mul_570[13] + kernel_img_mul_570[14] + 
                kernel_img_mul_570[15] + kernel_img_mul_570[16] + kernel_img_mul_570[17] + 
                kernel_img_mul_570[18] + kernel_img_mul_570[19] + kernel_img_mul_570[20] + 
                kernel_img_mul_570[21] + kernel_img_mul_570[22] + kernel_img_mul_570[23] + 
                kernel_img_mul_570[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4567:4560] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4567:4560] <= kernel_img_sum_570[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4567:4560] <= 'd0;
end

wire  [39:0]  kernel_img_mul_571[0:24];
assign kernel_img_mul_571[0] = buffer_data_4[4559:4552] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_571[1] = buffer_data_4[4567:4560] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_571[2] = buffer_data_4[4575:4568] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_571[3] = buffer_data_4[4583:4576] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_571[4] = buffer_data_4[4591:4584] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_571[5] = buffer_data_3[4559:4552] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_571[6] = buffer_data_3[4567:4560] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_571[7] = buffer_data_3[4575:4568] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_571[8] = buffer_data_3[4583:4576] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_571[9] = buffer_data_3[4591:4584] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_571[10] = buffer_data_2[4559:4552] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_571[11] = buffer_data_2[4567:4560] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_571[12] = buffer_data_2[4575:4568] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_571[13] = buffer_data_2[4583:4576] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_571[14] = buffer_data_2[4591:4584] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_571[15] = buffer_data_1[4559:4552] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_571[16] = buffer_data_1[4567:4560] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_571[17] = buffer_data_1[4575:4568] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_571[18] = buffer_data_1[4583:4576] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_571[19] = buffer_data_1[4591:4584] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_571[20] = buffer_data_0[4559:4552] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_571[21] = buffer_data_0[4567:4560] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_571[22] = buffer_data_0[4575:4568] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_571[23] = buffer_data_0[4583:4576] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_571[24] = buffer_data_0[4591:4584] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_571 = kernel_img_mul_571[0] + kernel_img_mul_571[1] + kernel_img_mul_571[2] + 
                kernel_img_mul_571[3] + kernel_img_mul_571[4] + kernel_img_mul_571[5] + 
                kernel_img_mul_571[6] + kernel_img_mul_571[7] + kernel_img_mul_571[8] + 
                kernel_img_mul_571[9] + kernel_img_mul_571[10] + kernel_img_mul_571[11] + 
                kernel_img_mul_571[12] + kernel_img_mul_571[13] + kernel_img_mul_571[14] + 
                kernel_img_mul_571[15] + kernel_img_mul_571[16] + kernel_img_mul_571[17] + 
                kernel_img_mul_571[18] + kernel_img_mul_571[19] + kernel_img_mul_571[20] + 
                kernel_img_mul_571[21] + kernel_img_mul_571[22] + kernel_img_mul_571[23] + 
                kernel_img_mul_571[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4575:4568] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4575:4568] <= kernel_img_sum_571[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4575:4568] <= 'd0;
end

wire  [39:0]  kernel_img_mul_572[0:24];
assign kernel_img_mul_572[0] = buffer_data_4[4567:4560] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_572[1] = buffer_data_4[4575:4568] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_572[2] = buffer_data_4[4583:4576] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_572[3] = buffer_data_4[4591:4584] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_572[4] = buffer_data_4[4599:4592] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_572[5] = buffer_data_3[4567:4560] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_572[6] = buffer_data_3[4575:4568] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_572[7] = buffer_data_3[4583:4576] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_572[8] = buffer_data_3[4591:4584] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_572[9] = buffer_data_3[4599:4592] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_572[10] = buffer_data_2[4567:4560] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_572[11] = buffer_data_2[4575:4568] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_572[12] = buffer_data_2[4583:4576] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_572[13] = buffer_data_2[4591:4584] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_572[14] = buffer_data_2[4599:4592] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_572[15] = buffer_data_1[4567:4560] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_572[16] = buffer_data_1[4575:4568] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_572[17] = buffer_data_1[4583:4576] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_572[18] = buffer_data_1[4591:4584] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_572[19] = buffer_data_1[4599:4592] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_572[20] = buffer_data_0[4567:4560] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_572[21] = buffer_data_0[4575:4568] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_572[22] = buffer_data_0[4583:4576] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_572[23] = buffer_data_0[4591:4584] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_572[24] = buffer_data_0[4599:4592] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_572 = kernel_img_mul_572[0] + kernel_img_mul_572[1] + kernel_img_mul_572[2] + 
                kernel_img_mul_572[3] + kernel_img_mul_572[4] + kernel_img_mul_572[5] + 
                kernel_img_mul_572[6] + kernel_img_mul_572[7] + kernel_img_mul_572[8] + 
                kernel_img_mul_572[9] + kernel_img_mul_572[10] + kernel_img_mul_572[11] + 
                kernel_img_mul_572[12] + kernel_img_mul_572[13] + kernel_img_mul_572[14] + 
                kernel_img_mul_572[15] + kernel_img_mul_572[16] + kernel_img_mul_572[17] + 
                kernel_img_mul_572[18] + kernel_img_mul_572[19] + kernel_img_mul_572[20] + 
                kernel_img_mul_572[21] + kernel_img_mul_572[22] + kernel_img_mul_572[23] + 
                kernel_img_mul_572[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4583:4576] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4583:4576] <= kernel_img_sum_572[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4583:4576] <= 'd0;
end

wire  [39:0]  kernel_img_mul_573[0:24];
assign kernel_img_mul_573[0] = buffer_data_4[4575:4568] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_573[1] = buffer_data_4[4583:4576] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_573[2] = buffer_data_4[4591:4584] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_573[3] = buffer_data_4[4599:4592] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_573[4] = buffer_data_4[4607:4600] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_573[5] = buffer_data_3[4575:4568] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_573[6] = buffer_data_3[4583:4576] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_573[7] = buffer_data_3[4591:4584] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_573[8] = buffer_data_3[4599:4592] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_573[9] = buffer_data_3[4607:4600] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_573[10] = buffer_data_2[4575:4568] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_573[11] = buffer_data_2[4583:4576] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_573[12] = buffer_data_2[4591:4584] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_573[13] = buffer_data_2[4599:4592] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_573[14] = buffer_data_2[4607:4600] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_573[15] = buffer_data_1[4575:4568] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_573[16] = buffer_data_1[4583:4576] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_573[17] = buffer_data_1[4591:4584] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_573[18] = buffer_data_1[4599:4592] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_573[19] = buffer_data_1[4607:4600] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_573[20] = buffer_data_0[4575:4568] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_573[21] = buffer_data_0[4583:4576] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_573[22] = buffer_data_0[4591:4584] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_573[23] = buffer_data_0[4599:4592] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_573[24] = buffer_data_0[4607:4600] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_573 = kernel_img_mul_573[0] + kernel_img_mul_573[1] + kernel_img_mul_573[2] + 
                kernel_img_mul_573[3] + kernel_img_mul_573[4] + kernel_img_mul_573[5] + 
                kernel_img_mul_573[6] + kernel_img_mul_573[7] + kernel_img_mul_573[8] + 
                kernel_img_mul_573[9] + kernel_img_mul_573[10] + kernel_img_mul_573[11] + 
                kernel_img_mul_573[12] + kernel_img_mul_573[13] + kernel_img_mul_573[14] + 
                kernel_img_mul_573[15] + kernel_img_mul_573[16] + kernel_img_mul_573[17] + 
                kernel_img_mul_573[18] + kernel_img_mul_573[19] + kernel_img_mul_573[20] + 
                kernel_img_mul_573[21] + kernel_img_mul_573[22] + kernel_img_mul_573[23] + 
                kernel_img_mul_573[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4591:4584] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4591:4584] <= kernel_img_sum_573[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4591:4584] <= 'd0;
end

wire  [39:0]  kernel_img_mul_574[0:24];
assign kernel_img_mul_574[0] = buffer_data_4[4583:4576] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_574[1] = buffer_data_4[4591:4584] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_574[2] = buffer_data_4[4599:4592] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_574[3] = buffer_data_4[4607:4600] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_574[4] = buffer_data_4[4615:4608] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_574[5] = buffer_data_3[4583:4576] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_574[6] = buffer_data_3[4591:4584] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_574[7] = buffer_data_3[4599:4592] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_574[8] = buffer_data_3[4607:4600] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_574[9] = buffer_data_3[4615:4608] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_574[10] = buffer_data_2[4583:4576] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_574[11] = buffer_data_2[4591:4584] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_574[12] = buffer_data_2[4599:4592] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_574[13] = buffer_data_2[4607:4600] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_574[14] = buffer_data_2[4615:4608] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_574[15] = buffer_data_1[4583:4576] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_574[16] = buffer_data_1[4591:4584] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_574[17] = buffer_data_1[4599:4592] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_574[18] = buffer_data_1[4607:4600] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_574[19] = buffer_data_1[4615:4608] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_574[20] = buffer_data_0[4583:4576] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_574[21] = buffer_data_0[4591:4584] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_574[22] = buffer_data_0[4599:4592] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_574[23] = buffer_data_0[4607:4600] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_574[24] = buffer_data_0[4615:4608] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_574 = kernel_img_mul_574[0] + kernel_img_mul_574[1] + kernel_img_mul_574[2] + 
                kernel_img_mul_574[3] + kernel_img_mul_574[4] + kernel_img_mul_574[5] + 
                kernel_img_mul_574[6] + kernel_img_mul_574[7] + kernel_img_mul_574[8] + 
                kernel_img_mul_574[9] + kernel_img_mul_574[10] + kernel_img_mul_574[11] + 
                kernel_img_mul_574[12] + kernel_img_mul_574[13] + kernel_img_mul_574[14] + 
                kernel_img_mul_574[15] + kernel_img_mul_574[16] + kernel_img_mul_574[17] + 
                kernel_img_mul_574[18] + kernel_img_mul_574[19] + kernel_img_mul_574[20] + 
                kernel_img_mul_574[21] + kernel_img_mul_574[22] + kernel_img_mul_574[23] + 
                kernel_img_mul_574[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4599:4592] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4599:4592] <= kernel_img_sum_574[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4599:4592] <= 'd0;
end

wire  [39:0]  kernel_img_mul_575[0:24];
assign kernel_img_mul_575[0] = buffer_data_4[4591:4584] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_575[1] = buffer_data_4[4599:4592] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_575[2] = buffer_data_4[4607:4600] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_575[3] = buffer_data_4[4615:4608] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_575[4] = buffer_data_4[4623:4616] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_575[5] = buffer_data_3[4591:4584] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_575[6] = buffer_data_3[4599:4592] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_575[7] = buffer_data_3[4607:4600] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_575[8] = buffer_data_3[4615:4608] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_575[9] = buffer_data_3[4623:4616] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_575[10] = buffer_data_2[4591:4584] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_575[11] = buffer_data_2[4599:4592] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_575[12] = buffer_data_2[4607:4600] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_575[13] = buffer_data_2[4615:4608] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_575[14] = buffer_data_2[4623:4616] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_575[15] = buffer_data_1[4591:4584] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_575[16] = buffer_data_1[4599:4592] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_575[17] = buffer_data_1[4607:4600] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_575[18] = buffer_data_1[4615:4608] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_575[19] = buffer_data_1[4623:4616] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_575[20] = buffer_data_0[4591:4584] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_575[21] = buffer_data_0[4599:4592] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_575[22] = buffer_data_0[4607:4600] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_575[23] = buffer_data_0[4615:4608] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_575[24] = buffer_data_0[4623:4616] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_575 = kernel_img_mul_575[0] + kernel_img_mul_575[1] + kernel_img_mul_575[2] + 
                kernel_img_mul_575[3] + kernel_img_mul_575[4] + kernel_img_mul_575[5] + 
                kernel_img_mul_575[6] + kernel_img_mul_575[7] + kernel_img_mul_575[8] + 
                kernel_img_mul_575[9] + kernel_img_mul_575[10] + kernel_img_mul_575[11] + 
                kernel_img_mul_575[12] + kernel_img_mul_575[13] + kernel_img_mul_575[14] + 
                kernel_img_mul_575[15] + kernel_img_mul_575[16] + kernel_img_mul_575[17] + 
                kernel_img_mul_575[18] + kernel_img_mul_575[19] + kernel_img_mul_575[20] + 
                kernel_img_mul_575[21] + kernel_img_mul_575[22] + kernel_img_mul_575[23] + 
                kernel_img_mul_575[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4607:4600] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4607:4600] <= kernel_img_sum_575[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4607:4600] <= 'd0;
end

wire  [39:0]  kernel_img_mul_576[0:24];
assign kernel_img_mul_576[0] = buffer_data_4[4599:4592] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_576[1] = buffer_data_4[4607:4600] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_576[2] = buffer_data_4[4615:4608] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_576[3] = buffer_data_4[4623:4616] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_576[4] = buffer_data_4[4631:4624] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_576[5] = buffer_data_3[4599:4592] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_576[6] = buffer_data_3[4607:4600] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_576[7] = buffer_data_3[4615:4608] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_576[8] = buffer_data_3[4623:4616] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_576[9] = buffer_data_3[4631:4624] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_576[10] = buffer_data_2[4599:4592] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_576[11] = buffer_data_2[4607:4600] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_576[12] = buffer_data_2[4615:4608] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_576[13] = buffer_data_2[4623:4616] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_576[14] = buffer_data_2[4631:4624] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_576[15] = buffer_data_1[4599:4592] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_576[16] = buffer_data_1[4607:4600] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_576[17] = buffer_data_1[4615:4608] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_576[18] = buffer_data_1[4623:4616] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_576[19] = buffer_data_1[4631:4624] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_576[20] = buffer_data_0[4599:4592] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_576[21] = buffer_data_0[4607:4600] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_576[22] = buffer_data_0[4615:4608] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_576[23] = buffer_data_0[4623:4616] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_576[24] = buffer_data_0[4631:4624] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_576 = kernel_img_mul_576[0] + kernel_img_mul_576[1] + kernel_img_mul_576[2] + 
                kernel_img_mul_576[3] + kernel_img_mul_576[4] + kernel_img_mul_576[5] + 
                kernel_img_mul_576[6] + kernel_img_mul_576[7] + kernel_img_mul_576[8] + 
                kernel_img_mul_576[9] + kernel_img_mul_576[10] + kernel_img_mul_576[11] + 
                kernel_img_mul_576[12] + kernel_img_mul_576[13] + kernel_img_mul_576[14] + 
                kernel_img_mul_576[15] + kernel_img_mul_576[16] + kernel_img_mul_576[17] + 
                kernel_img_mul_576[18] + kernel_img_mul_576[19] + kernel_img_mul_576[20] + 
                kernel_img_mul_576[21] + kernel_img_mul_576[22] + kernel_img_mul_576[23] + 
                kernel_img_mul_576[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4615:4608] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4615:4608] <= kernel_img_sum_576[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4615:4608] <= 'd0;
end

wire  [39:0]  kernel_img_mul_577[0:24];
assign kernel_img_mul_577[0] = buffer_data_4[4607:4600] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_577[1] = buffer_data_4[4615:4608] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_577[2] = buffer_data_4[4623:4616] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_577[3] = buffer_data_4[4631:4624] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_577[4] = buffer_data_4[4639:4632] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_577[5] = buffer_data_3[4607:4600] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_577[6] = buffer_data_3[4615:4608] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_577[7] = buffer_data_3[4623:4616] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_577[8] = buffer_data_3[4631:4624] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_577[9] = buffer_data_3[4639:4632] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_577[10] = buffer_data_2[4607:4600] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_577[11] = buffer_data_2[4615:4608] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_577[12] = buffer_data_2[4623:4616] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_577[13] = buffer_data_2[4631:4624] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_577[14] = buffer_data_2[4639:4632] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_577[15] = buffer_data_1[4607:4600] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_577[16] = buffer_data_1[4615:4608] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_577[17] = buffer_data_1[4623:4616] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_577[18] = buffer_data_1[4631:4624] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_577[19] = buffer_data_1[4639:4632] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_577[20] = buffer_data_0[4607:4600] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_577[21] = buffer_data_0[4615:4608] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_577[22] = buffer_data_0[4623:4616] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_577[23] = buffer_data_0[4631:4624] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_577[24] = buffer_data_0[4639:4632] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_577 = kernel_img_mul_577[0] + kernel_img_mul_577[1] + kernel_img_mul_577[2] + 
                kernel_img_mul_577[3] + kernel_img_mul_577[4] + kernel_img_mul_577[5] + 
                kernel_img_mul_577[6] + kernel_img_mul_577[7] + kernel_img_mul_577[8] + 
                kernel_img_mul_577[9] + kernel_img_mul_577[10] + kernel_img_mul_577[11] + 
                kernel_img_mul_577[12] + kernel_img_mul_577[13] + kernel_img_mul_577[14] + 
                kernel_img_mul_577[15] + kernel_img_mul_577[16] + kernel_img_mul_577[17] + 
                kernel_img_mul_577[18] + kernel_img_mul_577[19] + kernel_img_mul_577[20] + 
                kernel_img_mul_577[21] + kernel_img_mul_577[22] + kernel_img_mul_577[23] + 
                kernel_img_mul_577[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4623:4616] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4623:4616] <= kernel_img_sum_577[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4623:4616] <= 'd0;
end

wire  [39:0]  kernel_img_mul_578[0:24];
assign kernel_img_mul_578[0] = buffer_data_4[4615:4608] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_578[1] = buffer_data_4[4623:4616] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_578[2] = buffer_data_4[4631:4624] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_578[3] = buffer_data_4[4639:4632] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_578[4] = buffer_data_4[4647:4640] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_578[5] = buffer_data_3[4615:4608] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_578[6] = buffer_data_3[4623:4616] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_578[7] = buffer_data_3[4631:4624] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_578[8] = buffer_data_3[4639:4632] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_578[9] = buffer_data_3[4647:4640] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_578[10] = buffer_data_2[4615:4608] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_578[11] = buffer_data_2[4623:4616] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_578[12] = buffer_data_2[4631:4624] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_578[13] = buffer_data_2[4639:4632] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_578[14] = buffer_data_2[4647:4640] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_578[15] = buffer_data_1[4615:4608] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_578[16] = buffer_data_1[4623:4616] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_578[17] = buffer_data_1[4631:4624] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_578[18] = buffer_data_1[4639:4632] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_578[19] = buffer_data_1[4647:4640] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_578[20] = buffer_data_0[4615:4608] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_578[21] = buffer_data_0[4623:4616] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_578[22] = buffer_data_0[4631:4624] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_578[23] = buffer_data_0[4639:4632] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_578[24] = buffer_data_0[4647:4640] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_578 = kernel_img_mul_578[0] + kernel_img_mul_578[1] + kernel_img_mul_578[2] + 
                kernel_img_mul_578[3] + kernel_img_mul_578[4] + kernel_img_mul_578[5] + 
                kernel_img_mul_578[6] + kernel_img_mul_578[7] + kernel_img_mul_578[8] + 
                kernel_img_mul_578[9] + kernel_img_mul_578[10] + kernel_img_mul_578[11] + 
                kernel_img_mul_578[12] + kernel_img_mul_578[13] + kernel_img_mul_578[14] + 
                kernel_img_mul_578[15] + kernel_img_mul_578[16] + kernel_img_mul_578[17] + 
                kernel_img_mul_578[18] + kernel_img_mul_578[19] + kernel_img_mul_578[20] + 
                kernel_img_mul_578[21] + kernel_img_mul_578[22] + kernel_img_mul_578[23] + 
                kernel_img_mul_578[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4631:4624] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4631:4624] <= kernel_img_sum_578[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4631:4624] <= 'd0;
end

wire  [39:0]  kernel_img_mul_579[0:24];
assign kernel_img_mul_579[0] = buffer_data_4[4623:4616] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_579[1] = buffer_data_4[4631:4624] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_579[2] = buffer_data_4[4639:4632] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_579[3] = buffer_data_4[4647:4640] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_579[4] = buffer_data_4[4655:4648] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_579[5] = buffer_data_3[4623:4616] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_579[6] = buffer_data_3[4631:4624] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_579[7] = buffer_data_3[4639:4632] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_579[8] = buffer_data_3[4647:4640] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_579[9] = buffer_data_3[4655:4648] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_579[10] = buffer_data_2[4623:4616] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_579[11] = buffer_data_2[4631:4624] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_579[12] = buffer_data_2[4639:4632] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_579[13] = buffer_data_2[4647:4640] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_579[14] = buffer_data_2[4655:4648] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_579[15] = buffer_data_1[4623:4616] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_579[16] = buffer_data_1[4631:4624] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_579[17] = buffer_data_1[4639:4632] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_579[18] = buffer_data_1[4647:4640] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_579[19] = buffer_data_1[4655:4648] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_579[20] = buffer_data_0[4623:4616] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_579[21] = buffer_data_0[4631:4624] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_579[22] = buffer_data_0[4639:4632] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_579[23] = buffer_data_0[4647:4640] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_579[24] = buffer_data_0[4655:4648] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_579 = kernel_img_mul_579[0] + kernel_img_mul_579[1] + kernel_img_mul_579[2] + 
                kernel_img_mul_579[3] + kernel_img_mul_579[4] + kernel_img_mul_579[5] + 
                kernel_img_mul_579[6] + kernel_img_mul_579[7] + kernel_img_mul_579[8] + 
                kernel_img_mul_579[9] + kernel_img_mul_579[10] + kernel_img_mul_579[11] + 
                kernel_img_mul_579[12] + kernel_img_mul_579[13] + kernel_img_mul_579[14] + 
                kernel_img_mul_579[15] + kernel_img_mul_579[16] + kernel_img_mul_579[17] + 
                kernel_img_mul_579[18] + kernel_img_mul_579[19] + kernel_img_mul_579[20] + 
                kernel_img_mul_579[21] + kernel_img_mul_579[22] + kernel_img_mul_579[23] + 
                kernel_img_mul_579[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4639:4632] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4639:4632] <= kernel_img_sum_579[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4639:4632] <= 'd0;
end

wire  [39:0]  kernel_img_mul_580[0:24];
assign kernel_img_mul_580[0] = buffer_data_4[4631:4624] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_580[1] = buffer_data_4[4639:4632] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_580[2] = buffer_data_4[4647:4640] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_580[3] = buffer_data_4[4655:4648] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_580[4] = buffer_data_4[4663:4656] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_580[5] = buffer_data_3[4631:4624] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_580[6] = buffer_data_3[4639:4632] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_580[7] = buffer_data_3[4647:4640] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_580[8] = buffer_data_3[4655:4648] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_580[9] = buffer_data_3[4663:4656] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_580[10] = buffer_data_2[4631:4624] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_580[11] = buffer_data_2[4639:4632] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_580[12] = buffer_data_2[4647:4640] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_580[13] = buffer_data_2[4655:4648] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_580[14] = buffer_data_2[4663:4656] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_580[15] = buffer_data_1[4631:4624] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_580[16] = buffer_data_1[4639:4632] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_580[17] = buffer_data_1[4647:4640] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_580[18] = buffer_data_1[4655:4648] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_580[19] = buffer_data_1[4663:4656] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_580[20] = buffer_data_0[4631:4624] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_580[21] = buffer_data_0[4639:4632] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_580[22] = buffer_data_0[4647:4640] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_580[23] = buffer_data_0[4655:4648] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_580[24] = buffer_data_0[4663:4656] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_580 = kernel_img_mul_580[0] + kernel_img_mul_580[1] + kernel_img_mul_580[2] + 
                kernel_img_mul_580[3] + kernel_img_mul_580[4] + kernel_img_mul_580[5] + 
                kernel_img_mul_580[6] + kernel_img_mul_580[7] + kernel_img_mul_580[8] + 
                kernel_img_mul_580[9] + kernel_img_mul_580[10] + kernel_img_mul_580[11] + 
                kernel_img_mul_580[12] + kernel_img_mul_580[13] + kernel_img_mul_580[14] + 
                kernel_img_mul_580[15] + kernel_img_mul_580[16] + kernel_img_mul_580[17] + 
                kernel_img_mul_580[18] + kernel_img_mul_580[19] + kernel_img_mul_580[20] + 
                kernel_img_mul_580[21] + kernel_img_mul_580[22] + kernel_img_mul_580[23] + 
                kernel_img_mul_580[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4647:4640] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4647:4640] <= kernel_img_sum_580[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4647:4640] <= 'd0;
end

wire  [39:0]  kernel_img_mul_581[0:24];
assign kernel_img_mul_581[0] = buffer_data_4[4639:4632] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_581[1] = buffer_data_4[4647:4640] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_581[2] = buffer_data_4[4655:4648] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_581[3] = buffer_data_4[4663:4656] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_581[4] = buffer_data_4[4671:4664] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_581[5] = buffer_data_3[4639:4632] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_581[6] = buffer_data_3[4647:4640] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_581[7] = buffer_data_3[4655:4648] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_581[8] = buffer_data_3[4663:4656] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_581[9] = buffer_data_3[4671:4664] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_581[10] = buffer_data_2[4639:4632] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_581[11] = buffer_data_2[4647:4640] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_581[12] = buffer_data_2[4655:4648] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_581[13] = buffer_data_2[4663:4656] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_581[14] = buffer_data_2[4671:4664] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_581[15] = buffer_data_1[4639:4632] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_581[16] = buffer_data_1[4647:4640] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_581[17] = buffer_data_1[4655:4648] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_581[18] = buffer_data_1[4663:4656] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_581[19] = buffer_data_1[4671:4664] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_581[20] = buffer_data_0[4639:4632] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_581[21] = buffer_data_0[4647:4640] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_581[22] = buffer_data_0[4655:4648] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_581[23] = buffer_data_0[4663:4656] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_581[24] = buffer_data_0[4671:4664] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_581 = kernel_img_mul_581[0] + kernel_img_mul_581[1] + kernel_img_mul_581[2] + 
                kernel_img_mul_581[3] + kernel_img_mul_581[4] + kernel_img_mul_581[5] + 
                kernel_img_mul_581[6] + kernel_img_mul_581[7] + kernel_img_mul_581[8] + 
                kernel_img_mul_581[9] + kernel_img_mul_581[10] + kernel_img_mul_581[11] + 
                kernel_img_mul_581[12] + kernel_img_mul_581[13] + kernel_img_mul_581[14] + 
                kernel_img_mul_581[15] + kernel_img_mul_581[16] + kernel_img_mul_581[17] + 
                kernel_img_mul_581[18] + kernel_img_mul_581[19] + kernel_img_mul_581[20] + 
                kernel_img_mul_581[21] + kernel_img_mul_581[22] + kernel_img_mul_581[23] + 
                kernel_img_mul_581[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4655:4648] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4655:4648] <= kernel_img_sum_581[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4655:4648] <= 'd0;
end

wire  [39:0]  kernel_img_mul_582[0:24];
assign kernel_img_mul_582[0] = buffer_data_4[4647:4640] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_582[1] = buffer_data_4[4655:4648] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_582[2] = buffer_data_4[4663:4656] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_582[3] = buffer_data_4[4671:4664] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_582[4] = buffer_data_4[4679:4672] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_582[5] = buffer_data_3[4647:4640] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_582[6] = buffer_data_3[4655:4648] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_582[7] = buffer_data_3[4663:4656] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_582[8] = buffer_data_3[4671:4664] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_582[9] = buffer_data_3[4679:4672] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_582[10] = buffer_data_2[4647:4640] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_582[11] = buffer_data_2[4655:4648] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_582[12] = buffer_data_2[4663:4656] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_582[13] = buffer_data_2[4671:4664] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_582[14] = buffer_data_2[4679:4672] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_582[15] = buffer_data_1[4647:4640] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_582[16] = buffer_data_1[4655:4648] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_582[17] = buffer_data_1[4663:4656] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_582[18] = buffer_data_1[4671:4664] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_582[19] = buffer_data_1[4679:4672] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_582[20] = buffer_data_0[4647:4640] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_582[21] = buffer_data_0[4655:4648] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_582[22] = buffer_data_0[4663:4656] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_582[23] = buffer_data_0[4671:4664] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_582[24] = buffer_data_0[4679:4672] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_582 = kernel_img_mul_582[0] + kernel_img_mul_582[1] + kernel_img_mul_582[2] + 
                kernel_img_mul_582[3] + kernel_img_mul_582[4] + kernel_img_mul_582[5] + 
                kernel_img_mul_582[6] + kernel_img_mul_582[7] + kernel_img_mul_582[8] + 
                kernel_img_mul_582[9] + kernel_img_mul_582[10] + kernel_img_mul_582[11] + 
                kernel_img_mul_582[12] + kernel_img_mul_582[13] + kernel_img_mul_582[14] + 
                kernel_img_mul_582[15] + kernel_img_mul_582[16] + kernel_img_mul_582[17] + 
                kernel_img_mul_582[18] + kernel_img_mul_582[19] + kernel_img_mul_582[20] + 
                kernel_img_mul_582[21] + kernel_img_mul_582[22] + kernel_img_mul_582[23] + 
                kernel_img_mul_582[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4663:4656] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4663:4656] <= kernel_img_sum_582[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4663:4656] <= 'd0;
end

wire  [39:0]  kernel_img_mul_583[0:24];
assign kernel_img_mul_583[0] = buffer_data_4[4655:4648] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_583[1] = buffer_data_4[4663:4656] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_583[2] = buffer_data_4[4671:4664] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_583[3] = buffer_data_4[4679:4672] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_583[4] = buffer_data_4[4687:4680] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_583[5] = buffer_data_3[4655:4648] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_583[6] = buffer_data_3[4663:4656] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_583[7] = buffer_data_3[4671:4664] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_583[8] = buffer_data_3[4679:4672] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_583[9] = buffer_data_3[4687:4680] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_583[10] = buffer_data_2[4655:4648] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_583[11] = buffer_data_2[4663:4656] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_583[12] = buffer_data_2[4671:4664] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_583[13] = buffer_data_2[4679:4672] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_583[14] = buffer_data_2[4687:4680] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_583[15] = buffer_data_1[4655:4648] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_583[16] = buffer_data_1[4663:4656] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_583[17] = buffer_data_1[4671:4664] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_583[18] = buffer_data_1[4679:4672] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_583[19] = buffer_data_1[4687:4680] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_583[20] = buffer_data_0[4655:4648] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_583[21] = buffer_data_0[4663:4656] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_583[22] = buffer_data_0[4671:4664] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_583[23] = buffer_data_0[4679:4672] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_583[24] = buffer_data_0[4687:4680] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_583 = kernel_img_mul_583[0] + kernel_img_mul_583[1] + kernel_img_mul_583[2] + 
                kernel_img_mul_583[3] + kernel_img_mul_583[4] + kernel_img_mul_583[5] + 
                kernel_img_mul_583[6] + kernel_img_mul_583[7] + kernel_img_mul_583[8] + 
                kernel_img_mul_583[9] + kernel_img_mul_583[10] + kernel_img_mul_583[11] + 
                kernel_img_mul_583[12] + kernel_img_mul_583[13] + kernel_img_mul_583[14] + 
                kernel_img_mul_583[15] + kernel_img_mul_583[16] + kernel_img_mul_583[17] + 
                kernel_img_mul_583[18] + kernel_img_mul_583[19] + kernel_img_mul_583[20] + 
                kernel_img_mul_583[21] + kernel_img_mul_583[22] + kernel_img_mul_583[23] + 
                kernel_img_mul_583[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4671:4664] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4671:4664] <= kernel_img_sum_583[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4671:4664] <= 'd0;
end

wire  [39:0]  kernel_img_mul_584[0:24];
assign kernel_img_mul_584[0] = buffer_data_4[4663:4656] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_584[1] = buffer_data_4[4671:4664] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_584[2] = buffer_data_4[4679:4672] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_584[3] = buffer_data_4[4687:4680] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_584[4] = buffer_data_4[4695:4688] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_584[5] = buffer_data_3[4663:4656] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_584[6] = buffer_data_3[4671:4664] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_584[7] = buffer_data_3[4679:4672] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_584[8] = buffer_data_3[4687:4680] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_584[9] = buffer_data_3[4695:4688] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_584[10] = buffer_data_2[4663:4656] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_584[11] = buffer_data_2[4671:4664] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_584[12] = buffer_data_2[4679:4672] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_584[13] = buffer_data_2[4687:4680] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_584[14] = buffer_data_2[4695:4688] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_584[15] = buffer_data_1[4663:4656] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_584[16] = buffer_data_1[4671:4664] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_584[17] = buffer_data_1[4679:4672] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_584[18] = buffer_data_1[4687:4680] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_584[19] = buffer_data_1[4695:4688] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_584[20] = buffer_data_0[4663:4656] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_584[21] = buffer_data_0[4671:4664] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_584[22] = buffer_data_0[4679:4672] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_584[23] = buffer_data_0[4687:4680] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_584[24] = buffer_data_0[4695:4688] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_584 = kernel_img_mul_584[0] + kernel_img_mul_584[1] + kernel_img_mul_584[2] + 
                kernel_img_mul_584[3] + kernel_img_mul_584[4] + kernel_img_mul_584[5] + 
                kernel_img_mul_584[6] + kernel_img_mul_584[7] + kernel_img_mul_584[8] + 
                kernel_img_mul_584[9] + kernel_img_mul_584[10] + kernel_img_mul_584[11] + 
                kernel_img_mul_584[12] + kernel_img_mul_584[13] + kernel_img_mul_584[14] + 
                kernel_img_mul_584[15] + kernel_img_mul_584[16] + kernel_img_mul_584[17] + 
                kernel_img_mul_584[18] + kernel_img_mul_584[19] + kernel_img_mul_584[20] + 
                kernel_img_mul_584[21] + kernel_img_mul_584[22] + kernel_img_mul_584[23] + 
                kernel_img_mul_584[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4679:4672] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4679:4672] <= kernel_img_sum_584[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4679:4672] <= 'd0;
end

wire  [39:0]  kernel_img_mul_585[0:24];
assign kernel_img_mul_585[0] = buffer_data_4[4671:4664] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_585[1] = buffer_data_4[4679:4672] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_585[2] = buffer_data_4[4687:4680] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_585[3] = buffer_data_4[4695:4688] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_585[4] = buffer_data_4[4703:4696] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_585[5] = buffer_data_3[4671:4664] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_585[6] = buffer_data_3[4679:4672] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_585[7] = buffer_data_3[4687:4680] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_585[8] = buffer_data_3[4695:4688] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_585[9] = buffer_data_3[4703:4696] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_585[10] = buffer_data_2[4671:4664] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_585[11] = buffer_data_2[4679:4672] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_585[12] = buffer_data_2[4687:4680] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_585[13] = buffer_data_2[4695:4688] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_585[14] = buffer_data_2[4703:4696] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_585[15] = buffer_data_1[4671:4664] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_585[16] = buffer_data_1[4679:4672] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_585[17] = buffer_data_1[4687:4680] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_585[18] = buffer_data_1[4695:4688] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_585[19] = buffer_data_1[4703:4696] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_585[20] = buffer_data_0[4671:4664] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_585[21] = buffer_data_0[4679:4672] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_585[22] = buffer_data_0[4687:4680] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_585[23] = buffer_data_0[4695:4688] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_585[24] = buffer_data_0[4703:4696] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_585 = kernel_img_mul_585[0] + kernel_img_mul_585[1] + kernel_img_mul_585[2] + 
                kernel_img_mul_585[3] + kernel_img_mul_585[4] + kernel_img_mul_585[5] + 
                kernel_img_mul_585[6] + kernel_img_mul_585[7] + kernel_img_mul_585[8] + 
                kernel_img_mul_585[9] + kernel_img_mul_585[10] + kernel_img_mul_585[11] + 
                kernel_img_mul_585[12] + kernel_img_mul_585[13] + kernel_img_mul_585[14] + 
                kernel_img_mul_585[15] + kernel_img_mul_585[16] + kernel_img_mul_585[17] + 
                kernel_img_mul_585[18] + kernel_img_mul_585[19] + kernel_img_mul_585[20] + 
                kernel_img_mul_585[21] + kernel_img_mul_585[22] + kernel_img_mul_585[23] + 
                kernel_img_mul_585[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4687:4680] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4687:4680] <= kernel_img_sum_585[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4687:4680] <= 'd0;
end

wire  [39:0]  kernel_img_mul_586[0:24];
assign kernel_img_mul_586[0] = buffer_data_4[4679:4672] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_586[1] = buffer_data_4[4687:4680] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_586[2] = buffer_data_4[4695:4688] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_586[3] = buffer_data_4[4703:4696] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_586[4] = buffer_data_4[4711:4704] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_586[5] = buffer_data_3[4679:4672] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_586[6] = buffer_data_3[4687:4680] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_586[7] = buffer_data_3[4695:4688] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_586[8] = buffer_data_3[4703:4696] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_586[9] = buffer_data_3[4711:4704] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_586[10] = buffer_data_2[4679:4672] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_586[11] = buffer_data_2[4687:4680] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_586[12] = buffer_data_2[4695:4688] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_586[13] = buffer_data_2[4703:4696] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_586[14] = buffer_data_2[4711:4704] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_586[15] = buffer_data_1[4679:4672] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_586[16] = buffer_data_1[4687:4680] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_586[17] = buffer_data_1[4695:4688] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_586[18] = buffer_data_1[4703:4696] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_586[19] = buffer_data_1[4711:4704] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_586[20] = buffer_data_0[4679:4672] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_586[21] = buffer_data_0[4687:4680] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_586[22] = buffer_data_0[4695:4688] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_586[23] = buffer_data_0[4703:4696] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_586[24] = buffer_data_0[4711:4704] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_586 = kernel_img_mul_586[0] + kernel_img_mul_586[1] + kernel_img_mul_586[2] + 
                kernel_img_mul_586[3] + kernel_img_mul_586[4] + kernel_img_mul_586[5] + 
                kernel_img_mul_586[6] + kernel_img_mul_586[7] + kernel_img_mul_586[8] + 
                kernel_img_mul_586[9] + kernel_img_mul_586[10] + kernel_img_mul_586[11] + 
                kernel_img_mul_586[12] + kernel_img_mul_586[13] + kernel_img_mul_586[14] + 
                kernel_img_mul_586[15] + kernel_img_mul_586[16] + kernel_img_mul_586[17] + 
                kernel_img_mul_586[18] + kernel_img_mul_586[19] + kernel_img_mul_586[20] + 
                kernel_img_mul_586[21] + kernel_img_mul_586[22] + kernel_img_mul_586[23] + 
                kernel_img_mul_586[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4695:4688] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4695:4688] <= kernel_img_sum_586[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4695:4688] <= 'd0;
end

wire  [39:0]  kernel_img_mul_587[0:24];
assign kernel_img_mul_587[0] = buffer_data_4[4687:4680] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_587[1] = buffer_data_4[4695:4688] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_587[2] = buffer_data_4[4703:4696] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_587[3] = buffer_data_4[4711:4704] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_587[4] = buffer_data_4[4719:4712] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_587[5] = buffer_data_3[4687:4680] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_587[6] = buffer_data_3[4695:4688] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_587[7] = buffer_data_3[4703:4696] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_587[8] = buffer_data_3[4711:4704] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_587[9] = buffer_data_3[4719:4712] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_587[10] = buffer_data_2[4687:4680] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_587[11] = buffer_data_2[4695:4688] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_587[12] = buffer_data_2[4703:4696] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_587[13] = buffer_data_2[4711:4704] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_587[14] = buffer_data_2[4719:4712] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_587[15] = buffer_data_1[4687:4680] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_587[16] = buffer_data_1[4695:4688] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_587[17] = buffer_data_1[4703:4696] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_587[18] = buffer_data_1[4711:4704] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_587[19] = buffer_data_1[4719:4712] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_587[20] = buffer_data_0[4687:4680] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_587[21] = buffer_data_0[4695:4688] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_587[22] = buffer_data_0[4703:4696] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_587[23] = buffer_data_0[4711:4704] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_587[24] = buffer_data_0[4719:4712] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_587 = kernel_img_mul_587[0] + kernel_img_mul_587[1] + kernel_img_mul_587[2] + 
                kernel_img_mul_587[3] + kernel_img_mul_587[4] + kernel_img_mul_587[5] + 
                kernel_img_mul_587[6] + kernel_img_mul_587[7] + kernel_img_mul_587[8] + 
                kernel_img_mul_587[9] + kernel_img_mul_587[10] + kernel_img_mul_587[11] + 
                kernel_img_mul_587[12] + kernel_img_mul_587[13] + kernel_img_mul_587[14] + 
                kernel_img_mul_587[15] + kernel_img_mul_587[16] + kernel_img_mul_587[17] + 
                kernel_img_mul_587[18] + kernel_img_mul_587[19] + kernel_img_mul_587[20] + 
                kernel_img_mul_587[21] + kernel_img_mul_587[22] + kernel_img_mul_587[23] + 
                kernel_img_mul_587[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4703:4696] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4703:4696] <= kernel_img_sum_587[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4703:4696] <= 'd0;
end

wire  [39:0]  kernel_img_mul_588[0:24];
assign kernel_img_mul_588[0] = buffer_data_4[4695:4688] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_588[1] = buffer_data_4[4703:4696] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_588[2] = buffer_data_4[4711:4704] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_588[3] = buffer_data_4[4719:4712] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_588[4] = buffer_data_4[4727:4720] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_588[5] = buffer_data_3[4695:4688] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_588[6] = buffer_data_3[4703:4696] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_588[7] = buffer_data_3[4711:4704] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_588[8] = buffer_data_3[4719:4712] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_588[9] = buffer_data_3[4727:4720] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_588[10] = buffer_data_2[4695:4688] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_588[11] = buffer_data_2[4703:4696] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_588[12] = buffer_data_2[4711:4704] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_588[13] = buffer_data_2[4719:4712] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_588[14] = buffer_data_2[4727:4720] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_588[15] = buffer_data_1[4695:4688] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_588[16] = buffer_data_1[4703:4696] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_588[17] = buffer_data_1[4711:4704] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_588[18] = buffer_data_1[4719:4712] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_588[19] = buffer_data_1[4727:4720] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_588[20] = buffer_data_0[4695:4688] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_588[21] = buffer_data_0[4703:4696] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_588[22] = buffer_data_0[4711:4704] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_588[23] = buffer_data_0[4719:4712] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_588[24] = buffer_data_0[4727:4720] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_588 = kernel_img_mul_588[0] + kernel_img_mul_588[1] + kernel_img_mul_588[2] + 
                kernel_img_mul_588[3] + kernel_img_mul_588[4] + kernel_img_mul_588[5] + 
                kernel_img_mul_588[6] + kernel_img_mul_588[7] + kernel_img_mul_588[8] + 
                kernel_img_mul_588[9] + kernel_img_mul_588[10] + kernel_img_mul_588[11] + 
                kernel_img_mul_588[12] + kernel_img_mul_588[13] + kernel_img_mul_588[14] + 
                kernel_img_mul_588[15] + kernel_img_mul_588[16] + kernel_img_mul_588[17] + 
                kernel_img_mul_588[18] + kernel_img_mul_588[19] + kernel_img_mul_588[20] + 
                kernel_img_mul_588[21] + kernel_img_mul_588[22] + kernel_img_mul_588[23] + 
                kernel_img_mul_588[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4711:4704] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4711:4704] <= kernel_img_sum_588[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4711:4704] <= 'd0;
end

wire  [39:0]  kernel_img_mul_589[0:24];
assign kernel_img_mul_589[0] = buffer_data_4[4703:4696] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_589[1] = buffer_data_4[4711:4704] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_589[2] = buffer_data_4[4719:4712] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_589[3] = buffer_data_4[4727:4720] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_589[4] = buffer_data_4[4735:4728] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_589[5] = buffer_data_3[4703:4696] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_589[6] = buffer_data_3[4711:4704] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_589[7] = buffer_data_3[4719:4712] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_589[8] = buffer_data_3[4727:4720] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_589[9] = buffer_data_3[4735:4728] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_589[10] = buffer_data_2[4703:4696] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_589[11] = buffer_data_2[4711:4704] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_589[12] = buffer_data_2[4719:4712] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_589[13] = buffer_data_2[4727:4720] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_589[14] = buffer_data_2[4735:4728] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_589[15] = buffer_data_1[4703:4696] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_589[16] = buffer_data_1[4711:4704] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_589[17] = buffer_data_1[4719:4712] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_589[18] = buffer_data_1[4727:4720] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_589[19] = buffer_data_1[4735:4728] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_589[20] = buffer_data_0[4703:4696] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_589[21] = buffer_data_0[4711:4704] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_589[22] = buffer_data_0[4719:4712] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_589[23] = buffer_data_0[4727:4720] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_589[24] = buffer_data_0[4735:4728] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_589 = kernel_img_mul_589[0] + kernel_img_mul_589[1] + kernel_img_mul_589[2] + 
                kernel_img_mul_589[3] + kernel_img_mul_589[4] + kernel_img_mul_589[5] + 
                kernel_img_mul_589[6] + kernel_img_mul_589[7] + kernel_img_mul_589[8] + 
                kernel_img_mul_589[9] + kernel_img_mul_589[10] + kernel_img_mul_589[11] + 
                kernel_img_mul_589[12] + kernel_img_mul_589[13] + kernel_img_mul_589[14] + 
                kernel_img_mul_589[15] + kernel_img_mul_589[16] + kernel_img_mul_589[17] + 
                kernel_img_mul_589[18] + kernel_img_mul_589[19] + kernel_img_mul_589[20] + 
                kernel_img_mul_589[21] + kernel_img_mul_589[22] + kernel_img_mul_589[23] + 
                kernel_img_mul_589[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4719:4712] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4719:4712] <= kernel_img_sum_589[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4719:4712] <= 'd0;
end

wire  [39:0]  kernel_img_mul_590[0:24];
assign kernel_img_mul_590[0] = buffer_data_4[4711:4704] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_590[1] = buffer_data_4[4719:4712] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_590[2] = buffer_data_4[4727:4720] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_590[3] = buffer_data_4[4735:4728] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_590[4] = buffer_data_4[4743:4736] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_590[5] = buffer_data_3[4711:4704] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_590[6] = buffer_data_3[4719:4712] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_590[7] = buffer_data_3[4727:4720] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_590[8] = buffer_data_3[4735:4728] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_590[9] = buffer_data_3[4743:4736] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_590[10] = buffer_data_2[4711:4704] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_590[11] = buffer_data_2[4719:4712] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_590[12] = buffer_data_2[4727:4720] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_590[13] = buffer_data_2[4735:4728] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_590[14] = buffer_data_2[4743:4736] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_590[15] = buffer_data_1[4711:4704] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_590[16] = buffer_data_1[4719:4712] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_590[17] = buffer_data_1[4727:4720] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_590[18] = buffer_data_1[4735:4728] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_590[19] = buffer_data_1[4743:4736] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_590[20] = buffer_data_0[4711:4704] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_590[21] = buffer_data_0[4719:4712] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_590[22] = buffer_data_0[4727:4720] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_590[23] = buffer_data_0[4735:4728] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_590[24] = buffer_data_0[4743:4736] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_590 = kernel_img_mul_590[0] + kernel_img_mul_590[1] + kernel_img_mul_590[2] + 
                kernel_img_mul_590[3] + kernel_img_mul_590[4] + kernel_img_mul_590[5] + 
                kernel_img_mul_590[6] + kernel_img_mul_590[7] + kernel_img_mul_590[8] + 
                kernel_img_mul_590[9] + kernel_img_mul_590[10] + kernel_img_mul_590[11] + 
                kernel_img_mul_590[12] + kernel_img_mul_590[13] + kernel_img_mul_590[14] + 
                kernel_img_mul_590[15] + kernel_img_mul_590[16] + kernel_img_mul_590[17] + 
                kernel_img_mul_590[18] + kernel_img_mul_590[19] + kernel_img_mul_590[20] + 
                kernel_img_mul_590[21] + kernel_img_mul_590[22] + kernel_img_mul_590[23] + 
                kernel_img_mul_590[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4727:4720] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4727:4720] <= kernel_img_sum_590[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4727:4720] <= 'd0;
end

wire  [39:0]  kernel_img_mul_591[0:24];
assign kernel_img_mul_591[0] = buffer_data_4[4719:4712] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_591[1] = buffer_data_4[4727:4720] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_591[2] = buffer_data_4[4735:4728] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_591[3] = buffer_data_4[4743:4736] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_591[4] = buffer_data_4[4751:4744] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_591[5] = buffer_data_3[4719:4712] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_591[6] = buffer_data_3[4727:4720] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_591[7] = buffer_data_3[4735:4728] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_591[8] = buffer_data_3[4743:4736] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_591[9] = buffer_data_3[4751:4744] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_591[10] = buffer_data_2[4719:4712] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_591[11] = buffer_data_2[4727:4720] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_591[12] = buffer_data_2[4735:4728] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_591[13] = buffer_data_2[4743:4736] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_591[14] = buffer_data_2[4751:4744] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_591[15] = buffer_data_1[4719:4712] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_591[16] = buffer_data_1[4727:4720] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_591[17] = buffer_data_1[4735:4728] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_591[18] = buffer_data_1[4743:4736] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_591[19] = buffer_data_1[4751:4744] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_591[20] = buffer_data_0[4719:4712] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_591[21] = buffer_data_0[4727:4720] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_591[22] = buffer_data_0[4735:4728] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_591[23] = buffer_data_0[4743:4736] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_591[24] = buffer_data_0[4751:4744] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_591 = kernel_img_mul_591[0] + kernel_img_mul_591[1] + kernel_img_mul_591[2] + 
                kernel_img_mul_591[3] + kernel_img_mul_591[4] + kernel_img_mul_591[5] + 
                kernel_img_mul_591[6] + kernel_img_mul_591[7] + kernel_img_mul_591[8] + 
                kernel_img_mul_591[9] + kernel_img_mul_591[10] + kernel_img_mul_591[11] + 
                kernel_img_mul_591[12] + kernel_img_mul_591[13] + kernel_img_mul_591[14] + 
                kernel_img_mul_591[15] + kernel_img_mul_591[16] + kernel_img_mul_591[17] + 
                kernel_img_mul_591[18] + kernel_img_mul_591[19] + kernel_img_mul_591[20] + 
                kernel_img_mul_591[21] + kernel_img_mul_591[22] + kernel_img_mul_591[23] + 
                kernel_img_mul_591[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4735:4728] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4735:4728] <= kernel_img_sum_591[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4735:4728] <= 'd0;
end

wire  [39:0]  kernel_img_mul_592[0:24];
assign kernel_img_mul_592[0] = buffer_data_4[4727:4720] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_592[1] = buffer_data_4[4735:4728] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_592[2] = buffer_data_4[4743:4736] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_592[3] = buffer_data_4[4751:4744] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_592[4] = buffer_data_4[4759:4752] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_592[5] = buffer_data_3[4727:4720] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_592[6] = buffer_data_3[4735:4728] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_592[7] = buffer_data_3[4743:4736] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_592[8] = buffer_data_3[4751:4744] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_592[9] = buffer_data_3[4759:4752] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_592[10] = buffer_data_2[4727:4720] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_592[11] = buffer_data_2[4735:4728] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_592[12] = buffer_data_2[4743:4736] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_592[13] = buffer_data_2[4751:4744] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_592[14] = buffer_data_2[4759:4752] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_592[15] = buffer_data_1[4727:4720] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_592[16] = buffer_data_1[4735:4728] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_592[17] = buffer_data_1[4743:4736] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_592[18] = buffer_data_1[4751:4744] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_592[19] = buffer_data_1[4759:4752] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_592[20] = buffer_data_0[4727:4720] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_592[21] = buffer_data_0[4735:4728] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_592[22] = buffer_data_0[4743:4736] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_592[23] = buffer_data_0[4751:4744] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_592[24] = buffer_data_0[4759:4752] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_592 = kernel_img_mul_592[0] + kernel_img_mul_592[1] + kernel_img_mul_592[2] + 
                kernel_img_mul_592[3] + kernel_img_mul_592[4] + kernel_img_mul_592[5] + 
                kernel_img_mul_592[6] + kernel_img_mul_592[7] + kernel_img_mul_592[8] + 
                kernel_img_mul_592[9] + kernel_img_mul_592[10] + kernel_img_mul_592[11] + 
                kernel_img_mul_592[12] + kernel_img_mul_592[13] + kernel_img_mul_592[14] + 
                kernel_img_mul_592[15] + kernel_img_mul_592[16] + kernel_img_mul_592[17] + 
                kernel_img_mul_592[18] + kernel_img_mul_592[19] + kernel_img_mul_592[20] + 
                kernel_img_mul_592[21] + kernel_img_mul_592[22] + kernel_img_mul_592[23] + 
                kernel_img_mul_592[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4743:4736] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4743:4736] <= kernel_img_sum_592[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4743:4736] <= 'd0;
end

wire  [39:0]  kernel_img_mul_593[0:24];
assign kernel_img_mul_593[0] = buffer_data_4[4735:4728] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_593[1] = buffer_data_4[4743:4736] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_593[2] = buffer_data_4[4751:4744] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_593[3] = buffer_data_4[4759:4752] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_593[4] = buffer_data_4[4767:4760] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_593[5] = buffer_data_3[4735:4728] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_593[6] = buffer_data_3[4743:4736] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_593[7] = buffer_data_3[4751:4744] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_593[8] = buffer_data_3[4759:4752] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_593[9] = buffer_data_3[4767:4760] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_593[10] = buffer_data_2[4735:4728] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_593[11] = buffer_data_2[4743:4736] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_593[12] = buffer_data_2[4751:4744] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_593[13] = buffer_data_2[4759:4752] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_593[14] = buffer_data_2[4767:4760] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_593[15] = buffer_data_1[4735:4728] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_593[16] = buffer_data_1[4743:4736] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_593[17] = buffer_data_1[4751:4744] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_593[18] = buffer_data_1[4759:4752] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_593[19] = buffer_data_1[4767:4760] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_593[20] = buffer_data_0[4735:4728] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_593[21] = buffer_data_0[4743:4736] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_593[22] = buffer_data_0[4751:4744] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_593[23] = buffer_data_0[4759:4752] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_593[24] = buffer_data_0[4767:4760] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_593 = kernel_img_mul_593[0] + kernel_img_mul_593[1] + kernel_img_mul_593[2] + 
                kernel_img_mul_593[3] + kernel_img_mul_593[4] + kernel_img_mul_593[5] + 
                kernel_img_mul_593[6] + kernel_img_mul_593[7] + kernel_img_mul_593[8] + 
                kernel_img_mul_593[9] + kernel_img_mul_593[10] + kernel_img_mul_593[11] + 
                kernel_img_mul_593[12] + kernel_img_mul_593[13] + kernel_img_mul_593[14] + 
                kernel_img_mul_593[15] + kernel_img_mul_593[16] + kernel_img_mul_593[17] + 
                kernel_img_mul_593[18] + kernel_img_mul_593[19] + kernel_img_mul_593[20] + 
                kernel_img_mul_593[21] + kernel_img_mul_593[22] + kernel_img_mul_593[23] + 
                kernel_img_mul_593[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4751:4744] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4751:4744] <= kernel_img_sum_593[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4751:4744] <= 'd0;
end

wire  [39:0]  kernel_img_mul_594[0:24];
assign kernel_img_mul_594[0] = buffer_data_4[4743:4736] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_594[1] = buffer_data_4[4751:4744] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_594[2] = buffer_data_4[4759:4752] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_594[3] = buffer_data_4[4767:4760] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_594[4] = buffer_data_4[4775:4768] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_594[5] = buffer_data_3[4743:4736] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_594[6] = buffer_data_3[4751:4744] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_594[7] = buffer_data_3[4759:4752] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_594[8] = buffer_data_3[4767:4760] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_594[9] = buffer_data_3[4775:4768] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_594[10] = buffer_data_2[4743:4736] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_594[11] = buffer_data_2[4751:4744] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_594[12] = buffer_data_2[4759:4752] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_594[13] = buffer_data_2[4767:4760] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_594[14] = buffer_data_2[4775:4768] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_594[15] = buffer_data_1[4743:4736] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_594[16] = buffer_data_1[4751:4744] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_594[17] = buffer_data_1[4759:4752] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_594[18] = buffer_data_1[4767:4760] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_594[19] = buffer_data_1[4775:4768] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_594[20] = buffer_data_0[4743:4736] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_594[21] = buffer_data_0[4751:4744] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_594[22] = buffer_data_0[4759:4752] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_594[23] = buffer_data_0[4767:4760] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_594[24] = buffer_data_0[4775:4768] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_594 = kernel_img_mul_594[0] + kernel_img_mul_594[1] + kernel_img_mul_594[2] + 
                kernel_img_mul_594[3] + kernel_img_mul_594[4] + kernel_img_mul_594[5] + 
                kernel_img_mul_594[6] + kernel_img_mul_594[7] + kernel_img_mul_594[8] + 
                kernel_img_mul_594[9] + kernel_img_mul_594[10] + kernel_img_mul_594[11] + 
                kernel_img_mul_594[12] + kernel_img_mul_594[13] + kernel_img_mul_594[14] + 
                kernel_img_mul_594[15] + kernel_img_mul_594[16] + kernel_img_mul_594[17] + 
                kernel_img_mul_594[18] + kernel_img_mul_594[19] + kernel_img_mul_594[20] + 
                kernel_img_mul_594[21] + kernel_img_mul_594[22] + kernel_img_mul_594[23] + 
                kernel_img_mul_594[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4759:4752] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4759:4752] <= kernel_img_sum_594[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4759:4752] <= 'd0;
end

wire  [39:0]  kernel_img_mul_595[0:24];
assign kernel_img_mul_595[0] = buffer_data_4[4751:4744] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_595[1] = buffer_data_4[4759:4752] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_595[2] = buffer_data_4[4767:4760] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_595[3] = buffer_data_4[4775:4768] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_595[4] = buffer_data_4[4783:4776] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_595[5] = buffer_data_3[4751:4744] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_595[6] = buffer_data_3[4759:4752] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_595[7] = buffer_data_3[4767:4760] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_595[8] = buffer_data_3[4775:4768] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_595[9] = buffer_data_3[4783:4776] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_595[10] = buffer_data_2[4751:4744] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_595[11] = buffer_data_2[4759:4752] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_595[12] = buffer_data_2[4767:4760] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_595[13] = buffer_data_2[4775:4768] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_595[14] = buffer_data_2[4783:4776] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_595[15] = buffer_data_1[4751:4744] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_595[16] = buffer_data_1[4759:4752] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_595[17] = buffer_data_1[4767:4760] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_595[18] = buffer_data_1[4775:4768] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_595[19] = buffer_data_1[4783:4776] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_595[20] = buffer_data_0[4751:4744] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_595[21] = buffer_data_0[4759:4752] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_595[22] = buffer_data_0[4767:4760] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_595[23] = buffer_data_0[4775:4768] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_595[24] = buffer_data_0[4783:4776] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_595 = kernel_img_mul_595[0] + kernel_img_mul_595[1] + kernel_img_mul_595[2] + 
                kernel_img_mul_595[3] + kernel_img_mul_595[4] + kernel_img_mul_595[5] + 
                kernel_img_mul_595[6] + kernel_img_mul_595[7] + kernel_img_mul_595[8] + 
                kernel_img_mul_595[9] + kernel_img_mul_595[10] + kernel_img_mul_595[11] + 
                kernel_img_mul_595[12] + kernel_img_mul_595[13] + kernel_img_mul_595[14] + 
                kernel_img_mul_595[15] + kernel_img_mul_595[16] + kernel_img_mul_595[17] + 
                kernel_img_mul_595[18] + kernel_img_mul_595[19] + kernel_img_mul_595[20] + 
                kernel_img_mul_595[21] + kernel_img_mul_595[22] + kernel_img_mul_595[23] + 
                kernel_img_mul_595[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4767:4760] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4767:4760] <= kernel_img_sum_595[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4767:4760] <= 'd0;
end

wire  [39:0]  kernel_img_mul_596[0:24];
assign kernel_img_mul_596[0] = buffer_data_4[4759:4752] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_596[1] = buffer_data_4[4767:4760] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_596[2] = buffer_data_4[4775:4768] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_596[3] = buffer_data_4[4783:4776] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_596[4] = buffer_data_4[4791:4784] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_596[5] = buffer_data_3[4759:4752] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_596[6] = buffer_data_3[4767:4760] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_596[7] = buffer_data_3[4775:4768] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_596[8] = buffer_data_3[4783:4776] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_596[9] = buffer_data_3[4791:4784] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_596[10] = buffer_data_2[4759:4752] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_596[11] = buffer_data_2[4767:4760] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_596[12] = buffer_data_2[4775:4768] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_596[13] = buffer_data_2[4783:4776] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_596[14] = buffer_data_2[4791:4784] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_596[15] = buffer_data_1[4759:4752] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_596[16] = buffer_data_1[4767:4760] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_596[17] = buffer_data_1[4775:4768] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_596[18] = buffer_data_1[4783:4776] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_596[19] = buffer_data_1[4791:4784] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_596[20] = buffer_data_0[4759:4752] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_596[21] = buffer_data_0[4767:4760] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_596[22] = buffer_data_0[4775:4768] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_596[23] = buffer_data_0[4783:4776] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_596[24] = buffer_data_0[4791:4784] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_596 = kernel_img_mul_596[0] + kernel_img_mul_596[1] + kernel_img_mul_596[2] + 
                kernel_img_mul_596[3] + kernel_img_mul_596[4] + kernel_img_mul_596[5] + 
                kernel_img_mul_596[6] + kernel_img_mul_596[7] + kernel_img_mul_596[8] + 
                kernel_img_mul_596[9] + kernel_img_mul_596[10] + kernel_img_mul_596[11] + 
                kernel_img_mul_596[12] + kernel_img_mul_596[13] + kernel_img_mul_596[14] + 
                kernel_img_mul_596[15] + kernel_img_mul_596[16] + kernel_img_mul_596[17] + 
                kernel_img_mul_596[18] + kernel_img_mul_596[19] + kernel_img_mul_596[20] + 
                kernel_img_mul_596[21] + kernel_img_mul_596[22] + kernel_img_mul_596[23] + 
                kernel_img_mul_596[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4775:4768] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4775:4768] <= kernel_img_sum_596[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4775:4768] <= 'd0;
end

wire  [39:0]  kernel_img_mul_597[0:24];
assign kernel_img_mul_597[0] = buffer_data_4[4767:4760] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_597[1] = buffer_data_4[4775:4768] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_597[2] = buffer_data_4[4783:4776] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_597[3] = buffer_data_4[4791:4784] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_597[4] = buffer_data_4[4799:4792] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_597[5] = buffer_data_3[4767:4760] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_597[6] = buffer_data_3[4775:4768] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_597[7] = buffer_data_3[4783:4776] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_597[8] = buffer_data_3[4791:4784] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_597[9] = buffer_data_3[4799:4792] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_597[10] = buffer_data_2[4767:4760] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_597[11] = buffer_data_2[4775:4768] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_597[12] = buffer_data_2[4783:4776] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_597[13] = buffer_data_2[4791:4784] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_597[14] = buffer_data_2[4799:4792] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_597[15] = buffer_data_1[4767:4760] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_597[16] = buffer_data_1[4775:4768] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_597[17] = buffer_data_1[4783:4776] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_597[18] = buffer_data_1[4791:4784] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_597[19] = buffer_data_1[4799:4792] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_597[20] = buffer_data_0[4767:4760] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_597[21] = buffer_data_0[4775:4768] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_597[22] = buffer_data_0[4783:4776] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_597[23] = buffer_data_0[4791:4784] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_597[24] = buffer_data_0[4799:4792] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_597 = kernel_img_mul_597[0] + kernel_img_mul_597[1] + kernel_img_mul_597[2] + 
                kernel_img_mul_597[3] + kernel_img_mul_597[4] + kernel_img_mul_597[5] + 
                kernel_img_mul_597[6] + kernel_img_mul_597[7] + kernel_img_mul_597[8] + 
                kernel_img_mul_597[9] + kernel_img_mul_597[10] + kernel_img_mul_597[11] + 
                kernel_img_mul_597[12] + kernel_img_mul_597[13] + kernel_img_mul_597[14] + 
                kernel_img_mul_597[15] + kernel_img_mul_597[16] + kernel_img_mul_597[17] + 
                kernel_img_mul_597[18] + kernel_img_mul_597[19] + kernel_img_mul_597[20] + 
                kernel_img_mul_597[21] + kernel_img_mul_597[22] + kernel_img_mul_597[23] + 
                kernel_img_mul_597[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4783:4776] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4783:4776] <= kernel_img_sum_597[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4783:4776] <= 'd0;
end

wire  [39:0]  kernel_img_mul_598[0:24];
assign kernel_img_mul_598[0] = buffer_data_4[4775:4768] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_598[1] = buffer_data_4[4783:4776] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_598[2] = buffer_data_4[4791:4784] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_598[3] = buffer_data_4[4799:4792] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_598[4] = buffer_data_4[4807:4800] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_598[5] = buffer_data_3[4775:4768] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_598[6] = buffer_data_3[4783:4776] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_598[7] = buffer_data_3[4791:4784] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_598[8] = buffer_data_3[4799:4792] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_598[9] = buffer_data_3[4807:4800] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_598[10] = buffer_data_2[4775:4768] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_598[11] = buffer_data_2[4783:4776] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_598[12] = buffer_data_2[4791:4784] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_598[13] = buffer_data_2[4799:4792] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_598[14] = buffer_data_2[4807:4800] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_598[15] = buffer_data_1[4775:4768] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_598[16] = buffer_data_1[4783:4776] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_598[17] = buffer_data_1[4791:4784] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_598[18] = buffer_data_1[4799:4792] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_598[19] = buffer_data_1[4807:4800] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_598[20] = buffer_data_0[4775:4768] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_598[21] = buffer_data_0[4783:4776] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_598[22] = buffer_data_0[4791:4784] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_598[23] = buffer_data_0[4799:4792] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_598[24] = buffer_data_0[4807:4800] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_598 = kernel_img_mul_598[0] + kernel_img_mul_598[1] + kernel_img_mul_598[2] + 
                kernel_img_mul_598[3] + kernel_img_mul_598[4] + kernel_img_mul_598[5] + 
                kernel_img_mul_598[6] + kernel_img_mul_598[7] + kernel_img_mul_598[8] + 
                kernel_img_mul_598[9] + kernel_img_mul_598[10] + kernel_img_mul_598[11] + 
                kernel_img_mul_598[12] + kernel_img_mul_598[13] + kernel_img_mul_598[14] + 
                kernel_img_mul_598[15] + kernel_img_mul_598[16] + kernel_img_mul_598[17] + 
                kernel_img_mul_598[18] + kernel_img_mul_598[19] + kernel_img_mul_598[20] + 
                kernel_img_mul_598[21] + kernel_img_mul_598[22] + kernel_img_mul_598[23] + 
                kernel_img_mul_598[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4791:4784] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4791:4784] <= kernel_img_sum_598[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4791:4784] <= 'd0;
end

wire  [39:0]  kernel_img_mul_599[0:24];
assign kernel_img_mul_599[0] = buffer_data_4[4783:4776] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_599[1] = buffer_data_4[4791:4784] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_599[2] = buffer_data_4[4799:4792] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_599[3] = buffer_data_4[4807:4800] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_599[4] = buffer_data_4[4815:4808] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_599[5] = buffer_data_3[4783:4776] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_599[6] = buffer_data_3[4791:4784] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_599[7] = buffer_data_3[4799:4792] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_599[8] = buffer_data_3[4807:4800] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_599[9] = buffer_data_3[4815:4808] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_599[10] = buffer_data_2[4783:4776] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_599[11] = buffer_data_2[4791:4784] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_599[12] = buffer_data_2[4799:4792] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_599[13] = buffer_data_2[4807:4800] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_599[14] = buffer_data_2[4815:4808] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_599[15] = buffer_data_1[4783:4776] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_599[16] = buffer_data_1[4791:4784] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_599[17] = buffer_data_1[4799:4792] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_599[18] = buffer_data_1[4807:4800] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_599[19] = buffer_data_1[4815:4808] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_599[20] = buffer_data_0[4783:4776] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_599[21] = buffer_data_0[4791:4784] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_599[22] = buffer_data_0[4799:4792] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_599[23] = buffer_data_0[4807:4800] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_599[24] = buffer_data_0[4815:4808] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_599 = kernel_img_mul_599[0] + kernel_img_mul_599[1] + kernel_img_mul_599[2] + 
                kernel_img_mul_599[3] + kernel_img_mul_599[4] + kernel_img_mul_599[5] + 
                kernel_img_mul_599[6] + kernel_img_mul_599[7] + kernel_img_mul_599[8] + 
                kernel_img_mul_599[9] + kernel_img_mul_599[10] + kernel_img_mul_599[11] + 
                kernel_img_mul_599[12] + kernel_img_mul_599[13] + kernel_img_mul_599[14] + 
                kernel_img_mul_599[15] + kernel_img_mul_599[16] + kernel_img_mul_599[17] + 
                kernel_img_mul_599[18] + kernel_img_mul_599[19] + kernel_img_mul_599[20] + 
                kernel_img_mul_599[21] + kernel_img_mul_599[22] + kernel_img_mul_599[23] + 
                kernel_img_mul_599[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4799:4792] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4799:4792] <= kernel_img_sum_599[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4799:4792] <= 'd0;
end

wire  [39:0]  kernel_img_mul_600[0:24];
assign kernel_img_mul_600[0] = buffer_data_4[4791:4784] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_600[1] = buffer_data_4[4799:4792] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_600[2] = buffer_data_4[4807:4800] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_600[3] = buffer_data_4[4815:4808] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_600[4] = buffer_data_4[4823:4816] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_600[5] = buffer_data_3[4791:4784] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_600[6] = buffer_data_3[4799:4792] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_600[7] = buffer_data_3[4807:4800] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_600[8] = buffer_data_3[4815:4808] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_600[9] = buffer_data_3[4823:4816] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_600[10] = buffer_data_2[4791:4784] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_600[11] = buffer_data_2[4799:4792] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_600[12] = buffer_data_2[4807:4800] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_600[13] = buffer_data_2[4815:4808] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_600[14] = buffer_data_2[4823:4816] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_600[15] = buffer_data_1[4791:4784] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_600[16] = buffer_data_1[4799:4792] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_600[17] = buffer_data_1[4807:4800] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_600[18] = buffer_data_1[4815:4808] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_600[19] = buffer_data_1[4823:4816] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_600[20] = buffer_data_0[4791:4784] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_600[21] = buffer_data_0[4799:4792] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_600[22] = buffer_data_0[4807:4800] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_600[23] = buffer_data_0[4815:4808] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_600[24] = buffer_data_0[4823:4816] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_600 = kernel_img_mul_600[0] + kernel_img_mul_600[1] + kernel_img_mul_600[2] + 
                kernel_img_mul_600[3] + kernel_img_mul_600[4] + kernel_img_mul_600[5] + 
                kernel_img_mul_600[6] + kernel_img_mul_600[7] + kernel_img_mul_600[8] + 
                kernel_img_mul_600[9] + kernel_img_mul_600[10] + kernel_img_mul_600[11] + 
                kernel_img_mul_600[12] + kernel_img_mul_600[13] + kernel_img_mul_600[14] + 
                kernel_img_mul_600[15] + kernel_img_mul_600[16] + kernel_img_mul_600[17] + 
                kernel_img_mul_600[18] + kernel_img_mul_600[19] + kernel_img_mul_600[20] + 
                kernel_img_mul_600[21] + kernel_img_mul_600[22] + kernel_img_mul_600[23] + 
                kernel_img_mul_600[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4807:4800] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4807:4800] <= kernel_img_sum_600[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4807:4800] <= 'd0;
end

wire  [39:0]  kernel_img_mul_601[0:24];
assign kernel_img_mul_601[0] = buffer_data_4[4799:4792] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_601[1] = buffer_data_4[4807:4800] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_601[2] = buffer_data_4[4815:4808] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_601[3] = buffer_data_4[4823:4816] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_601[4] = buffer_data_4[4831:4824] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_601[5] = buffer_data_3[4799:4792] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_601[6] = buffer_data_3[4807:4800] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_601[7] = buffer_data_3[4815:4808] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_601[8] = buffer_data_3[4823:4816] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_601[9] = buffer_data_3[4831:4824] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_601[10] = buffer_data_2[4799:4792] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_601[11] = buffer_data_2[4807:4800] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_601[12] = buffer_data_2[4815:4808] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_601[13] = buffer_data_2[4823:4816] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_601[14] = buffer_data_2[4831:4824] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_601[15] = buffer_data_1[4799:4792] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_601[16] = buffer_data_1[4807:4800] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_601[17] = buffer_data_1[4815:4808] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_601[18] = buffer_data_1[4823:4816] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_601[19] = buffer_data_1[4831:4824] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_601[20] = buffer_data_0[4799:4792] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_601[21] = buffer_data_0[4807:4800] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_601[22] = buffer_data_0[4815:4808] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_601[23] = buffer_data_0[4823:4816] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_601[24] = buffer_data_0[4831:4824] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_601 = kernel_img_mul_601[0] + kernel_img_mul_601[1] + kernel_img_mul_601[2] + 
                kernel_img_mul_601[3] + kernel_img_mul_601[4] + kernel_img_mul_601[5] + 
                kernel_img_mul_601[6] + kernel_img_mul_601[7] + kernel_img_mul_601[8] + 
                kernel_img_mul_601[9] + kernel_img_mul_601[10] + kernel_img_mul_601[11] + 
                kernel_img_mul_601[12] + kernel_img_mul_601[13] + kernel_img_mul_601[14] + 
                kernel_img_mul_601[15] + kernel_img_mul_601[16] + kernel_img_mul_601[17] + 
                kernel_img_mul_601[18] + kernel_img_mul_601[19] + kernel_img_mul_601[20] + 
                kernel_img_mul_601[21] + kernel_img_mul_601[22] + kernel_img_mul_601[23] + 
                kernel_img_mul_601[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4815:4808] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4815:4808] <= kernel_img_sum_601[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4815:4808] <= 'd0;
end

wire  [39:0]  kernel_img_mul_602[0:24];
assign kernel_img_mul_602[0] = buffer_data_4[4807:4800] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_602[1] = buffer_data_4[4815:4808] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_602[2] = buffer_data_4[4823:4816] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_602[3] = buffer_data_4[4831:4824] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_602[4] = buffer_data_4[4839:4832] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_602[5] = buffer_data_3[4807:4800] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_602[6] = buffer_data_3[4815:4808] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_602[7] = buffer_data_3[4823:4816] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_602[8] = buffer_data_3[4831:4824] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_602[9] = buffer_data_3[4839:4832] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_602[10] = buffer_data_2[4807:4800] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_602[11] = buffer_data_2[4815:4808] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_602[12] = buffer_data_2[4823:4816] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_602[13] = buffer_data_2[4831:4824] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_602[14] = buffer_data_2[4839:4832] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_602[15] = buffer_data_1[4807:4800] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_602[16] = buffer_data_1[4815:4808] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_602[17] = buffer_data_1[4823:4816] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_602[18] = buffer_data_1[4831:4824] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_602[19] = buffer_data_1[4839:4832] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_602[20] = buffer_data_0[4807:4800] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_602[21] = buffer_data_0[4815:4808] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_602[22] = buffer_data_0[4823:4816] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_602[23] = buffer_data_0[4831:4824] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_602[24] = buffer_data_0[4839:4832] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_602 = kernel_img_mul_602[0] + kernel_img_mul_602[1] + kernel_img_mul_602[2] + 
                kernel_img_mul_602[3] + kernel_img_mul_602[4] + kernel_img_mul_602[5] + 
                kernel_img_mul_602[6] + kernel_img_mul_602[7] + kernel_img_mul_602[8] + 
                kernel_img_mul_602[9] + kernel_img_mul_602[10] + kernel_img_mul_602[11] + 
                kernel_img_mul_602[12] + kernel_img_mul_602[13] + kernel_img_mul_602[14] + 
                kernel_img_mul_602[15] + kernel_img_mul_602[16] + kernel_img_mul_602[17] + 
                kernel_img_mul_602[18] + kernel_img_mul_602[19] + kernel_img_mul_602[20] + 
                kernel_img_mul_602[21] + kernel_img_mul_602[22] + kernel_img_mul_602[23] + 
                kernel_img_mul_602[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4823:4816] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4823:4816] <= kernel_img_sum_602[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4823:4816] <= 'd0;
end

wire  [39:0]  kernel_img_mul_603[0:24];
assign kernel_img_mul_603[0] = buffer_data_4[4815:4808] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_603[1] = buffer_data_4[4823:4816] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_603[2] = buffer_data_4[4831:4824] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_603[3] = buffer_data_4[4839:4832] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_603[4] = buffer_data_4[4847:4840] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_603[5] = buffer_data_3[4815:4808] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_603[6] = buffer_data_3[4823:4816] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_603[7] = buffer_data_3[4831:4824] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_603[8] = buffer_data_3[4839:4832] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_603[9] = buffer_data_3[4847:4840] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_603[10] = buffer_data_2[4815:4808] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_603[11] = buffer_data_2[4823:4816] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_603[12] = buffer_data_2[4831:4824] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_603[13] = buffer_data_2[4839:4832] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_603[14] = buffer_data_2[4847:4840] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_603[15] = buffer_data_1[4815:4808] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_603[16] = buffer_data_1[4823:4816] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_603[17] = buffer_data_1[4831:4824] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_603[18] = buffer_data_1[4839:4832] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_603[19] = buffer_data_1[4847:4840] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_603[20] = buffer_data_0[4815:4808] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_603[21] = buffer_data_0[4823:4816] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_603[22] = buffer_data_0[4831:4824] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_603[23] = buffer_data_0[4839:4832] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_603[24] = buffer_data_0[4847:4840] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_603 = kernel_img_mul_603[0] + kernel_img_mul_603[1] + kernel_img_mul_603[2] + 
                kernel_img_mul_603[3] + kernel_img_mul_603[4] + kernel_img_mul_603[5] + 
                kernel_img_mul_603[6] + kernel_img_mul_603[7] + kernel_img_mul_603[8] + 
                kernel_img_mul_603[9] + kernel_img_mul_603[10] + kernel_img_mul_603[11] + 
                kernel_img_mul_603[12] + kernel_img_mul_603[13] + kernel_img_mul_603[14] + 
                kernel_img_mul_603[15] + kernel_img_mul_603[16] + kernel_img_mul_603[17] + 
                kernel_img_mul_603[18] + kernel_img_mul_603[19] + kernel_img_mul_603[20] + 
                kernel_img_mul_603[21] + kernel_img_mul_603[22] + kernel_img_mul_603[23] + 
                kernel_img_mul_603[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4831:4824] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4831:4824] <= kernel_img_sum_603[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4831:4824] <= 'd0;
end

wire  [39:0]  kernel_img_mul_604[0:24];
assign kernel_img_mul_604[0] = buffer_data_4[4823:4816] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_604[1] = buffer_data_4[4831:4824] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_604[2] = buffer_data_4[4839:4832] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_604[3] = buffer_data_4[4847:4840] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_604[4] = buffer_data_4[4855:4848] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_604[5] = buffer_data_3[4823:4816] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_604[6] = buffer_data_3[4831:4824] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_604[7] = buffer_data_3[4839:4832] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_604[8] = buffer_data_3[4847:4840] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_604[9] = buffer_data_3[4855:4848] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_604[10] = buffer_data_2[4823:4816] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_604[11] = buffer_data_2[4831:4824] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_604[12] = buffer_data_2[4839:4832] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_604[13] = buffer_data_2[4847:4840] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_604[14] = buffer_data_2[4855:4848] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_604[15] = buffer_data_1[4823:4816] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_604[16] = buffer_data_1[4831:4824] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_604[17] = buffer_data_1[4839:4832] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_604[18] = buffer_data_1[4847:4840] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_604[19] = buffer_data_1[4855:4848] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_604[20] = buffer_data_0[4823:4816] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_604[21] = buffer_data_0[4831:4824] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_604[22] = buffer_data_0[4839:4832] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_604[23] = buffer_data_0[4847:4840] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_604[24] = buffer_data_0[4855:4848] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_604 = kernel_img_mul_604[0] + kernel_img_mul_604[1] + kernel_img_mul_604[2] + 
                kernel_img_mul_604[3] + kernel_img_mul_604[4] + kernel_img_mul_604[5] + 
                kernel_img_mul_604[6] + kernel_img_mul_604[7] + kernel_img_mul_604[8] + 
                kernel_img_mul_604[9] + kernel_img_mul_604[10] + kernel_img_mul_604[11] + 
                kernel_img_mul_604[12] + kernel_img_mul_604[13] + kernel_img_mul_604[14] + 
                kernel_img_mul_604[15] + kernel_img_mul_604[16] + kernel_img_mul_604[17] + 
                kernel_img_mul_604[18] + kernel_img_mul_604[19] + kernel_img_mul_604[20] + 
                kernel_img_mul_604[21] + kernel_img_mul_604[22] + kernel_img_mul_604[23] + 
                kernel_img_mul_604[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4839:4832] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4839:4832] <= kernel_img_sum_604[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4839:4832] <= 'd0;
end

wire  [39:0]  kernel_img_mul_605[0:24];
assign kernel_img_mul_605[0] = buffer_data_4[4831:4824] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_605[1] = buffer_data_4[4839:4832] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_605[2] = buffer_data_4[4847:4840] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_605[3] = buffer_data_4[4855:4848] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_605[4] = buffer_data_4[4863:4856] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_605[5] = buffer_data_3[4831:4824] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_605[6] = buffer_data_3[4839:4832] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_605[7] = buffer_data_3[4847:4840] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_605[8] = buffer_data_3[4855:4848] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_605[9] = buffer_data_3[4863:4856] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_605[10] = buffer_data_2[4831:4824] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_605[11] = buffer_data_2[4839:4832] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_605[12] = buffer_data_2[4847:4840] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_605[13] = buffer_data_2[4855:4848] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_605[14] = buffer_data_2[4863:4856] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_605[15] = buffer_data_1[4831:4824] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_605[16] = buffer_data_1[4839:4832] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_605[17] = buffer_data_1[4847:4840] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_605[18] = buffer_data_1[4855:4848] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_605[19] = buffer_data_1[4863:4856] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_605[20] = buffer_data_0[4831:4824] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_605[21] = buffer_data_0[4839:4832] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_605[22] = buffer_data_0[4847:4840] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_605[23] = buffer_data_0[4855:4848] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_605[24] = buffer_data_0[4863:4856] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_605 = kernel_img_mul_605[0] + kernel_img_mul_605[1] + kernel_img_mul_605[2] + 
                kernel_img_mul_605[3] + kernel_img_mul_605[4] + kernel_img_mul_605[5] + 
                kernel_img_mul_605[6] + kernel_img_mul_605[7] + kernel_img_mul_605[8] + 
                kernel_img_mul_605[9] + kernel_img_mul_605[10] + kernel_img_mul_605[11] + 
                kernel_img_mul_605[12] + kernel_img_mul_605[13] + kernel_img_mul_605[14] + 
                kernel_img_mul_605[15] + kernel_img_mul_605[16] + kernel_img_mul_605[17] + 
                kernel_img_mul_605[18] + kernel_img_mul_605[19] + kernel_img_mul_605[20] + 
                kernel_img_mul_605[21] + kernel_img_mul_605[22] + kernel_img_mul_605[23] + 
                kernel_img_mul_605[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4847:4840] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4847:4840] <= kernel_img_sum_605[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4847:4840] <= 'd0;
end

wire  [39:0]  kernel_img_mul_606[0:24];
assign kernel_img_mul_606[0] = buffer_data_4[4839:4832] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_606[1] = buffer_data_4[4847:4840] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_606[2] = buffer_data_4[4855:4848] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_606[3] = buffer_data_4[4863:4856] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_606[4] = buffer_data_4[4871:4864] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_606[5] = buffer_data_3[4839:4832] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_606[6] = buffer_data_3[4847:4840] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_606[7] = buffer_data_3[4855:4848] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_606[8] = buffer_data_3[4863:4856] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_606[9] = buffer_data_3[4871:4864] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_606[10] = buffer_data_2[4839:4832] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_606[11] = buffer_data_2[4847:4840] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_606[12] = buffer_data_2[4855:4848] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_606[13] = buffer_data_2[4863:4856] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_606[14] = buffer_data_2[4871:4864] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_606[15] = buffer_data_1[4839:4832] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_606[16] = buffer_data_1[4847:4840] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_606[17] = buffer_data_1[4855:4848] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_606[18] = buffer_data_1[4863:4856] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_606[19] = buffer_data_1[4871:4864] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_606[20] = buffer_data_0[4839:4832] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_606[21] = buffer_data_0[4847:4840] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_606[22] = buffer_data_0[4855:4848] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_606[23] = buffer_data_0[4863:4856] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_606[24] = buffer_data_0[4871:4864] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_606 = kernel_img_mul_606[0] + kernel_img_mul_606[1] + kernel_img_mul_606[2] + 
                kernel_img_mul_606[3] + kernel_img_mul_606[4] + kernel_img_mul_606[5] + 
                kernel_img_mul_606[6] + kernel_img_mul_606[7] + kernel_img_mul_606[8] + 
                kernel_img_mul_606[9] + kernel_img_mul_606[10] + kernel_img_mul_606[11] + 
                kernel_img_mul_606[12] + kernel_img_mul_606[13] + kernel_img_mul_606[14] + 
                kernel_img_mul_606[15] + kernel_img_mul_606[16] + kernel_img_mul_606[17] + 
                kernel_img_mul_606[18] + kernel_img_mul_606[19] + kernel_img_mul_606[20] + 
                kernel_img_mul_606[21] + kernel_img_mul_606[22] + kernel_img_mul_606[23] + 
                kernel_img_mul_606[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4855:4848] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4855:4848] <= kernel_img_sum_606[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4855:4848] <= 'd0;
end

wire  [39:0]  kernel_img_mul_607[0:24];
assign kernel_img_mul_607[0] = buffer_data_4[4847:4840] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_607[1] = buffer_data_4[4855:4848] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_607[2] = buffer_data_4[4863:4856] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_607[3] = buffer_data_4[4871:4864] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_607[4] = buffer_data_4[4879:4872] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_607[5] = buffer_data_3[4847:4840] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_607[6] = buffer_data_3[4855:4848] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_607[7] = buffer_data_3[4863:4856] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_607[8] = buffer_data_3[4871:4864] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_607[9] = buffer_data_3[4879:4872] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_607[10] = buffer_data_2[4847:4840] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_607[11] = buffer_data_2[4855:4848] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_607[12] = buffer_data_2[4863:4856] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_607[13] = buffer_data_2[4871:4864] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_607[14] = buffer_data_2[4879:4872] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_607[15] = buffer_data_1[4847:4840] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_607[16] = buffer_data_1[4855:4848] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_607[17] = buffer_data_1[4863:4856] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_607[18] = buffer_data_1[4871:4864] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_607[19] = buffer_data_1[4879:4872] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_607[20] = buffer_data_0[4847:4840] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_607[21] = buffer_data_0[4855:4848] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_607[22] = buffer_data_0[4863:4856] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_607[23] = buffer_data_0[4871:4864] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_607[24] = buffer_data_0[4879:4872] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_607 = kernel_img_mul_607[0] + kernel_img_mul_607[1] + kernel_img_mul_607[2] + 
                kernel_img_mul_607[3] + kernel_img_mul_607[4] + kernel_img_mul_607[5] + 
                kernel_img_mul_607[6] + kernel_img_mul_607[7] + kernel_img_mul_607[8] + 
                kernel_img_mul_607[9] + kernel_img_mul_607[10] + kernel_img_mul_607[11] + 
                kernel_img_mul_607[12] + kernel_img_mul_607[13] + kernel_img_mul_607[14] + 
                kernel_img_mul_607[15] + kernel_img_mul_607[16] + kernel_img_mul_607[17] + 
                kernel_img_mul_607[18] + kernel_img_mul_607[19] + kernel_img_mul_607[20] + 
                kernel_img_mul_607[21] + kernel_img_mul_607[22] + kernel_img_mul_607[23] + 
                kernel_img_mul_607[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4863:4856] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4863:4856] <= kernel_img_sum_607[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4863:4856] <= 'd0;
end

wire  [39:0]  kernel_img_mul_608[0:24];
assign kernel_img_mul_608[0] = buffer_data_4[4855:4848] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_608[1] = buffer_data_4[4863:4856] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_608[2] = buffer_data_4[4871:4864] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_608[3] = buffer_data_4[4879:4872] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_608[4] = buffer_data_4[4887:4880] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_608[5] = buffer_data_3[4855:4848] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_608[6] = buffer_data_3[4863:4856] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_608[7] = buffer_data_3[4871:4864] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_608[8] = buffer_data_3[4879:4872] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_608[9] = buffer_data_3[4887:4880] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_608[10] = buffer_data_2[4855:4848] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_608[11] = buffer_data_2[4863:4856] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_608[12] = buffer_data_2[4871:4864] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_608[13] = buffer_data_2[4879:4872] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_608[14] = buffer_data_2[4887:4880] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_608[15] = buffer_data_1[4855:4848] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_608[16] = buffer_data_1[4863:4856] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_608[17] = buffer_data_1[4871:4864] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_608[18] = buffer_data_1[4879:4872] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_608[19] = buffer_data_1[4887:4880] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_608[20] = buffer_data_0[4855:4848] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_608[21] = buffer_data_0[4863:4856] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_608[22] = buffer_data_0[4871:4864] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_608[23] = buffer_data_0[4879:4872] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_608[24] = buffer_data_0[4887:4880] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_608 = kernel_img_mul_608[0] + kernel_img_mul_608[1] + kernel_img_mul_608[2] + 
                kernel_img_mul_608[3] + kernel_img_mul_608[4] + kernel_img_mul_608[5] + 
                kernel_img_mul_608[6] + kernel_img_mul_608[7] + kernel_img_mul_608[8] + 
                kernel_img_mul_608[9] + kernel_img_mul_608[10] + kernel_img_mul_608[11] + 
                kernel_img_mul_608[12] + kernel_img_mul_608[13] + kernel_img_mul_608[14] + 
                kernel_img_mul_608[15] + kernel_img_mul_608[16] + kernel_img_mul_608[17] + 
                kernel_img_mul_608[18] + kernel_img_mul_608[19] + kernel_img_mul_608[20] + 
                kernel_img_mul_608[21] + kernel_img_mul_608[22] + kernel_img_mul_608[23] + 
                kernel_img_mul_608[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4871:4864] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4871:4864] <= kernel_img_sum_608[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4871:4864] <= 'd0;
end

wire  [39:0]  kernel_img_mul_609[0:24];
assign kernel_img_mul_609[0] = buffer_data_4[4863:4856] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_609[1] = buffer_data_4[4871:4864] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_609[2] = buffer_data_4[4879:4872] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_609[3] = buffer_data_4[4887:4880] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_609[4] = buffer_data_4[4895:4888] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_609[5] = buffer_data_3[4863:4856] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_609[6] = buffer_data_3[4871:4864] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_609[7] = buffer_data_3[4879:4872] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_609[8] = buffer_data_3[4887:4880] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_609[9] = buffer_data_3[4895:4888] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_609[10] = buffer_data_2[4863:4856] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_609[11] = buffer_data_2[4871:4864] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_609[12] = buffer_data_2[4879:4872] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_609[13] = buffer_data_2[4887:4880] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_609[14] = buffer_data_2[4895:4888] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_609[15] = buffer_data_1[4863:4856] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_609[16] = buffer_data_1[4871:4864] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_609[17] = buffer_data_1[4879:4872] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_609[18] = buffer_data_1[4887:4880] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_609[19] = buffer_data_1[4895:4888] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_609[20] = buffer_data_0[4863:4856] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_609[21] = buffer_data_0[4871:4864] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_609[22] = buffer_data_0[4879:4872] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_609[23] = buffer_data_0[4887:4880] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_609[24] = buffer_data_0[4895:4888] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_609 = kernel_img_mul_609[0] + kernel_img_mul_609[1] + kernel_img_mul_609[2] + 
                kernel_img_mul_609[3] + kernel_img_mul_609[4] + kernel_img_mul_609[5] + 
                kernel_img_mul_609[6] + kernel_img_mul_609[7] + kernel_img_mul_609[8] + 
                kernel_img_mul_609[9] + kernel_img_mul_609[10] + kernel_img_mul_609[11] + 
                kernel_img_mul_609[12] + kernel_img_mul_609[13] + kernel_img_mul_609[14] + 
                kernel_img_mul_609[15] + kernel_img_mul_609[16] + kernel_img_mul_609[17] + 
                kernel_img_mul_609[18] + kernel_img_mul_609[19] + kernel_img_mul_609[20] + 
                kernel_img_mul_609[21] + kernel_img_mul_609[22] + kernel_img_mul_609[23] + 
                kernel_img_mul_609[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4879:4872] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4879:4872] <= kernel_img_sum_609[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4879:4872] <= 'd0;
end

wire  [39:0]  kernel_img_mul_610[0:24];
assign kernel_img_mul_610[0] = buffer_data_4[4871:4864] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_610[1] = buffer_data_4[4879:4872] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_610[2] = buffer_data_4[4887:4880] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_610[3] = buffer_data_4[4895:4888] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_610[4] = buffer_data_4[4903:4896] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_610[5] = buffer_data_3[4871:4864] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_610[6] = buffer_data_3[4879:4872] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_610[7] = buffer_data_3[4887:4880] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_610[8] = buffer_data_3[4895:4888] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_610[9] = buffer_data_3[4903:4896] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_610[10] = buffer_data_2[4871:4864] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_610[11] = buffer_data_2[4879:4872] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_610[12] = buffer_data_2[4887:4880] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_610[13] = buffer_data_2[4895:4888] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_610[14] = buffer_data_2[4903:4896] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_610[15] = buffer_data_1[4871:4864] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_610[16] = buffer_data_1[4879:4872] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_610[17] = buffer_data_1[4887:4880] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_610[18] = buffer_data_1[4895:4888] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_610[19] = buffer_data_1[4903:4896] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_610[20] = buffer_data_0[4871:4864] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_610[21] = buffer_data_0[4879:4872] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_610[22] = buffer_data_0[4887:4880] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_610[23] = buffer_data_0[4895:4888] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_610[24] = buffer_data_0[4903:4896] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_610 = kernel_img_mul_610[0] + kernel_img_mul_610[1] + kernel_img_mul_610[2] + 
                kernel_img_mul_610[3] + kernel_img_mul_610[4] + kernel_img_mul_610[5] + 
                kernel_img_mul_610[6] + kernel_img_mul_610[7] + kernel_img_mul_610[8] + 
                kernel_img_mul_610[9] + kernel_img_mul_610[10] + kernel_img_mul_610[11] + 
                kernel_img_mul_610[12] + kernel_img_mul_610[13] + kernel_img_mul_610[14] + 
                kernel_img_mul_610[15] + kernel_img_mul_610[16] + kernel_img_mul_610[17] + 
                kernel_img_mul_610[18] + kernel_img_mul_610[19] + kernel_img_mul_610[20] + 
                kernel_img_mul_610[21] + kernel_img_mul_610[22] + kernel_img_mul_610[23] + 
                kernel_img_mul_610[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4887:4880] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4887:4880] <= kernel_img_sum_610[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4887:4880] <= 'd0;
end

wire  [39:0]  kernel_img_mul_611[0:24];
assign kernel_img_mul_611[0] = buffer_data_4[4879:4872] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_611[1] = buffer_data_4[4887:4880] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_611[2] = buffer_data_4[4895:4888] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_611[3] = buffer_data_4[4903:4896] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_611[4] = buffer_data_4[4911:4904] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_611[5] = buffer_data_3[4879:4872] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_611[6] = buffer_data_3[4887:4880] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_611[7] = buffer_data_3[4895:4888] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_611[8] = buffer_data_3[4903:4896] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_611[9] = buffer_data_3[4911:4904] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_611[10] = buffer_data_2[4879:4872] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_611[11] = buffer_data_2[4887:4880] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_611[12] = buffer_data_2[4895:4888] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_611[13] = buffer_data_2[4903:4896] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_611[14] = buffer_data_2[4911:4904] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_611[15] = buffer_data_1[4879:4872] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_611[16] = buffer_data_1[4887:4880] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_611[17] = buffer_data_1[4895:4888] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_611[18] = buffer_data_1[4903:4896] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_611[19] = buffer_data_1[4911:4904] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_611[20] = buffer_data_0[4879:4872] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_611[21] = buffer_data_0[4887:4880] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_611[22] = buffer_data_0[4895:4888] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_611[23] = buffer_data_0[4903:4896] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_611[24] = buffer_data_0[4911:4904] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_611 = kernel_img_mul_611[0] + kernel_img_mul_611[1] + kernel_img_mul_611[2] + 
                kernel_img_mul_611[3] + kernel_img_mul_611[4] + kernel_img_mul_611[5] + 
                kernel_img_mul_611[6] + kernel_img_mul_611[7] + kernel_img_mul_611[8] + 
                kernel_img_mul_611[9] + kernel_img_mul_611[10] + kernel_img_mul_611[11] + 
                kernel_img_mul_611[12] + kernel_img_mul_611[13] + kernel_img_mul_611[14] + 
                kernel_img_mul_611[15] + kernel_img_mul_611[16] + kernel_img_mul_611[17] + 
                kernel_img_mul_611[18] + kernel_img_mul_611[19] + kernel_img_mul_611[20] + 
                kernel_img_mul_611[21] + kernel_img_mul_611[22] + kernel_img_mul_611[23] + 
                kernel_img_mul_611[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4895:4888] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4895:4888] <= kernel_img_sum_611[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4895:4888] <= 'd0;
end

wire  [39:0]  kernel_img_mul_612[0:24];
assign kernel_img_mul_612[0] = buffer_data_4[4887:4880] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_612[1] = buffer_data_4[4895:4888] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_612[2] = buffer_data_4[4903:4896] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_612[3] = buffer_data_4[4911:4904] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_612[4] = buffer_data_4[4919:4912] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_612[5] = buffer_data_3[4887:4880] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_612[6] = buffer_data_3[4895:4888] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_612[7] = buffer_data_3[4903:4896] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_612[8] = buffer_data_3[4911:4904] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_612[9] = buffer_data_3[4919:4912] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_612[10] = buffer_data_2[4887:4880] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_612[11] = buffer_data_2[4895:4888] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_612[12] = buffer_data_2[4903:4896] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_612[13] = buffer_data_2[4911:4904] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_612[14] = buffer_data_2[4919:4912] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_612[15] = buffer_data_1[4887:4880] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_612[16] = buffer_data_1[4895:4888] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_612[17] = buffer_data_1[4903:4896] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_612[18] = buffer_data_1[4911:4904] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_612[19] = buffer_data_1[4919:4912] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_612[20] = buffer_data_0[4887:4880] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_612[21] = buffer_data_0[4895:4888] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_612[22] = buffer_data_0[4903:4896] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_612[23] = buffer_data_0[4911:4904] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_612[24] = buffer_data_0[4919:4912] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_612 = kernel_img_mul_612[0] + kernel_img_mul_612[1] + kernel_img_mul_612[2] + 
                kernel_img_mul_612[3] + kernel_img_mul_612[4] + kernel_img_mul_612[5] + 
                kernel_img_mul_612[6] + kernel_img_mul_612[7] + kernel_img_mul_612[8] + 
                kernel_img_mul_612[9] + kernel_img_mul_612[10] + kernel_img_mul_612[11] + 
                kernel_img_mul_612[12] + kernel_img_mul_612[13] + kernel_img_mul_612[14] + 
                kernel_img_mul_612[15] + kernel_img_mul_612[16] + kernel_img_mul_612[17] + 
                kernel_img_mul_612[18] + kernel_img_mul_612[19] + kernel_img_mul_612[20] + 
                kernel_img_mul_612[21] + kernel_img_mul_612[22] + kernel_img_mul_612[23] + 
                kernel_img_mul_612[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4903:4896] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4903:4896] <= kernel_img_sum_612[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4903:4896] <= 'd0;
end

wire  [39:0]  kernel_img_mul_613[0:24];
assign kernel_img_mul_613[0] = buffer_data_4[4895:4888] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_613[1] = buffer_data_4[4903:4896] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_613[2] = buffer_data_4[4911:4904] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_613[3] = buffer_data_4[4919:4912] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_613[4] = buffer_data_4[4927:4920] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_613[5] = buffer_data_3[4895:4888] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_613[6] = buffer_data_3[4903:4896] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_613[7] = buffer_data_3[4911:4904] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_613[8] = buffer_data_3[4919:4912] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_613[9] = buffer_data_3[4927:4920] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_613[10] = buffer_data_2[4895:4888] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_613[11] = buffer_data_2[4903:4896] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_613[12] = buffer_data_2[4911:4904] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_613[13] = buffer_data_2[4919:4912] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_613[14] = buffer_data_2[4927:4920] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_613[15] = buffer_data_1[4895:4888] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_613[16] = buffer_data_1[4903:4896] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_613[17] = buffer_data_1[4911:4904] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_613[18] = buffer_data_1[4919:4912] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_613[19] = buffer_data_1[4927:4920] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_613[20] = buffer_data_0[4895:4888] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_613[21] = buffer_data_0[4903:4896] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_613[22] = buffer_data_0[4911:4904] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_613[23] = buffer_data_0[4919:4912] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_613[24] = buffer_data_0[4927:4920] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_613 = kernel_img_mul_613[0] + kernel_img_mul_613[1] + kernel_img_mul_613[2] + 
                kernel_img_mul_613[3] + kernel_img_mul_613[4] + kernel_img_mul_613[5] + 
                kernel_img_mul_613[6] + kernel_img_mul_613[7] + kernel_img_mul_613[8] + 
                kernel_img_mul_613[9] + kernel_img_mul_613[10] + kernel_img_mul_613[11] + 
                kernel_img_mul_613[12] + kernel_img_mul_613[13] + kernel_img_mul_613[14] + 
                kernel_img_mul_613[15] + kernel_img_mul_613[16] + kernel_img_mul_613[17] + 
                kernel_img_mul_613[18] + kernel_img_mul_613[19] + kernel_img_mul_613[20] + 
                kernel_img_mul_613[21] + kernel_img_mul_613[22] + kernel_img_mul_613[23] + 
                kernel_img_mul_613[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4911:4904] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4911:4904] <= kernel_img_sum_613[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4911:4904] <= 'd0;
end

wire  [39:0]  kernel_img_mul_614[0:24];
assign kernel_img_mul_614[0] = buffer_data_4[4903:4896] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_614[1] = buffer_data_4[4911:4904] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_614[2] = buffer_data_4[4919:4912] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_614[3] = buffer_data_4[4927:4920] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_614[4] = buffer_data_4[4935:4928] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_614[5] = buffer_data_3[4903:4896] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_614[6] = buffer_data_3[4911:4904] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_614[7] = buffer_data_3[4919:4912] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_614[8] = buffer_data_3[4927:4920] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_614[9] = buffer_data_3[4935:4928] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_614[10] = buffer_data_2[4903:4896] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_614[11] = buffer_data_2[4911:4904] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_614[12] = buffer_data_2[4919:4912] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_614[13] = buffer_data_2[4927:4920] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_614[14] = buffer_data_2[4935:4928] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_614[15] = buffer_data_1[4903:4896] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_614[16] = buffer_data_1[4911:4904] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_614[17] = buffer_data_1[4919:4912] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_614[18] = buffer_data_1[4927:4920] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_614[19] = buffer_data_1[4935:4928] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_614[20] = buffer_data_0[4903:4896] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_614[21] = buffer_data_0[4911:4904] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_614[22] = buffer_data_0[4919:4912] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_614[23] = buffer_data_0[4927:4920] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_614[24] = buffer_data_0[4935:4928] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_614 = kernel_img_mul_614[0] + kernel_img_mul_614[1] + kernel_img_mul_614[2] + 
                kernel_img_mul_614[3] + kernel_img_mul_614[4] + kernel_img_mul_614[5] + 
                kernel_img_mul_614[6] + kernel_img_mul_614[7] + kernel_img_mul_614[8] + 
                kernel_img_mul_614[9] + kernel_img_mul_614[10] + kernel_img_mul_614[11] + 
                kernel_img_mul_614[12] + kernel_img_mul_614[13] + kernel_img_mul_614[14] + 
                kernel_img_mul_614[15] + kernel_img_mul_614[16] + kernel_img_mul_614[17] + 
                kernel_img_mul_614[18] + kernel_img_mul_614[19] + kernel_img_mul_614[20] + 
                kernel_img_mul_614[21] + kernel_img_mul_614[22] + kernel_img_mul_614[23] + 
                kernel_img_mul_614[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4919:4912] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4919:4912] <= kernel_img_sum_614[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4919:4912] <= 'd0;
end

wire  [39:0]  kernel_img_mul_615[0:24];
assign kernel_img_mul_615[0] = buffer_data_4[4911:4904] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_615[1] = buffer_data_4[4919:4912] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_615[2] = buffer_data_4[4927:4920] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_615[3] = buffer_data_4[4935:4928] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_615[4] = buffer_data_4[4943:4936] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_615[5] = buffer_data_3[4911:4904] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_615[6] = buffer_data_3[4919:4912] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_615[7] = buffer_data_3[4927:4920] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_615[8] = buffer_data_3[4935:4928] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_615[9] = buffer_data_3[4943:4936] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_615[10] = buffer_data_2[4911:4904] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_615[11] = buffer_data_2[4919:4912] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_615[12] = buffer_data_2[4927:4920] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_615[13] = buffer_data_2[4935:4928] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_615[14] = buffer_data_2[4943:4936] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_615[15] = buffer_data_1[4911:4904] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_615[16] = buffer_data_1[4919:4912] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_615[17] = buffer_data_1[4927:4920] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_615[18] = buffer_data_1[4935:4928] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_615[19] = buffer_data_1[4943:4936] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_615[20] = buffer_data_0[4911:4904] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_615[21] = buffer_data_0[4919:4912] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_615[22] = buffer_data_0[4927:4920] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_615[23] = buffer_data_0[4935:4928] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_615[24] = buffer_data_0[4943:4936] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_615 = kernel_img_mul_615[0] + kernel_img_mul_615[1] + kernel_img_mul_615[2] + 
                kernel_img_mul_615[3] + kernel_img_mul_615[4] + kernel_img_mul_615[5] + 
                kernel_img_mul_615[6] + kernel_img_mul_615[7] + kernel_img_mul_615[8] + 
                kernel_img_mul_615[9] + kernel_img_mul_615[10] + kernel_img_mul_615[11] + 
                kernel_img_mul_615[12] + kernel_img_mul_615[13] + kernel_img_mul_615[14] + 
                kernel_img_mul_615[15] + kernel_img_mul_615[16] + kernel_img_mul_615[17] + 
                kernel_img_mul_615[18] + kernel_img_mul_615[19] + kernel_img_mul_615[20] + 
                kernel_img_mul_615[21] + kernel_img_mul_615[22] + kernel_img_mul_615[23] + 
                kernel_img_mul_615[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4927:4920] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4927:4920] <= kernel_img_sum_615[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4927:4920] <= 'd0;
end

wire  [39:0]  kernel_img_mul_616[0:24];
assign kernel_img_mul_616[0] = buffer_data_4[4919:4912] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_616[1] = buffer_data_4[4927:4920] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_616[2] = buffer_data_4[4935:4928] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_616[3] = buffer_data_4[4943:4936] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_616[4] = buffer_data_4[4951:4944] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_616[5] = buffer_data_3[4919:4912] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_616[6] = buffer_data_3[4927:4920] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_616[7] = buffer_data_3[4935:4928] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_616[8] = buffer_data_3[4943:4936] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_616[9] = buffer_data_3[4951:4944] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_616[10] = buffer_data_2[4919:4912] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_616[11] = buffer_data_2[4927:4920] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_616[12] = buffer_data_2[4935:4928] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_616[13] = buffer_data_2[4943:4936] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_616[14] = buffer_data_2[4951:4944] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_616[15] = buffer_data_1[4919:4912] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_616[16] = buffer_data_1[4927:4920] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_616[17] = buffer_data_1[4935:4928] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_616[18] = buffer_data_1[4943:4936] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_616[19] = buffer_data_1[4951:4944] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_616[20] = buffer_data_0[4919:4912] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_616[21] = buffer_data_0[4927:4920] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_616[22] = buffer_data_0[4935:4928] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_616[23] = buffer_data_0[4943:4936] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_616[24] = buffer_data_0[4951:4944] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_616 = kernel_img_mul_616[0] + kernel_img_mul_616[1] + kernel_img_mul_616[2] + 
                kernel_img_mul_616[3] + kernel_img_mul_616[4] + kernel_img_mul_616[5] + 
                kernel_img_mul_616[6] + kernel_img_mul_616[7] + kernel_img_mul_616[8] + 
                kernel_img_mul_616[9] + kernel_img_mul_616[10] + kernel_img_mul_616[11] + 
                kernel_img_mul_616[12] + kernel_img_mul_616[13] + kernel_img_mul_616[14] + 
                kernel_img_mul_616[15] + kernel_img_mul_616[16] + kernel_img_mul_616[17] + 
                kernel_img_mul_616[18] + kernel_img_mul_616[19] + kernel_img_mul_616[20] + 
                kernel_img_mul_616[21] + kernel_img_mul_616[22] + kernel_img_mul_616[23] + 
                kernel_img_mul_616[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4935:4928] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4935:4928] <= kernel_img_sum_616[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4935:4928] <= 'd0;
end

wire  [39:0]  kernel_img_mul_617[0:24];
assign kernel_img_mul_617[0] = buffer_data_4[4927:4920] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_617[1] = buffer_data_4[4935:4928] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_617[2] = buffer_data_4[4943:4936] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_617[3] = buffer_data_4[4951:4944] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_617[4] = buffer_data_4[4959:4952] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_617[5] = buffer_data_3[4927:4920] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_617[6] = buffer_data_3[4935:4928] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_617[7] = buffer_data_3[4943:4936] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_617[8] = buffer_data_3[4951:4944] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_617[9] = buffer_data_3[4959:4952] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_617[10] = buffer_data_2[4927:4920] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_617[11] = buffer_data_2[4935:4928] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_617[12] = buffer_data_2[4943:4936] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_617[13] = buffer_data_2[4951:4944] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_617[14] = buffer_data_2[4959:4952] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_617[15] = buffer_data_1[4927:4920] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_617[16] = buffer_data_1[4935:4928] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_617[17] = buffer_data_1[4943:4936] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_617[18] = buffer_data_1[4951:4944] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_617[19] = buffer_data_1[4959:4952] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_617[20] = buffer_data_0[4927:4920] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_617[21] = buffer_data_0[4935:4928] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_617[22] = buffer_data_0[4943:4936] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_617[23] = buffer_data_0[4951:4944] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_617[24] = buffer_data_0[4959:4952] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_617 = kernel_img_mul_617[0] + kernel_img_mul_617[1] + kernel_img_mul_617[2] + 
                kernel_img_mul_617[3] + kernel_img_mul_617[4] + kernel_img_mul_617[5] + 
                kernel_img_mul_617[6] + kernel_img_mul_617[7] + kernel_img_mul_617[8] + 
                kernel_img_mul_617[9] + kernel_img_mul_617[10] + kernel_img_mul_617[11] + 
                kernel_img_mul_617[12] + kernel_img_mul_617[13] + kernel_img_mul_617[14] + 
                kernel_img_mul_617[15] + kernel_img_mul_617[16] + kernel_img_mul_617[17] + 
                kernel_img_mul_617[18] + kernel_img_mul_617[19] + kernel_img_mul_617[20] + 
                kernel_img_mul_617[21] + kernel_img_mul_617[22] + kernel_img_mul_617[23] + 
                kernel_img_mul_617[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4943:4936] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4943:4936] <= kernel_img_sum_617[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4943:4936] <= 'd0;
end

wire  [39:0]  kernel_img_mul_618[0:24];
assign kernel_img_mul_618[0] = buffer_data_4[4935:4928] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_618[1] = buffer_data_4[4943:4936] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_618[2] = buffer_data_4[4951:4944] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_618[3] = buffer_data_4[4959:4952] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_618[4] = buffer_data_4[4967:4960] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_618[5] = buffer_data_3[4935:4928] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_618[6] = buffer_data_3[4943:4936] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_618[7] = buffer_data_3[4951:4944] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_618[8] = buffer_data_3[4959:4952] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_618[9] = buffer_data_3[4967:4960] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_618[10] = buffer_data_2[4935:4928] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_618[11] = buffer_data_2[4943:4936] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_618[12] = buffer_data_2[4951:4944] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_618[13] = buffer_data_2[4959:4952] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_618[14] = buffer_data_2[4967:4960] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_618[15] = buffer_data_1[4935:4928] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_618[16] = buffer_data_1[4943:4936] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_618[17] = buffer_data_1[4951:4944] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_618[18] = buffer_data_1[4959:4952] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_618[19] = buffer_data_1[4967:4960] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_618[20] = buffer_data_0[4935:4928] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_618[21] = buffer_data_0[4943:4936] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_618[22] = buffer_data_0[4951:4944] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_618[23] = buffer_data_0[4959:4952] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_618[24] = buffer_data_0[4967:4960] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_618 = kernel_img_mul_618[0] + kernel_img_mul_618[1] + kernel_img_mul_618[2] + 
                kernel_img_mul_618[3] + kernel_img_mul_618[4] + kernel_img_mul_618[5] + 
                kernel_img_mul_618[6] + kernel_img_mul_618[7] + kernel_img_mul_618[8] + 
                kernel_img_mul_618[9] + kernel_img_mul_618[10] + kernel_img_mul_618[11] + 
                kernel_img_mul_618[12] + kernel_img_mul_618[13] + kernel_img_mul_618[14] + 
                kernel_img_mul_618[15] + kernel_img_mul_618[16] + kernel_img_mul_618[17] + 
                kernel_img_mul_618[18] + kernel_img_mul_618[19] + kernel_img_mul_618[20] + 
                kernel_img_mul_618[21] + kernel_img_mul_618[22] + kernel_img_mul_618[23] + 
                kernel_img_mul_618[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4951:4944] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4951:4944] <= kernel_img_sum_618[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4951:4944] <= 'd0;
end

wire  [39:0]  kernel_img_mul_619[0:24];
assign kernel_img_mul_619[0] = buffer_data_4[4943:4936] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_619[1] = buffer_data_4[4951:4944] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_619[2] = buffer_data_4[4959:4952] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_619[3] = buffer_data_4[4967:4960] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_619[4] = buffer_data_4[4975:4968] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_619[5] = buffer_data_3[4943:4936] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_619[6] = buffer_data_3[4951:4944] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_619[7] = buffer_data_3[4959:4952] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_619[8] = buffer_data_3[4967:4960] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_619[9] = buffer_data_3[4975:4968] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_619[10] = buffer_data_2[4943:4936] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_619[11] = buffer_data_2[4951:4944] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_619[12] = buffer_data_2[4959:4952] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_619[13] = buffer_data_2[4967:4960] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_619[14] = buffer_data_2[4975:4968] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_619[15] = buffer_data_1[4943:4936] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_619[16] = buffer_data_1[4951:4944] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_619[17] = buffer_data_1[4959:4952] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_619[18] = buffer_data_1[4967:4960] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_619[19] = buffer_data_1[4975:4968] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_619[20] = buffer_data_0[4943:4936] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_619[21] = buffer_data_0[4951:4944] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_619[22] = buffer_data_0[4959:4952] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_619[23] = buffer_data_0[4967:4960] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_619[24] = buffer_data_0[4975:4968] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_619 = kernel_img_mul_619[0] + kernel_img_mul_619[1] + kernel_img_mul_619[2] + 
                kernel_img_mul_619[3] + kernel_img_mul_619[4] + kernel_img_mul_619[5] + 
                kernel_img_mul_619[6] + kernel_img_mul_619[7] + kernel_img_mul_619[8] + 
                kernel_img_mul_619[9] + kernel_img_mul_619[10] + kernel_img_mul_619[11] + 
                kernel_img_mul_619[12] + kernel_img_mul_619[13] + kernel_img_mul_619[14] + 
                kernel_img_mul_619[15] + kernel_img_mul_619[16] + kernel_img_mul_619[17] + 
                kernel_img_mul_619[18] + kernel_img_mul_619[19] + kernel_img_mul_619[20] + 
                kernel_img_mul_619[21] + kernel_img_mul_619[22] + kernel_img_mul_619[23] + 
                kernel_img_mul_619[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4959:4952] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4959:4952] <= kernel_img_sum_619[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4959:4952] <= 'd0;
end

wire  [39:0]  kernel_img_mul_620[0:24];
assign kernel_img_mul_620[0] = buffer_data_4[4951:4944] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_620[1] = buffer_data_4[4959:4952] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_620[2] = buffer_data_4[4967:4960] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_620[3] = buffer_data_4[4975:4968] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_620[4] = buffer_data_4[4983:4976] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_620[5] = buffer_data_3[4951:4944] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_620[6] = buffer_data_3[4959:4952] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_620[7] = buffer_data_3[4967:4960] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_620[8] = buffer_data_3[4975:4968] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_620[9] = buffer_data_3[4983:4976] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_620[10] = buffer_data_2[4951:4944] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_620[11] = buffer_data_2[4959:4952] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_620[12] = buffer_data_2[4967:4960] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_620[13] = buffer_data_2[4975:4968] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_620[14] = buffer_data_2[4983:4976] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_620[15] = buffer_data_1[4951:4944] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_620[16] = buffer_data_1[4959:4952] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_620[17] = buffer_data_1[4967:4960] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_620[18] = buffer_data_1[4975:4968] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_620[19] = buffer_data_1[4983:4976] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_620[20] = buffer_data_0[4951:4944] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_620[21] = buffer_data_0[4959:4952] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_620[22] = buffer_data_0[4967:4960] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_620[23] = buffer_data_0[4975:4968] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_620[24] = buffer_data_0[4983:4976] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_620 = kernel_img_mul_620[0] + kernel_img_mul_620[1] + kernel_img_mul_620[2] + 
                kernel_img_mul_620[3] + kernel_img_mul_620[4] + kernel_img_mul_620[5] + 
                kernel_img_mul_620[6] + kernel_img_mul_620[7] + kernel_img_mul_620[8] + 
                kernel_img_mul_620[9] + kernel_img_mul_620[10] + kernel_img_mul_620[11] + 
                kernel_img_mul_620[12] + kernel_img_mul_620[13] + kernel_img_mul_620[14] + 
                kernel_img_mul_620[15] + kernel_img_mul_620[16] + kernel_img_mul_620[17] + 
                kernel_img_mul_620[18] + kernel_img_mul_620[19] + kernel_img_mul_620[20] + 
                kernel_img_mul_620[21] + kernel_img_mul_620[22] + kernel_img_mul_620[23] + 
                kernel_img_mul_620[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4967:4960] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4967:4960] <= kernel_img_sum_620[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4967:4960] <= 'd0;
end

wire  [39:0]  kernel_img_mul_621[0:24];
assign kernel_img_mul_621[0] = buffer_data_4[4959:4952] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_621[1] = buffer_data_4[4967:4960] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_621[2] = buffer_data_4[4975:4968] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_621[3] = buffer_data_4[4983:4976] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_621[4] = buffer_data_4[4991:4984] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_621[5] = buffer_data_3[4959:4952] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_621[6] = buffer_data_3[4967:4960] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_621[7] = buffer_data_3[4975:4968] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_621[8] = buffer_data_3[4983:4976] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_621[9] = buffer_data_3[4991:4984] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_621[10] = buffer_data_2[4959:4952] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_621[11] = buffer_data_2[4967:4960] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_621[12] = buffer_data_2[4975:4968] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_621[13] = buffer_data_2[4983:4976] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_621[14] = buffer_data_2[4991:4984] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_621[15] = buffer_data_1[4959:4952] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_621[16] = buffer_data_1[4967:4960] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_621[17] = buffer_data_1[4975:4968] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_621[18] = buffer_data_1[4983:4976] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_621[19] = buffer_data_1[4991:4984] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_621[20] = buffer_data_0[4959:4952] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_621[21] = buffer_data_0[4967:4960] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_621[22] = buffer_data_0[4975:4968] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_621[23] = buffer_data_0[4983:4976] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_621[24] = buffer_data_0[4991:4984] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_621 = kernel_img_mul_621[0] + kernel_img_mul_621[1] + kernel_img_mul_621[2] + 
                kernel_img_mul_621[3] + kernel_img_mul_621[4] + kernel_img_mul_621[5] + 
                kernel_img_mul_621[6] + kernel_img_mul_621[7] + kernel_img_mul_621[8] + 
                kernel_img_mul_621[9] + kernel_img_mul_621[10] + kernel_img_mul_621[11] + 
                kernel_img_mul_621[12] + kernel_img_mul_621[13] + kernel_img_mul_621[14] + 
                kernel_img_mul_621[15] + kernel_img_mul_621[16] + kernel_img_mul_621[17] + 
                kernel_img_mul_621[18] + kernel_img_mul_621[19] + kernel_img_mul_621[20] + 
                kernel_img_mul_621[21] + kernel_img_mul_621[22] + kernel_img_mul_621[23] + 
                kernel_img_mul_621[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4975:4968] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4975:4968] <= kernel_img_sum_621[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4975:4968] <= 'd0;
end

wire  [39:0]  kernel_img_mul_622[0:24];
assign kernel_img_mul_622[0] = buffer_data_4[4967:4960] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_622[1] = buffer_data_4[4975:4968] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_622[2] = buffer_data_4[4983:4976] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_622[3] = buffer_data_4[4991:4984] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_622[4] = buffer_data_4[4999:4992] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_622[5] = buffer_data_3[4967:4960] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_622[6] = buffer_data_3[4975:4968] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_622[7] = buffer_data_3[4983:4976] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_622[8] = buffer_data_3[4991:4984] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_622[9] = buffer_data_3[4999:4992] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_622[10] = buffer_data_2[4967:4960] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_622[11] = buffer_data_2[4975:4968] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_622[12] = buffer_data_2[4983:4976] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_622[13] = buffer_data_2[4991:4984] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_622[14] = buffer_data_2[4999:4992] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_622[15] = buffer_data_1[4967:4960] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_622[16] = buffer_data_1[4975:4968] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_622[17] = buffer_data_1[4983:4976] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_622[18] = buffer_data_1[4991:4984] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_622[19] = buffer_data_1[4999:4992] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_622[20] = buffer_data_0[4967:4960] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_622[21] = buffer_data_0[4975:4968] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_622[22] = buffer_data_0[4983:4976] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_622[23] = buffer_data_0[4991:4984] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_622[24] = buffer_data_0[4999:4992] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_622 = kernel_img_mul_622[0] + kernel_img_mul_622[1] + kernel_img_mul_622[2] + 
                kernel_img_mul_622[3] + kernel_img_mul_622[4] + kernel_img_mul_622[5] + 
                kernel_img_mul_622[6] + kernel_img_mul_622[7] + kernel_img_mul_622[8] + 
                kernel_img_mul_622[9] + kernel_img_mul_622[10] + kernel_img_mul_622[11] + 
                kernel_img_mul_622[12] + kernel_img_mul_622[13] + kernel_img_mul_622[14] + 
                kernel_img_mul_622[15] + kernel_img_mul_622[16] + kernel_img_mul_622[17] + 
                kernel_img_mul_622[18] + kernel_img_mul_622[19] + kernel_img_mul_622[20] + 
                kernel_img_mul_622[21] + kernel_img_mul_622[22] + kernel_img_mul_622[23] + 
                kernel_img_mul_622[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4983:4976] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4983:4976] <= kernel_img_sum_622[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4983:4976] <= 'd0;
end

wire  [39:0]  kernel_img_mul_623[0:24];
assign kernel_img_mul_623[0] = buffer_data_4[4975:4968] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_623[1] = buffer_data_4[4983:4976] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_623[2] = buffer_data_4[4991:4984] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_623[3] = buffer_data_4[4999:4992] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_623[4] = buffer_data_4[5007:5000] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_623[5] = buffer_data_3[4975:4968] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_623[6] = buffer_data_3[4983:4976] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_623[7] = buffer_data_3[4991:4984] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_623[8] = buffer_data_3[4999:4992] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_623[9] = buffer_data_3[5007:5000] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_623[10] = buffer_data_2[4975:4968] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_623[11] = buffer_data_2[4983:4976] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_623[12] = buffer_data_2[4991:4984] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_623[13] = buffer_data_2[4999:4992] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_623[14] = buffer_data_2[5007:5000] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_623[15] = buffer_data_1[4975:4968] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_623[16] = buffer_data_1[4983:4976] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_623[17] = buffer_data_1[4991:4984] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_623[18] = buffer_data_1[4999:4992] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_623[19] = buffer_data_1[5007:5000] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_623[20] = buffer_data_0[4975:4968] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_623[21] = buffer_data_0[4983:4976] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_623[22] = buffer_data_0[4991:4984] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_623[23] = buffer_data_0[4999:4992] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_623[24] = buffer_data_0[5007:5000] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_623 = kernel_img_mul_623[0] + kernel_img_mul_623[1] + kernel_img_mul_623[2] + 
                kernel_img_mul_623[3] + kernel_img_mul_623[4] + kernel_img_mul_623[5] + 
                kernel_img_mul_623[6] + kernel_img_mul_623[7] + kernel_img_mul_623[8] + 
                kernel_img_mul_623[9] + kernel_img_mul_623[10] + kernel_img_mul_623[11] + 
                kernel_img_mul_623[12] + kernel_img_mul_623[13] + kernel_img_mul_623[14] + 
                kernel_img_mul_623[15] + kernel_img_mul_623[16] + kernel_img_mul_623[17] + 
                kernel_img_mul_623[18] + kernel_img_mul_623[19] + kernel_img_mul_623[20] + 
                kernel_img_mul_623[21] + kernel_img_mul_623[22] + kernel_img_mul_623[23] + 
                kernel_img_mul_623[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4991:4984] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4991:4984] <= kernel_img_sum_623[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4991:4984] <= 'd0;
end

wire  [39:0]  kernel_img_mul_624[0:24];
assign kernel_img_mul_624[0] = buffer_data_4[4983:4976] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_624[1] = buffer_data_4[4991:4984] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_624[2] = buffer_data_4[4999:4992] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_624[3] = buffer_data_4[5007:5000] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_624[4] = buffer_data_4[5015:5008] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_624[5] = buffer_data_3[4983:4976] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_624[6] = buffer_data_3[4991:4984] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_624[7] = buffer_data_3[4999:4992] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_624[8] = buffer_data_3[5007:5000] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_624[9] = buffer_data_3[5015:5008] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_624[10] = buffer_data_2[4983:4976] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_624[11] = buffer_data_2[4991:4984] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_624[12] = buffer_data_2[4999:4992] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_624[13] = buffer_data_2[5007:5000] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_624[14] = buffer_data_2[5015:5008] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_624[15] = buffer_data_1[4983:4976] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_624[16] = buffer_data_1[4991:4984] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_624[17] = buffer_data_1[4999:4992] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_624[18] = buffer_data_1[5007:5000] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_624[19] = buffer_data_1[5015:5008] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_624[20] = buffer_data_0[4983:4976] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_624[21] = buffer_data_0[4991:4984] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_624[22] = buffer_data_0[4999:4992] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_624[23] = buffer_data_0[5007:5000] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_624[24] = buffer_data_0[5015:5008] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_624 = kernel_img_mul_624[0] + kernel_img_mul_624[1] + kernel_img_mul_624[2] + 
                kernel_img_mul_624[3] + kernel_img_mul_624[4] + kernel_img_mul_624[5] + 
                kernel_img_mul_624[6] + kernel_img_mul_624[7] + kernel_img_mul_624[8] + 
                kernel_img_mul_624[9] + kernel_img_mul_624[10] + kernel_img_mul_624[11] + 
                kernel_img_mul_624[12] + kernel_img_mul_624[13] + kernel_img_mul_624[14] + 
                kernel_img_mul_624[15] + kernel_img_mul_624[16] + kernel_img_mul_624[17] + 
                kernel_img_mul_624[18] + kernel_img_mul_624[19] + kernel_img_mul_624[20] + 
                kernel_img_mul_624[21] + kernel_img_mul_624[22] + kernel_img_mul_624[23] + 
                kernel_img_mul_624[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[4999:4992] <= 'd0;
  else if (current_state==ST_START)
    blur_din[4999:4992] <= kernel_img_sum_624[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4999:4992] <= 'd0;
end

wire  [39:0]  kernel_img_mul_625[0:24];
assign kernel_img_mul_625[0] = buffer_data_4[4991:4984] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_625[1] = buffer_data_4[4999:4992] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_625[2] = buffer_data_4[5007:5000] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_625[3] = buffer_data_4[5015:5008] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_625[4] = buffer_data_4[5023:5016] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_625[5] = buffer_data_3[4991:4984] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_625[6] = buffer_data_3[4999:4992] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_625[7] = buffer_data_3[5007:5000] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_625[8] = buffer_data_3[5015:5008] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_625[9] = buffer_data_3[5023:5016] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_625[10] = buffer_data_2[4991:4984] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_625[11] = buffer_data_2[4999:4992] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_625[12] = buffer_data_2[5007:5000] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_625[13] = buffer_data_2[5015:5008] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_625[14] = buffer_data_2[5023:5016] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_625[15] = buffer_data_1[4991:4984] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_625[16] = buffer_data_1[4999:4992] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_625[17] = buffer_data_1[5007:5000] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_625[18] = buffer_data_1[5015:5008] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_625[19] = buffer_data_1[5023:5016] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_625[20] = buffer_data_0[4991:4984] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_625[21] = buffer_data_0[4999:4992] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_625[22] = buffer_data_0[5007:5000] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_625[23] = buffer_data_0[5015:5008] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_625[24] = buffer_data_0[5023:5016] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_625 = kernel_img_mul_625[0] + kernel_img_mul_625[1] + kernel_img_mul_625[2] + 
                kernel_img_mul_625[3] + kernel_img_mul_625[4] + kernel_img_mul_625[5] + 
                kernel_img_mul_625[6] + kernel_img_mul_625[7] + kernel_img_mul_625[8] + 
                kernel_img_mul_625[9] + kernel_img_mul_625[10] + kernel_img_mul_625[11] + 
                kernel_img_mul_625[12] + kernel_img_mul_625[13] + kernel_img_mul_625[14] + 
                kernel_img_mul_625[15] + kernel_img_mul_625[16] + kernel_img_mul_625[17] + 
                kernel_img_mul_625[18] + kernel_img_mul_625[19] + kernel_img_mul_625[20] + 
                kernel_img_mul_625[21] + kernel_img_mul_625[22] + kernel_img_mul_625[23] + 
                kernel_img_mul_625[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[5007:5000] <= 'd0;
  else if (current_state==ST_START)
    blur_din[5007:5000] <= kernel_img_sum_625[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5007:5000] <= 'd0;
end

wire  [39:0]  kernel_img_mul_626[0:24];
assign kernel_img_mul_626[0] = buffer_data_4[4999:4992] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_626[1] = buffer_data_4[5007:5000] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_626[2] = buffer_data_4[5015:5008] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_626[3] = buffer_data_4[5023:5016] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_626[4] = buffer_data_4[5031:5024] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_626[5] = buffer_data_3[4999:4992] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_626[6] = buffer_data_3[5007:5000] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_626[7] = buffer_data_3[5015:5008] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_626[8] = buffer_data_3[5023:5016] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_626[9] = buffer_data_3[5031:5024] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_626[10] = buffer_data_2[4999:4992] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_626[11] = buffer_data_2[5007:5000] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_626[12] = buffer_data_2[5015:5008] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_626[13] = buffer_data_2[5023:5016] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_626[14] = buffer_data_2[5031:5024] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_626[15] = buffer_data_1[4999:4992] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_626[16] = buffer_data_1[5007:5000] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_626[17] = buffer_data_1[5015:5008] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_626[18] = buffer_data_1[5023:5016] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_626[19] = buffer_data_1[5031:5024] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_626[20] = buffer_data_0[4999:4992] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_626[21] = buffer_data_0[5007:5000] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_626[22] = buffer_data_0[5015:5008] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_626[23] = buffer_data_0[5023:5016] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_626[24] = buffer_data_0[5031:5024] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_626 = kernel_img_mul_626[0] + kernel_img_mul_626[1] + kernel_img_mul_626[2] + 
                kernel_img_mul_626[3] + kernel_img_mul_626[4] + kernel_img_mul_626[5] + 
                kernel_img_mul_626[6] + kernel_img_mul_626[7] + kernel_img_mul_626[8] + 
                kernel_img_mul_626[9] + kernel_img_mul_626[10] + kernel_img_mul_626[11] + 
                kernel_img_mul_626[12] + kernel_img_mul_626[13] + kernel_img_mul_626[14] + 
                kernel_img_mul_626[15] + kernel_img_mul_626[16] + kernel_img_mul_626[17] + 
                kernel_img_mul_626[18] + kernel_img_mul_626[19] + kernel_img_mul_626[20] + 
                kernel_img_mul_626[21] + kernel_img_mul_626[22] + kernel_img_mul_626[23] + 
                kernel_img_mul_626[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[5015:5008] <= 'd0;
  else if (current_state==ST_START)
    blur_din[5015:5008] <= kernel_img_sum_626[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5015:5008] <= 'd0;
end

wire  [39:0]  kernel_img_mul_627[0:24];
assign kernel_img_mul_627[0] = buffer_data_4[5007:5000] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_627[1] = buffer_data_4[5015:5008] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_627[2] = buffer_data_4[5023:5016] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_627[3] = buffer_data_4[5031:5024] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_627[4] = buffer_data_4[5039:5032] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_627[5] = buffer_data_3[5007:5000] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_627[6] = buffer_data_3[5015:5008] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_627[7] = buffer_data_3[5023:5016] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_627[8] = buffer_data_3[5031:5024] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_627[9] = buffer_data_3[5039:5032] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_627[10] = buffer_data_2[5007:5000] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_627[11] = buffer_data_2[5015:5008] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_627[12] = buffer_data_2[5023:5016] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_627[13] = buffer_data_2[5031:5024] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_627[14] = buffer_data_2[5039:5032] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_627[15] = buffer_data_1[5007:5000] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_627[16] = buffer_data_1[5015:5008] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_627[17] = buffer_data_1[5023:5016] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_627[18] = buffer_data_1[5031:5024] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_627[19] = buffer_data_1[5039:5032] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_627[20] = buffer_data_0[5007:5000] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_627[21] = buffer_data_0[5015:5008] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_627[22] = buffer_data_0[5023:5016] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_627[23] = buffer_data_0[5031:5024] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_627[24] = buffer_data_0[5039:5032] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_627 = kernel_img_mul_627[0] + kernel_img_mul_627[1] + kernel_img_mul_627[2] + 
                kernel_img_mul_627[3] + kernel_img_mul_627[4] + kernel_img_mul_627[5] + 
                kernel_img_mul_627[6] + kernel_img_mul_627[7] + kernel_img_mul_627[8] + 
                kernel_img_mul_627[9] + kernel_img_mul_627[10] + kernel_img_mul_627[11] + 
                kernel_img_mul_627[12] + kernel_img_mul_627[13] + kernel_img_mul_627[14] + 
                kernel_img_mul_627[15] + kernel_img_mul_627[16] + kernel_img_mul_627[17] + 
                kernel_img_mul_627[18] + kernel_img_mul_627[19] + kernel_img_mul_627[20] + 
                kernel_img_mul_627[21] + kernel_img_mul_627[22] + kernel_img_mul_627[23] + 
                kernel_img_mul_627[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[5023:5016] <= 'd0;
  else if (current_state==ST_START)
    blur_din[5023:5016] <= kernel_img_sum_627[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5023:5016] <= 'd0;
end

wire  [39:0]  kernel_img_mul_628[0:24];
assign kernel_img_mul_628[0] = buffer_data_4[5015:5008] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_628[1] = buffer_data_4[5023:5016] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_628[2] = buffer_data_4[5031:5024] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_628[3] = buffer_data_4[5039:5032] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_628[4] = buffer_data_4[5047:5040] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_628[5] = buffer_data_3[5015:5008] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_628[6] = buffer_data_3[5023:5016] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_628[7] = buffer_data_3[5031:5024] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_628[8] = buffer_data_3[5039:5032] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_628[9] = buffer_data_3[5047:5040] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_628[10] = buffer_data_2[5015:5008] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_628[11] = buffer_data_2[5023:5016] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_628[12] = buffer_data_2[5031:5024] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_628[13] = buffer_data_2[5039:5032] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_628[14] = buffer_data_2[5047:5040] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_628[15] = buffer_data_1[5015:5008] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_628[16] = buffer_data_1[5023:5016] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_628[17] = buffer_data_1[5031:5024] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_628[18] = buffer_data_1[5039:5032] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_628[19] = buffer_data_1[5047:5040] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_628[20] = buffer_data_0[5015:5008] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_628[21] = buffer_data_0[5023:5016] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_628[22] = buffer_data_0[5031:5024] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_628[23] = buffer_data_0[5039:5032] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_628[24] = buffer_data_0[5047:5040] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_628 = kernel_img_mul_628[0] + kernel_img_mul_628[1] + kernel_img_mul_628[2] + 
                kernel_img_mul_628[3] + kernel_img_mul_628[4] + kernel_img_mul_628[5] + 
                kernel_img_mul_628[6] + kernel_img_mul_628[7] + kernel_img_mul_628[8] + 
                kernel_img_mul_628[9] + kernel_img_mul_628[10] + kernel_img_mul_628[11] + 
                kernel_img_mul_628[12] + kernel_img_mul_628[13] + kernel_img_mul_628[14] + 
                kernel_img_mul_628[15] + kernel_img_mul_628[16] + kernel_img_mul_628[17] + 
                kernel_img_mul_628[18] + kernel_img_mul_628[19] + kernel_img_mul_628[20] + 
                kernel_img_mul_628[21] + kernel_img_mul_628[22] + kernel_img_mul_628[23] + 
                kernel_img_mul_628[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[5031:5024] <= 'd0;
  else if (current_state==ST_START)
    blur_din[5031:5024] <= kernel_img_sum_628[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5031:5024] <= 'd0;
end

wire  [39:0]  kernel_img_mul_629[0:24];
assign kernel_img_mul_629[0] = buffer_data_4[5023:5016] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_629[1] = buffer_data_4[5031:5024] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_629[2] = buffer_data_4[5039:5032] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_629[3] = buffer_data_4[5047:5040] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_629[4] = buffer_data_4[5055:5048] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_629[5] = buffer_data_3[5023:5016] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_629[6] = buffer_data_3[5031:5024] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_629[7] = buffer_data_3[5039:5032] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_629[8] = buffer_data_3[5047:5040] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_629[9] = buffer_data_3[5055:5048] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_629[10] = buffer_data_2[5023:5016] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_629[11] = buffer_data_2[5031:5024] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_629[12] = buffer_data_2[5039:5032] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_629[13] = buffer_data_2[5047:5040] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_629[14] = buffer_data_2[5055:5048] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_629[15] = buffer_data_1[5023:5016] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_629[16] = buffer_data_1[5031:5024] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_629[17] = buffer_data_1[5039:5032] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_629[18] = buffer_data_1[5047:5040] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_629[19] = buffer_data_1[5055:5048] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_629[20] = buffer_data_0[5023:5016] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_629[21] = buffer_data_0[5031:5024] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_629[22] = buffer_data_0[5039:5032] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_629[23] = buffer_data_0[5047:5040] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_629[24] = buffer_data_0[5055:5048] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_629 = kernel_img_mul_629[0] + kernel_img_mul_629[1] + kernel_img_mul_629[2] + 
                kernel_img_mul_629[3] + kernel_img_mul_629[4] + kernel_img_mul_629[5] + 
                kernel_img_mul_629[6] + kernel_img_mul_629[7] + kernel_img_mul_629[8] + 
                kernel_img_mul_629[9] + kernel_img_mul_629[10] + kernel_img_mul_629[11] + 
                kernel_img_mul_629[12] + kernel_img_mul_629[13] + kernel_img_mul_629[14] + 
                kernel_img_mul_629[15] + kernel_img_mul_629[16] + kernel_img_mul_629[17] + 
                kernel_img_mul_629[18] + kernel_img_mul_629[19] + kernel_img_mul_629[20] + 
                kernel_img_mul_629[21] + kernel_img_mul_629[22] + kernel_img_mul_629[23] + 
                kernel_img_mul_629[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[5039:5032] <= 'd0;
  else if (current_state==ST_START)
    blur_din[5039:5032] <= kernel_img_sum_629[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5039:5032] <= 'd0;
end

wire  [39:0]  kernel_img_mul_630[0:24];
assign kernel_img_mul_630[0] = buffer_data_4[5031:5024] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_630[1] = buffer_data_4[5039:5032] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_630[2] = buffer_data_4[5047:5040] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_630[3] = buffer_data_4[5055:5048] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_630[4] = buffer_data_4[5063:5056] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_630[5] = buffer_data_3[5031:5024] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_630[6] = buffer_data_3[5039:5032] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_630[7] = buffer_data_3[5047:5040] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_630[8] = buffer_data_3[5055:5048] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_630[9] = buffer_data_3[5063:5056] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_630[10] = buffer_data_2[5031:5024] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_630[11] = buffer_data_2[5039:5032] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_630[12] = buffer_data_2[5047:5040] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_630[13] = buffer_data_2[5055:5048] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_630[14] = buffer_data_2[5063:5056] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_630[15] = buffer_data_1[5031:5024] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_630[16] = buffer_data_1[5039:5032] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_630[17] = buffer_data_1[5047:5040] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_630[18] = buffer_data_1[5055:5048] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_630[19] = buffer_data_1[5063:5056] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_630[20] = buffer_data_0[5031:5024] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_630[21] = buffer_data_0[5039:5032] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_630[22] = buffer_data_0[5047:5040] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_630[23] = buffer_data_0[5055:5048] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_630[24] = buffer_data_0[5063:5056] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_630 = kernel_img_mul_630[0] + kernel_img_mul_630[1] + kernel_img_mul_630[2] + 
                kernel_img_mul_630[3] + kernel_img_mul_630[4] + kernel_img_mul_630[5] + 
                kernel_img_mul_630[6] + kernel_img_mul_630[7] + kernel_img_mul_630[8] + 
                kernel_img_mul_630[9] + kernel_img_mul_630[10] + kernel_img_mul_630[11] + 
                kernel_img_mul_630[12] + kernel_img_mul_630[13] + kernel_img_mul_630[14] + 
                kernel_img_mul_630[15] + kernel_img_mul_630[16] + kernel_img_mul_630[17] + 
                kernel_img_mul_630[18] + kernel_img_mul_630[19] + kernel_img_mul_630[20] + 
                kernel_img_mul_630[21] + kernel_img_mul_630[22] + kernel_img_mul_630[23] + 
                kernel_img_mul_630[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[5047:5040] <= 'd0;
  else if (current_state==ST_START)
    blur_din[5047:5040] <= kernel_img_sum_630[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5047:5040] <= 'd0;
end

wire  [39:0]  kernel_img_mul_631[0:24];
assign kernel_img_mul_631[0] = buffer_data_4[5039:5032] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_631[1] = buffer_data_4[5047:5040] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_631[2] = buffer_data_4[5055:5048] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_631[3] = buffer_data_4[5063:5056] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_631[4] = buffer_data_4[5071:5064] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_631[5] = buffer_data_3[5039:5032] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_631[6] = buffer_data_3[5047:5040] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_631[7] = buffer_data_3[5055:5048] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_631[8] = buffer_data_3[5063:5056] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_631[9] = buffer_data_3[5071:5064] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_631[10] = buffer_data_2[5039:5032] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_631[11] = buffer_data_2[5047:5040] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_631[12] = buffer_data_2[5055:5048] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_631[13] = buffer_data_2[5063:5056] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_631[14] = buffer_data_2[5071:5064] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_631[15] = buffer_data_1[5039:5032] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_631[16] = buffer_data_1[5047:5040] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_631[17] = buffer_data_1[5055:5048] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_631[18] = buffer_data_1[5063:5056] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_631[19] = buffer_data_1[5071:5064] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_631[20] = buffer_data_0[5039:5032] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_631[21] = buffer_data_0[5047:5040] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_631[22] = buffer_data_0[5055:5048] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_631[23] = buffer_data_0[5063:5056] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_631[24] = buffer_data_0[5071:5064] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_631 = kernel_img_mul_631[0] + kernel_img_mul_631[1] + kernel_img_mul_631[2] + 
                kernel_img_mul_631[3] + kernel_img_mul_631[4] + kernel_img_mul_631[5] + 
                kernel_img_mul_631[6] + kernel_img_mul_631[7] + kernel_img_mul_631[8] + 
                kernel_img_mul_631[9] + kernel_img_mul_631[10] + kernel_img_mul_631[11] + 
                kernel_img_mul_631[12] + kernel_img_mul_631[13] + kernel_img_mul_631[14] + 
                kernel_img_mul_631[15] + kernel_img_mul_631[16] + kernel_img_mul_631[17] + 
                kernel_img_mul_631[18] + kernel_img_mul_631[19] + kernel_img_mul_631[20] + 
                kernel_img_mul_631[21] + kernel_img_mul_631[22] + kernel_img_mul_631[23] + 
                kernel_img_mul_631[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[5055:5048] <= 'd0;
  else if (current_state==ST_START)
    blur_din[5055:5048] <= kernel_img_sum_631[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5055:5048] <= 'd0;
end

wire  [39:0]  kernel_img_mul_632[0:24];
assign kernel_img_mul_632[0] = buffer_data_4[5047:5040] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_632[1] = buffer_data_4[5055:5048] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_632[2] = buffer_data_4[5063:5056] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_632[3] = buffer_data_4[5071:5064] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_632[4] = buffer_data_4[5079:5072] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_632[5] = buffer_data_3[5047:5040] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_632[6] = buffer_data_3[5055:5048] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_632[7] = buffer_data_3[5063:5056] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_632[8] = buffer_data_3[5071:5064] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_632[9] = buffer_data_3[5079:5072] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_632[10] = buffer_data_2[5047:5040] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_632[11] = buffer_data_2[5055:5048] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_632[12] = buffer_data_2[5063:5056] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_632[13] = buffer_data_2[5071:5064] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_632[14] = buffer_data_2[5079:5072] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_632[15] = buffer_data_1[5047:5040] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_632[16] = buffer_data_1[5055:5048] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_632[17] = buffer_data_1[5063:5056] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_632[18] = buffer_data_1[5071:5064] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_632[19] = buffer_data_1[5079:5072] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_632[20] = buffer_data_0[5047:5040] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_632[21] = buffer_data_0[5055:5048] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_632[22] = buffer_data_0[5063:5056] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_632[23] = buffer_data_0[5071:5064] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_632[24] = buffer_data_0[5079:5072] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_632 = kernel_img_mul_632[0] + kernel_img_mul_632[1] + kernel_img_mul_632[2] + 
                kernel_img_mul_632[3] + kernel_img_mul_632[4] + kernel_img_mul_632[5] + 
                kernel_img_mul_632[6] + kernel_img_mul_632[7] + kernel_img_mul_632[8] + 
                kernel_img_mul_632[9] + kernel_img_mul_632[10] + kernel_img_mul_632[11] + 
                kernel_img_mul_632[12] + kernel_img_mul_632[13] + kernel_img_mul_632[14] + 
                kernel_img_mul_632[15] + kernel_img_mul_632[16] + kernel_img_mul_632[17] + 
                kernel_img_mul_632[18] + kernel_img_mul_632[19] + kernel_img_mul_632[20] + 
                kernel_img_mul_632[21] + kernel_img_mul_632[22] + kernel_img_mul_632[23] + 
                kernel_img_mul_632[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[5063:5056] <= 'd0;
  else if (current_state==ST_START)
    blur_din[5063:5056] <= kernel_img_sum_632[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5063:5056] <= 'd0;
end

wire  [39:0]  kernel_img_mul_633[0:24];
assign kernel_img_mul_633[0] = buffer_data_4[5055:5048] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_633[1] = buffer_data_4[5063:5056] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_633[2] = buffer_data_4[5071:5064] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_633[3] = buffer_data_4[5079:5072] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_633[4] = buffer_data_4[5087:5080] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_633[5] = buffer_data_3[5055:5048] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_633[6] = buffer_data_3[5063:5056] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_633[7] = buffer_data_3[5071:5064] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_633[8] = buffer_data_3[5079:5072] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_633[9] = buffer_data_3[5087:5080] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_633[10] = buffer_data_2[5055:5048] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_633[11] = buffer_data_2[5063:5056] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_633[12] = buffer_data_2[5071:5064] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_633[13] = buffer_data_2[5079:5072] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_633[14] = buffer_data_2[5087:5080] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_633[15] = buffer_data_1[5055:5048] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_633[16] = buffer_data_1[5063:5056] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_633[17] = buffer_data_1[5071:5064] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_633[18] = buffer_data_1[5079:5072] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_633[19] = buffer_data_1[5087:5080] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_633[20] = buffer_data_0[5055:5048] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_633[21] = buffer_data_0[5063:5056] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_633[22] = buffer_data_0[5071:5064] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_633[23] = buffer_data_0[5079:5072] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_633[24] = buffer_data_0[5087:5080] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_633 = kernel_img_mul_633[0] + kernel_img_mul_633[1] + kernel_img_mul_633[2] + 
                kernel_img_mul_633[3] + kernel_img_mul_633[4] + kernel_img_mul_633[5] + 
                kernel_img_mul_633[6] + kernel_img_mul_633[7] + kernel_img_mul_633[8] + 
                kernel_img_mul_633[9] + kernel_img_mul_633[10] + kernel_img_mul_633[11] + 
                kernel_img_mul_633[12] + kernel_img_mul_633[13] + kernel_img_mul_633[14] + 
                kernel_img_mul_633[15] + kernel_img_mul_633[16] + kernel_img_mul_633[17] + 
                kernel_img_mul_633[18] + kernel_img_mul_633[19] + kernel_img_mul_633[20] + 
                kernel_img_mul_633[21] + kernel_img_mul_633[22] + kernel_img_mul_633[23] + 
                kernel_img_mul_633[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[5071:5064] <= 'd0;
  else if (current_state==ST_START)
    blur_din[5071:5064] <= kernel_img_sum_633[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5071:5064] <= 'd0;
end

wire  [39:0]  kernel_img_mul_634[0:24];
assign kernel_img_mul_634[0] = buffer_data_4[5063:5056] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_634[1] = buffer_data_4[5071:5064] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_634[2] = buffer_data_4[5079:5072] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_634[3] = buffer_data_4[5087:5080] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_634[4] = buffer_data_4[5095:5088] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_634[5] = buffer_data_3[5063:5056] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_634[6] = buffer_data_3[5071:5064] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_634[7] = buffer_data_3[5079:5072] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_634[8] = buffer_data_3[5087:5080] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_634[9] = buffer_data_3[5095:5088] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_634[10] = buffer_data_2[5063:5056] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_634[11] = buffer_data_2[5071:5064] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_634[12] = buffer_data_2[5079:5072] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_634[13] = buffer_data_2[5087:5080] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_634[14] = buffer_data_2[5095:5088] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_634[15] = buffer_data_1[5063:5056] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_634[16] = buffer_data_1[5071:5064] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_634[17] = buffer_data_1[5079:5072] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_634[18] = buffer_data_1[5087:5080] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_634[19] = buffer_data_1[5095:5088] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_634[20] = buffer_data_0[5063:5056] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_634[21] = buffer_data_0[5071:5064] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_634[22] = buffer_data_0[5079:5072] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_634[23] = buffer_data_0[5087:5080] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_634[24] = buffer_data_0[5095:5088] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_634 = kernel_img_mul_634[0] + kernel_img_mul_634[1] + kernel_img_mul_634[2] + 
                kernel_img_mul_634[3] + kernel_img_mul_634[4] + kernel_img_mul_634[5] + 
                kernel_img_mul_634[6] + kernel_img_mul_634[7] + kernel_img_mul_634[8] + 
                kernel_img_mul_634[9] + kernel_img_mul_634[10] + kernel_img_mul_634[11] + 
                kernel_img_mul_634[12] + kernel_img_mul_634[13] + kernel_img_mul_634[14] + 
                kernel_img_mul_634[15] + kernel_img_mul_634[16] + kernel_img_mul_634[17] + 
                kernel_img_mul_634[18] + kernel_img_mul_634[19] + kernel_img_mul_634[20] + 
                kernel_img_mul_634[21] + kernel_img_mul_634[22] + kernel_img_mul_634[23] + 
                kernel_img_mul_634[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[5079:5072] <= 'd0;
  else if (current_state==ST_START)
    blur_din[5079:5072] <= kernel_img_sum_634[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5079:5072] <= 'd0;
end

wire  [39:0]  kernel_img_mul_635[0:24];
assign kernel_img_mul_635[0] = buffer_data_4[5071:5064] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_635[1] = buffer_data_4[5079:5072] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_635[2] = buffer_data_4[5087:5080] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_635[3] = buffer_data_4[5095:5088] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_635[4] = buffer_data_4[5103:5096] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_635[5] = buffer_data_3[5071:5064] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_635[6] = buffer_data_3[5079:5072] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_635[7] = buffer_data_3[5087:5080] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_635[8] = buffer_data_3[5095:5088] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_635[9] = buffer_data_3[5103:5096] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_635[10] = buffer_data_2[5071:5064] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_635[11] = buffer_data_2[5079:5072] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_635[12] = buffer_data_2[5087:5080] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_635[13] = buffer_data_2[5095:5088] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_635[14] = buffer_data_2[5103:5096] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_635[15] = buffer_data_1[5071:5064] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_635[16] = buffer_data_1[5079:5072] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_635[17] = buffer_data_1[5087:5080] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_635[18] = buffer_data_1[5095:5088] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_635[19] = buffer_data_1[5103:5096] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_635[20] = buffer_data_0[5071:5064] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_635[21] = buffer_data_0[5079:5072] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_635[22] = buffer_data_0[5087:5080] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_635[23] = buffer_data_0[5095:5088] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_635[24] = buffer_data_0[5103:5096] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_635 = kernel_img_mul_635[0] + kernel_img_mul_635[1] + kernel_img_mul_635[2] + 
                kernel_img_mul_635[3] + kernel_img_mul_635[4] + kernel_img_mul_635[5] + 
                kernel_img_mul_635[6] + kernel_img_mul_635[7] + kernel_img_mul_635[8] + 
                kernel_img_mul_635[9] + kernel_img_mul_635[10] + kernel_img_mul_635[11] + 
                kernel_img_mul_635[12] + kernel_img_mul_635[13] + kernel_img_mul_635[14] + 
                kernel_img_mul_635[15] + kernel_img_mul_635[16] + kernel_img_mul_635[17] + 
                kernel_img_mul_635[18] + kernel_img_mul_635[19] + kernel_img_mul_635[20] + 
                kernel_img_mul_635[21] + kernel_img_mul_635[22] + kernel_img_mul_635[23] + 
                kernel_img_mul_635[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[5087:5080] <= 'd0;
  else if (current_state==ST_START)
    blur_din[5087:5080] <= kernel_img_sum_635[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5087:5080] <= 'd0;
end

wire  [39:0]  kernel_img_mul_636[0:24];
assign kernel_img_mul_636[0] = buffer_data_4[5079:5072] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_636[1] = buffer_data_4[5087:5080] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_636[2] = buffer_data_4[5095:5088] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_636[3] = buffer_data_4[5103:5096] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_636[4] = buffer_data_4[5111:5104] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_636[5] = buffer_data_3[5079:5072] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_636[6] = buffer_data_3[5087:5080] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_636[7] = buffer_data_3[5095:5088] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_636[8] = buffer_data_3[5103:5096] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_636[9] = buffer_data_3[5111:5104] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_636[10] = buffer_data_2[5079:5072] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_636[11] = buffer_data_2[5087:5080] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_636[12] = buffer_data_2[5095:5088] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_636[13] = buffer_data_2[5103:5096] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_636[14] = buffer_data_2[5111:5104] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_636[15] = buffer_data_1[5079:5072] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_636[16] = buffer_data_1[5087:5080] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_636[17] = buffer_data_1[5095:5088] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_636[18] = buffer_data_1[5103:5096] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_636[19] = buffer_data_1[5111:5104] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_636[20] = buffer_data_0[5079:5072] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_636[21] = buffer_data_0[5087:5080] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_636[22] = buffer_data_0[5095:5088] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_636[23] = buffer_data_0[5103:5096] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_636[24] = buffer_data_0[5111:5104] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_636 = kernel_img_mul_636[0] + kernel_img_mul_636[1] + kernel_img_mul_636[2] + 
                kernel_img_mul_636[3] + kernel_img_mul_636[4] + kernel_img_mul_636[5] + 
                kernel_img_mul_636[6] + kernel_img_mul_636[7] + kernel_img_mul_636[8] + 
                kernel_img_mul_636[9] + kernel_img_mul_636[10] + kernel_img_mul_636[11] + 
                kernel_img_mul_636[12] + kernel_img_mul_636[13] + kernel_img_mul_636[14] + 
                kernel_img_mul_636[15] + kernel_img_mul_636[16] + kernel_img_mul_636[17] + 
                kernel_img_mul_636[18] + kernel_img_mul_636[19] + kernel_img_mul_636[20] + 
                kernel_img_mul_636[21] + kernel_img_mul_636[22] + kernel_img_mul_636[23] + 
                kernel_img_mul_636[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[5095:5088] <= 'd0;
  else if (current_state==ST_START)
    blur_din[5095:5088] <= kernel_img_sum_636[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5095:5088] <= 'd0;
end

wire  [39:0]  kernel_img_mul_637[0:24];
assign kernel_img_mul_637[0] = buffer_data_4[5087:5080] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_637[1] = buffer_data_4[5095:5088] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_637[2] = buffer_data_4[5103:5096] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_637[3] = buffer_data_4[5111:5104] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_637[4] = buffer_data_4[5119:5112] * G_Kernel_5x5[0][159:128];
assign kernel_img_mul_637[5] = buffer_data_3[5087:5080] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_637[6] = buffer_data_3[5095:5088] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_637[7] = buffer_data_3[5103:5096] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_637[8] = buffer_data_3[5111:5104] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_637[9] = buffer_data_3[5119:5112] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_637[10] = buffer_data_2[5087:5080] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_637[11] = buffer_data_2[5095:5088] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_637[12] = buffer_data_2[5103:5096] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_637[13] = buffer_data_2[5111:5104] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_637[14] = buffer_data_2[5119:5112] * G_Kernel_5x5[2][159:128];
assign kernel_img_mul_637[15] = buffer_data_1[5087:5080] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_637[16] = buffer_data_1[5095:5088] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_637[17] = buffer_data_1[5103:5096] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_637[18] = buffer_data_1[5111:5104] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_637[19] = buffer_data_1[5119:5112] * G_Kernel_5x5[1][159:128];
assign kernel_img_mul_637[20] = buffer_data_0[5087:5080] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_637[21] = buffer_data_0[5095:5088] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_637[22] = buffer_data_0[5103:5096] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_637[23] = buffer_data_0[5111:5104] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_637[24] = buffer_data_0[5119:5112] * G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_637 = kernel_img_mul_637[0] + kernel_img_mul_637[1] + kernel_img_mul_637[2] + 
                kernel_img_mul_637[3] + kernel_img_mul_637[4] + kernel_img_mul_637[5] + 
                kernel_img_mul_637[6] + kernel_img_mul_637[7] + kernel_img_mul_637[8] + 
                kernel_img_mul_637[9] + kernel_img_mul_637[10] + kernel_img_mul_637[11] + 
                kernel_img_mul_637[12] + kernel_img_mul_637[13] + kernel_img_mul_637[14] + 
                kernel_img_mul_637[15] + kernel_img_mul_637[16] + kernel_img_mul_637[17] + 
                kernel_img_mul_637[18] + kernel_img_mul_637[19] + kernel_img_mul_637[20] + 
                kernel_img_mul_637[21] + kernel_img_mul_637[22] + kernel_img_mul_637[23] + 
                kernel_img_mul_637[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[5103:5096] <= 'd0;
  else if (current_state==ST_START)
    blur_din[5103:5096] <= kernel_img_sum_637[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5103:5096] <= 'd0;
end

wire  [39:0]  kernel_img_mul_638[0:24];
assign kernel_img_mul_638[0] = buffer_data_4[5095:5088] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_638[1] = buffer_data_4[5103:5096] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_638[2] = buffer_data_4[5111:5104] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_638[3] = buffer_data_4[5119:5112] * G_Kernel_5x5[0][127:96];
assign kernel_img_mul_638[5] = buffer_data_3[5095:5088] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_638[6] = buffer_data_3[5103:5096] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_638[7] = buffer_data_3[5111:5104] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_638[8] = buffer_data_3[5119:5112] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_638[10] = buffer_data_2[5095:5088] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_638[11] = buffer_data_2[5103:5096] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_638[12] = buffer_data_2[5111:5104] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_638[13] = buffer_data_2[5119:5112] * G_Kernel_5x5[2][127:96];
assign kernel_img_mul_638[15] = buffer_data_1[5095:5088] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_638[16] = buffer_data_1[5103:5096] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_638[17] = buffer_data_1[5111:5104] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_638[18] = buffer_data_1[5119:5112] * G_Kernel_5x5[1][127:96];
assign kernel_img_mul_638[20] = buffer_data_0[5095:5088] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_638[21] = buffer_data_0[5103:5096] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_638[22] = buffer_data_0[5111:5104] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_638[23] = buffer_data_0[5119:5112] * G_Kernel_5x5[0][127:96];
wire  [39:0]  kernel_img_sum_638 = kernel_img_mul_638[0] + kernel_img_mul_638[1] + kernel_img_mul_638[2] + 
                kernel_img_mul_638[3] + kernel_img_mul_638[5] + kernel_img_mul_638[6] + 
                kernel_img_mul_638[7] + kernel_img_mul_638[8] + kernel_img_mul_638[10] + 
                kernel_img_mul_638[11] + kernel_img_mul_638[12] + kernel_img_mul_638[13] + 
                kernel_img_mul_638[15] + kernel_img_mul_638[16] + kernel_img_mul_638[17] + 
                kernel_img_mul_638[18] + kernel_img_mul_638[20] + kernel_img_mul_638[21] + 
                kernel_img_mul_638[22] + kernel_img_mul_638[23] + 'd0;
always @(posedge clk) begin
  if (!rst_n)
    blur_din[5111:5104] <= 'd0;
  else if (current_state==ST_START)
    blur_din[5111:5104] <= kernel_img_sum_638[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5111:5104] <= 'd0;
end

wire  [39:0]  kernel_img_mul_639[0:24];
assign kernel_img_mul_639[0] = buffer_data_4[5103:5096] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_639[1] = buffer_data_4[5111:5104] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_639[2] = buffer_data_4[5119:5112] * G_Kernel_5x5[0][95:64];
assign kernel_img_mul_639[5] = buffer_data_3[5103:5096] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_639[6] = buffer_data_3[5111:5104] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_639[7] = buffer_data_3[5119:5112] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_639[10] = buffer_data_2[5103:5096] * G_Kernel_5x5[2][31:0];
assign kernel_img_mul_639[11] = buffer_data_2[5111:5104] * G_Kernel_5x5[2][63:32];
assign kernel_img_mul_639[12] = buffer_data_2[5119:5112] * G_Kernel_5x5[2][95:64];
assign kernel_img_mul_639[15] = buffer_data_1[5103:5096] * G_Kernel_5x5[1][31:0];
assign kernel_img_mul_639[16] = buffer_data_1[5111:5104] * G_Kernel_5x5[1][63:32];
assign kernel_img_mul_639[17] = buffer_data_1[5119:5112] * G_Kernel_5x5[1][95:64];
assign kernel_img_mul_639[20] = buffer_data_0[5103:5096] * G_Kernel_5x5[0][31:0];
assign kernel_img_mul_639[21] = buffer_data_0[5111:5104] * G_Kernel_5x5[0][63:32];
assign kernel_img_mul_639[22] = buffer_data_0[5119:5112] * G_Kernel_5x5[0][95:64];
wire  [39:0]  kernel_img_sum_639 = kernel_img_mul_639[0] + kernel_img_mul_639[1] + kernel_img_mul_639[2] + 
                kernel_img_mul_639[5] + kernel_img_mul_639[6] + kernel_img_mul_639[7] + 
                kernel_img_mul_639[10] + kernel_img_mul_639[11] + kernel_img_mul_639[12] + 
                kernel_img_mul_639[15] + kernel_img_mul_639[16] + kernel_img_mul_639[17] + 
                kernel_img_mul_639[20] + kernel_img_mul_639[21] + kernel_img_mul_639[22] + 
                'd0;
always @(posedge clk) begin
  if (!rst_n)
    blur_din[5119:5112] <= 'd0;
  else if (current_state==ST_START)
    blur_din[5119:5112] <= kernel_img_sum_639[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5119:5112] <= 'd0;
end




/*
 *  FSM
 *
 */

always @(posedge clk) begin
  if (!rst_n) begin
    current_state <= ST_IDLE;    
  end
  else begin
    current_state <= next_state;
  end
end

always @(*) begin
  case(current_state)
    ST_IDLE: begin
      if(start)
        next_state = ST_READY;
      else
        next_state = ST_IDLE;
    end
    ST_READY: begin
      if(ready_start_relay)
        next_state = ST_START;
      else 
        next_state = ST_READY;
    end
    ST_START: begin
      if(done)//CHANGE LATER
        next_state = ST_IDLE;
      else
        next_state = ST_START;
    end
    default:
      next_state = ST_IDLE;
  endcase
end



endmodule 