module bus_partition(
    img0,
    img1,
    img2,
    img3,
    img4,
    img_out0,
    img_out1,
    img_out2,
    img_out3,
    img_out4,
    buffer_col
);

input[5119:0]   img0,
                img1,
                img2,
                img3,
                img4;
output[175:0]   img_out0,
                img_out1,
                img_out2,
                img_out3,
                img_out4;
input[5:0]      buffer_col;

always @(*) begin
  case(buffer_col)
    'd0: begin
      img_out0[7:0] = 'd0;
      img_out0[15:8] = 'd0;
      img_out0[23:16] = 'd0;
      img_out0[31:24] = img0[7:0];
      img_out0[39:32] = img0[15:8];
      img_out0[47:40] = img0[23:16];
      img_out0[55:48] = img0[31:24];
      img_out0[63:56] = img0[39:32];
      img_out0[71:64] = img0[47:40];
      img_out0[79:72] = img0[55:48];
      img_out0[87:80] = img0[63:56];
      img_out0[95:88] = img0[71:64];
      img_out0[103:96] = img0[79:72];
      img_out0[111:104] = img0[87:80];
      img_out0[119:112] = img0[95:88];
      img_out0[127:120] = img0[103:96];
      img_out0[135:128] = img0[111:104];
      img_out0[143:136] = img0[119:112];
      img_out0[151:144] = img0[127:120];
      img_out0[159:152] = img0[135:128];
      img_out0[167:160] = img0[143:136];
      img_out0[175:168] = img0[151:144];
      img_out1[7:0] = 'd0;
      img_out1[15:8] = 'd0;
      img_out1[23:16] = 'd0;
      img_out1[31:24] = img1[7:0];
      img_out1[39:32] = img1[15:8];
      img_out1[47:40] = img1[23:16];
      img_out1[55:48] = img1[31:24];
      img_out1[63:56] = img1[39:32];
      img_out1[71:64] = img1[47:40];
      img_out1[79:72] = img1[55:48];
      img_out1[87:80] = img1[63:56];
      img_out1[95:88] = img1[71:64];
      img_out1[103:96] = img1[79:72];
      img_out1[111:104] = img1[87:80];
      img_out1[119:112] = img1[95:88];
      img_out1[127:120] = img1[103:96];
      img_out1[135:128] = img1[111:104];
      img_out1[143:136] = img1[119:112];
      img_out1[151:144] = img1[127:120];
      img_out1[159:152] = img1[135:128];
      img_out1[167:160] = img1[143:136];
      img_out1[175:168] = img1[151:144];
      img_out2[7:0] = 'd0;
      img_out2[15:8] = 'd0;
      img_out2[23:16] = 'd0;
      img_out2[31:24] = img2[7:0];
      img_out2[39:32] = img2[15:8];
      img_out2[47:40] = img2[23:16];
      img_out2[55:48] = img2[31:24];
      img_out2[63:56] = img2[39:32];
      img_out2[71:64] = img2[47:40];
      img_out2[79:72] = img2[55:48];
      img_out2[87:80] = img2[63:56];
      img_out2[95:88] = img2[71:64];
      img_out2[103:96] = img2[79:72];
      img_out2[111:104] = img2[87:80];
      img_out2[119:112] = img2[95:88];
      img_out2[127:120] = img2[103:96];
      img_out2[135:128] = img2[111:104];
      img_out2[143:136] = img2[119:112];
      img_out2[151:144] = img2[127:120];
      img_out2[159:152] = img2[135:128];
      img_out2[167:160] = img2[143:136];
      img_out2[175:168] = img2[151:144];
      img_out3[7:0] = 'd0;
      img_out3[15:8] = 'd0;
      img_out3[23:16] = 'd0;
      img_out3[31:24] = img3[7:0];
      img_out3[39:32] = img3[15:8];
      img_out3[47:40] = img3[23:16];
      img_out3[55:48] = img3[31:24];
      img_out3[63:56] = img3[39:32];
      img_out3[71:64] = img3[47:40];
      img_out3[79:72] = img3[55:48];
      img_out3[87:80] = img3[63:56];
      img_out3[95:88] = img3[71:64];
      img_out3[103:96] = img3[79:72];
      img_out3[111:104] = img3[87:80];
      img_out3[119:112] = img3[95:88];
      img_out3[127:120] = img3[103:96];
      img_out3[135:128] = img3[111:104];
      img_out3[143:136] = img3[119:112];
      img_out3[151:144] = img3[127:120];
      img_out3[159:152] = img3[135:128];
      img_out3[167:160] = img3[143:136];
      img_out3[175:168] = img3[151:144];
      img_out4[7:0] = 'd0;
      img_out4[15:8] = 'd0;
      img_out4[23:16] = 'd0;
      img_out4[31:24] = img4[7:0];
      img_out4[39:32] = img4[15:8];
      img_out4[47:40] = img4[23:16];
      img_out4[55:48] = img4[31:24];
      img_out4[63:56] = img4[39:32];
      img_out4[71:64] = img4[47:40];
      img_out4[79:72] = img4[55:48];
      img_out4[87:80] = img4[63:56];
      img_out4[95:88] = img4[71:64];
      img_out4[103:96] = img4[79:72];
      img_out4[111:104] = img4[87:80];
      img_out4[119:112] = img4[95:88];
      img_out4[127:120] = img4[103:96];
      img_out4[135:128] = img4[111:104];
      img_out4[143:136] = img4[119:112];
      img_out4[151:144] = img4[127:120];
      img_out4[159:152] = img4[135:128];
      img_out4[167:160] = img4[143:136];
      img_out4[175:168] = img4[151:144];
    end
    'd1: begin
      img_out0[7:0] = img0[111:104];
      img_out0[15:8] = img0[119:112];
      img_out0[23:16] = img0[127:120];
      img_out0[31:24] = img0[135:128];
      img_out0[39:32] = img0[143:136];
      img_out0[47:40] = img0[151:144];
      img_out0[55:48] = img0[159:152];
      img_out0[63:56] = img0[167:160];
      img_out0[71:64] = img0[175:168];
      img_out0[79:72] = img0[183:176];
      img_out0[87:80] = img0[191:184];
      img_out0[95:88] = img0[199:192];
      img_out0[103:96] = img0[207:200];
      img_out0[111:104] = img0[215:208];
      img_out0[119:112] = img0[223:216];
      img_out0[127:120] = img0[231:224];
      img_out0[135:128] = img0[239:232];
      img_out0[143:136] = img0[247:240];
      img_out0[151:144] = img0[255:248];
      img_out0[159:152] = img0[263:256];
      img_out0[167:160] = img0[271:264];
      img_out0[175:168] = img0[279:272];
      img_out1[7:0] = img1[111:104];
      img_out1[15:8] = img1[119:112];
      img_out1[23:16] = img1[127:120];
      img_out1[31:24] = img1[135:128];
      img_out1[39:32] = img1[143:136];
      img_out1[47:40] = img1[151:144];
      img_out1[55:48] = img1[159:152];
      img_out1[63:56] = img1[167:160];
      img_out1[71:64] = img1[175:168];
      img_out1[79:72] = img1[183:176];
      img_out1[87:80] = img1[191:184];
      img_out1[95:88] = img1[199:192];
      img_out1[103:96] = img1[207:200];
      img_out1[111:104] = img1[215:208];
      img_out1[119:112] = img1[223:216];
      img_out1[127:120] = img1[231:224];
      img_out1[135:128] = img1[239:232];
      img_out1[143:136] = img1[247:240];
      img_out1[151:144] = img1[255:248];
      img_out1[159:152] = img1[263:256];
      img_out1[167:160] = img1[271:264];
      img_out1[175:168] = img1[279:272];
      img_out2[7:0] = img2[111:104];
      img_out2[15:8] = img2[119:112];
      img_out2[23:16] = img2[127:120];
      img_out2[31:24] = img2[135:128];
      img_out2[39:32] = img2[143:136];
      img_out2[47:40] = img2[151:144];
      img_out2[55:48] = img2[159:152];
      img_out2[63:56] = img2[167:160];
      img_out2[71:64] = img2[175:168];
      img_out2[79:72] = img2[183:176];
      img_out2[87:80] = img2[191:184];
      img_out2[95:88] = img2[199:192];
      img_out2[103:96] = img2[207:200];
      img_out2[111:104] = img2[215:208];
      img_out2[119:112] = img2[223:216];
      img_out2[127:120] = img2[231:224];
      img_out2[135:128] = img2[239:232];
      img_out2[143:136] = img2[247:240];
      img_out2[151:144] = img2[255:248];
      img_out2[159:152] = img2[263:256];
      img_out2[167:160] = img2[271:264];
      img_out2[175:168] = img2[279:272];
      img_out3[7:0] = img3[111:104];
      img_out3[15:8] = img3[119:112];
      img_out3[23:16] = img3[127:120];
      img_out3[31:24] = img3[135:128];
      img_out3[39:32] = img3[143:136];
      img_out3[47:40] = img3[151:144];
      img_out3[55:48] = img3[159:152];
      img_out3[63:56] = img3[167:160];
      img_out3[71:64] = img3[175:168];
      img_out3[79:72] = img3[183:176];
      img_out3[87:80] = img3[191:184];
      img_out3[95:88] = img3[199:192];
      img_out3[103:96] = img3[207:200];
      img_out3[111:104] = img3[215:208];
      img_out3[119:112] = img3[223:216];
      img_out3[127:120] = img3[231:224];
      img_out3[135:128] = img3[239:232];
      img_out3[143:136] = img3[247:240];
      img_out3[151:144] = img3[255:248];
      img_out3[159:152] = img3[263:256];
      img_out3[167:160] = img3[271:264];
      img_out3[175:168] = img3[279:272];
      img_out4[7:0] = img4[111:104];
      img_out4[15:8] = img4[119:112];
      img_out4[23:16] = img4[127:120];
      img_out4[31:24] = img4[135:128];
      img_out4[39:32] = img4[143:136];
      img_out4[47:40] = img4[151:144];
      img_out4[55:48] = img4[159:152];
      img_out4[63:56] = img4[167:160];
      img_out4[71:64] = img4[175:168];
      img_out4[79:72] = img4[183:176];
      img_out4[87:80] = img4[191:184];
      img_out4[95:88] = img4[199:192];
      img_out4[103:96] = img4[207:200];
      img_out4[111:104] = img4[215:208];
      img_out4[119:112] = img4[223:216];
      img_out4[127:120] = img4[231:224];
      img_out4[135:128] = img4[239:232];
      img_out4[143:136] = img4[247:240];
      img_out4[151:144] = img4[255:248];
      img_out4[159:152] = img4[263:256];
      img_out4[167:160] = img4[271:264];
      img_out4[175:168] = img4[279:272];
    end
    'd2: begin
      img_out0[7:0] = img0[239:232];
      img_out0[15:8] = img0[247:240];
      img_out0[23:16] = img0[255:248];
      img_out0[31:24] = img0[263:256];
      img_out0[39:32] = img0[271:264];
      img_out0[47:40] = img0[279:272];
      img_out0[55:48] = img0[287:280];
      img_out0[63:56] = img0[295:288];
      img_out0[71:64] = img0[303:296];
      img_out0[79:72] = img0[311:304];
      img_out0[87:80] = img0[319:312];
      img_out0[95:88] = img0[327:320];
      img_out0[103:96] = img0[335:328];
      img_out0[111:104] = img0[343:336];
      img_out0[119:112] = img0[351:344];
      img_out0[127:120] = img0[359:352];
      img_out0[135:128] = img0[367:360];
      img_out0[143:136] = img0[375:368];
      img_out0[151:144] = img0[383:376];
      img_out0[159:152] = img0[391:384];
      img_out0[167:160] = img0[399:392];
      img_out0[175:168] = img0[407:400];
      img_out1[7:0] = img1[239:232];
      img_out1[15:8] = img1[247:240];
      img_out1[23:16] = img1[255:248];
      img_out1[31:24] = img1[263:256];
      img_out1[39:32] = img1[271:264];
      img_out1[47:40] = img1[279:272];
      img_out1[55:48] = img1[287:280];
      img_out1[63:56] = img1[295:288];
      img_out1[71:64] = img1[303:296];
      img_out1[79:72] = img1[311:304];
      img_out1[87:80] = img1[319:312];
      img_out1[95:88] = img1[327:320];
      img_out1[103:96] = img1[335:328];
      img_out1[111:104] = img1[343:336];
      img_out1[119:112] = img1[351:344];
      img_out1[127:120] = img1[359:352];
      img_out1[135:128] = img1[367:360];
      img_out1[143:136] = img1[375:368];
      img_out1[151:144] = img1[383:376];
      img_out1[159:152] = img1[391:384];
      img_out1[167:160] = img1[399:392];
      img_out1[175:168] = img1[407:400];
      img_out2[7:0] = img2[239:232];
      img_out2[15:8] = img2[247:240];
      img_out2[23:16] = img2[255:248];
      img_out2[31:24] = img2[263:256];
      img_out2[39:32] = img2[271:264];
      img_out2[47:40] = img2[279:272];
      img_out2[55:48] = img2[287:280];
      img_out2[63:56] = img2[295:288];
      img_out2[71:64] = img2[303:296];
      img_out2[79:72] = img2[311:304];
      img_out2[87:80] = img2[319:312];
      img_out2[95:88] = img2[327:320];
      img_out2[103:96] = img2[335:328];
      img_out2[111:104] = img2[343:336];
      img_out2[119:112] = img2[351:344];
      img_out2[127:120] = img2[359:352];
      img_out2[135:128] = img2[367:360];
      img_out2[143:136] = img2[375:368];
      img_out2[151:144] = img2[383:376];
      img_out2[159:152] = img2[391:384];
      img_out2[167:160] = img2[399:392];
      img_out2[175:168] = img2[407:400];
      img_out3[7:0] = img3[239:232];
      img_out3[15:8] = img3[247:240];
      img_out3[23:16] = img3[255:248];
      img_out3[31:24] = img3[263:256];
      img_out3[39:32] = img3[271:264];
      img_out3[47:40] = img3[279:272];
      img_out3[55:48] = img3[287:280];
      img_out3[63:56] = img3[295:288];
      img_out3[71:64] = img3[303:296];
      img_out3[79:72] = img3[311:304];
      img_out3[87:80] = img3[319:312];
      img_out3[95:88] = img3[327:320];
      img_out3[103:96] = img3[335:328];
      img_out3[111:104] = img3[343:336];
      img_out3[119:112] = img3[351:344];
      img_out3[127:120] = img3[359:352];
      img_out3[135:128] = img3[367:360];
      img_out3[143:136] = img3[375:368];
      img_out3[151:144] = img3[383:376];
      img_out3[159:152] = img3[391:384];
      img_out3[167:160] = img3[399:392];
      img_out3[175:168] = img3[407:400];
      img_out4[7:0] = img4[239:232];
      img_out4[15:8] = img4[247:240];
      img_out4[23:16] = img4[255:248];
      img_out4[31:24] = img4[263:256];
      img_out4[39:32] = img4[271:264];
      img_out4[47:40] = img4[279:272];
      img_out4[55:48] = img4[287:280];
      img_out4[63:56] = img4[295:288];
      img_out4[71:64] = img4[303:296];
      img_out4[79:72] = img4[311:304];
      img_out4[87:80] = img4[319:312];
      img_out4[95:88] = img4[327:320];
      img_out4[103:96] = img4[335:328];
      img_out4[111:104] = img4[343:336];
      img_out4[119:112] = img4[351:344];
      img_out4[127:120] = img4[359:352];
      img_out4[135:128] = img4[367:360];
      img_out4[143:136] = img4[375:368];
      img_out4[151:144] = img4[383:376];
      img_out4[159:152] = img4[391:384];
      img_out4[167:160] = img4[399:392];
      img_out4[175:168] = img4[407:400];
    end
    'd3: begin
      img_out0[7:0] = img0[367:360];
      img_out0[15:8] = img0[375:368];
      img_out0[23:16] = img0[383:376];
      img_out0[31:24] = img0[391:384];
      img_out0[39:32] = img0[399:392];
      img_out0[47:40] = img0[407:400];
      img_out0[55:48] = img0[415:408];
      img_out0[63:56] = img0[423:416];
      img_out0[71:64] = img0[431:424];
      img_out0[79:72] = img0[439:432];
      img_out0[87:80] = img0[447:440];
      img_out0[95:88] = img0[455:448];
      img_out0[103:96] = img0[463:456];
      img_out0[111:104] = img0[471:464];
      img_out0[119:112] = img0[479:472];
      img_out0[127:120] = img0[487:480];
      img_out0[135:128] = img0[495:488];
      img_out0[143:136] = img0[503:496];
      img_out0[151:144] = img0[511:504];
      img_out0[159:152] = img0[519:512];
      img_out0[167:160] = img0[527:520];
      img_out0[175:168] = img0[535:528];
      img_out1[7:0] = img1[367:360];
      img_out1[15:8] = img1[375:368];
      img_out1[23:16] = img1[383:376];
      img_out1[31:24] = img1[391:384];
      img_out1[39:32] = img1[399:392];
      img_out1[47:40] = img1[407:400];
      img_out1[55:48] = img1[415:408];
      img_out1[63:56] = img1[423:416];
      img_out1[71:64] = img1[431:424];
      img_out1[79:72] = img1[439:432];
      img_out1[87:80] = img1[447:440];
      img_out1[95:88] = img1[455:448];
      img_out1[103:96] = img1[463:456];
      img_out1[111:104] = img1[471:464];
      img_out1[119:112] = img1[479:472];
      img_out1[127:120] = img1[487:480];
      img_out1[135:128] = img1[495:488];
      img_out1[143:136] = img1[503:496];
      img_out1[151:144] = img1[511:504];
      img_out1[159:152] = img1[519:512];
      img_out1[167:160] = img1[527:520];
      img_out1[175:168] = img1[535:528];
      img_out2[7:0] = img2[367:360];
      img_out2[15:8] = img2[375:368];
      img_out2[23:16] = img2[383:376];
      img_out2[31:24] = img2[391:384];
      img_out2[39:32] = img2[399:392];
      img_out2[47:40] = img2[407:400];
      img_out2[55:48] = img2[415:408];
      img_out2[63:56] = img2[423:416];
      img_out2[71:64] = img2[431:424];
      img_out2[79:72] = img2[439:432];
      img_out2[87:80] = img2[447:440];
      img_out2[95:88] = img2[455:448];
      img_out2[103:96] = img2[463:456];
      img_out2[111:104] = img2[471:464];
      img_out2[119:112] = img2[479:472];
      img_out2[127:120] = img2[487:480];
      img_out2[135:128] = img2[495:488];
      img_out2[143:136] = img2[503:496];
      img_out2[151:144] = img2[511:504];
      img_out2[159:152] = img2[519:512];
      img_out2[167:160] = img2[527:520];
      img_out2[175:168] = img2[535:528];
      img_out3[7:0] = img3[367:360];
      img_out3[15:8] = img3[375:368];
      img_out3[23:16] = img3[383:376];
      img_out3[31:24] = img3[391:384];
      img_out3[39:32] = img3[399:392];
      img_out3[47:40] = img3[407:400];
      img_out3[55:48] = img3[415:408];
      img_out3[63:56] = img3[423:416];
      img_out3[71:64] = img3[431:424];
      img_out3[79:72] = img3[439:432];
      img_out3[87:80] = img3[447:440];
      img_out3[95:88] = img3[455:448];
      img_out3[103:96] = img3[463:456];
      img_out3[111:104] = img3[471:464];
      img_out3[119:112] = img3[479:472];
      img_out3[127:120] = img3[487:480];
      img_out3[135:128] = img3[495:488];
      img_out3[143:136] = img3[503:496];
      img_out3[151:144] = img3[511:504];
      img_out3[159:152] = img3[519:512];
      img_out3[167:160] = img3[527:520];
      img_out3[175:168] = img3[535:528];
      img_out4[7:0] = img4[367:360];
      img_out4[15:8] = img4[375:368];
      img_out4[23:16] = img4[383:376];
      img_out4[31:24] = img4[391:384];
      img_out4[39:32] = img4[399:392];
      img_out4[47:40] = img4[407:400];
      img_out4[55:48] = img4[415:408];
      img_out4[63:56] = img4[423:416];
      img_out4[71:64] = img4[431:424];
      img_out4[79:72] = img4[439:432];
      img_out4[87:80] = img4[447:440];
      img_out4[95:88] = img4[455:448];
      img_out4[103:96] = img4[463:456];
      img_out4[111:104] = img4[471:464];
      img_out4[119:112] = img4[479:472];
      img_out4[127:120] = img4[487:480];
      img_out4[135:128] = img4[495:488];
      img_out4[143:136] = img4[503:496];
      img_out4[151:144] = img4[511:504];
      img_out4[159:152] = img4[519:512];
      img_out4[167:160] = img4[527:520];
      img_out4[175:168] = img4[535:528];
    end
    'd4: begin
      img_out0[7:0] = img0[495:488];
      img_out0[15:8] = img0[503:496];
      img_out0[23:16] = img0[511:504];
      img_out0[31:24] = img0[519:512];
      img_out0[39:32] = img0[527:520];
      img_out0[47:40] = img0[535:528];
      img_out0[55:48] = img0[543:536];
      img_out0[63:56] = img0[551:544];
      img_out0[71:64] = img0[559:552];
      img_out0[79:72] = img0[567:560];
      img_out0[87:80] = img0[575:568];
      img_out0[95:88] = img0[583:576];
      img_out0[103:96] = img0[591:584];
      img_out0[111:104] = img0[599:592];
      img_out0[119:112] = img0[607:600];
      img_out0[127:120] = img0[615:608];
      img_out0[135:128] = img0[623:616];
      img_out0[143:136] = img0[631:624];
      img_out0[151:144] = img0[639:632];
      img_out0[159:152] = img0[647:640];
      img_out0[167:160] = img0[655:648];
      img_out0[175:168] = img0[663:656];
      img_out1[7:0] = img1[495:488];
      img_out1[15:8] = img1[503:496];
      img_out1[23:16] = img1[511:504];
      img_out1[31:24] = img1[519:512];
      img_out1[39:32] = img1[527:520];
      img_out1[47:40] = img1[535:528];
      img_out1[55:48] = img1[543:536];
      img_out1[63:56] = img1[551:544];
      img_out1[71:64] = img1[559:552];
      img_out1[79:72] = img1[567:560];
      img_out1[87:80] = img1[575:568];
      img_out1[95:88] = img1[583:576];
      img_out1[103:96] = img1[591:584];
      img_out1[111:104] = img1[599:592];
      img_out1[119:112] = img1[607:600];
      img_out1[127:120] = img1[615:608];
      img_out1[135:128] = img1[623:616];
      img_out1[143:136] = img1[631:624];
      img_out1[151:144] = img1[639:632];
      img_out1[159:152] = img1[647:640];
      img_out1[167:160] = img1[655:648];
      img_out1[175:168] = img1[663:656];
      img_out2[7:0] = img2[495:488];
      img_out2[15:8] = img2[503:496];
      img_out2[23:16] = img2[511:504];
      img_out2[31:24] = img2[519:512];
      img_out2[39:32] = img2[527:520];
      img_out2[47:40] = img2[535:528];
      img_out2[55:48] = img2[543:536];
      img_out2[63:56] = img2[551:544];
      img_out2[71:64] = img2[559:552];
      img_out2[79:72] = img2[567:560];
      img_out2[87:80] = img2[575:568];
      img_out2[95:88] = img2[583:576];
      img_out2[103:96] = img2[591:584];
      img_out2[111:104] = img2[599:592];
      img_out2[119:112] = img2[607:600];
      img_out2[127:120] = img2[615:608];
      img_out2[135:128] = img2[623:616];
      img_out2[143:136] = img2[631:624];
      img_out2[151:144] = img2[639:632];
      img_out2[159:152] = img2[647:640];
      img_out2[167:160] = img2[655:648];
      img_out2[175:168] = img2[663:656];
      img_out3[7:0] = img3[495:488];
      img_out3[15:8] = img3[503:496];
      img_out3[23:16] = img3[511:504];
      img_out3[31:24] = img3[519:512];
      img_out3[39:32] = img3[527:520];
      img_out3[47:40] = img3[535:528];
      img_out3[55:48] = img3[543:536];
      img_out3[63:56] = img3[551:544];
      img_out3[71:64] = img3[559:552];
      img_out3[79:72] = img3[567:560];
      img_out3[87:80] = img3[575:568];
      img_out3[95:88] = img3[583:576];
      img_out3[103:96] = img3[591:584];
      img_out3[111:104] = img3[599:592];
      img_out3[119:112] = img3[607:600];
      img_out3[127:120] = img3[615:608];
      img_out3[135:128] = img3[623:616];
      img_out3[143:136] = img3[631:624];
      img_out3[151:144] = img3[639:632];
      img_out3[159:152] = img3[647:640];
      img_out3[167:160] = img3[655:648];
      img_out3[175:168] = img3[663:656];
      img_out4[7:0] = img4[495:488];
      img_out4[15:8] = img4[503:496];
      img_out4[23:16] = img4[511:504];
      img_out4[31:24] = img4[519:512];
      img_out4[39:32] = img4[527:520];
      img_out4[47:40] = img4[535:528];
      img_out4[55:48] = img4[543:536];
      img_out4[63:56] = img4[551:544];
      img_out4[71:64] = img4[559:552];
      img_out4[79:72] = img4[567:560];
      img_out4[87:80] = img4[575:568];
      img_out4[95:88] = img4[583:576];
      img_out4[103:96] = img4[591:584];
      img_out4[111:104] = img4[599:592];
      img_out4[119:112] = img4[607:600];
      img_out4[127:120] = img4[615:608];
      img_out4[135:128] = img4[623:616];
      img_out4[143:136] = img4[631:624];
      img_out4[151:144] = img4[639:632];
      img_out4[159:152] = img4[647:640];
      img_out4[167:160] = img4[655:648];
      img_out4[175:168] = img4[663:656];
    end
    'd5: begin
      img_out0[7:0] = img0[623:616];
      img_out0[15:8] = img0[631:624];
      img_out0[23:16] = img0[639:632];
      img_out0[31:24] = img0[647:640];
      img_out0[39:32] = img0[655:648];
      img_out0[47:40] = img0[663:656];
      img_out0[55:48] = img0[671:664];
      img_out0[63:56] = img0[679:672];
      img_out0[71:64] = img0[687:680];
      img_out0[79:72] = img0[695:688];
      img_out0[87:80] = img0[703:696];
      img_out0[95:88] = img0[711:704];
      img_out0[103:96] = img0[719:712];
      img_out0[111:104] = img0[727:720];
      img_out0[119:112] = img0[735:728];
      img_out0[127:120] = img0[743:736];
      img_out0[135:128] = img0[751:744];
      img_out0[143:136] = img0[759:752];
      img_out0[151:144] = img0[767:760];
      img_out0[159:152] = img0[775:768];
      img_out0[167:160] = img0[783:776];
      img_out0[175:168] = img0[791:784];
      img_out1[7:0] = img1[623:616];
      img_out1[15:8] = img1[631:624];
      img_out1[23:16] = img1[639:632];
      img_out1[31:24] = img1[647:640];
      img_out1[39:32] = img1[655:648];
      img_out1[47:40] = img1[663:656];
      img_out1[55:48] = img1[671:664];
      img_out1[63:56] = img1[679:672];
      img_out1[71:64] = img1[687:680];
      img_out1[79:72] = img1[695:688];
      img_out1[87:80] = img1[703:696];
      img_out1[95:88] = img1[711:704];
      img_out1[103:96] = img1[719:712];
      img_out1[111:104] = img1[727:720];
      img_out1[119:112] = img1[735:728];
      img_out1[127:120] = img1[743:736];
      img_out1[135:128] = img1[751:744];
      img_out1[143:136] = img1[759:752];
      img_out1[151:144] = img1[767:760];
      img_out1[159:152] = img1[775:768];
      img_out1[167:160] = img1[783:776];
      img_out1[175:168] = img1[791:784];
      img_out2[7:0] = img2[623:616];
      img_out2[15:8] = img2[631:624];
      img_out2[23:16] = img2[639:632];
      img_out2[31:24] = img2[647:640];
      img_out2[39:32] = img2[655:648];
      img_out2[47:40] = img2[663:656];
      img_out2[55:48] = img2[671:664];
      img_out2[63:56] = img2[679:672];
      img_out2[71:64] = img2[687:680];
      img_out2[79:72] = img2[695:688];
      img_out2[87:80] = img2[703:696];
      img_out2[95:88] = img2[711:704];
      img_out2[103:96] = img2[719:712];
      img_out2[111:104] = img2[727:720];
      img_out2[119:112] = img2[735:728];
      img_out2[127:120] = img2[743:736];
      img_out2[135:128] = img2[751:744];
      img_out2[143:136] = img2[759:752];
      img_out2[151:144] = img2[767:760];
      img_out2[159:152] = img2[775:768];
      img_out2[167:160] = img2[783:776];
      img_out2[175:168] = img2[791:784];
      img_out3[7:0] = img3[623:616];
      img_out3[15:8] = img3[631:624];
      img_out3[23:16] = img3[639:632];
      img_out3[31:24] = img3[647:640];
      img_out3[39:32] = img3[655:648];
      img_out3[47:40] = img3[663:656];
      img_out3[55:48] = img3[671:664];
      img_out3[63:56] = img3[679:672];
      img_out3[71:64] = img3[687:680];
      img_out3[79:72] = img3[695:688];
      img_out3[87:80] = img3[703:696];
      img_out3[95:88] = img3[711:704];
      img_out3[103:96] = img3[719:712];
      img_out3[111:104] = img3[727:720];
      img_out3[119:112] = img3[735:728];
      img_out3[127:120] = img3[743:736];
      img_out3[135:128] = img3[751:744];
      img_out3[143:136] = img3[759:752];
      img_out3[151:144] = img3[767:760];
      img_out3[159:152] = img3[775:768];
      img_out3[167:160] = img3[783:776];
      img_out3[175:168] = img3[791:784];
      img_out4[7:0] = img4[623:616];
      img_out4[15:8] = img4[631:624];
      img_out4[23:16] = img4[639:632];
      img_out4[31:24] = img4[647:640];
      img_out4[39:32] = img4[655:648];
      img_out4[47:40] = img4[663:656];
      img_out4[55:48] = img4[671:664];
      img_out4[63:56] = img4[679:672];
      img_out4[71:64] = img4[687:680];
      img_out4[79:72] = img4[695:688];
      img_out4[87:80] = img4[703:696];
      img_out4[95:88] = img4[711:704];
      img_out4[103:96] = img4[719:712];
      img_out4[111:104] = img4[727:720];
      img_out4[119:112] = img4[735:728];
      img_out4[127:120] = img4[743:736];
      img_out4[135:128] = img4[751:744];
      img_out4[143:136] = img4[759:752];
      img_out4[151:144] = img4[767:760];
      img_out4[159:152] = img4[775:768];
      img_out4[167:160] = img4[783:776];
      img_out4[175:168] = img4[791:784];
    end
    'd6: begin
      img_out0[7:0] = img0[751:744];
      img_out0[15:8] = img0[759:752];
      img_out0[23:16] = img0[767:760];
      img_out0[31:24] = img0[775:768];
      img_out0[39:32] = img0[783:776];
      img_out0[47:40] = img0[791:784];
      img_out0[55:48] = img0[799:792];
      img_out0[63:56] = img0[807:800];
      img_out0[71:64] = img0[815:808];
      img_out0[79:72] = img0[823:816];
      img_out0[87:80] = img0[831:824];
      img_out0[95:88] = img0[839:832];
      img_out0[103:96] = img0[847:840];
      img_out0[111:104] = img0[855:848];
      img_out0[119:112] = img0[863:856];
      img_out0[127:120] = img0[871:864];
      img_out0[135:128] = img0[879:872];
      img_out0[143:136] = img0[887:880];
      img_out0[151:144] = img0[895:888];
      img_out0[159:152] = img0[903:896];
      img_out0[167:160] = img0[911:904];
      img_out0[175:168] = img0[919:912];
      img_out1[7:0] = img1[751:744];
      img_out1[15:8] = img1[759:752];
      img_out1[23:16] = img1[767:760];
      img_out1[31:24] = img1[775:768];
      img_out1[39:32] = img1[783:776];
      img_out1[47:40] = img1[791:784];
      img_out1[55:48] = img1[799:792];
      img_out1[63:56] = img1[807:800];
      img_out1[71:64] = img1[815:808];
      img_out1[79:72] = img1[823:816];
      img_out1[87:80] = img1[831:824];
      img_out1[95:88] = img1[839:832];
      img_out1[103:96] = img1[847:840];
      img_out1[111:104] = img1[855:848];
      img_out1[119:112] = img1[863:856];
      img_out1[127:120] = img1[871:864];
      img_out1[135:128] = img1[879:872];
      img_out1[143:136] = img1[887:880];
      img_out1[151:144] = img1[895:888];
      img_out1[159:152] = img1[903:896];
      img_out1[167:160] = img1[911:904];
      img_out1[175:168] = img1[919:912];
      img_out2[7:0] = img2[751:744];
      img_out2[15:8] = img2[759:752];
      img_out2[23:16] = img2[767:760];
      img_out2[31:24] = img2[775:768];
      img_out2[39:32] = img2[783:776];
      img_out2[47:40] = img2[791:784];
      img_out2[55:48] = img2[799:792];
      img_out2[63:56] = img2[807:800];
      img_out2[71:64] = img2[815:808];
      img_out2[79:72] = img2[823:816];
      img_out2[87:80] = img2[831:824];
      img_out2[95:88] = img2[839:832];
      img_out2[103:96] = img2[847:840];
      img_out2[111:104] = img2[855:848];
      img_out2[119:112] = img2[863:856];
      img_out2[127:120] = img2[871:864];
      img_out2[135:128] = img2[879:872];
      img_out2[143:136] = img2[887:880];
      img_out2[151:144] = img2[895:888];
      img_out2[159:152] = img2[903:896];
      img_out2[167:160] = img2[911:904];
      img_out2[175:168] = img2[919:912];
      img_out3[7:0] = img3[751:744];
      img_out3[15:8] = img3[759:752];
      img_out3[23:16] = img3[767:760];
      img_out3[31:24] = img3[775:768];
      img_out3[39:32] = img3[783:776];
      img_out3[47:40] = img3[791:784];
      img_out3[55:48] = img3[799:792];
      img_out3[63:56] = img3[807:800];
      img_out3[71:64] = img3[815:808];
      img_out3[79:72] = img3[823:816];
      img_out3[87:80] = img3[831:824];
      img_out3[95:88] = img3[839:832];
      img_out3[103:96] = img3[847:840];
      img_out3[111:104] = img3[855:848];
      img_out3[119:112] = img3[863:856];
      img_out3[127:120] = img3[871:864];
      img_out3[135:128] = img3[879:872];
      img_out3[143:136] = img3[887:880];
      img_out3[151:144] = img3[895:888];
      img_out3[159:152] = img3[903:896];
      img_out3[167:160] = img3[911:904];
      img_out3[175:168] = img3[919:912];
      img_out4[7:0] = img4[751:744];
      img_out4[15:8] = img4[759:752];
      img_out4[23:16] = img4[767:760];
      img_out4[31:24] = img4[775:768];
      img_out4[39:32] = img4[783:776];
      img_out4[47:40] = img4[791:784];
      img_out4[55:48] = img4[799:792];
      img_out4[63:56] = img4[807:800];
      img_out4[71:64] = img4[815:808];
      img_out4[79:72] = img4[823:816];
      img_out4[87:80] = img4[831:824];
      img_out4[95:88] = img4[839:832];
      img_out4[103:96] = img4[847:840];
      img_out4[111:104] = img4[855:848];
      img_out4[119:112] = img4[863:856];
      img_out4[127:120] = img4[871:864];
      img_out4[135:128] = img4[879:872];
      img_out4[143:136] = img4[887:880];
      img_out4[151:144] = img4[895:888];
      img_out4[159:152] = img4[903:896];
      img_out4[167:160] = img4[911:904];
      img_out4[175:168] = img4[919:912];
    end
    'd7: begin
      img_out0[7:0] = img0[879:872];
      img_out0[15:8] = img0[887:880];
      img_out0[23:16] = img0[895:888];
      img_out0[31:24] = img0[903:896];
      img_out0[39:32] = img0[911:904];
      img_out0[47:40] = img0[919:912];
      img_out0[55:48] = img0[927:920];
      img_out0[63:56] = img0[935:928];
      img_out0[71:64] = img0[943:936];
      img_out0[79:72] = img0[951:944];
      img_out0[87:80] = img0[959:952];
      img_out0[95:88] = img0[967:960];
      img_out0[103:96] = img0[975:968];
      img_out0[111:104] = img0[983:976];
      img_out0[119:112] = img0[991:984];
      img_out0[127:120] = img0[999:992];
      img_out0[135:128] = img0[1007:1000];
      img_out0[143:136] = img0[1015:1008];
      img_out0[151:144] = img0[1023:1016];
      img_out0[159:152] = img0[1031:1024];
      img_out0[167:160] = img0[1039:1032];
      img_out0[175:168] = img0[1047:1040];
      img_out1[7:0] = img1[879:872];
      img_out1[15:8] = img1[887:880];
      img_out1[23:16] = img1[895:888];
      img_out1[31:24] = img1[903:896];
      img_out1[39:32] = img1[911:904];
      img_out1[47:40] = img1[919:912];
      img_out1[55:48] = img1[927:920];
      img_out1[63:56] = img1[935:928];
      img_out1[71:64] = img1[943:936];
      img_out1[79:72] = img1[951:944];
      img_out1[87:80] = img1[959:952];
      img_out1[95:88] = img1[967:960];
      img_out1[103:96] = img1[975:968];
      img_out1[111:104] = img1[983:976];
      img_out1[119:112] = img1[991:984];
      img_out1[127:120] = img1[999:992];
      img_out1[135:128] = img1[1007:1000];
      img_out1[143:136] = img1[1015:1008];
      img_out1[151:144] = img1[1023:1016];
      img_out1[159:152] = img1[1031:1024];
      img_out1[167:160] = img1[1039:1032];
      img_out1[175:168] = img1[1047:1040];
      img_out2[7:0] = img2[879:872];
      img_out2[15:8] = img2[887:880];
      img_out2[23:16] = img2[895:888];
      img_out2[31:24] = img2[903:896];
      img_out2[39:32] = img2[911:904];
      img_out2[47:40] = img2[919:912];
      img_out2[55:48] = img2[927:920];
      img_out2[63:56] = img2[935:928];
      img_out2[71:64] = img2[943:936];
      img_out2[79:72] = img2[951:944];
      img_out2[87:80] = img2[959:952];
      img_out2[95:88] = img2[967:960];
      img_out2[103:96] = img2[975:968];
      img_out2[111:104] = img2[983:976];
      img_out2[119:112] = img2[991:984];
      img_out2[127:120] = img2[999:992];
      img_out2[135:128] = img2[1007:1000];
      img_out2[143:136] = img2[1015:1008];
      img_out2[151:144] = img2[1023:1016];
      img_out2[159:152] = img2[1031:1024];
      img_out2[167:160] = img2[1039:1032];
      img_out2[175:168] = img2[1047:1040];
      img_out3[7:0] = img3[879:872];
      img_out3[15:8] = img3[887:880];
      img_out3[23:16] = img3[895:888];
      img_out3[31:24] = img3[903:896];
      img_out3[39:32] = img3[911:904];
      img_out3[47:40] = img3[919:912];
      img_out3[55:48] = img3[927:920];
      img_out3[63:56] = img3[935:928];
      img_out3[71:64] = img3[943:936];
      img_out3[79:72] = img3[951:944];
      img_out3[87:80] = img3[959:952];
      img_out3[95:88] = img3[967:960];
      img_out3[103:96] = img3[975:968];
      img_out3[111:104] = img3[983:976];
      img_out3[119:112] = img3[991:984];
      img_out3[127:120] = img3[999:992];
      img_out3[135:128] = img3[1007:1000];
      img_out3[143:136] = img3[1015:1008];
      img_out3[151:144] = img3[1023:1016];
      img_out3[159:152] = img3[1031:1024];
      img_out3[167:160] = img3[1039:1032];
      img_out3[175:168] = img3[1047:1040];
      img_out4[7:0] = img4[879:872];
      img_out4[15:8] = img4[887:880];
      img_out4[23:16] = img4[895:888];
      img_out4[31:24] = img4[903:896];
      img_out4[39:32] = img4[911:904];
      img_out4[47:40] = img4[919:912];
      img_out4[55:48] = img4[927:920];
      img_out4[63:56] = img4[935:928];
      img_out4[71:64] = img4[943:936];
      img_out4[79:72] = img4[951:944];
      img_out4[87:80] = img4[959:952];
      img_out4[95:88] = img4[967:960];
      img_out4[103:96] = img4[975:968];
      img_out4[111:104] = img4[983:976];
      img_out4[119:112] = img4[991:984];
      img_out4[127:120] = img4[999:992];
      img_out4[135:128] = img4[1007:1000];
      img_out4[143:136] = img4[1015:1008];
      img_out4[151:144] = img4[1023:1016];
      img_out4[159:152] = img4[1031:1024];
      img_out4[167:160] = img4[1039:1032];
      img_out4[175:168] = img4[1047:1040];
    end
    'd8: begin
      img_out0[7:0] = img0[1007:1000];
      img_out0[15:8] = img0[1015:1008];
      img_out0[23:16] = img0[1023:1016];
      img_out0[31:24] = img0[1031:1024];
      img_out0[39:32] = img0[1039:1032];
      img_out0[47:40] = img0[1047:1040];
      img_out0[55:48] = img0[1055:1048];
      img_out0[63:56] = img0[1063:1056];
      img_out0[71:64] = img0[1071:1064];
      img_out0[79:72] = img0[1079:1072];
      img_out0[87:80] = img0[1087:1080];
      img_out0[95:88] = img0[1095:1088];
      img_out0[103:96] = img0[1103:1096];
      img_out0[111:104] = img0[1111:1104];
      img_out0[119:112] = img0[1119:1112];
      img_out0[127:120] = img0[1127:1120];
      img_out0[135:128] = img0[1135:1128];
      img_out0[143:136] = img0[1143:1136];
      img_out0[151:144] = img0[1151:1144];
      img_out0[159:152] = img0[1159:1152];
      img_out0[167:160] = img0[1167:1160];
      img_out0[175:168] = img0[1175:1168];
      img_out1[7:0] = img1[1007:1000];
      img_out1[15:8] = img1[1015:1008];
      img_out1[23:16] = img1[1023:1016];
      img_out1[31:24] = img1[1031:1024];
      img_out1[39:32] = img1[1039:1032];
      img_out1[47:40] = img1[1047:1040];
      img_out1[55:48] = img1[1055:1048];
      img_out1[63:56] = img1[1063:1056];
      img_out1[71:64] = img1[1071:1064];
      img_out1[79:72] = img1[1079:1072];
      img_out1[87:80] = img1[1087:1080];
      img_out1[95:88] = img1[1095:1088];
      img_out1[103:96] = img1[1103:1096];
      img_out1[111:104] = img1[1111:1104];
      img_out1[119:112] = img1[1119:1112];
      img_out1[127:120] = img1[1127:1120];
      img_out1[135:128] = img1[1135:1128];
      img_out1[143:136] = img1[1143:1136];
      img_out1[151:144] = img1[1151:1144];
      img_out1[159:152] = img1[1159:1152];
      img_out1[167:160] = img1[1167:1160];
      img_out1[175:168] = img1[1175:1168];
      img_out2[7:0] = img2[1007:1000];
      img_out2[15:8] = img2[1015:1008];
      img_out2[23:16] = img2[1023:1016];
      img_out2[31:24] = img2[1031:1024];
      img_out2[39:32] = img2[1039:1032];
      img_out2[47:40] = img2[1047:1040];
      img_out2[55:48] = img2[1055:1048];
      img_out2[63:56] = img2[1063:1056];
      img_out2[71:64] = img2[1071:1064];
      img_out2[79:72] = img2[1079:1072];
      img_out2[87:80] = img2[1087:1080];
      img_out2[95:88] = img2[1095:1088];
      img_out2[103:96] = img2[1103:1096];
      img_out2[111:104] = img2[1111:1104];
      img_out2[119:112] = img2[1119:1112];
      img_out2[127:120] = img2[1127:1120];
      img_out2[135:128] = img2[1135:1128];
      img_out2[143:136] = img2[1143:1136];
      img_out2[151:144] = img2[1151:1144];
      img_out2[159:152] = img2[1159:1152];
      img_out2[167:160] = img2[1167:1160];
      img_out2[175:168] = img2[1175:1168];
      img_out3[7:0] = img3[1007:1000];
      img_out3[15:8] = img3[1015:1008];
      img_out3[23:16] = img3[1023:1016];
      img_out3[31:24] = img3[1031:1024];
      img_out3[39:32] = img3[1039:1032];
      img_out3[47:40] = img3[1047:1040];
      img_out3[55:48] = img3[1055:1048];
      img_out3[63:56] = img3[1063:1056];
      img_out3[71:64] = img3[1071:1064];
      img_out3[79:72] = img3[1079:1072];
      img_out3[87:80] = img3[1087:1080];
      img_out3[95:88] = img3[1095:1088];
      img_out3[103:96] = img3[1103:1096];
      img_out3[111:104] = img3[1111:1104];
      img_out3[119:112] = img3[1119:1112];
      img_out3[127:120] = img3[1127:1120];
      img_out3[135:128] = img3[1135:1128];
      img_out3[143:136] = img3[1143:1136];
      img_out3[151:144] = img3[1151:1144];
      img_out3[159:152] = img3[1159:1152];
      img_out3[167:160] = img3[1167:1160];
      img_out3[175:168] = img3[1175:1168];
      img_out4[7:0] = img4[1007:1000];
      img_out4[15:8] = img4[1015:1008];
      img_out4[23:16] = img4[1023:1016];
      img_out4[31:24] = img4[1031:1024];
      img_out4[39:32] = img4[1039:1032];
      img_out4[47:40] = img4[1047:1040];
      img_out4[55:48] = img4[1055:1048];
      img_out4[63:56] = img4[1063:1056];
      img_out4[71:64] = img4[1071:1064];
      img_out4[79:72] = img4[1079:1072];
      img_out4[87:80] = img4[1087:1080];
      img_out4[95:88] = img4[1095:1088];
      img_out4[103:96] = img4[1103:1096];
      img_out4[111:104] = img4[1111:1104];
      img_out4[119:112] = img4[1119:1112];
      img_out4[127:120] = img4[1127:1120];
      img_out4[135:128] = img4[1135:1128];
      img_out4[143:136] = img4[1143:1136];
      img_out4[151:144] = img4[1151:1144];
      img_out4[159:152] = img4[1159:1152];
      img_out4[167:160] = img4[1167:1160];
      img_out4[175:168] = img4[1175:1168];
    end
    'd9: begin
      img_out0[7:0] = img0[1135:1128];
      img_out0[15:8] = img0[1143:1136];
      img_out0[23:16] = img0[1151:1144];
      img_out0[31:24] = img0[1159:1152];
      img_out0[39:32] = img0[1167:1160];
      img_out0[47:40] = img0[1175:1168];
      img_out0[55:48] = img0[1183:1176];
      img_out0[63:56] = img0[1191:1184];
      img_out0[71:64] = img0[1199:1192];
      img_out0[79:72] = img0[1207:1200];
      img_out0[87:80] = img0[1215:1208];
      img_out0[95:88] = img0[1223:1216];
      img_out0[103:96] = img0[1231:1224];
      img_out0[111:104] = img0[1239:1232];
      img_out0[119:112] = img0[1247:1240];
      img_out0[127:120] = img0[1255:1248];
      img_out0[135:128] = img0[1263:1256];
      img_out0[143:136] = img0[1271:1264];
      img_out0[151:144] = img0[1279:1272];
      img_out0[159:152] = img0[1287:1280];
      img_out0[167:160] = img0[1295:1288];
      img_out0[175:168] = img0[1303:1296];
      img_out1[7:0] = img1[1135:1128];
      img_out1[15:8] = img1[1143:1136];
      img_out1[23:16] = img1[1151:1144];
      img_out1[31:24] = img1[1159:1152];
      img_out1[39:32] = img1[1167:1160];
      img_out1[47:40] = img1[1175:1168];
      img_out1[55:48] = img1[1183:1176];
      img_out1[63:56] = img1[1191:1184];
      img_out1[71:64] = img1[1199:1192];
      img_out1[79:72] = img1[1207:1200];
      img_out1[87:80] = img1[1215:1208];
      img_out1[95:88] = img1[1223:1216];
      img_out1[103:96] = img1[1231:1224];
      img_out1[111:104] = img1[1239:1232];
      img_out1[119:112] = img1[1247:1240];
      img_out1[127:120] = img1[1255:1248];
      img_out1[135:128] = img1[1263:1256];
      img_out1[143:136] = img1[1271:1264];
      img_out1[151:144] = img1[1279:1272];
      img_out1[159:152] = img1[1287:1280];
      img_out1[167:160] = img1[1295:1288];
      img_out1[175:168] = img1[1303:1296];
      img_out2[7:0] = img2[1135:1128];
      img_out2[15:8] = img2[1143:1136];
      img_out2[23:16] = img2[1151:1144];
      img_out2[31:24] = img2[1159:1152];
      img_out2[39:32] = img2[1167:1160];
      img_out2[47:40] = img2[1175:1168];
      img_out2[55:48] = img2[1183:1176];
      img_out2[63:56] = img2[1191:1184];
      img_out2[71:64] = img2[1199:1192];
      img_out2[79:72] = img2[1207:1200];
      img_out2[87:80] = img2[1215:1208];
      img_out2[95:88] = img2[1223:1216];
      img_out2[103:96] = img2[1231:1224];
      img_out2[111:104] = img2[1239:1232];
      img_out2[119:112] = img2[1247:1240];
      img_out2[127:120] = img2[1255:1248];
      img_out2[135:128] = img2[1263:1256];
      img_out2[143:136] = img2[1271:1264];
      img_out2[151:144] = img2[1279:1272];
      img_out2[159:152] = img2[1287:1280];
      img_out2[167:160] = img2[1295:1288];
      img_out2[175:168] = img2[1303:1296];
      img_out3[7:0] = img3[1135:1128];
      img_out3[15:8] = img3[1143:1136];
      img_out3[23:16] = img3[1151:1144];
      img_out3[31:24] = img3[1159:1152];
      img_out3[39:32] = img3[1167:1160];
      img_out3[47:40] = img3[1175:1168];
      img_out3[55:48] = img3[1183:1176];
      img_out3[63:56] = img3[1191:1184];
      img_out3[71:64] = img3[1199:1192];
      img_out3[79:72] = img3[1207:1200];
      img_out3[87:80] = img3[1215:1208];
      img_out3[95:88] = img3[1223:1216];
      img_out3[103:96] = img3[1231:1224];
      img_out3[111:104] = img3[1239:1232];
      img_out3[119:112] = img3[1247:1240];
      img_out3[127:120] = img3[1255:1248];
      img_out3[135:128] = img3[1263:1256];
      img_out3[143:136] = img3[1271:1264];
      img_out3[151:144] = img3[1279:1272];
      img_out3[159:152] = img3[1287:1280];
      img_out3[167:160] = img3[1295:1288];
      img_out3[175:168] = img3[1303:1296];
      img_out4[7:0] = img4[1135:1128];
      img_out4[15:8] = img4[1143:1136];
      img_out4[23:16] = img4[1151:1144];
      img_out4[31:24] = img4[1159:1152];
      img_out4[39:32] = img4[1167:1160];
      img_out4[47:40] = img4[1175:1168];
      img_out4[55:48] = img4[1183:1176];
      img_out4[63:56] = img4[1191:1184];
      img_out4[71:64] = img4[1199:1192];
      img_out4[79:72] = img4[1207:1200];
      img_out4[87:80] = img4[1215:1208];
      img_out4[95:88] = img4[1223:1216];
      img_out4[103:96] = img4[1231:1224];
      img_out4[111:104] = img4[1239:1232];
      img_out4[119:112] = img4[1247:1240];
      img_out4[127:120] = img4[1255:1248];
      img_out4[135:128] = img4[1263:1256];
      img_out4[143:136] = img4[1271:1264];
      img_out4[151:144] = img4[1279:1272];
      img_out4[159:152] = img4[1287:1280];
      img_out4[167:160] = img4[1295:1288];
      img_out4[175:168] = img4[1303:1296];
    end
    'd10: begin
      img_out0[7:0] = img0[1263:1256];
      img_out0[15:8] = img0[1271:1264];
      img_out0[23:16] = img0[1279:1272];
      img_out0[31:24] = img0[1287:1280];
      img_out0[39:32] = img0[1295:1288];
      img_out0[47:40] = img0[1303:1296];
      img_out0[55:48] = img0[1311:1304];
      img_out0[63:56] = img0[1319:1312];
      img_out0[71:64] = img0[1327:1320];
      img_out0[79:72] = img0[1335:1328];
      img_out0[87:80] = img0[1343:1336];
      img_out0[95:88] = img0[1351:1344];
      img_out0[103:96] = img0[1359:1352];
      img_out0[111:104] = img0[1367:1360];
      img_out0[119:112] = img0[1375:1368];
      img_out0[127:120] = img0[1383:1376];
      img_out0[135:128] = img0[1391:1384];
      img_out0[143:136] = img0[1399:1392];
      img_out0[151:144] = img0[1407:1400];
      img_out0[159:152] = img0[1415:1408];
      img_out0[167:160] = img0[1423:1416];
      img_out0[175:168] = img0[1431:1424];
      img_out1[7:0] = img1[1263:1256];
      img_out1[15:8] = img1[1271:1264];
      img_out1[23:16] = img1[1279:1272];
      img_out1[31:24] = img1[1287:1280];
      img_out1[39:32] = img1[1295:1288];
      img_out1[47:40] = img1[1303:1296];
      img_out1[55:48] = img1[1311:1304];
      img_out1[63:56] = img1[1319:1312];
      img_out1[71:64] = img1[1327:1320];
      img_out1[79:72] = img1[1335:1328];
      img_out1[87:80] = img1[1343:1336];
      img_out1[95:88] = img1[1351:1344];
      img_out1[103:96] = img1[1359:1352];
      img_out1[111:104] = img1[1367:1360];
      img_out1[119:112] = img1[1375:1368];
      img_out1[127:120] = img1[1383:1376];
      img_out1[135:128] = img1[1391:1384];
      img_out1[143:136] = img1[1399:1392];
      img_out1[151:144] = img1[1407:1400];
      img_out1[159:152] = img1[1415:1408];
      img_out1[167:160] = img1[1423:1416];
      img_out1[175:168] = img1[1431:1424];
      img_out2[7:0] = img2[1263:1256];
      img_out2[15:8] = img2[1271:1264];
      img_out2[23:16] = img2[1279:1272];
      img_out2[31:24] = img2[1287:1280];
      img_out2[39:32] = img2[1295:1288];
      img_out2[47:40] = img2[1303:1296];
      img_out2[55:48] = img2[1311:1304];
      img_out2[63:56] = img2[1319:1312];
      img_out2[71:64] = img2[1327:1320];
      img_out2[79:72] = img2[1335:1328];
      img_out2[87:80] = img2[1343:1336];
      img_out2[95:88] = img2[1351:1344];
      img_out2[103:96] = img2[1359:1352];
      img_out2[111:104] = img2[1367:1360];
      img_out2[119:112] = img2[1375:1368];
      img_out2[127:120] = img2[1383:1376];
      img_out2[135:128] = img2[1391:1384];
      img_out2[143:136] = img2[1399:1392];
      img_out2[151:144] = img2[1407:1400];
      img_out2[159:152] = img2[1415:1408];
      img_out2[167:160] = img2[1423:1416];
      img_out2[175:168] = img2[1431:1424];
      img_out3[7:0] = img3[1263:1256];
      img_out3[15:8] = img3[1271:1264];
      img_out3[23:16] = img3[1279:1272];
      img_out3[31:24] = img3[1287:1280];
      img_out3[39:32] = img3[1295:1288];
      img_out3[47:40] = img3[1303:1296];
      img_out3[55:48] = img3[1311:1304];
      img_out3[63:56] = img3[1319:1312];
      img_out3[71:64] = img3[1327:1320];
      img_out3[79:72] = img3[1335:1328];
      img_out3[87:80] = img3[1343:1336];
      img_out3[95:88] = img3[1351:1344];
      img_out3[103:96] = img3[1359:1352];
      img_out3[111:104] = img3[1367:1360];
      img_out3[119:112] = img3[1375:1368];
      img_out3[127:120] = img3[1383:1376];
      img_out3[135:128] = img3[1391:1384];
      img_out3[143:136] = img3[1399:1392];
      img_out3[151:144] = img3[1407:1400];
      img_out3[159:152] = img3[1415:1408];
      img_out3[167:160] = img3[1423:1416];
      img_out3[175:168] = img3[1431:1424];
      img_out4[7:0] = img4[1263:1256];
      img_out4[15:8] = img4[1271:1264];
      img_out4[23:16] = img4[1279:1272];
      img_out4[31:24] = img4[1287:1280];
      img_out4[39:32] = img4[1295:1288];
      img_out4[47:40] = img4[1303:1296];
      img_out4[55:48] = img4[1311:1304];
      img_out4[63:56] = img4[1319:1312];
      img_out4[71:64] = img4[1327:1320];
      img_out4[79:72] = img4[1335:1328];
      img_out4[87:80] = img4[1343:1336];
      img_out4[95:88] = img4[1351:1344];
      img_out4[103:96] = img4[1359:1352];
      img_out4[111:104] = img4[1367:1360];
      img_out4[119:112] = img4[1375:1368];
      img_out4[127:120] = img4[1383:1376];
      img_out4[135:128] = img4[1391:1384];
      img_out4[143:136] = img4[1399:1392];
      img_out4[151:144] = img4[1407:1400];
      img_out4[159:152] = img4[1415:1408];
      img_out4[167:160] = img4[1423:1416];
      img_out4[175:168] = img4[1431:1424];
    end
    'd11: begin
      img_out0[7:0] = img0[1391:1384];
      img_out0[15:8] = img0[1399:1392];
      img_out0[23:16] = img0[1407:1400];
      img_out0[31:24] = img0[1415:1408];
      img_out0[39:32] = img0[1423:1416];
      img_out0[47:40] = img0[1431:1424];
      img_out0[55:48] = img0[1439:1432];
      img_out0[63:56] = img0[1447:1440];
      img_out0[71:64] = img0[1455:1448];
      img_out0[79:72] = img0[1463:1456];
      img_out0[87:80] = img0[1471:1464];
      img_out0[95:88] = img0[1479:1472];
      img_out0[103:96] = img0[1487:1480];
      img_out0[111:104] = img0[1495:1488];
      img_out0[119:112] = img0[1503:1496];
      img_out0[127:120] = img0[1511:1504];
      img_out0[135:128] = img0[1519:1512];
      img_out0[143:136] = img0[1527:1520];
      img_out0[151:144] = img0[1535:1528];
      img_out0[159:152] = img0[1543:1536];
      img_out0[167:160] = img0[1551:1544];
      img_out0[175:168] = img0[1559:1552];
      img_out1[7:0] = img1[1391:1384];
      img_out1[15:8] = img1[1399:1392];
      img_out1[23:16] = img1[1407:1400];
      img_out1[31:24] = img1[1415:1408];
      img_out1[39:32] = img1[1423:1416];
      img_out1[47:40] = img1[1431:1424];
      img_out1[55:48] = img1[1439:1432];
      img_out1[63:56] = img1[1447:1440];
      img_out1[71:64] = img1[1455:1448];
      img_out1[79:72] = img1[1463:1456];
      img_out1[87:80] = img1[1471:1464];
      img_out1[95:88] = img1[1479:1472];
      img_out1[103:96] = img1[1487:1480];
      img_out1[111:104] = img1[1495:1488];
      img_out1[119:112] = img1[1503:1496];
      img_out1[127:120] = img1[1511:1504];
      img_out1[135:128] = img1[1519:1512];
      img_out1[143:136] = img1[1527:1520];
      img_out1[151:144] = img1[1535:1528];
      img_out1[159:152] = img1[1543:1536];
      img_out1[167:160] = img1[1551:1544];
      img_out1[175:168] = img1[1559:1552];
      img_out2[7:0] = img2[1391:1384];
      img_out2[15:8] = img2[1399:1392];
      img_out2[23:16] = img2[1407:1400];
      img_out2[31:24] = img2[1415:1408];
      img_out2[39:32] = img2[1423:1416];
      img_out2[47:40] = img2[1431:1424];
      img_out2[55:48] = img2[1439:1432];
      img_out2[63:56] = img2[1447:1440];
      img_out2[71:64] = img2[1455:1448];
      img_out2[79:72] = img2[1463:1456];
      img_out2[87:80] = img2[1471:1464];
      img_out2[95:88] = img2[1479:1472];
      img_out2[103:96] = img2[1487:1480];
      img_out2[111:104] = img2[1495:1488];
      img_out2[119:112] = img2[1503:1496];
      img_out2[127:120] = img2[1511:1504];
      img_out2[135:128] = img2[1519:1512];
      img_out2[143:136] = img2[1527:1520];
      img_out2[151:144] = img2[1535:1528];
      img_out2[159:152] = img2[1543:1536];
      img_out2[167:160] = img2[1551:1544];
      img_out2[175:168] = img2[1559:1552];
      img_out3[7:0] = img3[1391:1384];
      img_out3[15:8] = img3[1399:1392];
      img_out3[23:16] = img3[1407:1400];
      img_out3[31:24] = img3[1415:1408];
      img_out3[39:32] = img3[1423:1416];
      img_out3[47:40] = img3[1431:1424];
      img_out3[55:48] = img3[1439:1432];
      img_out3[63:56] = img3[1447:1440];
      img_out3[71:64] = img3[1455:1448];
      img_out3[79:72] = img3[1463:1456];
      img_out3[87:80] = img3[1471:1464];
      img_out3[95:88] = img3[1479:1472];
      img_out3[103:96] = img3[1487:1480];
      img_out3[111:104] = img3[1495:1488];
      img_out3[119:112] = img3[1503:1496];
      img_out3[127:120] = img3[1511:1504];
      img_out3[135:128] = img3[1519:1512];
      img_out3[143:136] = img3[1527:1520];
      img_out3[151:144] = img3[1535:1528];
      img_out3[159:152] = img3[1543:1536];
      img_out3[167:160] = img3[1551:1544];
      img_out3[175:168] = img3[1559:1552];
      img_out4[7:0] = img4[1391:1384];
      img_out4[15:8] = img4[1399:1392];
      img_out4[23:16] = img4[1407:1400];
      img_out4[31:24] = img4[1415:1408];
      img_out4[39:32] = img4[1423:1416];
      img_out4[47:40] = img4[1431:1424];
      img_out4[55:48] = img4[1439:1432];
      img_out4[63:56] = img4[1447:1440];
      img_out4[71:64] = img4[1455:1448];
      img_out4[79:72] = img4[1463:1456];
      img_out4[87:80] = img4[1471:1464];
      img_out4[95:88] = img4[1479:1472];
      img_out4[103:96] = img4[1487:1480];
      img_out4[111:104] = img4[1495:1488];
      img_out4[119:112] = img4[1503:1496];
      img_out4[127:120] = img4[1511:1504];
      img_out4[135:128] = img4[1519:1512];
      img_out4[143:136] = img4[1527:1520];
      img_out4[151:144] = img4[1535:1528];
      img_out4[159:152] = img4[1543:1536];
      img_out4[167:160] = img4[1551:1544];
      img_out4[175:168] = img4[1559:1552];
    end
    'd12: begin
      img_out0[7:0] = img0[1519:1512];
      img_out0[15:8] = img0[1527:1520];
      img_out0[23:16] = img0[1535:1528];
      img_out0[31:24] = img0[1543:1536];
      img_out0[39:32] = img0[1551:1544];
      img_out0[47:40] = img0[1559:1552];
      img_out0[55:48] = img0[1567:1560];
      img_out0[63:56] = img0[1575:1568];
      img_out0[71:64] = img0[1583:1576];
      img_out0[79:72] = img0[1591:1584];
      img_out0[87:80] = img0[1599:1592];
      img_out0[95:88] = img0[1607:1600];
      img_out0[103:96] = img0[1615:1608];
      img_out0[111:104] = img0[1623:1616];
      img_out0[119:112] = img0[1631:1624];
      img_out0[127:120] = img0[1639:1632];
      img_out0[135:128] = img0[1647:1640];
      img_out0[143:136] = img0[1655:1648];
      img_out0[151:144] = img0[1663:1656];
      img_out0[159:152] = img0[1671:1664];
      img_out0[167:160] = img0[1679:1672];
      img_out0[175:168] = img0[1687:1680];
      img_out1[7:0] = img1[1519:1512];
      img_out1[15:8] = img1[1527:1520];
      img_out1[23:16] = img1[1535:1528];
      img_out1[31:24] = img1[1543:1536];
      img_out1[39:32] = img1[1551:1544];
      img_out1[47:40] = img1[1559:1552];
      img_out1[55:48] = img1[1567:1560];
      img_out1[63:56] = img1[1575:1568];
      img_out1[71:64] = img1[1583:1576];
      img_out1[79:72] = img1[1591:1584];
      img_out1[87:80] = img1[1599:1592];
      img_out1[95:88] = img1[1607:1600];
      img_out1[103:96] = img1[1615:1608];
      img_out1[111:104] = img1[1623:1616];
      img_out1[119:112] = img1[1631:1624];
      img_out1[127:120] = img1[1639:1632];
      img_out1[135:128] = img1[1647:1640];
      img_out1[143:136] = img1[1655:1648];
      img_out1[151:144] = img1[1663:1656];
      img_out1[159:152] = img1[1671:1664];
      img_out1[167:160] = img1[1679:1672];
      img_out1[175:168] = img1[1687:1680];
      img_out2[7:0] = img2[1519:1512];
      img_out2[15:8] = img2[1527:1520];
      img_out2[23:16] = img2[1535:1528];
      img_out2[31:24] = img2[1543:1536];
      img_out2[39:32] = img2[1551:1544];
      img_out2[47:40] = img2[1559:1552];
      img_out2[55:48] = img2[1567:1560];
      img_out2[63:56] = img2[1575:1568];
      img_out2[71:64] = img2[1583:1576];
      img_out2[79:72] = img2[1591:1584];
      img_out2[87:80] = img2[1599:1592];
      img_out2[95:88] = img2[1607:1600];
      img_out2[103:96] = img2[1615:1608];
      img_out2[111:104] = img2[1623:1616];
      img_out2[119:112] = img2[1631:1624];
      img_out2[127:120] = img2[1639:1632];
      img_out2[135:128] = img2[1647:1640];
      img_out2[143:136] = img2[1655:1648];
      img_out2[151:144] = img2[1663:1656];
      img_out2[159:152] = img2[1671:1664];
      img_out2[167:160] = img2[1679:1672];
      img_out2[175:168] = img2[1687:1680];
      img_out3[7:0] = img3[1519:1512];
      img_out3[15:8] = img3[1527:1520];
      img_out3[23:16] = img3[1535:1528];
      img_out3[31:24] = img3[1543:1536];
      img_out3[39:32] = img3[1551:1544];
      img_out3[47:40] = img3[1559:1552];
      img_out3[55:48] = img3[1567:1560];
      img_out3[63:56] = img3[1575:1568];
      img_out3[71:64] = img3[1583:1576];
      img_out3[79:72] = img3[1591:1584];
      img_out3[87:80] = img3[1599:1592];
      img_out3[95:88] = img3[1607:1600];
      img_out3[103:96] = img3[1615:1608];
      img_out3[111:104] = img3[1623:1616];
      img_out3[119:112] = img3[1631:1624];
      img_out3[127:120] = img3[1639:1632];
      img_out3[135:128] = img3[1647:1640];
      img_out3[143:136] = img3[1655:1648];
      img_out3[151:144] = img3[1663:1656];
      img_out3[159:152] = img3[1671:1664];
      img_out3[167:160] = img3[1679:1672];
      img_out3[175:168] = img3[1687:1680];
      img_out4[7:0] = img4[1519:1512];
      img_out4[15:8] = img4[1527:1520];
      img_out4[23:16] = img4[1535:1528];
      img_out4[31:24] = img4[1543:1536];
      img_out4[39:32] = img4[1551:1544];
      img_out4[47:40] = img4[1559:1552];
      img_out4[55:48] = img4[1567:1560];
      img_out4[63:56] = img4[1575:1568];
      img_out4[71:64] = img4[1583:1576];
      img_out4[79:72] = img4[1591:1584];
      img_out4[87:80] = img4[1599:1592];
      img_out4[95:88] = img4[1607:1600];
      img_out4[103:96] = img4[1615:1608];
      img_out4[111:104] = img4[1623:1616];
      img_out4[119:112] = img4[1631:1624];
      img_out4[127:120] = img4[1639:1632];
      img_out4[135:128] = img4[1647:1640];
      img_out4[143:136] = img4[1655:1648];
      img_out4[151:144] = img4[1663:1656];
      img_out4[159:152] = img4[1671:1664];
      img_out4[167:160] = img4[1679:1672];
      img_out4[175:168] = img4[1687:1680];
    end
    'd13: begin
      img_out0[7:0] = img0[1647:1640];
      img_out0[15:8] = img0[1655:1648];
      img_out0[23:16] = img0[1663:1656];
      img_out0[31:24] = img0[1671:1664];
      img_out0[39:32] = img0[1679:1672];
      img_out0[47:40] = img0[1687:1680];
      img_out0[55:48] = img0[1695:1688];
      img_out0[63:56] = img0[1703:1696];
      img_out0[71:64] = img0[1711:1704];
      img_out0[79:72] = img0[1719:1712];
      img_out0[87:80] = img0[1727:1720];
      img_out0[95:88] = img0[1735:1728];
      img_out0[103:96] = img0[1743:1736];
      img_out0[111:104] = img0[1751:1744];
      img_out0[119:112] = img0[1759:1752];
      img_out0[127:120] = img0[1767:1760];
      img_out0[135:128] = img0[1775:1768];
      img_out0[143:136] = img0[1783:1776];
      img_out0[151:144] = img0[1791:1784];
      img_out0[159:152] = img0[1799:1792];
      img_out0[167:160] = img0[1807:1800];
      img_out0[175:168] = img0[1815:1808];
      img_out1[7:0] = img1[1647:1640];
      img_out1[15:8] = img1[1655:1648];
      img_out1[23:16] = img1[1663:1656];
      img_out1[31:24] = img1[1671:1664];
      img_out1[39:32] = img1[1679:1672];
      img_out1[47:40] = img1[1687:1680];
      img_out1[55:48] = img1[1695:1688];
      img_out1[63:56] = img1[1703:1696];
      img_out1[71:64] = img1[1711:1704];
      img_out1[79:72] = img1[1719:1712];
      img_out1[87:80] = img1[1727:1720];
      img_out1[95:88] = img1[1735:1728];
      img_out1[103:96] = img1[1743:1736];
      img_out1[111:104] = img1[1751:1744];
      img_out1[119:112] = img1[1759:1752];
      img_out1[127:120] = img1[1767:1760];
      img_out1[135:128] = img1[1775:1768];
      img_out1[143:136] = img1[1783:1776];
      img_out1[151:144] = img1[1791:1784];
      img_out1[159:152] = img1[1799:1792];
      img_out1[167:160] = img1[1807:1800];
      img_out1[175:168] = img1[1815:1808];
      img_out2[7:0] = img2[1647:1640];
      img_out2[15:8] = img2[1655:1648];
      img_out2[23:16] = img2[1663:1656];
      img_out2[31:24] = img2[1671:1664];
      img_out2[39:32] = img2[1679:1672];
      img_out2[47:40] = img2[1687:1680];
      img_out2[55:48] = img2[1695:1688];
      img_out2[63:56] = img2[1703:1696];
      img_out2[71:64] = img2[1711:1704];
      img_out2[79:72] = img2[1719:1712];
      img_out2[87:80] = img2[1727:1720];
      img_out2[95:88] = img2[1735:1728];
      img_out2[103:96] = img2[1743:1736];
      img_out2[111:104] = img2[1751:1744];
      img_out2[119:112] = img2[1759:1752];
      img_out2[127:120] = img2[1767:1760];
      img_out2[135:128] = img2[1775:1768];
      img_out2[143:136] = img2[1783:1776];
      img_out2[151:144] = img2[1791:1784];
      img_out2[159:152] = img2[1799:1792];
      img_out2[167:160] = img2[1807:1800];
      img_out2[175:168] = img2[1815:1808];
      img_out3[7:0] = img3[1647:1640];
      img_out3[15:8] = img3[1655:1648];
      img_out3[23:16] = img3[1663:1656];
      img_out3[31:24] = img3[1671:1664];
      img_out3[39:32] = img3[1679:1672];
      img_out3[47:40] = img3[1687:1680];
      img_out3[55:48] = img3[1695:1688];
      img_out3[63:56] = img3[1703:1696];
      img_out3[71:64] = img3[1711:1704];
      img_out3[79:72] = img3[1719:1712];
      img_out3[87:80] = img3[1727:1720];
      img_out3[95:88] = img3[1735:1728];
      img_out3[103:96] = img3[1743:1736];
      img_out3[111:104] = img3[1751:1744];
      img_out3[119:112] = img3[1759:1752];
      img_out3[127:120] = img3[1767:1760];
      img_out3[135:128] = img3[1775:1768];
      img_out3[143:136] = img3[1783:1776];
      img_out3[151:144] = img3[1791:1784];
      img_out3[159:152] = img3[1799:1792];
      img_out3[167:160] = img3[1807:1800];
      img_out3[175:168] = img3[1815:1808];
      img_out4[7:0] = img4[1647:1640];
      img_out4[15:8] = img4[1655:1648];
      img_out4[23:16] = img4[1663:1656];
      img_out4[31:24] = img4[1671:1664];
      img_out4[39:32] = img4[1679:1672];
      img_out4[47:40] = img4[1687:1680];
      img_out4[55:48] = img4[1695:1688];
      img_out4[63:56] = img4[1703:1696];
      img_out4[71:64] = img4[1711:1704];
      img_out4[79:72] = img4[1719:1712];
      img_out4[87:80] = img4[1727:1720];
      img_out4[95:88] = img4[1735:1728];
      img_out4[103:96] = img4[1743:1736];
      img_out4[111:104] = img4[1751:1744];
      img_out4[119:112] = img4[1759:1752];
      img_out4[127:120] = img4[1767:1760];
      img_out4[135:128] = img4[1775:1768];
      img_out4[143:136] = img4[1783:1776];
      img_out4[151:144] = img4[1791:1784];
      img_out4[159:152] = img4[1799:1792];
      img_out4[167:160] = img4[1807:1800];
      img_out4[175:168] = img4[1815:1808];
    end
    'd14: begin
      img_out0[7:0] = img0[1775:1768];
      img_out0[15:8] = img0[1783:1776];
      img_out0[23:16] = img0[1791:1784];
      img_out0[31:24] = img0[1799:1792];
      img_out0[39:32] = img0[1807:1800];
      img_out0[47:40] = img0[1815:1808];
      img_out0[55:48] = img0[1823:1816];
      img_out0[63:56] = img0[1831:1824];
      img_out0[71:64] = img0[1839:1832];
      img_out0[79:72] = img0[1847:1840];
      img_out0[87:80] = img0[1855:1848];
      img_out0[95:88] = img0[1863:1856];
      img_out0[103:96] = img0[1871:1864];
      img_out0[111:104] = img0[1879:1872];
      img_out0[119:112] = img0[1887:1880];
      img_out0[127:120] = img0[1895:1888];
      img_out0[135:128] = img0[1903:1896];
      img_out0[143:136] = img0[1911:1904];
      img_out0[151:144] = img0[1919:1912];
      img_out0[159:152] = img0[1927:1920];
      img_out0[167:160] = img0[1935:1928];
      img_out0[175:168] = img0[1943:1936];
      img_out1[7:0] = img1[1775:1768];
      img_out1[15:8] = img1[1783:1776];
      img_out1[23:16] = img1[1791:1784];
      img_out1[31:24] = img1[1799:1792];
      img_out1[39:32] = img1[1807:1800];
      img_out1[47:40] = img1[1815:1808];
      img_out1[55:48] = img1[1823:1816];
      img_out1[63:56] = img1[1831:1824];
      img_out1[71:64] = img1[1839:1832];
      img_out1[79:72] = img1[1847:1840];
      img_out1[87:80] = img1[1855:1848];
      img_out1[95:88] = img1[1863:1856];
      img_out1[103:96] = img1[1871:1864];
      img_out1[111:104] = img1[1879:1872];
      img_out1[119:112] = img1[1887:1880];
      img_out1[127:120] = img1[1895:1888];
      img_out1[135:128] = img1[1903:1896];
      img_out1[143:136] = img1[1911:1904];
      img_out1[151:144] = img1[1919:1912];
      img_out1[159:152] = img1[1927:1920];
      img_out1[167:160] = img1[1935:1928];
      img_out1[175:168] = img1[1943:1936];
      img_out2[7:0] = img2[1775:1768];
      img_out2[15:8] = img2[1783:1776];
      img_out2[23:16] = img2[1791:1784];
      img_out2[31:24] = img2[1799:1792];
      img_out2[39:32] = img2[1807:1800];
      img_out2[47:40] = img2[1815:1808];
      img_out2[55:48] = img2[1823:1816];
      img_out2[63:56] = img2[1831:1824];
      img_out2[71:64] = img2[1839:1832];
      img_out2[79:72] = img2[1847:1840];
      img_out2[87:80] = img2[1855:1848];
      img_out2[95:88] = img2[1863:1856];
      img_out2[103:96] = img2[1871:1864];
      img_out2[111:104] = img2[1879:1872];
      img_out2[119:112] = img2[1887:1880];
      img_out2[127:120] = img2[1895:1888];
      img_out2[135:128] = img2[1903:1896];
      img_out2[143:136] = img2[1911:1904];
      img_out2[151:144] = img2[1919:1912];
      img_out2[159:152] = img2[1927:1920];
      img_out2[167:160] = img2[1935:1928];
      img_out2[175:168] = img2[1943:1936];
      img_out3[7:0] = img3[1775:1768];
      img_out3[15:8] = img3[1783:1776];
      img_out3[23:16] = img3[1791:1784];
      img_out3[31:24] = img3[1799:1792];
      img_out3[39:32] = img3[1807:1800];
      img_out3[47:40] = img3[1815:1808];
      img_out3[55:48] = img3[1823:1816];
      img_out3[63:56] = img3[1831:1824];
      img_out3[71:64] = img3[1839:1832];
      img_out3[79:72] = img3[1847:1840];
      img_out3[87:80] = img3[1855:1848];
      img_out3[95:88] = img3[1863:1856];
      img_out3[103:96] = img3[1871:1864];
      img_out3[111:104] = img3[1879:1872];
      img_out3[119:112] = img3[1887:1880];
      img_out3[127:120] = img3[1895:1888];
      img_out3[135:128] = img3[1903:1896];
      img_out3[143:136] = img3[1911:1904];
      img_out3[151:144] = img3[1919:1912];
      img_out3[159:152] = img3[1927:1920];
      img_out3[167:160] = img3[1935:1928];
      img_out3[175:168] = img3[1943:1936];
      img_out4[7:0] = img4[1775:1768];
      img_out4[15:8] = img4[1783:1776];
      img_out4[23:16] = img4[1791:1784];
      img_out4[31:24] = img4[1799:1792];
      img_out4[39:32] = img4[1807:1800];
      img_out4[47:40] = img4[1815:1808];
      img_out4[55:48] = img4[1823:1816];
      img_out4[63:56] = img4[1831:1824];
      img_out4[71:64] = img4[1839:1832];
      img_out4[79:72] = img4[1847:1840];
      img_out4[87:80] = img4[1855:1848];
      img_out4[95:88] = img4[1863:1856];
      img_out4[103:96] = img4[1871:1864];
      img_out4[111:104] = img4[1879:1872];
      img_out4[119:112] = img4[1887:1880];
      img_out4[127:120] = img4[1895:1888];
      img_out4[135:128] = img4[1903:1896];
      img_out4[143:136] = img4[1911:1904];
      img_out4[151:144] = img4[1919:1912];
      img_out4[159:152] = img4[1927:1920];
      img_out4[167:160] = img4[1935:1928];
      img_out4[175:168] = img4[1943:1936];
    end
    'd15: begin
      img_out0[7:0] = img0[1903:1896];
      img_out0[15:8] = img0[1911:1904];
      img_out0[23:16] = img0[1919:1912];
      img_out0[31:24] = img0[1927:1920];
      img_out0[39:32] = img0[1935:1928];
      img_out0[47:40] = img0[1943:1936];
      img_out0[55:48] = img0[1951:1944];
      img_out0[63:56] = img0[1959:1952];
      img_out0[71:64] = img0[1967:1960];
      img_out0[79:72] = img0[1975:1968];
      img_out0[87:80] = img0[1983:1976];
      img_out0[95:88] = img0[1991:1984];
      img_out0[103:96] = img0[1999:1992];
      img_out0[111:104] = img0[2007:2000];
      img_out0[119:112] = img0[2015:2008];
      img_out0[127:120] = img0[2023:2016];
      img_out0[135:128] = img0[2031:2024];
      img_out0[143:136] = img0[2039:2032];
      img_out0[151:144] = img0[2047:2040];
      img_out0[159:152] = img0[2055:2048];
      img_out0[167:160] = img0[2063:2056];
      img_out0[175:168] = img0[2071:2064];
      img_out1[7:0] = img1[1903:1896];
      img_out1[15:8] = img1[1911:1904];
      img_out1[23:16] = img1[1919:1912];
      img_out1[31:24] = img1[1927:1920];
      img_out1[39:32] = img1[1935:1928];
      img_out1[47:40] = img1[1943:1936];
      img_out1[55:48] = img1[1951:1944];
      img_out1[63:56] = img1[1959:1952];
      img_out1[71:64] = img1[1967:1960];
      img_out1[79:72] = img1[1975:1968];
      img_out1[87:80] = img1[1983:1976];
      img_out1[95:88] = img1[1991:1984];
      img_out1[103:96] = img1[1999:1992];
      img_out1[111:104] = img1[2007:2000];
      img_out1[119:112] = img1[2015:2008];
      img_out1[127:120] = img1[2023:2016];
      img_out1[135:128] = img1[2031:2024];
      img_out1[143:136] = img1[2039:2032];
      img_out1[151:144] = img1[2047:2040];
      img_out1[159:152] = img1[2055:2048];
      img_out1[167:160] = img1[2063:2056];
      img_out1[175:168] = img1[2071:2064];
      img_out2[7:0] = img2[1903:1896];
      img_out2[15:8] = img2[1911:1904];
      img_out2[23:16] = img2[1919:1912];
      img_out2[31:24] = img2[1927:1920];
      img_out2[39:32] = img2[1935:1928];
      img_out2[47:40] = img2[1943:1936];
      img_out2[55:48] = img2[1951:1944];
      img_out2[63:56] = img2[1959:1952];
      img_out2[71:64] = img2[1967:1960];
      img_out2[79:72] = img2[1975:1968];
      img_out2[87:80] = img2[1983:1976];
      img_out2[95:88] = img2[1991:1984];
      img_out2[103:96] = img2[1999:1992];
      img_out2[111:104] = img2[2007:2000];
      img_out2[119:112] = img2[2015:2008];
      img_out2[127:120] = img2[2023:2016];
      img_out2[135:128] = img2[2031:2024];
      img_out2[143:136] = img2[2039:2032];
      img_out2[151:144] = img2[2047:2040];
      img_out2[159:152] = img2[2055:2048];
      img_out2[167:160] = img2[2063:2056];
      img_out2[175:168] = img2[2071:2064];
      img_out3[7:0] = img3[1903:1896];
      img_out3[15:8] = img3[1911:1904];
      img_out3[23:16] = img3[1919:1912];
      img_out3[31:24] = img3[1927:1920];
      img_out3[39:32] = img3[1935:1928];
      img_out3[47:40] = img3[1943:1936];
      img_out3[55:48] = img3[1951:1944];
      img_out3[63:56] = img3[1959:1952];
      img_out3[71:64] = img3[1967:1960];
      img_out3[79:72] = img3[1975:1968];
      img_out3[87:80] = img3[1983:1976];
      img_out3[95:88] = img3[1991:1984];
      img_out3[103:96] = img3[1999:1992];
      img_out3[111:104] = img3[2007:2000];
      img_out3[119:112] = img3[2015:2008];
      img_out3[127:120] = img3[2023:2016];
      img_out3[135:128] = img3[2031:2024];
      img_out3[143:136] = img3[2039:2032];
      img_out3[151:144] = img3[2047:2040];
      img_out3[159:152] = img3[2055:2048];
      img_out3[167:160] = img3[2063:2056];
      img_out3[175:168] = img3[2071:2064];
      img_out4[7:0] = img4[1903:1896];
      img_out4[15:8] = img4[1911:1904];
      img_out4[23:16] = img4[1919:1912];
      img_out4[31:24] = img4[1927:1920];
      img_out4[39:32] = img4[1935:1928];
      img_out4[47:40] = img4[1943:1936];
      img_out4[55:48] = img4[1951:1944];
      img_out4[63:56] = img4[1959:1952];
      img_out4[71:64] = img4[1967:1960];
      img_out4[79:72] = img4[1975:1968];
      img_out4[87:80] = img4[1983:1976];
      img_out4[95:88] = img4[1991:1984];
      img_out4[103:96] = img4[1999:1992];
      img_out4[111:104] = img4[2007:2000];
      img_out4[119:112] = img4[2015:2008];
      img_out4[127:120] = img4[2023:2016];
      img_out4[135:128] = img4[2031:2024];
      img_out4[143:136] = img4[2039:2032];
      img_out4[151:144] = img4[2047:2040];
      img_out4[159:152] = img4[2055:2048];
      img_out4[167:160] = img4[2063:2056];
      img_out4[175:168] = img4[2071:2064];
    end
    'd16: begin
      img_out0[7:0] = img0[2031:2024];
      img_out0[15:8] = img0[2039:2032];
      img_out0[23:16] = img0[2047:2040];
      img_out0[31:24] = img0[2055:2048];
      img_out0[39:32] = img0[2063:2056];
      img_out0[47:40] = img0[2071:2064];
      img_out0[55:48] = img0[2079:2072];
      img_out0[63:56] = img0[2087:2080];
      img_out0[71:64] = img0[2095:2088];
      img_out0[79:72] = img0[2103:2096];
      img_out0[87:80] = img0[2111:2104];
      img_out0[95:88] = img0[2119:2112];
      img_out0[103:96] = img0[2127:2120];
      img_out0[111:104] = img0[2135:2128];
      img_out0[119:112] = img0[2143:2136];
      img_out0[127:120] = img0[2151:2144];
      img_out0[135:128] = img0[2159:2152];
      img_out0[143:136] = img0[2167:2160];
      img_out0[151:144] = img0[2175:2168];
      img_out0[159:152] = img0[2183:2176];
      img_out0[167:160] = img0[2191:2184];
      img_out0[175:168] = img0[2199:2192];
      img_out1[7:0] = img1[2031:2024];
      img_out1[15:8] = img1[2039:2032];
      img_out1[23:16] = img1[2047:2040];
      img_out1[31:24] = img1[2055:2048];
      img_out1[39:32] = img1[2063:2056];
      img_out1[47:40] = img1[2071:2064];
      img_out1[55:48] = img1[2079:2072];
      img_out1[63:56] = img1[2087:2080];
      img_out1[71:64] = img1[2095:2088];
      img_out1[79:72] = img1[2103:2096];
      img_out1[87:80] = img1[2111:2104];
      img_out1[95:88] = img1[2119:2112];
      img_out1[103:96] = img1[2127:2120];
      img_out1[111:104] = img1[2135:2128];
      img_out1[119:112] = img1[2143:2136];
      img_out1[127:120] = img1[2151:2144];
      img_out1[135:128] = img1[2159:2152];
      img_out1[143:136] = img1[2167:2160];
      img_out1[151:144] = img1[2175:2168];
      img_out1[159:152] = img1[2183:2176];
      img_out1[167:160] = img1[2191:2184];
      img_out1[175:168] = img1[2199:2192];
      img_out2[7:0] = img2[2031:2024];
      img_out2[15:8] = img2[2039:2032];
      img_out2[23:16] = img2[2047:2040];
      img_out2[31:24] = img2[2055:2048];
      img_out2[39:32] = img2[2063:2056];
      img_out2[47:40] = img2[2071:2064];
      img_out2[55:48] = img2[2079:2072];
      img_out2[63:56] = img2[2087:2080];
      img_out2[71:64] = img2[2095:2088];
      img_out2[79:72] = img2[2103:2096];
      img_out2[87:80] = img2[2111:2104];
      img_out2[95:88] = img2[2119:2112];
      img_out2[103:96] = img2[2127:2120];
      img_out2[111:104] = img2[2135:2128];
      img_out2[119:112] = img2[2143:2136];
      img_out2[127:120] = img2[2151:2144];
      img_out2[135:128] = img2[2159:2152];
      img_out2[143:136] = img2[2167:2160];
      img_out2[151:144] = img2[2175:2168];
      img_out2[159:152] = img2[2183:2176];
      img_out2[167:160] = img2[2191:2184];
      img_out2[175:168] = img2[2199:2192];
      img_out3[7:0] = img3[2031:2024];
      img_out3[15:8] = img3[2039:2032];
      img_out3[23:16] = img3[2047:2040];
      img_out3[31:24] = img3[2055:2048];
      img_out3[39:32] = img3[2063:2056];
      img_out3[47:40] = img3[2071:2064];
      img_out3[55:48] = img3[2079:2072];
      img_out3[63:56] = img3[2087:2080];
      img_out3[71:64] = img3[2095:2088];
      img_out3[79:72] = img3[2103:2096];
      img_out3[87:80] = img3[2111:2104];
      img_out3[95:88] = img3[2119:2112];
      img_out3[103:96] = img3[2127:2120];
      img_out3[111:104] = img3[2135:2128];
      img_out3[119:112] = img3[2143:2136];
      img_out3[127:120] = img3[2151:2144];
      img_out3[135:128] = img3[2159:2152];
      img_out3[143:136] = img3[2167:2160];
      img_out3[151:144] = img3[2175:2168];
      img_out3[159:152] = img3[2183:2176];
      img_out3[167:160] = img3[2191:2184];
      img_out3[175:168] = img3[2199:2192];
      img_out4[7:0] = img4[2031:2024];
      img_out4[15:8] = img4[2039:2032];
      img_out4[23:16] = img4[2047:2040];
      img_out4[31:24] = img4[2055:2048];
      img_out4[39:32] = img4[2063:2056];
      img_out4[47:40] = img4[2071:2064];
      img_out4[55:48] = img4[2079:2072];
      img_out4[63:56] = img4[2087:2080];
      img_out4[71:64] = img4[2095:2088];
      img_out4[79:72] = img4[2103:2096];
      img_out4[87:80] = img4[2111:2104];
      img_out4[95:88] = img4[2119:2112];
      img_out4[103:96] = img4[2127:2120];
      img_out4[111:104] = img4[2135:2128];
      img_out4[119:112] = img4[2143:2136];
      img_out4[127:120] = img4[2151:2144];
      img_out4[135:128] = img4[2159:2152];
      img_out4[143:136] = img4[2167:2160];
      img_out4[151:144] = img4[2175:2168];
      img_out4[159:152] = img4[2183:2176];
      img_out4[167:160] = img4[2191:2184];
      img_out4[175:168] = img4[2199:2192];
    end
    'd17: begin
      img_out0[7:0] = img0[2159:2152];
      img_out0[15:8] = img0[2167:2160];
      img_out0[23:16] = img0[2175:2168];
      img_out0[31:24] = img0[2183:2176];
      img_out0[39:32] = img0[2191:2184];
      img_out0[47:40] = img0[2199:2192];
      img_out0[55:48] = img0[2207:2200];
      img_out0[63:56] = img0[2215:2208];
      img_out0[71:64] = img0[2223:2216];
      img_out0[79:72] = img0[2231:2224];
      img_out0[87:80] = img0[2239:2232];
      img_out0[95:88] = img0[2247:2240];
      img_out0[103:96] = img0[2255:2248];
      img_out0[111:104] = img0[2263:2256];
      img_out0[119:112] = img0[2271:2264];
      img_out0[127:120] = img0[2279:2272];
      img_out0[135:128] = img0[2287:2280];
      img_out0[143:136] = img0[2295:2288];
      img_out0[151:144] = img0[2303:2296];
      img_out0[159:152] = img0[2311:2304];
      img_out0[167:160] = img0[2319:2312];
      img_out0[175:168] = img0[2327:2320];
      img_out1[7:0] = img1[2159:2152];
      img_out1[15:8] = img1[2167:2160];
      img_out1[23:16] = img1[2175:2168];
      img_out1[31:24] = img1[2183:2176];
      img_out1[39:32] = img1[2191:2184];
      img_out1[47:40] = img1[2199:2192];
      img_out1[55:48] = img1[2207:2200];
      img_out1[63:56] = img1[2215:2208];
      img_out1[71:64] = img1[2223:2216];
      img_out1[79:72] = img1[2231:2224];
      img_out1[87:80] = img1[2239:2232];
      img_out1[95:88] = img1[2247:2240];
      img_out1[103:96] = img1[2255:2248];
      img_out1[111:104] = img1[2263:2256];
      img_out1[119:112] = img1[2271:2264];
      img_out1[127:120] = img1[2279:2272];
      img_out1[135:128] = img1[2287:2280];
      img_out1[143:136] = img1[2295:2288];
      img_out1[151:144] = img1[2303:2296];
      img_out1[159:152] = img1[2311:2304];
      img_out1[167:160] = img1[2319:2312];
      img_out1[175:168] = img1[2327:2320];
      img_out2[7:0] = img2[2159:2152];
      img_out2[15:8] = img2[2167:2160];
      img_out2[23:16] = img2[2175:2168];
      img_out2[31:24] = img2[2183:2176];
      img_out2[39:32] = img2[2191:2184];
      img_out2[47:40] = img2[2199:2192];
      img_out2[55:48] = img2[2207:2200];
      img_out2[63:56] = img2[2215:2208];
      img_out2[71:64] = img2[2223:2216];
      img_out2[79:72] = img2[2231:2224];
      img_out2[87:80] = img2[2239:2232];
      img_out2[95:88] = img2[2247:2240];
      img_out2[103:96] = img2[2255:2248];
      img_out2[111:104] = img2[2263:2256];
      img_out2[119:112] = img2[2271:2264];
      img_out2[127:120] = img2[2279:2272];
      img_out2[135:128] = img2[2287:2280];
      img_out2[143:136] = img2[2295:2288];
      img_out2[151:144] = img2[2303:2296];
      img_out2[159:152] = img2[2311:2304];
      img_out2[167:160] = img2[2319:2312];
      img_out2[175:168] = img2[2327:2320];
      img_out3[7:0] = img3[2159:2152];
      img_out3[15:8] = img3[2167:2160];
      img_out3[23:16] = img3[2175:2168];
      img_out3[31:24] = img3[2183:2176];
      img_out3[39:32] = img3[2191:2184];
      img_out3[47:40] = img3[2199:2192];
      img_out3[55:48] = img3[2207:2200];
      img_out3[63:56] = img3[2215:2208];
      img_out3[71:64] = img3[2223:2216];
      img_out3[79:72] = img3[2231:2224];
      img_out3[87:80] = img3[2239:2232];
      img_out3[95:88] = img3[2247:2240];
      img_out3[103:96] = img3[2255:2248];
      img_out3[111:104] = img3[2263:2256];
      img_out3[119:112] = img3[2271:2264];
      img_out3[127:120] = img3[2279:2272];
      img_out3[135:128] = img3[2287:2280];
      img_out3[143:136] = img3[2295:2288];
      img_out3[151:144] = img3[2303:2296];
      img_out3[159:152] = img3[2311:2304];
      img_out3[167:160] = img3[2319:2312];
      img_out3[175:168] = img3[2327:2320];
      img_out4[7:0] = img4[2159:2152];
      img_out4[15:8] = img4[2167:2160];
      img_out4[23:16] = img4[2175:2168];
      img_out4[31:24] = img4[2183:2176];
      img_out4[39:32] = img4[2191:2184];
      img_out4[47:40] = img4[2199:2192];
      img_out4[55:48] = img4[2207:2200];
      img_out4[63:56] = img4[2215:2208];
      img_out4[71:64] = img4[2223:2216];
      img_out4[79:72] = img4[2231:2224];
      img_out4[87:80] = img4[2239:2232];
      img_out4[95:88] = img4[2247:2240];
      img_out4[103:96] = img4[2255:2248];
      img_out4[111:104] = img4[2263:2256];
      img_out4[119:112] = img4[2271:2264];
      img_out4[127:120] = img4[2279:2272];
      img_out4[135:128] = img4[2287:2280];
      img_out4[143:136] = img4[2295:2288];
      img_out4[151:144] = img4[2303:2296];
      img_out4[159:152] = img4[2311:2304];
      img_out4[167:160] = img4[2319:2312];
      img_out4[175:168] = img4[2327:2320];
    end
    'd18: begin
      img_out0[7:0] = img0[2287:2280];
      img_out0[15:8] = img0[2295:2288];
      img_out0[23:16] = img0[2303:2296];
      img_out0[31:24] = img0[2311:2304];
      img_out0[39:32] = img0[2319:2312];
      img_out0[47:40] = img0[2327:2320];
      img_out0[55:48] = img0[2335:2328];
      img_out0[63:56] = img0[2343:2336];
      img_out0[71:64] = img0[2351:2344];
      img_out0[79:72] = img0[2359:2352];
      img_out0[87:80] = img0[2367:2360];
      img_out0[95:88] = img0[2375:2368];
      img_out0[103:96] = img0[2383:2376];
      img_out0[111:104] = img0[2391:2384];
      img_out0[119:112] = img0[2399:2392];
      img_out0[127:120] = img0[2407:2400];
      img_out0[135:128] = img0[2415:2408];
      img_out0[143:136] = img0[2423:2416];
      img_out0[151:144] = img0[2431:2424];
      img_out0[159:152] = img0[2439:2432];
      img_out0[167:160] = img0[2447:2440];
      img_out0[175:168] = img0[2455:2448];
      img_out1[7:0] = img1[2287:2280];
      img_out1[15:8] = img1[2295:2288];
      img_out1[23:16] = img1[2303:2296];
      img_out1[31:24] = img1[2311:2304];
      img_out1[39:32] = img1[2319:2312];
      img_out1[47:40] = img1[2327:2320];
      img_out1[55:48] = img1[2335:2328];
      img_out1[63:56] = img1[2343:2336];
      img_out1[71:64] = img1[2351:2344];
      img_out1[79:72] = img1[2359:2352];
      img_out1[87:80] = img1[2367:2360];
      img_out1[95:88] = img1[2375:2368];
      img_out1[103:96] = img1[2383:2376];
      img_out1[111:104] = img1[2391:2384];
      img_out1[119:112] = img1[2399:2392];
      img_out1[127:120] = img1[2407:2400];
      img_out1[135:128] = img1[2415:2408];
      img_out1[143:136] = img1[2423:2416];
      img_out1[151:144] = img1[2431:2424];
      img_out1[159:152] = img1[2439:2432];
      img_out1[167:160] = img1[2447:2440];
      img_out1[175:168] = img1[2455:2448];
      img_out2[7:0] = img2[2287:2280];
      img_out2[15:8] = img2[2295:2288];
      img_out2[23:16] = img2[2303:2296];
      img_out2[31:24] = img2[2311:2304];
      img_out2[39:32] = img2[2319:2312];
      img_out2[47:40] = img2[2327:2320];
      img_out2[55:48] = img2[2335:2328];
      img_out2[63:56] = img2[2343:2336];
      img_out2[71:64] = img2[2351:2344];
      img_out2[79:72] = img2[2359:2352];
      img_out2[87:80] = img2[2367:2360];
      img_out2[95:88] = img2[2375:2368];
      img_out2[103:96] = img2[2383:2376];
      img_out2[111:104] = img2[2391:2384];
      img_out2[119:112] = img2[2399:2392];
      img_out2[127:120] = img2[2407:2400];
      img_out2[135:128] = img2[2415:2408];
      img_out2[143:136] = img2[2423:2416];
      img_out2[151:144] = img2[2431:2424];
      img_out2[159:152] = img2[2439:2432];
      img_out2[167:160] = img2[2447:2440];
      img_out2[175:168] = img2[2455:2448];
      img_out3[7:0] = img3[2287:2280];
      img_out3[15:8] = img3[2295:2288];
      img_out3[23:16] = img3[2303:2296];
      img_out3[31:24] = img3[2311:2304];
      img_out3[39:32] = img3[2319:2312];
      img_out3[47:40] = img3[2327:2320];
      img_out3[55:48] = img3[2335:2328];
      img_out3[63:56] = img3[2343:2336];
      img_out3[71:64] = img3[2351:2344];
      img_out3[79:72] = img3[2359:2352];
      img_out3[87:80] = img3[2367:2360];
      img_out3[95:88] = img3[2375:2368];
      img_out3[103:96] = img3[2383:2376];
      img_out3[111:104] = img3[2391:2384];
      img_out3[119:112] = img3[2399:2392];
      img_out3[127:120] = img3[2407:2400];
      img_out3[135:128] = img3[2415:2408];
      img_out3[143:136] = img3[2423:2416];
      img_out3[151:144] = img3[2431:2424];
      img_out3[159:152] = img3[2439:2432];
      img_out3[167:160] = img3[2447:2440];
      img_out3[175:168] = img3[2455:2448];
      img_out4[7:0] = img4[2287:2280];
      img_out4[15:8] = img4[2295:2288];
      img_out4[23:16] = img4[2303:2296];
      img_out4[31:24] = img4[2311:2304];
      img_out4[39:32] = img4[2319:2312];
      img_out4[47:40] = img4[2327:2320];
      img_out4[55:48] = img4[2335:2328];
      img_out4[63:56] = img4[2343:2336];
      img_out4[71:64] = img4[2351:2344];
      img_out4[79:72] = img4[2359:2352];
      img_out4[87:80] = img4[2367:2360];
      img_out4[95:88] = img4[2375:2368];
      img_out4[103:96] = img4[2383:2376];
      img_out4[111:104] = img4[2391:2384];
      img_out4[119:112] = img4[2399:2392];
      img_out4[127:120] = img4[2407:2400];
      img_out4[135:128] = img4[2415:2408];
      img_out4[143:136] = img4[2423:2416];
      img_out4[151:144] = img4[2431:2424];
      img_out4[159:152] = img4[2439:2432];
      img_out4[167:160] = img4[2447:2440];
      img_out4[175:168] = img4[2455:2448];
    end
    'd19: begin
      img_out0[7:0] = img0[2415:2408];
      img_out0[15:8] = img0[2423:2416];
      img_out0[23:16] = img0[2431:2424];
      img_out0[31:24] = img0[2439:2432];
      img_out0[39:32] = img0[2447:2440];
      img_out0[47:40] = img0[2455:2448];
      img_out0[55:48] = img0[2463:2456];
      img_out0[63:56] = img0[2471:2464];
      img_out0[71:64] = img0[2479:2472];
      img_out0[79:72] = img0[2487:2480];
      img_out0[87:80] = img0[2495:2488];
      img_out0[95:88] = img0[2503:2496];
      img_out0[103:96] = img0[2511:2504];
      img_out0[111:104] = img0[2519:2512];
      img_out0[119:112] = img0[2527:2520];
      img_out0[127:120] = img0[2535:2528];
      img_out0[135:128] = img0[2543:2536];
      img_out0[143:136] = img0[2551:2544];
      img_out0[151:144] = img0[2559:2552];
      img_out0[159:152] = img0[2567:2560];
      img_out0[167:160] = img0[2575:2568];
      img_out0[175:168] = img0[2583:2576];
      img_out1[7:0] = img1[2415:2408];
      img_out1[15:8] = img1[2423:2416];
      img_out1[23:16] = img1[2431:2424];
      img_out1[31:24] = img1[2439:2432];
      img_out1[39:32] = img1[2447:2440];
      img_out1[47:40] = img1[2455:2448];
      img_out1[55:48] = img1[2463:2456];
      img_out1[63:56] = img1[2471:2464];
      img_out1[71:64] = img1[2479:2472];
      img_out1[79:72] = img1[2487:2480];
      img_out1[87:80] = img1[2495:2488];
      img_out1[95:88] = img1[2503:2496];
      img_out1[103:96] = img1[2511:2504];
      img_out1[111:104] = img1[2519:2512];
      img_out1[119:112] = img1[2527:2520];
      img_out1[127:120] = img1[2535:2528];
      img_out1[135:128] = img1[2543:2536];
      img_out1[143:136] = img1[2551:2544];
      img_out1[151:144] = img1[2559:2552];
      img_out1[159:152] = img1[2567:2560];
      img_out1[167:160] = img1[2575:2568];
      img_out1[175:168] = img1[2583:2576];
      img_out2[7:0] = img2[2415:2408];
      img_out2[15:8] = img2[2423:2416];
      img_out2[23:16] = img2[2431:2424];
      img_out2[31:24] = img2[2439:2432];
      img_out2[39:32] = img2[2447:2440];
      img_out2[47:40] = img2[2455:2448];
      img_out2[55:48] = img2[2463:2456];
      img_out2[63:56] = img2[2471:2464];
      img_out2[71:64] = img2[2479:2472];
      img_out2[79:72] = img2[2487:2480];
      img_out2[87:80] = img2[2495:2488];
      img_out2[95:88] = img2[2503:2496];
      img_out2[103:96] = img2[2511:2504];
      img_out2[111:104] = img2[2519:2512];
      img_out2[119:112] = img2[2527:2520];
      img_out2[127:120] = img2[2535:2528];
      img_out2[135:128] = img2[2543:2536];
      img_out2[143:136] = img2[2551:2544];
      img_out2[151:144] = img2[2559:2552];
      img_out2[159:152] = img2[2567:2560];
      img_out2[167:160] = img2[2575:2568];
      img_out2[175:168] = img2[2583:2576];
      img_out3[7:0] = img3[2415:2408];
      img_out3[15:8] = img3[2423:2416];
      img_out3[23:16] = img3[2431:2424];
      img_out3[31:24] = img3[2439:2432];
      img_out3[39:32] = img3[2447:2440];
      img_out3[47:40] = img3[2455:2448];
      img_out3[55:48] = img3[2463:2456];
      img_out3[63:56] = img3[2471:2464];
      img_out3[71:64] = img3[2479:2472];
      img_out3[79:72] = img3[2487:2480];
      img_out3[87:80] = img3[2495:2488];
      img_out3[95:88] = img3[2503:2496];
      img_out3[103:96] = img3[2511:2504];
      img_out3[111:104] = img3[2519:2512];
      img_out3[119:112] = img3[2527:2520];
      img_out3[127:120] = img3[2535:2528];
      img_out3[135:128] = img3[2543:2536];
      img_out3[143:136] = img3[2551:2544];
      img_out3[151:144] = img3[2559:2552];
      img_out3[159:152] = img3[2567:2560];
      img_out3[167:160] = img3[2575:2568];
      img_out3[175:168] = img3[2583:2576];
      img_out4[7:0] = img4[2415:2408];
      img_out4[15:8] = img4[2423:2416];
      img_out4[23:16] = img4[2431:2424];
      img_out4[31:24] = img4[2439:2432];
      img_out4[39:32] = img4[2447:2440];
      img_out4[47:40] = img4[2455:2448];
      img_out4[55:48] = img4[2463:2456];
      img_out4[63:56] = img4[2471:2464];
      img_out4[71:64] = img4[2479:2472];
      img_out4[79:72] = img4[2487:2480];
      img_out4[87:80] = img4[2495:2488];
      img_out4[95:88] = img4[2503:2496];
      img_out4[103:96] = img4[2511:2504];
      img_out4[111:104] = img4[2519:2512];
      img_out4[119:112] = img4[2527:2520];
      img_out4[127:120] = img4[2535:2528];
      img_out4[135:128] = img4[2543:2536];
      img_out4[143:136] = img4[2551:2544];
      img_out4[151:144] = img4[2559:2552];
      img_out4[159:152] = img4[2567:2560];
      img_out4[167:160] = img4[2575:2568];
      img_out4[175:168] = img4[2583:2576];
    end
    'd20: begin
      img_out0[7:0] = img0[2543:2536];
      img_out0[15:8] = img0[2551:2544];
      img_out0[23:16] = img0[2559:2552];
      img_out0[31:24] = img0[2567:2560];
      img_out0[39:32] = img0[2575:2568];
      img_out0[47:40] = img0[2583:2576];
      img_out0[55:48] = img0[2591:2584];
      img_out0[63:56] = img0[2599:2592];
      img_out0[71:64] = img0[2607:2600];
      img_out0[79:72] = img0[2615:2608];
      img_out0[87:80] = img0[2623:2616];
      img_out0[95:88] = img0[2631:2624];
      img_out0[103:96] = img0[2639:2632];
      img_out0[111:104] = img0[2647:2640];
      img_out0[119:112] = img0[2655:2648];
      img_out0[127:120] = img0[2663:2656];
      img_out0[135:128] = img0[2671:2664];
      img_out0[143:136] = img0[2679:2672];
      img_out0[151:144] = img0[2687:2680];
      img_out0[159:152] = img0[2695:2688];
      img_out0[167:160] = img0[2703:2696];
      img_out0[175:168] = img0[2711:2704];
      img_out1[7:0] = img1[2543:2536];
      img_out1[15:8] = img1[2551:2544];
      img_out1[23:16] = img1[2559:2552];
      img_out1[31:24] = img1[2567:2560];
      img_out1[39:32] = img1[2575:2568];
      img_out1[47:40] = img1[2583:2576];
      img_out1[55:48] = img1[2591:2584];
      img_out1[63:56] = img1[2599:2592];
      img_out1[71:64] = img1[2607:2600];
      img_out1[79:72] = img1[2615:2608];
      img_out1[87:80] = img1[2623:2616];
      img_out1[95:88] = img1[2631:2624];
      img_out1[103:96] = img1[2639:2632];
      img_out1[111:104] = img1[2647:2640];
      img_out1[119:112] = img1[2655:2648];
      img_out1[127:120] = img1[2663:2656];
      img_out1[135:128] = img1[2671:2664];
      img_out1[143:136] = img1[2679:2672];
      img_out1[151:144] = img1[2687:2680];
      img_out1[159:152] = img1[2695:2688];
      img_out1[167:160] = img1[2703:2696];
      img_out1[175:168] = img1[2711:2704];
      img_out2[7:0] = img2[2543:2536];
      img_out2[15:8] = img2[2551:2544];
      img_out2[23:16] = img2[2559:2552];
      img_out2[31:24] = img2[2567:2560];
      img_out2[39:32] = img2[2575:2568];
      img_out2[47:40] = img2[2583:2576];
      img_out2[55:48] = img2[2591:2584];
      img_out2[63:56] = img2[2599:2592];
      img_out2[71:64] = img2[2607:2600];
      img_out2[79:72] = img2[2615:2608];
      img_out2[87:80] = img2[2623:2616];
      img_out2[95:88] = img2[2631:2624];
      img_out2[103:96] = img2[2639:2632];
      img_out2[111:104] = img2[2647:2640];
      img_out2[119:112] = img2[2655:2648];
      img_out2[127:120] = img2[2663:2656];
      img_out2[135:128] = img2[2671:2664];
      img_out2[143:136] = img2[2679:2672];
      img_out2[151:144] = img2[2687:2680];
      img_out2[159:152] = img2[2695:2688];
      img_out2[167:160] = img2[2703:2696];
      img_out2[175:168] = img2[2711:2704];
      img_out3[7:0] = img3[2543:2536];
      img_out3[15:8] = img3[2551:2544];
      img_out3[23:16] = img3[2559:2552];
      img_out3[31:24] = img3[2567:2560];
      img_out3[39:32] = img3[2575:2568];
      img_out3[47:40] = img3[2583:2576];
      img_out3[55:48] = img3[2591:2584];
      img_out3[63:56] = img3[2599:2592];
      img_out3[71:64] = img3[2607:2600];
      img_out3[79:72] = img3[2615:2608];
      img_out3[87:80] = img3[2623:2616];
      img_out3[95:88] = img3[2631:2624];
      img_out3[103:96] = img3[2639:2632];
      img_out3[111:104] = img3[2647:2640];
      img_out3[119:112] = img3[2655:2648];
      img_out3[127:120] = img3[2663:2656];
      img_out3[135:128] = img3[2671:2664];
      img_out3[143:136] = img3[2679:2672];
      img_out3[151:144] = img3[2687:2680];
      img_out3[159:152] = img3[2695:2688];
      img_out3[167:160] = img3[2703:2696];
      img_out3[175:168] = img3[2711:2704];
      img_out4[7:0] = img4[2543:2536];
      img_out4[15:8] = img4[2551:2544];
      img_out4[23:16] = img4[2559:2552];
      img_out4[31:24] = img4[2567:2560];
      img_out4[39:32] = img4[2575:2568];
      img_out4[47:40] = img4[2583:2576];
      img_out4[55:48] = img4[2591:2584];
      img_out4[63:56] = img4[2599:2592];
      img_out4[71:64] = img4[2607:2600];
      img_out4[79:72] = img4[2615:2608];
      img_out4[87:80] = img4[2623:2616];
      img_out4[95:88] = img4[2631:2624];
      img_out4[103:96] = img4[2639:2632];
      img_out4[111:104] = img4[2647:2640];
      img_out4[119:112] = img4[2655:2648];
      img_out4[127:120] = img4[2663:2656];
      img_out4[135:128] = img4[2671:2664];
      img_out4[143:136] = img4[2679:2672];
      img_out4[151:144] = img4[2687:2680];
      img_out4[159:152] = img4[2695:2688];
      img_out4[167:160] = img4[2703:2696];
      img_out4[175:168] = img4[2711:2704];
    end
    'd21: begin
      img_out0[7:0] = img0[2671:2664];
      img_out0[15:8] = img0[2679:2672];
      img_out0[23:16] = img0[2687:2680];
      img_out0[31:24] = img0[2695:2688];
      img_out0[39:32] = img0[2703:2696];
      img_out0[47:40] = img0[2711:2704];
      img_out0[55:48] = img0[2719:2712];
      img_out0[63:56] = img0[2727:2720];
      img_out0[71:64] = img0[2735:2728];
      img_out0[79:72] = img0[2743:2736];
      img_out0[87:80] = img0[2751:2744];
      img_out0[95:88] = img0[2759:2752];
      img_out0[103:96] = img0[2767:2760];
      img_out0[111:104] = img0[2775:2768];
      img_out0[119:112] = img0[2783:2776];
      img_out0[127:120] = img0[2791:2784];
      img_out0[135:128] = img0[2799:2792];
      img_out0[143:136] = img0[2807:2800];
      img_out0[151:144] = img0[2815:2808];
      img_out0[159:152] = img0[2823:2816];
      img_out0[167:160] = img0[2831:2824];
      img_out0[175:168] = img0[2839:2832];
      img_out1[7:0] = img1[2671:2664];
      img_out1[15:8] = img1[2679:2672];
      img_out1[23:16] = img1[2687:2680];
      img_out1[31:24] = img1[2695:2688];
      img_out1[39:32] = img1[2703:2696];
      img_out1[47:40] = img1[2711:2704];
      img_out1[55:48] = img1[2719:2712];
      img_out1[63:56] = img1[2727:2720];
      img_out1[71:64] = img1[2735:2728];
      img_out1[79:72] = img1[2743:2736];
      img_out1[87:80] = img1[2751:2744];
      img_out1[95:88] = img1[2759:2752];
      img_out1[103:96] = img1[2767:2760];
      img_out1[111:104] = img1[2775:2768];
      img_out1[119:112] = img1[2783:2776];
      img_out1[127:120] = img1[2791:2784];
      img_out1[135:128] = img1[2799:2792];
      img_out1[143:136] = img1[2807:2800];
      img_out1[151:144] = img1[2815:2808];
      img_out1[159:152] = img1[2823:2816];
      img_out1[167:160] = img1[2831:2824];
      img_out1[175:168] = img1[2839:2832];
      img_out2[7:0] = img2[2671:2664];
      img_out2[15:8] = img2[2679:2672];
      img_out2[23:16] = img2[2687:2680];
      img_out2[31:24] = img2[2695:2688];
      img_out2[39:32] = img2[2703:2696];
      img_out2[47:40] = img2[2711:2704];
      img_out2[55:48] = img2[2719:2712];
      img_out2[63:56] = img2[2727:2720];
      img_out2[71:64] = img2[2735:2728];
      img_out2[79:72] = img2[2743:2736];
      img_out2[87:80] = img2[2751:2744];
      img_out2[95:88] = img2[2759:2752];
      img_out2[103:96] = img2[2767:2760];
      img_out2[111:104] = img2[2775:2768];
      img_out2[119:112] = img2[2783:2776];
      img_out2[127:120] = img2[2791:2784];
      img_out2[135:128] = img2[2799:2792];
      img_out2[143:136] = img2[2807:2800];
      img_out2[151:144] = img2[2815:2808];
      img_out2[159:152] = img2[2823:2816];
      img_out2[167:160] = img2[2831:2824];
      img_out2[175:168] = img2[2839:2832];
      img_out3[7:0] = img3[2671:2664];
      img_out3[15:8] = img3[2679:2672];
      img_out3[23:16] = img3[2687:2680];
      img_out3[31:24] = img3[2695:2688];
      img_out3[39:32] = img3[2703:2696];
      img_out3[47:40] = img3[2711:2704];
      img_out3[55:48] = img3[2719:2712];
      img_out3[63:56] = img3[2727:2720];
      img_out3[71:64] = img3[2735:2728];
      img_out3[79:72] = img3[2743:2736];
      img_out3[87:80] = img3[2751:2744];
      img_out3[95:88] = img3[2759:2752];
      img_out3[103:96] = img3[2767:2760];
      img_out3[111:104] = img3[2775:2768];
      img_out3[119:112] = img3[2783:2776];
      img_out3[127:120] = img3[2791:2784];
      img_out3[135:128] = img3[2799:2792];
      img_out3[143:136] = img3[2807:2800];
      img_out3[151:144] = img3[2815:2808];
      img_out3[159:152] = img3[2823:2816];
      img_out3[167:160] = img3[2831:2824];
      img_out3[175:168] = img3[2839:2832];
      img_out4[7:0] = img4[2671:2664];
      img_out4[15:8] = img4[2679:2672];
      img_out4[23:16] = img4[2687:2680];
      img_out4[31:24] = img4[2695:2688];
      img_out4[39:32] = img4[2703:2696];
      img_out4[47:40] = img4[2711:2704];
      img_out4[55:48] = img4[2719:2712];
      img_out4[63:56] = img4[2727:2720];
      img_out4[71:64] = img4[2735:2728];
      img_out4[79:72] = img4[2743:2736];
      img_out4[87:80] = img4[2751:2744];
      img_out4[95:88] = img4[2759:2752];
      img_out4[103:96] = img4[2767:2760];
      img_out4[111:104] = img4[2775:2768];
      img_out4[119:112] = img4[2783:2776];
      img_out4[127:120] = img4[2791:2784];
      img_out4[135:128] = img4[2799:2792];
      img_out4[143:136] = img4[2807:2800];
      img_out4[151:144] = img4[2815:2808];
      img_out4[159:152] = img4[2823:2816];
      img_out4[167:160] = img4[2831:2824];
      img_out4[175:168] = img4[2839:2832];
    end
    'd22: begin
      img_out0[7:0] = img0[2799:2792];
      img_out0[15:8] = img0[2807:2800];
      img_out0[23:16] = img0[2815:2808];
      img_out0[31:24] = img0[2823:2816];
      img_out0[39:32] = img0[2831:2824];
      img_out0[47:40] = img0[2839:2832];
      img_out0[55:48] = img0[2847:2840];
      img_out0[63:56] = img0[2855:2848];
      img_out0[71:64] = img0[2863:2856];
      img_out0[79:72] = img0[2871:2864];
      img_out0[87:80] = img0[2879:2872];
      img_out0[95:88] = img0[2887:2880];
      img_out0[103:96] = img0[2895:2888];
      img_out0[111:104] = img0[2903:2896];
      img_out0[119:112] = img0[2911:2904];
      img_out0[127:120] = img0[2919:2912];
      img_out0[135:128] = img0[2927:2920];
      img_out0[143:136] = img0[2935:2928];
      img_out0[151:144] = img0[2943:2936];
      img_out0[159:152] = img0[2951:2944];
      img_out0[167:160] = img0[2959:2952];
      img_out0[175:168] = img0[2967:2960];
      img_out1[7:0] = img1[2799:2792];
      img_out1[15:8] = img1[2807:2800];
      img_out1[23:16] = img1[2815:2808];
      img_out1[31:24] = img1[2823:2816];
      img_out1[39:32] = img1[2831:2824];
      img_out1[47:40] = img1[2839:2832];
      img_out1[55:48] = img1[2847:2840];
      img_out1[63:56] = img1[2855:2848];
      img_out1[71:64] = img1[2863:2856];
      img_out1[79:72] = img1[2871:2864];
      img_out1[87:80] = img1[2879:2872];
      img_out1[95:88] = img1[2887:2880];
      img_out1[103:96] = img1[2895:2888];
      img_out1[111:104] = img1[2903:2896];
      img_out1[119:112] = img1[2911:2904];
      img_out1[127:120] = img1[2919:2912];
      img_out1[135:128] = img1[2927:2920];
      img_out1[143:136] = img1[2935:2928];
      img_out1[151:144] = img1[2943:2936];
      img_out1[159:152] = img1[2951:2944];
      img_out1[167:160] = img1[2959:2952];
      img_out1[175:168] = img1[2967:2960];
      img_out2[7:0] = img2[2799:2792];
      img_out2[15:8] = img2[2807:2800];
      img_out2[23:16] = img2[2815:2808];
      img_out2[31:24] = img2[2823:2816];
      img_out2[39:32] = img2[2831:2824];
      img_out2[47:40] = img2[2839:2832];
      img_out2[55:48] = img2[2847:2840];
      img_out2[63:56] = img2[2855:2848];
      img_out2[71:64] = img2[2863:2856];
      img_out2[79:72] = img2[2871:2864];
      img_out2[87:80] = img2[2879:2872];
      img_out2[95:88] = img2[2887:2880];
      img_out2[103:96] = img2[2895:2888];
      img_out2[111:104] = img2[2903:2896];
      img_out2[119:112] = img2[2911:2904];
      img_out2[127:120] = img2[2919:2912];
      img_out2[135:128] = img2[2927:2920];
      img_out2[143:136] = img2[2935:2928];
      img_out2[151:144] = img2[2943:2936];
      img_out2[159:152] = img2[2951:2944];
      img_out2[167:160] = img2[2959:2952];
      img_out2[175:168] = img2[2967:2960];
      img_out3[7:0] = img3[2799:2792];
      img_out3[15:8] = img3[2807:2800];
      img_out3[23:16] = img3[2815:2808];
      img_out3[31:24] = img3[2823:2816];
      img_out3[39:32] = img3[2831:2824];
      img_out3[47:40] = img3[2839:2832];
      img_out3[55:48] = img3[2847:2840];
      img_out3[63:56] = img3[2855:2848];
      img_out3[71:64] = img3[2863:2856];
      img_out3[79:72] = img3[2871:2864];
      img_out3[87:80] = img3[2879:2872];
      img_out3[95:88] = img3[2887:2880];
      img_out3[103:96] = img3[2895:2888];
      img_out3[111:104] = img3[2903:2896];
      img_out3[119:112] = img3[2911:2904];
      img_out3[127:120] = img3[2919:2912];
      img_out3[135:128] = img3[2927:2920];
      img_out3[143:136] = img3[2935:2928];
      img_out3[151:144] = img3[2943:2936];
      img_out3[159:152] = img3[2951:2944];
      img_out3[167:160] = img3[2959:2952];
      img_out3[175:168] = img3[2967:2960];
      img_out4[7:0] = img4[2799:2792];
      img_out4[15:8] = img4[2807:2800];
      img_out4[23:16] = img4[2815:2808];
      img_out4[31:24] = img4[2823:2816];
      img_out4[39:32] = img4[2831:2824];
      img_out4[47:40] = img4[2839:2832];
      img_out4[55:48] = img4[2847:2840];
      img_out4[63:56] = img4[2855:2848];
      img_out4[71:64] = img4[2863:2856];
      img_out4[79:72] = img4[2871:2864];
      img_out4[87:80] = img4[2879:2872];
      img_out4[95:88] = img4[2887:2880];
      img_out4[103:96] = img4[2895:2888];
      img_out4[111:104] = img4[2903:2896];
      img_out4[119:112] = img4[2911:2904];
      img_out4[127:120] = img4[2919:2912];
      img_out4[135:128] = img4[2927:2920];
      img_out4[143:136] = img4[2935:2928];
      img_out4[151:144] = img4[2943:2936];
      img_out4[159:152] = img4[2951:2944];
      img_out4[167:160] = img4[2959:2952];
      img_out4[175:168] = img4[2967:2960];
    end
    'd23: begin
      img_out0[7:0] = img0[2927:2920];
      img_out0[15:8] = img0[2935:2928];
      img_out0[23:16] = img0[2943:2936];
      img_out0[31:24] = img0[2951:2944];
      img_out0[39:32] = img0[2959:2952];
      img_out0[47:40] = img0[2967:2960];
      img_out0[55:48] = img0[2975:2968];
      img_out0[63:56] = img0[2983:2976];
      img_out0[71:64] = img0[2991:2984];
      img_out0[79:72] = img0[2999:2992];
      img_out0[87:80] = img0[3007:3000];
      img_out0[95:88] = img0[3015:3008];
      img_out0[103:96] = img0[3023:3016];
      img_out0[111:104] = img0[3031:3024];
      img_out0[119:112] = img0[3039:3032];
      img_out0[127:120] = img0[3047:3040];
      img_out0[135:128] = img0[3055:3048];
      img_out0[143:136] = img0[3063:3056];
      img_out0[151:144] = img0[3071:3064];
      img_out0[159:152] = img0[3079:3072];
      img_out0[167:160] = img0[3087:3080];
      img_out0[175:168] = img0[3095:3088];
      img_out1[7:0] = img1[2927:2920];
      img_out1[15:8] = img1[2935:2928];
      img_out1[23:16] = img1[2943:2936];
      img_out1[31:24] = img1[2951:2944];
      img_out1[39:32] = img1[2959:2952];
      img_out1[47:40] = img1[2967:2960];
      img_out1[55:48] = img1[2975:2968];
      img_out1[63:56] = img1[2983:2976];
      img_out1[71:64] = img1[2991:2984];
      img_out1[79:72] = img1[2999:2992];
      img_out1[87:80] = img1[3007:3000];
      img_out1[95:88] = img1[3015:3008];
      img_out1[103:96] = img1[3023:3016];
      img_out1[111:104] = img1[3031:3024];
      img_out1[119:112] = img1[3039:3032];
      img_out1[127:120] = img1[3047:3040];
      img_out1[135:128] = img1[3055:3048];
      img_out1[143:136] = img1[3063:3056];
      img_out1[151:144] = img1[3071:3064];
      img_out1[159:152] = img1[3079:3072];
      img_out1[167:160] = img1[3087:3080];
      img_out1[175:168] = img1[3095:3088];
      img_out2[7:0] = img2[2927:2920];
      img_out2[15:8] = img2[2935:2928];
      img_out2[23:16] = img2[2943:2936];
      img_out2[31:24] = img2[2951:2944];
      img_out2[39:32] = img2[2959:2952];
      img_out2[47:40] = img2[2967:2960];
      img_out2[55:48] = img2[2975:2968];
      img_out2[63:56] = img2[2983:2976];
      img_out2[71:64] = img2[2991:2984];
      img_out2[79:72] = img2[2999:2992];
      img_out2[87:80] = img2[3007:3000];
      img_out2[95:88] = img2[3015:3008];
      img_out2[103:96] = img2[3023:3016];
      img_out2[111:104] = img2[3031:3024];
      img_out2[119:112] = img2[3039:3032];
      img_out2[127:120] = img2[3047:3040];
      img_out2[135:128] = img2[3055:3048];
      img_out2[143:136] = img2[3063:3056];
      img_out2[151:144] = img2[3071:3064];
      img_out2[159:152] = img2[3079:3072];
      img_out2[167:160] = img2[3087:3080];
      img_out2[175:168] = img2[3095:3088];
      img_out3[7:0] = img3[2927:2920];
      img_out3[15:8] = img3[2935:2928];
      img_out3[23:16] = img3[2943:2936];
      img_out3[31:24] = img3[2951:2944];
      img_out3[39:32] = img3[2959:2952];
      img_out3[47:40] = img3[2967:2960];
      img_out3[55:48] = img3[2975:2968];
      img_out3[63:56] = img3[2983:2976];
      img_out3[71:64] = img3[2991:2984];
      img_out3[79:72] = img3[2999:2992];
      img_out3[87:80] = img3[3007:3000];
      img_out3[95:88] = img3[3015:3008];
      img_out3[103:96] = img3[3023:3016];
      img_out3[111:104] = img3[3031:3024];
      img_out3[119:112] = img3[3039:3032];
      img_out3[127:120] = img3[3047:3040];
      img_out3[135:128] = img3[3055:3048];
      img_out3[143:136] = img3[3063:3056];
      img_out3[151:144] = img3[3071:3064];
      img_out3[159:152] = img3[3079:3072];
      img_out3[167:160] = img3[3087:3080];
      img_out3[175:168] = img3[3095:3088];
      img_out4[7:0] = img4[2927:2920];
      img_out4[15:8] = img4[2935:2928];
      img_out4[23:16] = img4[2943:2936];
      img_out4[31:24] = img4[2951:2944];
      img_out4[39:32] = img4[2959:2952];
      img_out4[47:40] = img4[2967:2960];
      img_out4[55:48] = img4[2975:2968];
      img_out4[63:56] = img4[2983:2976];
      img_out4[71:64] = img4[2991:2984];
      img_out4[79:72] = img4[2999:2992];
      img_out4[87:80] = img4[3007:3000];
      img_out4[95:88] = img4[3015:3008];
      img_out4[103:96] = img4[3023:3016];
      img_out4[111:104] = img4[3031:3024];
      img_out4[119:112] = img4[3039:3032];
      img_out4[127:120] = img4[3047:3040];
      img_out4[135:128] = img4[3055:3048];
      img_out4[143:136] = img4[3063:3056];
      img_out4[151:144] = img4[3071:3064];
      img_out4[159:152] = img4[3079:3072];
      img_out4[167:160] = img4[3087:3080];
      img_out4[175:168] = img4[3095:3088];
    end
    'd24: begin
      img_out0[7:0] = img0[3055:3048];
      img_out0[15:8] = img0[3063:3056];
      img_out0[23:16] = img0[3071:3064];
      img_out0[31:24] = img0[3079:3072];
      img_out0[39:32] = img0[3087:3080];
      img_out0[47:40] = img0[3095:3088];
      img_out0[55:48] = img0[3103:3096];
      img_out0[63:56] = img0[3111:3104];
      img_out0[71:64] = img0[3119:3112];
      img_out0[79:72] = img0[3127:3120];
      img_out0[87:80] = img0[3135:3128];
      img_out0[95:88] = img0[3143:3136];
      img_out0[103:96] = img0[3151:3144];
      img_out0[111:104] = img0[3159:3152];
      img_out0[119:112] = img0[3167:3160];
      img_out0[127:120] = img0[3175:3168];
      img_out0[135:128] = img0[3183:3176];
      img_out0[143:136] = img0[3191:3184];
      img_out0[151:144] = img0[3199:3192];
      img_out0[159:152] = img0[3207:3200];
      img_out0[167:160] = img0[3215:3208];
      img_out0[175:168] = img0[3223:3216];
      img_out1[7:0] = img1[3055:3048];
      img_out1[15:8] = img1[3063:3056];
      img_out1[23:16] = img1[3071:3064];
      img_out1[31:24] = img1[3079:3072];
      img_out1[39:32] = img1[3087:3080];
      img_out1[47:40] = img1[3095:3088];
      img_out1[55:48] = img1[3103:3096];
      img_out1[63:56] = img1[3111:3104];
      img_out1[71:64] = img1[3119:3112];
      img_out1[79:72] = img1[3127:3120];
      img_out1[87:80] = img1[3135:3128];
      img_out1[95:88] = img1[3143:3136];
      img_out1[103:96] = img1[3151:3144];
      img_out1[111:104] = img1[3159:3152];
      img_out1[119:112] = img1[3167:3160];
      img_out1[127:120] = img1[3175:3168];
      img_out1[135:128] = img1[3183:3176];
      img_out1[143:136] = img1[3191:3184];
      img_out1[151:144] = img1[3199:3192];
      img_out1[159:152] = img1[3207:3200];
      img_out1[167:160] = img1[3215:3208];
      img_out1[175:168] = img1[3223:3216];
      img_out2[7:0] = img2[3055:3048];
      img_out2[15:8] = img2[3063:3056];
      img_out2[23:16] = img2[3071:3064];
      img_out2[31:24] = img2[3079:3072];
      img_out2[39:32] = img2[3087:3080];
      img_out2[47:40] = img2[3095:3088];
      img_out2[55:48] = img2[3103:3096];
      img_out2[63:56] = img2[3111:3104];
      img_out2[71:64] = img2[3119:3112];
      img_out2[79:72] = img2[3127:3120];
      img_out2[87:80] = img2[3135:3128];
      img_out2[95:88] = img2[3143:3136];
      img_out2[103:96] = img2[3151:3144];
      img_out2[111:104] = img2[3159:3152];
      img_out2[119:112] = img2[3167:3160];
      img_out2[127:120] = img2[3175:3168];
      img_out2[135:128] = img2[3183:3176];
      img_out2[143:136] = img2[3191:3184];
      img_out2[151:144] = img2[3199:3192];
      img_out2[159:152] = img2[3207:3200];
      img_out2[167:160] = img2[3215:3208];
      img_out2[175:168] = img2[3223:3216];
      img_out3[7:0] = img3[3055:3048];
      img_out3[15:8] = img3[3063:3056];
      img_out3[23:16] = img3[3071:3064];
      img_out3[31:24] = img3[3079:3072];
      img_out3[39:32] = img3[3087:3080];
      img_out3[47:40] = img3[3095:3088];
      img_out3[55:48] = img3[3103:3096];
      img_out3[63:56] = img3[3111:3104];
      img_out3[71:64] = img3[3119:3112];
      img_out3[79:72] = img3[3127:3120];
      img_out3[87:80] = img3[3135:3128];
      img_out3[95:88] = img3[3143:3136];
      img_out3[103:96] = img3[3151:3144];
      img_out3[111:104] = img3[3159:3152];
      img_out3[119:112] = img3[3167:3160];
      img_out3[127:120] = img3[3175:3168];
      img_out3[135:128] = img3[3183:3176];
      img_out3[143:136] = img3[3191:3184];
      img_out3[151:144] = img3[3199:3192];
      img_out3[159:152] = img3[3207:3200];
      img_out3[167:160] = img3[3215:3208];
      img_out3[175:168] = img3[3223:3216];
      img_out4[7:0] = img4[3055:3048];
      img_out4[15:8] = img4[3063:3056];
      img_out4[23:16] = img4[3071:3064];
      img_out4[31:24] = img4[3079:3072];
      img_out4[39:32] = img4[3087:3080];
      img_out4[47:40] = img4[3095:3088];
      img_out4[55:48] = img4[3103:3096];
      img_out4[63:56] = img4[3111:3104];
      img_out4[71:64] = img4[3119:3112];
      img_out4[79:72] = img4[3127:3120];
      img_out4[87:80] = img4[3135:3128];
      img_out4[95:88] = img4[3143:3136];
      img_out4[103:96] = img4[3151:3144];
      img_out4[111:104] = img4[3159:3152];
      img_out4[119:112] = img4[3167:3160];
      img_out4[127:120] = img4[3175:3168];
      img_out4[135:128] = img4[3183:3176];
      img_out4[143:136] = img4[3191:3184];
      img_out4[151:144] = img4[3199:3192];
      img_out4[159:152] = img4[3207:3200];
      img_out4[167:160] = img4[3215:3208];
      img_out4[175:168] = img4[3223:3216];
    end
    'd25: begin
      img_out0[7:0] = img0[3183:3176];
      img_out0[15:8] = img0[3191:3184];
      img_out0[23:16] = img0[3199:3192];
      img_out0[31:24] = img0[3207:3200];
      img_out0[39:32] = img0[3215:3208];
      img_out0[47:40] = img0[3223:3216];
      img_out0[55:48] = img0[3231:3224];
      img_out0[63:56] = img0[3239:3232];
      img_out0[71:64] = img0[3247:3240];
      img_out0[79:72] = img0[3255:3248];
      img_out0[87:80] = img0[3263:3256];
      img_out0[95:88] = img0[3271:3264];
      img_out0[103:96] = img0[3279:3272];
      img_out0[111:104] = img0[3287:3280];
      img_out0[119:112] = img0[3295:3288];
      img_out0[127:120] = img0[3303:3296];
      img_out0[135:128] = img0[3311:3304];
      img_out0[143:136] = img0[3319:3312];
      img_out0[151:144] = img0[3327:3320];
      img_out0[159:152] = img0[3335:3328];
      img_out0[167:160] = img0[3343:3336];
      img_out0[175:168] = img0[3351:3344];
      img_out1[7:0] = img1[3183:3176];
      img_out1[15:8] = img1[3191:3184];
      img_out1[23:16] = img1[3199:3192];
      img_out1[31:24] = img1[3207:3200];
      img_out1[39:32] = img1[3215:3208];
      img_out1[47:40] = img1[3223:3216];
      img_out1[55:48] = img1[3231:3224];
      img_out1[63:56] = img1[3239:3232];
      img_out1[71:64] = img1[3247:3240];
      img_out1[79:72] = img1[3255:3248];
      img_out1[87:80] = img1[3263:3256];
      img_out1[95:88] = img1[3271:3264];
      img_out1[103:96] = img1[3279:3272];
      img_out1[111:104] = img1[3287:3280];
      img_out1[119:112] = img1[3295:3288];
      img_out1[127:120] = img1[3303:3296];
      img_out1[135:128] = img1[3311:3304];
      img_out1[143:136] = img1[3319:3312];
      img_out1[151:144] = img1[3327:3320];
      img_out1[159:152] = img1[3335:3328];
      img_out1[167:160] = img1[3343:3336];
      img_out1[175:168] = img1[3351:3344];
      img_out2[7:0] = img2[3183:3176];
      img_out2[15:8] = img2[3191:3184];
      img_out2[23:16] = img2[3199:3192];
      img_out2[31:24] = img2[3207:3200];
      img_out2[39:32] = img2[3215:3208];
      img_out2[47:40] = img2[3223:3216];
      img_out2[55:48] = img2[3231:3224];
      img_out2[63:56] = img2[3239:3232];
      img_out2[71:64] = img2[3247:3240];
      img_out2[79:72] = img2[3255:3248];
      img_out2[87:80] = img2[3263:3256];
      img_out2[95:88] = img2[3271:3264];
      img_out2[103:96] = img2[3279:3272];
      img_out2[111:104] = img2[3287:3280];
      img_out2[119:112] = img2[3295:3288];
      img_out2[127:120] = img2[3303:3296];
      img_out2[135:128] = img2[3311:3304];
      img_out2[143:136] = img2[3319:3312];
      img_out2[151:144] = img2[3327:3320];
      img_out2[159:152] = img2[3335:3328];
      img_out2[167:160] = img2[3343:3336];
      img_out2[175:168] = img2[3351:3344];
      img_out3[7:0] = img3[3183:3176];
      img_out3[15:8] = img3[3191:3184];
      img_out3[23:16] = img3[3199:3192];
      img_out3[31:24] = img3[3207:3200];
      img_out3[39:32] = img3[3215:3208];
      img_out3[47:40] = img3[3223:3216];
      img_out3[55:48] = img3[3231:3224];
      img_out3[63:56] = img3[3239:3232];
      img_out3[71:64] = img3[3247:3240];
      img_out3[79:72] = img3[3255:3248];
      img_out3[87:80] = img3[3263:3256];
      img_out3[95:88] = img3[3271:3264];
      img_out3[103:96] = img3[3279:3272];
      img_out3[111:104] = img3[3287:3280];
      img_out3[119:112] = img3[3295:3288];
      img_out3[127:120] = img3[3303:3296];
      img_out3[135:128] = img3[3311:3304];
      img_out3[143:136] = img3[3319:3312];
      img_out3[151:144] = img3[3327:3320];
      img_out3[159:152] = img3[3335:3328];
      img_out3[167:160] = img3[3343:3336];
      img_out3[175:168] = img3[3351:3344];
      img_out4[7:0] = img4[3183:3176];
      img_out4[15:8] = img4[3191:3184];
      img_out4[23:16] = img4[3199:3192];
      img_out4[31:24] = img4[3207:3200];
      img_out4[39:32] = img4[3215:3208];
      img_out4[47:40] = img4[3223:3216];
      img_out4[55:48] = img4[3231:3224];
      img_out4[63:56] = img4[3239:3232];
      img_out4[71:64] = img4[3247:3240];
      img_out4[79:72] = img4[3255:3248];
      img_out4[87:80] = img4[3263:3256];
      img_out4[95:88] = img4[3271:3264];
      img_out4[103:96] = img4[3279:3272];
      img_out4[111:104] = img4[3287:3280];
      img_out4[119:112] = img4[3295:3288];
      img_out4[127:120] = img4[3303:3296];
      img_out4[135:128] = img4[3311:3304];
      img_out4[143:136] = img4[3319:3312];
      img_out4[151:144] = img4[3327:3320];
      img_out4[159:152] = img4[3335:3328];
      img_out4[167:160] = img4[3343:3336];
      img_out4[175:168] = img4[3351:3344];
    end
    'd26: begin
      img_out0[7:0] = img0[3311:3304];
      img_out0[15:8] = img0[3319:3312];
      img_out0[23:16] = img0[3327:3320];
      img_out0[31:24] = img0[3335:3328];
      img_out0[39:32] = img0[3343:3336];
      img_out0[47:40] = img0[3351:3344];
      img_out0[55:48] = img0[3359:3352];
      img_out0[63:56] = img0[3367:3360];
      img_out0[71:64] = img0[3375:3368];
      img_out0[79:72] = img0[3383:3376];
      img_out0[87:80] = img0[3391:3384];
      img_out0[95:88] = img0[3399:3392];
      img_out0[103:96] = img0[3407:3400];
      img_out0[111:104] = img0[3415:3408];
      img_out0[119:112] = img0[3423:3416];
      img_out0[127:120] = img0[3431:3424];
      img_out0[135:128] = img0[3439:3432];
      img_out0[143:136] = img0[3447:3440];
      img_out0[151:144] = img0[3455:3448];
      img_out0[159:152] = img0[3463:3456];
      img_out0[167:160] = img0[3471:3464];
      img_out0[175:168] = img0[3479:3472];
      img_out1[7:0] = img1[3311:3304];
      img_out1[15:8] = img1[3319:3312];
      img_out1[23:16] = img1[3327:3320];
      img_out1[31:24] = img1[3335:3328];
      img_out1[39:32] = img1[3343:3336];
      img_out1[47:40] = img1[3351:3344];
      img_out1[55:48] = img1[3359:3352];
      img_out1[63:56] = img1[3367:3360];
      img_out1[71:64] = img1[3375:3368];
      img_out1[79:72] = img1[3383:3376];
      img_out1[87:80] = img1[3391:3384];
      img_out1[95:88] = img1[3399:3392];
      img_out1[103:96] = img1[3407:3400];
      img_out1[111:104] = img1[3415:3408];
      img_out1[119:112] = img1[3423:3416];
      img_out1[127:120] = img1[3431:3424];
      img_out1[135:128] = img1[3439:3432];
      img_out1[143:136] = img1[3447:3440];
      img_out1[151:144] = img1[3455:3448];
      img_out1[159:152] = img1[3463:3456];
      img_out1[167:160] = img1[3471:3464];
      img_out1[175:168] = img1[3479:3472];
      img_out2[7:0] = img2[3311:3304];
      img_out2[15:8] = img2[3319:3312];
      img_out2[23:16] = img2[3327:3320];
      img_out2[31:24] = img2[3335:3328];
      img_out2[39:32] = img2[3343:3336];
      img_out2[47:40] = img2[3351:3344];
      img_out2[55:48] = img2[3359:3352];
      img_out2[63:56] = img2[3367:3360];
      img_out2[71:64] = img2[3375:3368];
      img_out2[79:72] = img2[3383:3376];
      img_out2[87:80] = img2[3391:3384];
      img_out2[95:88] = img2[3399:3392];
      img_out2[103:96] = img2[3407:3400];
      img_out2[111:104] = img2[3415:3408];
      img_out2[119:112] = img2[3423:3416];
      img_out2[127:120] = img2[3431:3424];
      img_out2[135:128] = img2[3439:3432];
      img_out2[143:136] = img2[3447:3440];
      img_out2[151:144] = img2[3455:3448];
      img_out2[159:152] = img2[3463:3456];
      img_out2[167:160] = img2[3471:3464];
      img_out2[175:168] = img2[3479:3472];
      img_out3[7:0] = img3[3311:3304];
      img_out3[15:8] = img3[3319:3312];
      img_out3[23:16] = img3[3327:3320];
      img_out3[31:24] = img3[3335:3328];
      img_out3[39:32] = img3[3343:3336];
      img_out3[47:40] = img3[3351:3344];
      img_out3[55:48] = img3[3359:3352];
      img_out3[63:56] = img3[3367:3360];
      img_out3[71:64] = img3[3375:3368];
      img_out3[79:72] = img3[3383:3376];
      img_out3[87:80] = img3[3391:3384];
      img_out3[95:88] = img3[3399:3392];
      img_out3[103:96] = img3[3407:3400];
      img_out3[111:104] = img3[3415:3408];
      img_out3[119:112] = img3[3423:3416];
      img_out3[127:120] = img3[3431:3424];
      img_out3[135:128] = img3[3439:3432];
      img_out3[143:136] = img3[3447:3440];
      img_out3[151:144] = img3[3455:3448];
      img_out3[159:152] = img3[3463:3456];
      img_out3[167:160] = img3[3471:3464];
      img_out3[175:168] = img3[3479:3472];
      img_out4[7:0] = img4[3311:3304];
      img_out4[15:8] = img4[3319:3312];
      img_out4[23:16] = img4[3327:3320];
      img_out4[31:24] = img4[3335:3328];
      img_out4[39:32] = img4[3343:3336];
      img_out4[47:40] = img4[3351:3344];
      img_out4[55:48] = img4[3359:3352];
      img_out4[63:56] = img4[3367:3360];
      img_out4[71:64] = img4[3375:3368];
      img_out4[79:72] = img4[3383:3376];
      img_out4[87:80] = img4[3391:3384];
      img_out4[95:88] = img4[3399:3392];
      img_out4[103:96] = img4[3407:3400];
      img_out4[111:104] = img4[3415:3408];
      img_out4[119:112] = img4[3423:3416];
      img_out4[127:120] = img4[3431:3424];
      img_out4[135:128] = img4[3439:3432];
      img_out4[143:136] = img4[3447:3440];
      img_out4[151:144] = img4[3455:3448];
      img_out4[159:152] = img4[3463:3456];
      img_out4[167:160] = img4[3471:3464];
      img_out4[175:168] = img4[3479:3472];
    end
    'd27: begin
      img_out0[7:0] = img0[3439:3432];
      img_out0[15:8] = img0[3447:3440];
      img_out0[23:16] = img0[3455:3448];
      img_out0[31:24] = img0[3463:3456];
      img_out0[39:32] = img0[3471:3464];
      img_out0[47:40] = img0[3479:3472];
      img_out0[55:48] = img0[3487:3480];
      img_out0[63:56] = img0[3495:3488];
      img_out0[71:64] = img0[3503:3496];
      img_out0[79:72] = img0[3511:3504];
      img_out0[87:80] = img0[3519:3512];
      img_out0[95:88] = img0[3527:3520];
      img_out0[103:96] = img0[3535:3528];
      img_out0[111:104] = img0[3543:3536];
      img_out0[119:112] = img0[3551:3544];
      img_out0[127:120] = img0[3559:3552];
      img_out0[135:128] = img0[3567:3560];
      img_out0[143:136] = img0[3575:3568];
      img_out0[151:144] = img0[3583:3576];
      img_out0[159:152] = img0[3591:3584];
      img_out0[167:160] = img0[3599:3592];
      img_out0[175:168] = img0[3607:3600];
      img_out1[7:0] = img1[3439:3432];
      img_out1[15:8] = img1[3447:3440];
      img_out1[23:16] = img1[3455:3448];
      img_out1[31:24] = img1[3463:3456];
      img_out1[39:32] = img1[3471:3464];
      img_out1[47:40] = img1[3479:3472];
      img_out1[55:48] = img1[3487:3480];
      img_out1[63:56] = img1[3495:3488];
      img_out1[71:64] = img1[3503:3496];
      img_out1[79:72] = img1[3511:3504];
      img_out1[87:80] = img1[3519:3512];
      img_out1[95:88] = img1[3527:3520];
      img_out1[103:96] = img1[3535:3528];
      img_out1[111:104] = img1[3543:3536];
      img_out1[119:112] = img1[3551:3544];
      img_out1[127:120] = img1[3559:3552];
      img_out1[135:128] = img1[3567:3560];
      img_out1[143:136] = img1[3575:3568];
      img_out1[151:144] = img1[3583:3576];
      img_out1[159:152] = img1[3591:3584];
      img_out1[167:160] = img1[3599:3592];
      img_out1[175:168] = img1[3607:3600];
      img_out2[7:0] = img2[3439:3432];
      img_out2[15:8] = img2[3447:3440];
      img_out2[23:16] = img2[3455:3448];
      img_out2[31:24] = img2[3463:3456];
      img_out2[39:32] = img2[3471:3464];
      img_out2[47:40] = img2[3479:3472];
      img_out2[55:48] = img2[3487:3480];
      img_out2[63:56] = img2[3495:3488];
      img_out2[71:64] = img2[3503:3496];
      img_out2[79:72] = img2[3511:3504];
      img_out2[87:80] = img2[3519:3512];
      img_out2[95:88] = img2[3527:3520];
      img_out2[103:96] = img2[3535:3528];
      img_out2[111:104] = img2[3543:3536];
      img_out2[119:112] = img2[3551:3544];
      img_out2[127:120] = img2[3559:3552];
      img_out2[135:128] = img2[3567:3560];
      img_out2[143:136] = img2[3575:3568];
      img_out2[151:144] = img2[3583:3576];
      img_out2[159:152] = img2[3591:3584];
      img_out2[167:160] = img2[3599:3592];
      img_out2[175:168] = img2[3607:3600];
      img_out3[7:0] = img3[3439:3432];
      img_out3[15:8] = img3[3447:3440];
      img_out3[23:16] = img3[3455:3448];
      img_out3[31:24] = img3[3463:3456];
      img_out3[39:32] = img3[3471:3464];
      img_out3[47:40] = img3[3479:3472];
      img_out3[55:48] = img3[3487:3480];
      img_out3[63:56] = img3[3495:3488];
      img_out3[71:64] = img3[3503:3496];
      img_out3[79:72] = img3[3511:3504];
      img_out3[87:80] = img3[3519:3512];
      img_out3[95:88] = img3[3527:3520];
      img_out3[103:96] = img3[3535:3528];
      img_out3[111:104] = img3[3543:3536];
      img_out3[119:112] = img3[3551:3544];
      img_out3[127:120] = img3[3559:3552];
      img_out3[135:128] = img3[3567:3560];
      img_out3[143:136] = img3[3575:3568];
      img_out3[151:144] = img3[3583:3576];
      img_out3[159:152] = img3[3591:3584];
      img_out3[167:160] = img3[3599:3592];
      img_out3[175:168] = img3[3607:3600];
      img_out4[7:0] = img4[3439:3432];
      img_out4[15:8] = img4[3447:3440];
      img_out4[23:16] = img4[3455:3448];
      img_out4[31:24] = img4[3463:3456];
      img_out4[39:32] = img4[3471:3464];
      img_out4[47:40] = img4[3479:3472];
      img_out4[55:48] = img4[3487:3480];
      img_out4[63:56] = img4[3495:3488];
      img_out4[71:64] = img4[3503:3496];
      img_out4[79:72] = img4[3511:3504];
      img_out4[87:80] = img4[3519:3512];
      img_out4[95:88] = img4[3527:3520];
      img_out4[103:96] = img4[3535:3528];
      img_out4[111:104] = img4[3543:3536];
      img_out4[119:112] = img4[3551:3544];
      img_out4[127:120] = img4[3559:3552];
      img_out4[135:128] = img4[3567:3560];
      img_out4[143:136] = img4[3575:3568];
      img_out4[151:144] = img4[3583:3576];
      img_out4[159:152] = img4[3591:3584];
      img_out4[167:160] = img4[3599:3592];
      img_out4[175:168] = img4[3607:3600];
    end
    'd28: begin
      img_out0[7:0] = img0[3567:3560];
      img_out0[15:8] = img0[3575:3568];
      img_out0[23:16] = img0[3583:3576];
      img_out0[31:24] = img0[3591:3584];
      img_out0[39:32] = img0[3599:3592];
      img_out0[47:40] = img0[3607:3600];
      img_out0[55:48] = img0[3615:3608];
      img_out0[63:56] = img0[3623:3616];
      img_out0[71:64] = img0[3631:3624];
      img_out0[79:72] = img0[3639:3632];
      img_out0[87:80] = img0[3647:3640];
      img_out0[95:88] = img0[3655:3648];
      img_out0[103:96] = img0[3663:3656];
      img_out0[111:104] = img0[3671:3664];
      img_out0[119:112] = img0[3679:3672];
      img_out0[127:120] = img0[3687:3680];
      img_out0[135:128] = img0[3695:3688];
      img_out0[143:136] = img0[3703:3696];
      img_out0[151:144] = img0[3711:3704];
      img_out0[159:152] = img0[3719:3712];
      img_out0[167:160] = img0[3727:3720];
      img_out0[175:168] = img0[3735:3728];
      img_out1[7:0] = img1[3567:3560];
      img_out1[15:8] = img1[3575:3568];
      img_out1[23:16] = img1[3583:3576];
      img_out1[31:24] = img1[3591:3584];
      img_out1[39:32] = img1[3599:3592];
      img_out1[47:40] = img1[3607:3600];
      img_out1[55:48] = img1[3615:3608];
      img_out1[63:56] = img1[3623:3616];
      img_out1[71:64] = img1[3631:3624];
      img_out1[79:72] = img1[3639:3632];
      img_out1[87:80] = img1[3647:3640];
      img_out1[95:88] = img1[3655:3648];
      img_out1[103:96] = img1[3663:3656];
      img_out1[111:104] = img1[3671:3664];
      img_out1[119:112] = img1[3679:3672];
      img_out1[127:120] = img1[3687:3680];
      img_out1[135:128] = img1[3695:3688];
      img_out1[143:136] = img1[3703:3696];
      img_out1[151:144] = img1[3711:3704];
      img_out1[159:152] = img1[3719:3712];
      img_out1[167:160] = img1[3727:3720];
      img_out1[175:168] = img1[3735:3728];
      img_out2[7:0] = img2[3567:3560];
      img_out2[15:8] = img2[3575:3568];
      img_out2[23:16] = img2[3583:3576];
      img_out2[31:24] = img2[3591:3584];
      img_out2[39:32] = img2[3599:3592];
      img_out2[47:40] = img2[3607:3600];
      img_out2[55:48] = img2[3615:3608];
      img_out2[63:56] = img2[3623:3616];
      img_out2[71:64] = img2[3631:3624];
      img_out2[79:72] = img2[3639:3632];
      img_out2[87:80] = img2[3647:3640];
      img_out2[95:88] = img2[3655:3648];
      img_out2[103:96] = img2[3663:3656];
      img_out2[111:104] = img2[3671:3664];
      img_out2[119:112] = img2[3679:3672];
      img_out2[127:120] = img2[3687:3680];
      img_out2[135:128] = img2[3695:3688];
      img_out2[143:136] = img2[3703:3696];
      img_out2[151:144] = img2[3711:3704];
      img_out2[159:152] = img2[3719:3712];
      img_out2[167:160] = img2[3727:3720];
      img_out2[175:168] = img2[3735:3728];
      img_out3[7:0] = img3[3567:3560];
      img_out3[15:8] = img3[3575:3568];
      img_out3[23:16] = img3[3583:3576];
      img_out3[31:24] = img3[3591:3584];
      img_out3[39:32] = img3[3599:3592];
      img_out3[47:40] = img3[3607:3600];
      img_out3[55:48] = img3[3615:3608];
      img_out3[63:56] = img3[3623:3616];
      img_out3[71:64] = img3[3631:3624];
      img_out3[79:72] = img3[3639:3632];
      img_out3[87:80] = img3[3647:3640];
      img_out3[95:88] = img3[3655:3648];
      img_out3[103:96] = img3[3663:3656];
      img_out3[111:104] = img3[3671:3664];
      img_out3[119:112] = img3[3679:3672];
      img_out3[127:120] = img3[3687:3680];
      img_out3[135:128] = img3[3695:3688];
      img_out3[143:136] = img3[3703:3696];
      img_out3[151:144] = img3[3711:3704];
      img_out3[159:152] = img3[3719:3712];
      img_out3[167:160] = img3[3727:3720];
      img_out3[175:168] = img3[3735:3728];
      img_out4[7:0] = img4[3567:3560];
      img_out4[15:8] = img4[3575:3568];
      img_out4[23:16] = img4[3583:3576];
      img_out4[31:24] = img4[3591:3584];
      img_out4[39:32] = img4[3599:3592];
      img_out4[47:40] = img4[3607:3600];
      img_out4[55:48] = img4[3615:3608];
      img_out4[63:56] = img4[3623:3616];
      img_out4[71:64] = img4[3631:3624];
      img_out4[79:72] = img4[3639:3632];
      img_out4[87:80] = img4[3647:3640];
      img_out4[95:88] = img4[3655:3648];
      img_out4[103:96] = img4[3663:3656];
      img_out4[111:104] = img4[3671:3664];
      img_out4[119:112] = img4[3679:3672];
      img_out4[127:120] = img4[3687:3680];
      img_out4[135:128] = img4[3695:3688];
      img_out4[143:136] = img4[3703:3696];
      img_out4[151:144] = img4[3711:3704];
      img_out4[159:152] = img4[3719:3712];
      img_out4[167:160] = img4[3727:3720];
      img_out4[175:168] = img4[3735:3728];
    end
    'd29: begin
      img_out0[7:0] = img0[3695:3688];
      img_out0[15:8] = img0[3703:3696];
      img_out0[23:16] = img0[3711:3704];
      img_out0[31:24] = img0[3719:3712];
      img_out0[39:32] = img0[3727:3720];
      img_out0[47:40] = img0[3735:3728];
      img_out0[55:48] = img0[3743:3736];
      img_out0[63:56] = img0[3751:3744];
      img_out0[71:64] = img0[3759:3752];
      img_out0[79:72] = img0[3767:3760];
      img_out0[87:80] = img0[3775:3768];
      img_out0[95:88] = img0[3783:3776];
      img_out0[103:96] = img0[3791:3784];
      img_out0[111:104] = img0[3799:3792];
      img_out0[119:112] = img0[3807:3800];
      img_out0[127:120] = img0[3815:3808];
      img_out0[135:128] = img0[3823:3816];
      img_out0[143:136] = img0[3831:3824];
      img_out0[151:144] = img0[3839:3832];
      img_out0[159:152] = img0[3847:3840];
      img_out0[167:160] = img0[3855:3848];
      img_out0[175:168] = img0[3863:3856];
      img_out1[7:0] = img1[3695:3688];
      img_out1[15:8] = img1[3703:3696];
      img_out1[23:16] = img1[3711:3704];
      img_out1[31:24] = img1[3719:3712];
      img_out1[39:32] = img1[3727:3720];
      img_out1[47:40] = img1[3735:3728];
      img_out1[55:48] = img1[3743:3736];
      img_out1[63:56] = img1[3751:3744];
      img_out1[71:64] = img1[3759:3752];
      img_out1[79:72] = img1[3767:3760];
      img_out1[87:80] = img1[3775:3768];
      img_out1[95:88] = img1[3783:3776];
      img_out1[103:96] = img1[3791:3784];
      img_out1[111:104] = img1[3799:3792];
      img_out1[119:112] = img1[3807:3800];
      img_out1[127:120] = img1[3815:3808];
      img_out1[135:128] = img1[3823:3816];
      img_out1[143:136] = img1[3831:3824];
      img_out1[151:144] = img1[3839:3832];
      img_out1[159:152] = img1[3847:3840];
      img_out1[167:160] = img1[3855:3848];
      img_out1[175:168] = img1[3863:3856];
      img_out2[7:0] = img2[3695:3688];
      img_out2[15:8] = img2[3703:3696];
      img_out2[23:16] = img2[3711:3704];
      img_out2[31:24] = img2[3719:3712];
      img_out2[39:32] = img2[3727:3720];
      img_out2[47:40] = img2[3735:3728];
      img_out2[55:48] = img2[3743:3736];
      img_out2[63:56] = img2[3751:3744];
      img_out2[71:64] = img2[3759:3752];
      img_out2[79:72] = img2[3767:3760];
      img_out2[87:80] = img2[3775:3768];
      img_out2[95:88] = img2[3783:3776];
      img_out2[103:96] = img2[3791:3784];
      img_out2[111:104] = img2[3799:3792];
      img_out2[119:112] = img2[3807:3800];
      img_out2[127:120] = img2[3815:3808];
      img_out2[135:128] = img2[3823:3816];
      img_out2[143:136] = img2[3831:3824];
      img_out2[151:144] = img2[3839:3832];
      img_out2[159:152] = img2[3847:3840];
      img_out2[167:160] = img2[3855:3848];
      img_out2[175:168] = img2[3863:3856];
      img_out3[7:0] = img3[3695:3688];
      img_out3[15:8] = img3[3703:3696];
      img_out3[23:16] = img3[3711:3704];
      img_out3[31:24] = img3[3719:3712];
      img_out3[39:32] = img3[3727:3720];
      img_out3[47:40] = img3[3735:3728];
      img_out3[55:48] = img3[3743:3736];
      img_out3[63:56] = img3[3751:3744];
      img_out3[71:64] = img3[3759:3752];
      img_out3[79:72] = img3[3767:3760];
      img_out3[87:80] = img3[3775:3768];
      img_out3[95:88] = img3[3783:3776];
      img_out3[103:96] = img3[3791:3784];
      img_out3[111:104] = img3[3799:3792];
      img_out3[119:112] = img3[3807:3800];
      img_out3[127:120] = img3[3815:3808];
      img_out3[135:128] = img3[3823:3816];
      img_out3[143:136] = img3[3831:3824];
      img_out3[151:144] = img3[3839:3832];
      img_out3[159:152] = img3[3847:3840];
      img_out3[167:160] = img3[3855:3848];
      img_out3[175:168] = img3[3863:3856];
      img_out4[7:0] = img4[3695:3688];
      img_out4[15:8] = img4[3703:3696];
      img_out4[23:16] = img4[3711:3704];
      img_out4[31:24] = img4[3719:3712];
      img_out4[39:32] = img4[3727:3720];
      img_out4[47:40] = img4[3735:3728];
      img_out4[55:48] = img4[3743:3736];
      img_out4[63:56] = img4[3751:3744];
      img_out4[71:64] = img4[3759:3752];
      img_out4[79:72] = img4[3767:3760];
      img_out4[87:80] = img4[3775:3768];
      img_out4[95:88] = img4[3783:3776];
      img_out4[103:96] = img4[3791:3784];
      img_out4[111:104] = img4[3799:3792];
      img_out4[119:112] = img4[3807:3800];
      img_out4[127:120] = img4[3815:3808];
      img_out4[135:128] = img4[3823:3816];
      img_out4[143:136] = img4[3831:3824];
      img_out4[151:144] = img4[3839:3832];
      img_out4[159:152] = img4[3847:3840];
      img_out4[167:160] = img4[3855:3848];
      img_out4[175:168] = img4[3863:3856];
    end
    'd30: begin
      img_out0[7:0] = img0[3823:3816];
      img_out0[15:8] = img0[3831:3824];
      img_out0[23:16] = img0[3839:3832];
      img_out0[31:24] = img0[3847:3840];
      img_out0[39:32] = img0[3855:3848];
      img_out0[47:40] = img0[3863:3856];
      img_out0[55:48] = img0[3871:3864];
      img_out0[63:56] = img0[3879:3872];
      img_out0[71:64] = img0[3887:3880];
      img_out0[79:72] = img0[3895:3888];
      img_out0[87:80] = img0[3903:3896];
      img_out0[95:88] = img0[3911:3904];
      img_out0[103:96] = img0[3919:3912];
      img_out0[111:104] = img0[3927:3920];
      img_out0[119:112] = img0[3935:3928];
      img_out0[127:120] = img0[3943:3936];
      img_out0[135:128] = img0[3951:3944];
      img_out0[143:136] = img0[3959:3952];
      img_out0[151:144] = img0[3967:3960];
      img_out0[159:152] = img0[3975:3968];
      img_out0[167:160] = img0[3983:3976];
      img_out0[175:168] = img0[3991:3984];
      img_out1[7:0] = img1[3823:3816];
      img_out1[15:8] = img1[3831:3824];
      img_out1[23:16] = img1[3839:3832];
      img_out1[31:24] = img1[3847:3840];
      img_out1[39:32] = img1[3855:3848];
      img_out1[47:40] = img1[3863:3856];
      img_out1[55:48] = img1[3871:3864];
      img_out1[63:56] = img1[3879:3872];
      img_out1[71:64] = img1[3887:3880];
      img_out1[79:72] = img1[3895:3888];
      img_out1[87:80] = img1[3903:3896];
      img_out1[95:88] = img1[3911:3904];
      img_out1[103:96] = img1[3919:3912];
      img_out1[111:104] = img1[3927:3920];
      img_out1[119:112] = img1[3935:3928];
      img_out1[127:120] = img1[3943:3936];
      img_out1[135:128] = img1[3951:3944];
      img_out1[143:136] = img1[3959:3952];
      img_out1[151:144] = img1[3967:3960];
      img_out1[159:152] = img1[3975:3968];
      img_out1[167:160] = img1[3983:3976];
      img_out1[175:168] = img1[3991:3984];
      img_out2[7:0] = img2[3823:3816];
      img_out2[15:8] = img2[3831:3824];
      img_out2[23:16] = img2[3839:3832];
      img_out2[31:24] = img2[3847:3840];
      img_out2[39:32] = img2[3855:3848];
      img_out2[47:40] = img2[3863:3856];
      img_out2[55:48] = img2[3871:3864];
      img_out2[63:56] = img2[3879:3872];
      img_out2[71:64] = img2[3887:3880];
      img_out2[79:72] = img2[3895:3888];
      img_out2[87:80] = img2[3903:3896];
      img_out2[95:88] = img2[3911:3904];
      img_out2[103:96] = img2[3919:3912];
      img_out2[111:104] = img2[3927:3920];
      img_out2[119:112] = img2[3935:3928];
      img_out2[127:120] = img2[3943:3936];
      img_out2[135:128] = img2[3951:3944];
      img_out2[143:136] = img2[3959:3952];
      img_out2[151:144] = img2[3967:3960];
      img_out2[159:152] = img2[3975:3968];
      img_out2[167:160] = img2[3983:3976];
      img_out2[175:168] = img2[3991:3984];
      img_out3[7:0] = img3[3823:3816];
      img_out3[15:8] = img3[3831:3824];
      img_out3[23:16] = img3[3839:3832];
      img_out3[31:24] = img3[3847:3840];
      img_out3[39:32] = img3[3855:3848];
      img_out3[47:40] = img3[3863:3856];
      img_out3[55:48] = img3[3871:3864];
      img_out3[63:56] = img3[3879:3872];
      img_out3[71:64] = img3[3887:3880];
      img_out3[79:72] = img3[3895:3888];
      img_out3[87:80] = img3[3903:3896];
      img_out3[95:88] = img3[3911:3904];
      img_out3[103:96] = img3[3919:3912];
      img_out3[111:104] = img3[3927:3920];
      img_out3[119:112] = img3[3935:3928];
      img_out3[127:120] = img3[3943:3936];
      img_out3[135:128] = img3[3951:3944];
      img_out3[143:136] = img3[3959:3952];
      img_out3[151:144] = img3[3967:3960];
      img_out3[159:152] = img3[3975:3968];
      img_out3[167:160] = img3[3983:3976];
      img_out3[175:168] = img3[3991:3984];
      img_out4[7:0] = img4[3823:3816];
      img_out4[15:8] = img4[3831:3824];
      img_out4[23:16] = img4[3839:3832];
      img_out4[31:24] = img4[3847:3840];
      img_out4[39:32] = img4[3855:3848];
      img_out4[47:40] = img4[3863:3856];
      img_out4[55:48] = img4[3871:3864];
      img_out4[63:56] = img4[3879:3872];
      img_out4[71:64] = img4[3887:3880];
      img_out4[79:72] = img4[3895:3888];
      img_out4[87:80] = img4[3903:3896];
      img_out4[95:88] = img4[3911:3904];
      img_out4[103:96] = img4[3919:3912];
      img_out4[111:104] = img4[3927:3920];
      img_out4[119:112] = img4[3935:3928];
      img_out4[127:120] = img4[3943:3936];
      img_out4[135:128] = img4[3951:3944];
      img_out4[143:136] = img4[3959:3952];
      img_out4[151:144] = img4[3967:3960];
      img_out4[159:152] = img4[3975:3968];
      img_out4[167:160] = img4[3983:3976];
      img_out4[175:168] = img4[3991:3984];
    end
    'd31: begin
      img_out0[7:0] = img0[3951:3944];
      img_out0[15:8] = img0[3959:3952];
      img_out0[23:16] = img0[3967:3960];
      img_out0[31:24] = img0[3975:3968];
      img_out0[39:32] = img0[3983:3976];
      img_out0[47:40] = img0[3991:3984];
      img_out0[55:48] = img0[3999:3992];
      img_out0[63:56] = img0[4007:4000];
      img_out0[71:64] = img0[4015:4008];
      img_out0[79:72] = img0[4023:4016];
      img_out0[87:80] = img0[4031:4024];
      img_out0[95:88] = img0[4039:4032];
      img_out0[103:96] = img0[4047:4040];
      img_out0[111:104] = img0[4055:4048];
      img_out0[119:112] = img0[4063:4056];
      img_out0[127:120] = img0[4071:4064];
      img_out0[135:128] = img0[4079:4072];
      img_out0[143:136] = img0[4087:4080];
      img_out0[151:144] = img0[4095:4088];
      img_out0[159:152] = img0[4103:4096];
      img_out0[167:160] = img0[4111:4104];
      img_out0[175:168] = img0[4119:4112];
      img_out1[7:0] = img1[3951:3944];
      img_out1[15:8] = img1[3959:3952];
      img_out1[23:16] = img1[3967:3960];
      img_out1[31:24] = img1[3975:3968];
      img_out1[39:32] = img1[3983:3976];
      img_out1[47:40] = img1[3991:3984];
      img_out1[55:48] = img1[3999:3992];
      img_out1[63:56] = img1[4007:4000];
      img_out1[71:64] = img1[4015:4008];
      img_out1[79:72] = img1[4023:4016];
      img_out1[87:80] = img1[4031:4024];
      img_out1[95:88] = img1[4039:4032];
      img_out1[103:96] = img1[4047:4040];
      img_out1[111:104] = img1[4055:4048];
      img_out1[119:112] = img1[4063:4056];
      img_out1[127:120] = img1[4071:4064];
      img_out1[135:128] = img1[4079:4072];
      img_out1[143:136] = img1[4087:4080];
      img_out1[151:144] = img1[4095:4088];
      img_out1[159:152] = img1[4103:4096];
      img_out1[167:160] = img1[4111:4104];
      img_out1[175:168] = img1[4119:4112];
      img_out2[7:0] = img2[3951:3944];
      img_out2[15:8] = img2[3959:3952];
      img_out2[23:16] = img2[3967:3960];
      img_out2[31:24] = img2[3975:3968];
      img_out2[39:32] = img2[3983:3976];
      img_out2[47:40] = img2[3991:3984];
      img_out2[55:48] = img2[3999:3992];
      img_out2[63:56] = img2[4007:4000];
      img_out2[71:64] = img2[4015:4008];
      img_out2[79:72] = img2[4023:4016];
      img_out2[87:80] = img2[4031:4024];
      img_out2[95:88] = img2[4039:4032];
      img_out2[103:96] = img2[4047:4040];
      img_out2[111:104] = img2[4055:4048];
      img_out2[119:112] = img2[4063:4056];
      img_out2[127:120] = img2[4071:4064];
      img_out2[135:128] = img2[4079:4072];
      img_out2[143:136] = img2[4087:4080];
      img_out2[151:144] = img2[4095:4088];
      img_out2[159:152] = img2[4103:4096];
      img_out2[167:160] = img2[4111:4104];
      img_out2[175:168] = img2[4119:4112];
      img_out3[7:0] = img3[3951:3944];
      img_out3[15:8] = img3[3959:3952];
      img_out3[23:16] = img3[3967:3960];
      img_out3[31:24] = img3[3975:3968];
      img_out3[39:32] = img3[3983:3976];
      img_out3[47:40] = img3[3991:3984];
      img_out3[55:48] = img3[3999:3992];
      img_out3[63:56] = img3[4007:4000];
      img_out3[71:64] = img3[4015:4008];
      img_out3[79:72] = img3[4023:4016];
      img_out3[87:80] = img3[4031:4024];
      img_out3[95:88] = img3[4039:4032];
      img_out3[103:96] = img3[4047:4040];
      img_out3[111:104] = img3[4055:4048];
      img_out3[119:112] = img3[4063:4056];
      img_out3[127:120] = img3[4071:4064];
      img_out3[135:128] = img3[4079:4072];
      img_out3[143:136] = img3[4087:4080];
      img_out3[151:144] = img3[4095:4088];
      img_out3[159:152] = img3[4103:4096];
      img_out3[167:160] = img3[4111:4104];
      img_out3[175:168] = img3[4119:4112];
      img_out4[7:0] = img4[3951:3944];
      img_out4[15:8] = img4[3959:3952];
      img_out4[23:16] = img4[3967:3960];
      img_out4[31:24] = img4[3975:3968];
      img_out4[39:32] = img4[3983:3976];
      img_out4[47:40] = img4[3991:3984];
      img_out4[55:48] = img4[3999:3992];
      img_out4[63:56] = img4[4007:4000];
      img_out4[71:64] = img4[4015:4008];
      img_out4[79:72] = img4[4023:4016];
      img_out4[87:80] = img4[4031:4024];
      img_out4[95:88] = img4[4039:4032];
      img_out4[103:96] = img4[4047:4040];
      img_out4[111:104] = img4[4055:4048];
      img_out4[119:112] = img4[4063:4056];
      img_out4[127:120] = img4[4071:4064];
      img_out4[135:128] = img4[4079:4072];
      img_out4[143:136] = img4[4087:4080];
      img_out4[151:144] = img4[4095:4088];
      img_out4[159:152] = img4[4103:4096];
      img_out4[167:160] = img4[4111:4104];
      img_out4[175:168] = img4[4119:4112];
    end
    'd32: begin
      img_out0[7:0] = img0[4079:4072];
      img_out0[15:8] = img0[4087:4080];
      img_out0[23:16] = img0[4095:4088];
      img_out0[31:24] = img0[4103:4096];
      img_out0[39:32] = img0[4111:4104];
      img_out0[47:40] = img0[4119:4112];
      img_out0[55:48] = img0[4127:4120];
      img_out0[63:56] = img0[4135:4128];
      img_out0[71:64] = img0[4143:4136];
      img_out0[79:72] = img0[4151:4144];
      img_out0[87:80] = img0[4159:4152];
      img_out0[95:88] = img0[4167:4160];
      img_out0[103:96] = img0[4175:4168];
      img_out0[111:104] = img0[4183:4176];
      img_out0[119:112] = img0[4191:4184];
      img_out0[127:120] = img0[4199:4192];
      img_out0[135:128] = img0[4207:4200];
      img_out0[143:136] = img0[4215:4208];
      img_out0[151:144] = img0[4223:4216];
      img_out0[159:152] = img0[4231:4224];
      img_out0[167:160] = img0[4239:4232];
      img_out0[175:168] = img0[4247:4240];
      img_out1[7:0] = img1[4079:4072];
      img_out1[15:8] = img1[4087:4080];
      img_out1[23:16] = img1[4095:4088];
      img_out1[31:24] = img1[4103:4096];
      img_out1[39:32] = img1[4111:4104];
      img_out1[47:40] = img1[4119:4112];
      img_out1[55:48] = img1[4127:4120];
      img_out1[63:56] = img1[4135:4128];
      img_out1[71:64] = img1[4143:4136];
      img_out1[79:72] = img1[4151:4144];
      img_out1[87:80] = img1[4159:4152];
      img_out1[95:88] = img1[4167:4160];
      img_out1[103:96] = img1[4175:4168];
      img_out1[111:104] = img1[4183:4176];
      img_out1[119:112] = img1[4191:4184];
      img_out1[127:120] = img1[4199:4192];
      img_out1[135:128] = img1[4207:4200];
      img_out1[143:136] = img1[4215:4208];
      img_out1[151:144] = img1[4223:4216];
      img_out1[159:152] = img1[4231:4224];
      img_out1[167:160] = img1[4239:4232];
      img_out1[175:168] = img1[4247:4240];
      img_out2[7:0] = img2[4079:4072];
      img_out2[15:8] = img2[4087:4080];
      img_out2[23:16] = img2[4095:4088];
      img_out2[31:24] = img2[4103:4096];
      img_out2[39:32] = img2[4111:4104];
      img_out2[47:40] = img2[4119:4112];
      img_out2[55:48] = img2[4127:4120];
      img_out2[63:56] = img2[4135:4128];
      img_out2[71:64] = img2[4143:4136];
      img_out2[79:72] = img2[4151:4144];
      img_out2[87:80] = img2[4159:4152];
      img_out2[95:88] = img2[4167:4160];
      img_out2[103:96] = img2[4175:4168];
      img_out2[111:104] = img2[4183:4176];
      img_out2[119:112] = img2[4191:4184];
      img_out2[127:120] = img2[4199:4192];
      img_out2[135:128] = img2[4207:4200];
      img_out2[143:136] = img2[4215:4208];
      img_out2[151:144] = img2[4223:4216];
      img_out2[159:152] = img2[4231:4224];
      img_out2[167:160] = img2[4239:4232];
      img_out2[175:168] = img2[4247:4240];
      img_out3[7:0] = img3[4079:4072];
      img_out3[15:8] = img3[4087:4080];
      img_out3[23:16] = img3[4095:4088];
      img_out3[31:24] = img3[4103:4096];
      img_out3[39:32] = img3[4111:4104];
      img_out3[47:40] = img3[4119:4112];
      img_out3[55:48] = img3[4127:4120];
      img_out3[63:56] = img3[4135:4128];
      img_out3[71:64] = img3[4143:4136];
      img_out3[79:72] = img3[4151:4144];
      img_out3[87:80] = img3[4159:4152];
      img_out3[95:88] = img3[4167:4160];
      img_out3[103:96] = img3[4175:4168];
      img_out3[111:104] = img3[4183:4176];
      img_out3[119:112] = img3[4191:4184];
      img_out3[127:120] = img3[4199:4192];
      img_out3[135:128] = img3[4207:4200];
      img_out3[143:136] = img3[4215:4208];
      img_out3[151:144] = img3[4223:4216];
      img_out3[159:152] = img3[4231:4224];
      img_out3[167:160] = img3[4239:4232];
      img_out3[175:168] = img3[4247:4240];
      img_out4[7:0] = img4[4079:4072];
      img_out4[15:8] = img4[4087:4080];
      img_out4[23:16] = img4[4095:4088];
      img_out4[31:24] = img4[4103:4096];
      img_out4[39:32] = img4[4111:4104];
      img_out4[47:40] = img4[4119:4112];
      img_out4[55:48] = img4[4127:4120];
      img_out4[63:56] = img4[4135:4128];
      img_out4[71:64] = img4[4143:4136];
      img_out4[79:72] = img4[4151:4144];
      img_out4[87:80] = img4[4159:4152];
      img_out4[95:88] = img4[4167:4160];
      img_out4[103:96] = img4[4175:4168];
      img_out4[111:104] = img4[4183:4176];
      img_out4[119:112] = img4[4191:4184];
      img_out4[127:120] = img4[4199:4192];
      img_out4[135:128] = img4[4207:4200];
      img_out4[143:136] = img4[4215:4208];
      img_out4[151:144] = img4[4223:4216];
      img_out4[159:152] = img4[4231:4224];
      img_out4[167:160] = img4[4239:4232];
      img_out4[175:168] = img4[4247:4240];
    end
    'd33: begin
      img_out0[7:0] = img0[4207:4200];
      img_out0[15:8] = img0[4215:4208];
      img_out0[23:16] = img0[4223:4216];
      img_out0[31:24] = img0[4231:4224];
      img_out0[39:32] = img0[4239:4232];
      img_out0[47:40] = img0[4247:4240];
      img_out0[55:48] = img0[4255:4248];
      img_out0[63:56] = img0[4263:4256];
      img_out0[71:64] = img0[4271:4264];
      img_out0[79:72] = img0[4279:4272];
      img_out0[87:80] = img0[4287:4280];
      img_out0[95:88] = img0[4295:4288];
      img_out0[103:96] = img0[4303:4296];
      img_out0[111:104] = img0[4311:4304];
      img_out0[119:112] = img0[4319:4312];
      img_out0[127:120] = img0[4327:4320];
      img_out0[135:128] = img0[4335:4328];
      img_out0[143:136] = img0[4343:4336];
      img_out0[151:144] = img0[4351:4344];
      img_out0[159:152] = img0[4359:4352];
      img_out0[167:160] = img0[4367:4360];
      img_out0[175:168] = img0[4375:4368];
      img_out1[7:0] = img1[4207:4200];
      img_out1[15:8] = img1[4215:4208];
      img_out1[23:16] = img1[4223:4216];
      img_out1[31:24] = img1[4231:4224];
      img_out1[39:32] = img1[4239:4232];
      img_out1[47:40] = img1[4247:4240];
      img_out1[55:48] = img1[4255:4248];
      img_out1[63:56] = img1[4263:4256];
      img_out1[71:64] = img1[4271:4264];
      img_out1[79:72] = img1[4279:4272];
      img_out1[87:80] = img1[4287:4280];
      img_out1[95:88] = img1[4295:4288];
      img_out1[103:96] = img1[4303:4296];
      img_out1[111:104] = img1[4311:4304];
      img_out1[119:112] = img1[4319:4312];
      img_out1[127:120] = img1[4327:4320];
      img_out1[135:128] = img1[4335:4328];
      img_out1[143:136] = img1[4343:4336];
      img_out1[151:144] = img1[4351:4344];
      img_out1[159:152] = img1[4359:4352];
      img_out1[167:160] = img1[4367:4360];
      img_out1[175:168] = img1[4375:4368];
      img_out2[7:0] = img2[4207:4200];
      img_out2[15:8] = img2[4215:4208];
      img_out2[23:16] = img2[4223:4216];
      img_out2[31:24] = img2[4231:4224];
      img_out2[39:32] = img2[4239:4232];
      img_out2[47:40] = img2[4247:4240];
      img_out2[55:48] = img2[4255:4248];
      img_out2[63:56] = img2[4263:4256];
      img_out2[71:64] = img2[4271:4264];
      img_out2[79:72] = img2[4279:4272];
      img_out2[87:80] = img2[4287:4280];
      img_out2[95:88] = img2[4295:4288];
      img_out2[103:96] = img2[4303:4296];
      img_out2[111:104] = img2[4311:4304];
      img_out2[119:112] = img2[4319:4312];
      img_out2[127:120] = img2[4327:4320];
      img_out2[135:128] = img2[4335:4328];
      img_out2[143:136] = img2[4343:4336];
      img_out2[151:144] = img2[4351:4344];
      img_out2[159:152] = img2[4359:4352];
      img_out2[167:160] = img2[4367:4360];
      img_out2[175:168] = img2[4375:4368];
      img_out3[7:0] = img3[4207:4200];
      img_out3[15:8] = img3[4215:4208];
      img_out3[23:16] = img3[4223:4216];
      img_out3[31:24] = img3[4231:4224];
      img_out3[39:32] = img3[4239:4232];
      img_out3[47:40] = img3[4247:4240];
      img_out3[55:48] = img3[4255:4248];
      img_out3[63:56] = img3[4263:4256];
      img_out3[71:64] = img3[4271:4264];
      img_out3[79:72] = img3[4279:4272];
      img_out3[87:80] = img3[4287:4280];
      img_out3[95:88] = img3[4295:4288];
      img_out3[103:96] = img3[4303:4296];
      img_out3[111:104] = img3[4311:4304];
      img_out3[119:112] = img3[4319:4312];
      img_out3[127:120] = img3[4327:4320];
      img_out3[135:128] = img3[4335:4328];
      img_out3[143:136] = img3[4343:4336];
      img_out3[151:144] = img3[4351:4344];
      img_out3[159:152] = img3[4359:4352];
      img_out3[167:160] = img3[4367:4360];
      img_out3[175:168] = img3[4375:4368];
      img_out4[7:0] = img4[4207:4200];
      img_out4[15:8] = img4[4215:4208];
      img_out4[23:16] = img4[4223:4216];
      img_out4[31:24] = img4[4231:4224];
      img_out4[39:32] = img4[4239:4232];
      img_out4[47:40] = img4[4247:4240];
      img_out4[55:48] = img4[4255:4248];
      img_out4[63:56] = img4[4263:4256];
      img_out4[71:64] = img4[4271:4264];
      img_out4[79:72] = img4[4279:4272];
      img_out4[87:80] = img4[4287:4280];
      img_out4[95:88] = img4[4295:4288];
      img_out4[103:96] = img4[4303:4296];
      img_out4[111:104] = img4[4311:4304];
      img_out4[119:112] = img4[4319:4312];
      img_out4[127:120] = img4[4327:4320];
      img_out4[135:128] = img4[4335:4328];
      img_out4[143:136] = img4[4343:4336];
      img_out4[151:144] = img4[4351:4344];
      img_out4[159:152] = img4[4359:4352];
      img_out4[167:160] = img4[4367:4360];
      img_out4[175:168] = img4[4375:4368];
    end
    'd34: begin
      img_out0[7:0] = img0[4335:4328];
      img_out0[15:8] = img0[4343:4336];
      img_out0[23:16] = img0[4351:4344];
      img_out0[31:24] = img0[4359:4352];
      img_out0[39:32] = img0[4367:4360];
      img_out0[47:40] = img0[4375:4368];
      img_out0[55:48] = img0[4383:4376];
      img_out0[63:56] = img0[4391:4384];
      img_out0[71:64] = img0[4399:4392];
      img_out0[79:72] = img0[4407:4400];
      img_out0[87:80] = img0[4415:4408];
      img_out0[95:88] = img0[4423:4416];
      img_out0[103:96] = img0[4431:4424];
      img_out0[111:104] = img0[4439:4432];
      img_out0[119:112] = img0[4447:4440];
      img_out0[127:120] = img0[4455:4448];
      img_out0[135:128] = img0[4463:4456];
      img_out0[143:136] = img0[4471:4464];
      img_out0[151:144] = img0[4479:4472];
      img_out0[159:152] = img0[4487:4480];
      img_out0[167:160] = img0[4495:4488];
      img_out0[175:168] = img0[4503:4496];
      img_out1[7:0] = img1[4335:4328];
      img_out1[15:8] = img1[4343:4336];
      img_out1[23:16] = img1[4351:4344];
      img_out1[31:24] = img1[4359:4352];
      img_out1[39:32] = img1[4367:4360];
      img_out1[47:40] = img1[4375:4368];
      img_out1[55:48] = img1[4383:4376];
      img_out1[63:56] = img1[4391:4384];
      img_out1[71:64] = img1[4399:4392];
      img_out1[79:72] = img1[4407:4400];
      img_out1[87:80] = img1[4415:4408];
      img_out1[95:88] = img1[4423:4416];
      img_out1[103:96] = img1[4431:4424];
      img_out1[111:104] = img1[4439:4432];
      img_out1[119:112] = img1[4447:4440];
      img_out1[127:120] = img1[4455:4448];
      img_out1[135:128] = img1[4463:4456];
      img_out1[143:136] = img1[4471:4464];
      img_out1[151:144] = img1[4479:4472];
      img_out1[159:152] = img1[4487:4480];
      img_out1[167:160] = img1[4495:4488];
      img_out1[175:168] = img1[4503:4496];
      img_out2[7:0] = img2[4335:4328];
      img_out2[15:8] = img2[4343:4336];
      img_out2[23:16] = img2[4351:4344];
      img_out2[31:24] = img2[4359:4352];
      img_out2[39:32] = img2[4367:4360];
      img_out2[47:40] = img2[4375:4368];
      img_out2[55:48] = img2[4383:4376];
      img_out2[63:56] = img2[4391:4384];
      img_out2[71:64] = img2[4399:4392];
      img_out2[79:72] = img2[4407:4400];
      img_out2[87:80] = img2[4415:4408];
      img_out2[95:88] = img2[4423:4416];
      img_out2[103:96] = img2[4431:4424];
      img_out2[111:104] = img2[4439:4432];
      img_out2[119:112] = img2[4447:4440];
      img_out2[127:120] = img2[4455:4448];
      img_out2[135:128] = img2[4463:4456];
      img_out2[143:136] = img2[4471:4464];
      img_out2[151:144] = img2[4479:4472];
      img_out2[159:152] = img2[4487:4480];
      img_out2[167:160] = img2[4495:4488];
      img_out2[175:168] = img2[4503:4496];
      img_out3[7:0] = img3[4335:4328];
      img_out3[15:8] = img3[4343:4336];
      img_out3[23:16] = img3[4351:4344];
      img_out3[31:24] = img3[4359:4352];
      img_out3[39:32] = img3[4367:4360];
      img_out3[47:40] = img3[4375:4368];
      img_out3[55:48] = img3[4383:4376];
      img_out3[63:56] = img3[4391:4384];
      img_out3[71:64] = img3[4399:4392];
      img_out3[79:72] = img3[4407:4400];
      img_out3[87:80] = img3[4415:4408];
      img_out3[95:88] = img3[4423:4416];
      img_out3[103:96] = img3[4431:4424];
      img_out3[111:104] = img3[4439:4432];
      img_out3[119:112] = img3[4447:4440];
      img_out3[127:120] = img3[4455:4448];
      img_out3[135:128] = img3[4463:4456];
      img_out3[143:136] = img3[4471:4464];
      img_out3[151:144] = img3[4479:4472];
      img_out3[159:152] = img3[4487:4480];
      img_out3[167:160] = img3[4495:4488];
      img_out3[175:168] = img3[4503:4496];
      img_out4[7:0] = img4[4335:4328];
      img_out4[15:8] = img4[4343:4336];
      img_out4[23:16] = img4[4351:4344];
      img_out4[31:24] = img4[4359:4352];
      img_out4[39:32] = img4[4367:4360];
      img_out4[47:40] = img4[4375:4368];
      img_out4[55:48] = img4[4383:4376];
      img_out4[63:56] = img4[4391:4384];
      img_out4[71:64] = img4[4399:4392];
      img_out4[79:72] = img4[4407:4400];
      img_out4[87:80] = img4[4415:4408];
      img_out4[95:88] = img4[4423:4416];
      img_out4[103:96] = img4[4431:4424];
      img_out4[111:104] = img4[4439:4432];
      img_out4[119:112] = img4[4447:4440];
      img_out4[127:120] = img4[4455:4448];
      img_out4[135:128] = img4[4463:4456];
      img_out4[143:136] = img4[4471:4464];
      img_out4[151:144] = img4[4479:4472];
      img_out4[159:152] = img4[4487:4480];
      img_out4[167:160] = img4[4495:4488];
      img_out4[175:168] = img4[4503:4496];
    end
    'd35: begin
      img_out0[7:0] = img0[4463:4456];
      img_out0[15:8] = img0[4471:4464];
      img_out0[23:16] = img0[4479:4472];
      img_out0[31:24] = img0[4487:4480];
      img_out0[39:32] = img0[4495:4488];
      img_out0[47:40] = img0[4503:4496];
      img_out0[55:48] = img0[4511:4504];
      img_out0[63:56] = img0[4519:4512];
      img_out0[71:64] = img0[4527:4520];
      img_out0[79:72] = img0[4535:4528];
      img_out0[87:80] = img0[4543:4536];
      img_out0[95:88] = img0[4551:4544];
      img_out0[103:96] = img0[4559:4552];
      img_out0[111:104] = img0[4567:4560];
      img_out0[119:112] = img0[4575:4568];
      img_out0[127:120] = img0[4583:4576];
      img_out0[135:128] = img0[4591:4584];
      img_out0[143:136] = img0[4599:4592];
      img_out0[151:144] = img0[4607:4600];
      img_out0[159:152] = img0[4615:4608];
      img_out0[167:160] = img0[4623:4616];
      img_out0[175:168] = img0[4631:4624];
      img_out1[7:0] = img1[4463:4456];
      img_out1[15:8] = img1[4471:4464];
      img_out1[23:16] = img1[4479:4472];
      img_out1[31:24] = img1[4487:4480];
      img_out1[39:32] = img1[4495:4488];
      img_out1[47:40] = img1[4503:4496];
      img_out1[55:48] = img1[4511:4504];
      img_out1[63:56] = img1[4519:4512];
      img_out1[71:64] = img1[4527:4520];
      img_out1[79:72] = img1[4535:4528];
      img_out1[87:80] = img1[4543:4536];
      img_out1[95:88] = img1[4551:4544];
      img_out1[103:96] = img1[4559:4552];
      img_out1[111:104] = img1[4567:4560];
      img_out1[119:112] = img1[4575:4568];
      img_out1[127:120] = img1[4583:4576];
      img_out1[135:128] = img1[4591:4584];
      img_out1[143:136] = img1[4599:4592];
      img_out1[151:144] = img1[4607:4600];
      img_out1[159:152] = img1[4615:4608];
      img_out1[167:160] = img1[4623:4616];
      img_out1[175:168] = img1[4631:4624];
      img_out2[7:0] = img2[4463:4456];
      img_out2[15:8] = img2[4471:4464];
      img_out2[23:16] = img2[4479:4472];
      img_out2[31:24] = img2[4487:4480];
      img_out2[39:32] = img2[4495:4488];
      img_out2[47:40] = img2[4503:4496];
      img_out2[55:48] = img2[4511:4504];
      img_out2[63:56] = img2[4519:4512];
      img_out2[71:64] = img2[4527:4520];
      img_out2[79:72] = img2[4535:4528];
      img_out2[87:80] = img2[4543:4536];
      img_out2[95:88] = img2[4551:4544];
      img_out2[103:96] = img2[4559:4552];
      img_out2[111:104] = img2[4567:4560];
      img_out2[119:112] = img2[4575:4568];
      img_out2[127:120] = img2[4583:4576];
      img_out2[135:128] = img2[4591:4584];
      img_out2[143:136] = img2[4599:4592];
      img_out2[151:144] = img2[4607:4600];
      img_out2[159:152] = img2[4615:4608];
      img_out2[167:160] = img2[4623:4616];
      img_out2[175:168] = img2[4631:4624];
      img_out3[7:0] = img3[4463:4456];
      img_out3[15:8] = img3[4471:4464];
      img_out3[23:16] = img3[4479:4472];
      img_out3[31:24] = img3[4487:4480];
      img_out3[39:32] = img3[4495:4488];
      img_out3[47:40] = img3[4503:4496];
      img_out3[55:48] = img3[4511:4504];
      img_out3[63:56] = img3[4519:4512];
      img_out3[71:64] = img3[4527:4520];
      img_out3[79:72] = img3[4535:4528];
      img_out3[87:80] = img3[4543:4536];
      img_out3[95:88] = img3[4551:4544];
      img_out3[103:96] = img3[4559:4552];
      img_out3[111:104] = img3[4567:4560];
      img_out3[119:112] = img3[4575:4568];
      img_out3[127:120] = img3[4583:4576];
      img_out3[135:128] = img3[4591:4584];
      img_out3[143:136] = img3[4599:4592];
      img_out3[151:144] = img3[4607:4600];
      img_out3[159:152] = img3[4615:4608];
      img_out3[167:160] = img3[4623:4616];
      img_out3[175:168] = img3[4631:4624];
      img_out4[7:0] = img4[4463:4456];
      img_out4[15:8] = img4[4471:4464];
      img_out4[23:16] = img4[4479:4472];
      img_out4[31:24] = img4[4487:4480];
      img_out4[39:32] = img4[4495:4488];
      img_out4[47:40] = img4[4503:4496];
      img_out4[55:48] = img4[4511:4504];
      img_out4[63:56] = img4[4519:4512];
      img_out4[71:64] = img4[4527:4520];
      img_out4[79:72] = img4[4535:4528];
      img_out4[87:80] = img4[4543:4536];
      img_out4[95:88] = img4[4551:4544];
      img_out4[103:96] = img4[4559:4552];
      img_out4[111:104] = img4[4567:4560];
      img_out4[119:112] = img4[4575:4568];
      img_out4[127:120] = img4[4583:4576];
      img_out4[135:128] = img4[4591:4584];
      img_out4[143:136] = img4[4599:4592];
      img_out4[151:144] = img4[4607:4600];
      img_out4[159:152] = img4[4615:4608];
      img_out4[167:160] = img4[4623:4616];
      img_out4[175:168] = img4[4631:4624];
    end
    'd36: begin
      img_out0[7:0] = img0[4591:4584];
      img_out0[15:8] = img0[4599:4592];
      img_out0[23:16] = img0[4607:4600];
      img_out0[31:24] = img0[4615:4608];
      img_out0[39:32] = img0[4623:4616];
      img_out0[47:40] = img0[4631:4624];
      img_out0[55:48] = img0[4639:4632];
      img_out0[63:56] = img0[4647:4640];
      img_out0[71:64] = img0[4655:4648];
      img_out0[79:72] = img0[4663:4656];
      img_out0[87:80] = img0[4671:4664];
      img_out0[95:88] = img0[4679:4672];
      img_out0[103:96] = img0[4687:4680];
      img_out0[111:104] = img0[4695:4688];
      img_out0[119:112] = img0[4703:4696];
      img_out0[127:120] = img0[4711:4704];
      img_out0[135:128] = img0[4719:4712];
      img_out0[143:136] = img0[4727:4720];
      img_out0[151:144] = img0[4735:4728];
      img_out0[159:152] = img0[4743:4736];
      img_out0[167:160] = img0[4751:4744];
      img_out0[175:168] = img0[4759:4752];
      img_out1[7:0] = img1[4591:4584];
      img_out1[15:8] = img1[4599:4592];
      img_out1[23:16] = img1[4607:4600];
      img_out1[31:24] = img1[4615:4608];
      img_out1[39:32] = img1[4623:4616];
      img_out1[47:40] = img1[4631:4624];
      img_out1[55:48] = img1[4639:4632];
      img_out1[63:56] = img1[4647:4640];
      img_out1[71:64] = img1[4655:4648];
      img_out1[79:72] = img1[4663:4656];
      img_out1[87:80] = img1[4671:4664];
      img_out1[95:88] = img1[4679:4672];
      img_out1[103:96] = img1[4687:4680];
      img_out1[111:104] = img1[4695:4688];
      img_out1[119:112] = img1[4703:4696];
      img_out1[127:120] = img1[4711:4704];
      img_out1[135:128] = img1[4719:4712];
      img_out1[143:136] = img1[4727:4720];
      img_out1[151:144] = img1[4735:4728];
      img_out1[159:152] = img1[4743:4736];
      img_out1[167:160] = img1[4751:4744];
      img_out1[175:168] = img1[4759:4752];
      img_out2[7:0] = img2[4591:4584];
      img_out2[15:8] = img2[4599:4592];
      img_out2[23:16] = img2[4607:4600];
      img_out2[31:24] = img2[4615:4608];
      img_out2[39:32] = img2[4623:4616];
      img_out2[47:40] = img2[4631:4624];
      img_out2[55:48] = img2[4639:4632];
      img_out2[63:56] = img2[4647:4640];
      img_out2[71:64] = img2[4655:4648];
      img_out2[79:72] = img2[4663:4656];
      img_out2[87:80] = img2[4671:4664];
      img_out2[95:88] = img2[4679:4672];
      img_out2[103:96] = img2[4687:4680];
      img_out2[111:104] = img2[4695:4688];
      img_out2[119:112] = img2[4703:4696];
      img_out2[127:120] = img2[4711:4704];
      img_out2[135:128] = img2[4719:4712];
      img_out2[143:136] = img2[4727:4720];
      img_out2[151:144] = img2[4735:4728];
      img_out2[159:152] = img2[4743:4736];
      img_out2[167:160] = img2[4751:4744];
      img_out2[175:168] = img2[4759:4752];
      img_out3[7:0] = img3[4591:4584];
      img_out3[15:8] = img3[4599:4592];
      img_out3[23:16] = img3[4607:4600];
      img_out3[31:24] = img3[4615:4608];
      img_out3[39:32] = img3[4623:4616];
      img_out3[47:40] = img3[4631:4624];
      img_out3[55:48] = img3[4639:4632];
      img_out3[63:56] = img3[4647:4640];
      img_out3[71:64] = img3[4655:4648];
      img_out3[79:72] = img3[4663:4656];
      img_out3[87:80] = img3[4671:4664];
      img_out3[95:88] = img3[4679:4672];
      img_out3[103:96] = img3[4687:4680];
      img_out3[111:104] = img3[4695:4688];
      img_out3[119:112] = img3[4703:4696];
      img_out3[127:120] = img3[4711:4704];
      img_out3[135:128] = img3[4719:4712];
      img_out3[143:136] = img3[4727:4720];
      img_out3[151:144] = img3[4735:4728];
      img_out3[159:152] = img3[4743:4736];
      img_out3[167:160] = img3[4751:4744];
      img_out3[175:168] = img3[4759:4752];
      img_out4[7:0] = img4[4591:4584];
      img_out4[15:8] = img4[4599:4592];
      img_out4[23:16] = img4[4607:4600];
      img_out4[31:24] = img4[4615:4608];
      img_out4[39:32] = img4[4623:4616];
      img_out4[47:40] = img4[4631:4624];
      img_out4[55:48] = img4[4639:4632];
      img_out4[63:56] = img4[4647:4640];
      img_out4[71:64] = img4[4655:4648];
      img_out4[79:72] = img4[4663:4656];
      img_out4[87:80] = img4[4671:4664];
      img_out4[95:88] = img4[4679:4672];
      img_out4[103:96] = img4[4687:4680];
      img_out4[111:104] = img4[4695:4688];
      img_out4[119:112] = img4[4703:4696];
      img_out4[127:120] = img4[4711:4704];
      img_out4[135:128] = img4[4719:4712];
      img_out4[143:136] = img4[4727:4720];
      img_out4[151:144] = img4[4735:4728];
      img_out4[159:152] = img4[4743:4736];
      img_out4[167:160] = img4[4751:4744];
      img_out4[175:168] = img4[4759:4752];
    end
    'd37: begin
      img_out0[7:0] = img0[4719:4712];
      img_out0[15:8] = img0[4727:4720];
      img_out0[23:16] = img0[4735:4728];
      img_out0[31:24] = img0[4743:4736];
      img_out0[39:32] = img0[4751:4744];
      img_out0[47:40] = img0[4759:4752];
      img_out0[55:48] = img0[4767:4760];
      img_out0[63:56] = img0[4775:4768];
      img_out0[71:64] = img0[4783:4776];
      img_out0[79:72] = img0[4791:4784];
      img_out0[87:80] = img0[4799:4792];
      img_out0[95:88] = img0[4807:4800];
      img_out0[103:96] = img0[4815:4808];
      img_out0[111:104] = img0[4823:4816];
      img_out0[119:112] = img0[4831:4824];
      img_out0[127:120] = img0[4839:4832];
      img_out0[135:128] = img0[4847:4840];
      img_out0[143:136] = img0[4855:4848];
      img_out0[151:144] = img0[4863:4856];
      img_out0[159:152] = img0[4871:4864];
      img_out0[167:160] = img0[4879:4872];
      img_out0[175:168] = img0[4887:4880];
      img_out1[7:0] = img1[4719:4712];
      img_out1[15:8] = img1[4727:4720];
      img_out1[23:16] = img1[4735:4728];
      img_out1[31:24] = img1[4743:4736];
      img_out1[39:32] = img1[4751:4744];
      img_out1[47:40] = img1[4759:4752];
      img_out1[55:48] = img1[4767:4760];
      img_out1[63:56] = img1[4775:4768];
      img_out1[71:64] = img1[4783:4776];
      img_out1[79:72] = img1[4791:4784];
      img_out1[87:80] = img1[4799:4792];
      img_out1[95:88] = img1[4807:4800];
      img_out1[103:96] = img1[4815:4808];
      img_out1[111:104] = img1[4823:4816];
      img_out1[119:112] = img1[4831:4824];
      img_out1[127:120] = img1[4839:4832];
      img_out1[135:128] = img1[4847:4840];
      img_out1[143:136] = img1[4855:4848];
      img_out1[151:144] = img1[4863:4856];
      img_out1[159:152] = img1[4871:4864];
      img_out1[167:160] = img1[4879:4872];
      img_out1[175:168] = img1[4887:4880];
      img_out2[7:0] = img2[4719:4712];
      img_out2[15:8] = img2[4727:4720];
      img_out2[23:16] = img2[4735:4728];
      img_out2[31:24] = img2[4743:4736];
      img_out2[39:32] = img2[4751:4744];
      img_out2[47:40] = img2[4759:4752];
      img_out2[55:48] = img2[4767:4760];
      img_out2[63:56] = img2[4775:4768];
      img_out2[71:64] = img2[4783:4776];
      img_out2[79:72] = img2[4791:4784];
      img_out2[87:80] = img2[4799:4792];
      img_out2[95:88] = img2[4807:4800];
      img_out2[103:96] = img2[4815:4808];
      img_out2[111:104] = img2[4823:4816];
      img_out2[119:112] = img2[4831:4824];
      img_out2[127:120] = img2[4839:4832];
      img_out2[135:128] = img2[4847:4840];
      img_out2[143:136] = img2[4855:4848];
      img_out2[151:144] = img2[4863:4856];
      img_out2[159:152] = img2[4871:4864];
      img_out2[167:160] = img2[4879:4872];
      img_out2[175:168] = img2[4887:4880];
      img_out3[7:0] = img3[4719:4712];
      img_out3[15:8] = img3[4727:4720];
      img_out3[23:16] = img3[4735:4728];
      img_out3[31:24] = img3[4743:4736];
      img_out3[39:32] = img3[4751:4744];
      img_out3[47:40] = img3[4759:4752];
      img_out3[55:48] = img3[4767:4760];
      img_out3[63:56] = img3[4775:4768];
      img_out3[71:64] = img3[4783:4776];
      img_out3[79:72] = img3[4791:4784];
      img_out3[87:80] = img3[4799:4792];
      img_out3[95:88] = img3[4807:4800];
      img_out3[103:96] = img3[4815:4808];
      img_out3[111:104] = img3[4823:4816];
      img_out3[119:112] = img3[4831:4824];
      img_out3[127:120] = img3[4839:4832];
      img_out3[135:128] = img3[4847:4840];
      img_out3[143:136] = img3[4855:4848];
      img_out3[151:144] = img3[4863:4856];
      img_out3[159:152] = img3[4871:4864];
      img_out3[167:160] = img3[4879:4872];
      img_out3[175:168] = img3[4887:4880];
      img_out4[7:0] = img4[4719:4712];
      img_out4[15:8] = img4[4727:4720];
      img_out4[23:16] = img4[4735:4728];
      img_out4[31:24] = img4[4743:4736];
      img_out4[39:32] = img4[4751:4744];
      img_out4[47:40] = img4[4759:4752];
      img_out4[55:48] = img4[4767:4760];
      img_out4[63:56] = img4[4775:4768];
      img_out4[71:64] = img4[4783:4776];
      img_out4[79:72] = img4[4791:4784];
      img_out4[87:80] = img4[4799:4792];
      img_out4[95:88] = img4[4807:4800];
      img_out4[103:96] = img4[4815:4808];
      img_out4[111:104] = img4[4823:4816];
      img_out4[119:112] = img4[4831:4824];
      img_out4[127:120] = img4[4839:4832];
      img_out4[135:128] = img4[4847:4840];
      img_out4[143:136] = img4[4855:4848];
      img_out4[151:144] = img4[4863:4856];
      img_out4[159:152] = img4[4871:4864];
      img_out4[167:160] = img4[4879:4872];
      img_out4[175:168] = img4[4887:4880];
    end
    'd38: begin
      img_out0[7:0] = img0[4847:4840];
      img_out0[15:8] = img0[4855:4848];
      img_out0[23:16] = img0[4863:4856];
      img_out0[31:24] = img0[4871:4864];
      img_out0[39:32] = img0[4879:4872];
      img_out0[47:40] = img0[4887:4880];
      img_out0[55:48] = img0[4895:4888];
      img_out0[63:56] = img0[4903:4896];
      img_out0[71:64] = img0[4911:4904];
      img_out0[79:72] = img0[4919:4912];
      img_out0[87:80] = img0[4927:4920];
      img_out0[95:88] = img0[4935:4928];
      img_out0[103:96] = img0[4943:4936];
      img_out0[111:104] = img0[4951:4944];
      img_out0[119:112] = img0[4959:4952];
      img_out0[127:120] = img0[4967:4960];
      img_out0[135:128] = img0[4975:4968];
      img_out0[143:136] = img0[4983:4976];
      img_out0[151:144] = img0[4991:4984];
      img_out0[159:152] = img0[4999:4992];
      img_out0[167:160] = img0[5007:5000];
      img_out0[175:168] = img0[5015:5008];
      img_out1[7:0] = img1[4847:4840];
      img_out1[15:8] = img1[4855:4848];
      img_out1[23:16] = img1[4863:4856];
      img_out1[31:24] = img1[4871:4864];
      img_out1[39:32] = img1[4879:4872];
      img_out1[47:40] = img1[4887:4880];
      img_out1[55:48] = img1[4895:4888];
      img_out1[63:56] = img1[4903:4896];
      img_out1[71:64] = img1[4911:4904];
      img_out1[79:72] = img1[4919:4912];
      img_out1[87:80] = img1[4927:4920];
      img_out1[95:88] = img1[4935:4928];
      img_out1[103:96] = img1[4943:4936];
      img_out1[111:104] = img1[4951:4944];
      img_out1[119:112] = img1[4959:4952];
      img_out1[127:120] = img1[4967:4960];
      img_out1[135:128] = img1[4975:4968];
      img_out1[143:136] = img1[4983:4976];
      img_out1[151:144] = img1[4991:4984];
      img_out1[159:152] = img1[4999:4992];
      img_out1[167:160] = img1[5007:5000];
      img_out1[175:168] = img1[5015:5008];
      img_out2[7:0] = img2[4847:4840];
      img_out2[15:8] = img2[4855:4848];
      img_out2[23:16] = img2[4863:4856];
      img_out2[31:24] = img2[4871:4864];
      img_out2[39:32] = img2[4879:4872];
      img_out2[47:40] = img2[4887:4880];
      img_out2[55:48] = img2[4895:4888];
      img_out2[63:56] = img2[4903:4896];
      img_out2[71:64] = img2[4911:4904];
      img_out2[79:72] = img2[4919:4912];
      img_out2[87:80] = img2[4927:4920];
      img_out2[95:88] = img2[4935:4928];
      img_out2[103:96] = img2[4943:4936];
      img_out2[111:104] = img2[4951:4944];
      img_out2[119:112] = img2[4959:4952];
      img_out2[127:120] = img2[4967:4960];
      img_out2[135:128] = img2[4975:4968];
      img_out2[143:136] = img2[4983:4976];
      img_out2[151:144] = img2[4991:4984];
      img_out2[159:152] = img2[4999:4992];
      img_out2[167:160] = img2[5007:5000];
      img_out2[175:168] = img2[5015:5008];
      img_out3[7:0] = img3[4847:4840];
      img_out3[15:8] = img3[4855:4848];
      img_out3[23:16] = img3[4863:4856];
      img_out3[31:24] = img3[4871:4864];
      img_out3[39:32] = img3[4879:4872];
      img_out3[47:40] = img3[4887:4880];
      img_out3[55:48] = img3[4895:4888];
      img_out3[63:56] = img3[4903:4896];
      img_out3[71:64] = img3[4911:4904];
      img_out3[79:72] = img3[4919:4912];
      img_out3[87:80] = img3[4927:4920];
      img_out3[95:88] = img3[4935:4928];
      img_out3[103:96] = img3[4943:4936];
      img_out3[111:104] = img3[4951:4944];
      img_out3[119:112] = img3[4959:4952];
      img_out3[127:120] = img3[4967:4960];
      img_out3[135:128] = img3[4975:4968];
      img_out3[143:136] = img3[4983:4976];
      img_out3[151:144] = img3[4991:4984];
      img_out3[159:152] = img3[4999:4992];
      img_out3[167:160] = img3[5007:5000];
      img_out3[175:168] = img3[5015:5008];
      img_out4[7:0] = img4[4847:4840];
      img_out4[15:8] = img4[4855:4848];
      img_out4[23:16] = img4[4863:4856];
      img_out4[31:24] = img4[4871:4864];
      img_out4[39:32] = img4[4879:4872];
      img_out4[47:40] = img4[4887:4880];
      img_out4[55:48] = img4[4895:4888];
      img_out4[63:56] = img4[4903:4896];
      img_out4[71:64] = img4[4911:4904];
      img_out4[79:72] = img4[4919:4912];
      img_out4[87:80] = img4[4927:4920];
      img_out4[95:88] = img4[4935:4928];
      img_out4[103:96] = img4[4943:4936];
      img_out4[111:104] = img4[4951:4944];
      img_out4[119:112] = img4[4959:4952];
      img_out4[127:120] = img4[4967:4960];
      img_out4[135:128] = img4[4975:4968];
      img_out4[143:136] = img4[4983:4976];
      img_out4[151:144] = img4[4991:4984];
      img_out4[159:152] = img4[4999:4992];
      img_out4[167:160] = img4[5007:5000];
      img_out4[175:168] = img4[5015:5008];
    end
    'd39: begin
      img_out0[7:0] = img0[4975:4968];
      img_out0[15:8] = img0[4983:4976];
      img_out0[23:16] = img0[4991:4984];
      img_out0[31:24] = img0[4999:4992];
      img_out0[39:32] = img0[5007:5000];
      img_out0[47:40] = img0[5015:5008];
      img_out0[55:48] = img0[5023:5016];
      img_out0[63:56] = img0[5031:5024];
      img_out0[71:64] = img0[5039:5032];
      img_out0[79:72] = img0[5047:5040];
      img_out0[87:80] = img0[5055:5048];
      img_out0[95:88] = img0[5063:5056];
      img_out0[103:96] = img0[5071:5064];
      img_out0[111:104] = img0[5079:5072];
      img_out0[119:112] = img0[5087:5080];
      img_out0[127:120] = img0[5095:5088];
      img_out0[135:128] = img0[5103:5096];
      img_out0[143:136] = img0[5111:5104];
      img_out0[151:144] = img0[5119:5112];
      img_out0[159:152] = 'd0;
      img_out0[167:160] = 'd0;
      img_out0[175:168] = 'd0;
      img_out1[7:0] = img1[4975:4968];
      img_out1[15:8] = img1[4983:4976];
      img_out1[23:16] = img1[4991:4984];
      img_out1[31:24] = img1[4999:4992];
      img_out1[39:32] = img1[5007:5000];
      img_out1[47:40] = img1[5015:5008];
      img_out1[55:48] = img1[5023:5016];
      img_out1[63:56] = img1[5031:5024];
      img_out1[71:64] = img1[5039:5032];
      img_out1[79:72] = img1[5047:5040];
      img_out1[87:80] = img1[5055:5048];
      img_out1[95:88] = img1[5063:5056];
      img_out1[103:96] = img1[5071:5064];
      img_out1[111:104] = img1[5079:5072];
      img_out1[119:112] = img1[5087:5080];
      img_out1[127:120] = img1[5095:5088];
      img_out1[135:128] = img1[5103:5096];
      img_out1[143:136] = img1[5111:5104];
      img_out1[151:144] = img1[5119:5112];
      img_out1[159:152] = 'd0;
      img_out1[167:160] = 'd0;
      img_out1[175:168] = 'd0;
      img_out2[7:0] = img2[4975:4968];
      img_out2[15:8] = img2[4983:4976];
      img_out2[23:16] = img2[4991:4984];
      img_out2[31:24] = img2[4999:4992];
      img_out2[39:32] = img2[5007:5000];
      img_out2[47:40] = img2[5015:5008];
      img_out2[55:48] = img2[5023:5016];
      img_out2[63:56] = img2[5031:5024];
      img_out2[71:64] = img2[5039:5032];
      img_out2[79:72] = img2[5047:5040];
      img_out2[87:80] = img2[5055:5048];
      img_out2[95:88] = img2[5063:5056];
      img_out2[103:96] = img2[5071:5064];
      img_out2[111:104] = img2[5079:5072];
      img_out2[119:112] = img2[5087:5080];
      img_out2[127:120] = img2[5095:5088];
      img_out2[135:128] = img2[5103:5096];
      img_out2[143:136] = img2[5111:5104];
      img_out2[151:144] = img2[5119:5112];
      img_out2[159:152] = 'd0;
      img_out2[167:160] = 'd0;
      img_out2[175:168] = 'd0;
      img_out3[7:0] = img3[4975:4968];
      img_out3[15:8] = img3[4983:4976];
      img_out3[23:16] = img3[4991:4984];
      img_out3[31:24] = img3[4999:4992];
      img_out3[39:32] = img3[5007:5000];
      img_out3[47:40] = img3[5015:5008];
      img_out3[55:48] = img3[5023:5016];
      img_out3[63:56] = img3[5031:5024];
      img_out3[71:64] = img3[5039:5032];
      img_out3[79:72] = img3[5047:5040];
      img_out3[87:80] = img3[5055:5048];
      img_out3[95:88] = img3[5063:5056];
      img_out3[103:96] = img3[5071:5064];
      img_out3[111:104] = img3[5079:5072];
      img_out3[119:112] = img3[5087:5080];
      img_out3[127:120] = img3[5095:5088];
      img_out3[135:128] = img3[5103:5096];
      img_out3[143:136] = img3[5111:5104];
      img_out3[151:144] = img3[5119:5112];
      img_out3[159:152] = 'd0;
      img_out3[167:160] = 'd0;
      img_out3[175:168] = 'd0;
      img_out4[7:0] = img4[4975:4968];
      img_out4[15:8] = img4[4983:4976];
      img_out4[23:16] = img4[4991:4984];
      img_out4[31:24] = img4[4999:4992];
      img_out4[39:32] = img4[5007:5000];
      img_out4[47:40] = img4[5015:5008];
      img_out4[55:48] = img4[5023:5016];
      img_out4[63:56] = img4[5031:5024];
      img_out4[71:64] = img4[5039:5032];
      img_out4[79:72] = img4[5047:5040];
      img_out4[87:80] = img4[5055:5048];
      img_out4[95:88] = img4[5063:5056];
      img_out4[103:96] = img4[5071:5064];
      img_out4[111:104] = img4[5079:5072];
      img_out4[119:112] = img4[5087:5080];
      img_out4[127:120] = img4[5095:5088];
      img_out4[135:128] = img4[5103:5096];
      img_out4[143:136] = img4[5111:5104];
      img_out4[151:144] = img4[5119:5112];
      img_out4[159:152] = 'd0;
      img_out4[167:160] = 'd0;
      img_out4[175:168] = 'd0;
    end
    default: begin
      img_out0[7:0] = 'd0;
      img_out0[15:8] = 'd0;
      img_out0[23:16] = 'd0;
      img_out0[31:24] = 'd0;
      img_out0[39:32] = 'd0;
      img_out0[47:40] = 'd0;
      img_out0[55:48] = 'd0;
      img_out0[63:56] = 'd0;
      img_out0[71:64] = 'd0;
      img_out0[79:72] = 'd0;
      img_out0[87:80] = 'd0;
      img_out0[95:88] = 'd0;
      img_out0[103:96] = 'd0;
      img_out0[111:104] = 'd0;
      img_out0[119:112] = 'd0;
      img_out0[127:120] = 'd0;
      img_out0[135:128] = 'd0;
      img_out0[143:136] = 'd0;
      img_out0[151:144] = 'd0;
      img_out0[159:152] = 'd0;
      img_out0[167:160] = 'd0;
      img_out0[175:168] = 'd0;
      img_out1[7:0] = 'd0;
      img_out1[15:8] = 'd0;
      img_out1[23:16] = 'd0;
      img_out1[31:24] = 'd0;
      img_out1[39:32] = 'd0;
      img_out1[47:40] = 'd0;
      img_out1[55:48] = 'd0;
      img_out1[63:56] = 'd0;
      img_out1[71:64] = 'd0;
      img_out1[79:72] = 'd0;
      img_out1[87:80] = 'd0;
      img_out1[95:88] = 'd0;
      img_out1[103:96] = 'd0;
      img_out1[111:104] = 'd0;
      img_out1[119:112] = 'd0;
      img_out1[127:120] = 'd0;
      img_out1[135:128] = 'd0;
      img_out1[143:136] = 'd0;
      img_out1[151:144] = 'd0;
      img_out1[159:152] = 'd0;
      img_out1[167:160] = 'd0;
      img_out1[175:168] = 'd0;
      img_out2[7:0] = 'd0;
      img_out2[15:8] = 'd0;
      img_out2[23:16] = 'd0;
      img_out2[31:24] = 'd0;
      img_out2[39:32] = 'd0;
      img_out2[47:40] = 'd0;
      img_out2[55:48] = 'd0;
      img_out2[63:56] = 'd0;
      img_out2[71:64] = 'd0;
      img_out2[79:72] = 'd0;
      img_out2[87:80] = 'd0;
      img_out2[95:88] = 'd0;
      img_out2[103:96] = 'd0;
      img_out2[111:104] = 'd0;
      img_out2[119:112] = 'd0;
      img_out2[127:120] = 'd0;
      img_out2[135:128] = 'd0;
      img_out2[143:136] = 'd0;
      img_out2[151:144] = 'd0;
      img_out2[159:152] = 'd0;
      img_out2[167:160] = 'd0;
      img_out2[175:168] = 'd0;
      img_out3[7:0] = 'd0;
      img_out3[15:8] = 'd0;
      img_out3[23:16] = 'd0;
      img_out3[31:24] = 'd0;
      img_out3[39:32] = 'd0;
      img_out3[47:40] = 'd0;
      img_out3[55:48] = 'd0;
      img_out3[63:56] = 'd0;
      img_out3[71:64] = 'd0;
      img_out3[79:72] = 'd0;
      img_out3[87:80] = 'd0;
      img_out3[95:88] = 'd0;
      img_out3[103:96] = 'd0;
      img_out3[111:104] = 'd0;
      img_out3[119:112] = 'd0;
      img_out3[127:120] = 'd0;
      img_out3[135:128] = 'd0;
      img_out3[143:136] = 'd0;
      img_out3[151:144] = 'd0;
      img_out3[159:152] = 'd0;
      img_out3[167:160] = 'd0;
      img_out3[175:168] = 'd0;
      img_out4[7:0] = 'd0;
      img_out4[15:8] = 'd0;
      img_out4[23:16] = 'd0;
      img_out4[31:24] = 'd0;
      img_out4[39:32] = 'd0;
      img_out4[47:40] = 'd0;
      img_out4[55:48] = 'd0;
      img_out4[63:56] = 'd0;
      img_out4[71:64] = 'd0;
      img_out4[79:72] = 'd0;
      img_out4[87:80] = 'd0;
      img_out4[95:88] = 'd0;
      img_out4[103:96] = 'd0;
      img_out4[111:104] = 'd0;
      img_out4[119:112] = 'd0;
      img_out4[127:120] = 'd0;
      img_out4[135:128] = 'd0;
      img_out4[143:136] = 'd0;
      img_out4[151:144] = 'd0;
      img_out4[159:152] = 'd0;
      img_out4[167:160] = 'd0;
      img_out4[175:168] = 'd0;
    end
  endcase
end

endmodule
