module Gaussian_Blur_7x7(
  clk,
  rst_n,
  buffer_data_0,
  buffer_data_1,
  buffer_data_2,
  buffer_data_3,
  buffer_data_4,
  buffer_data_5,
  buffer_data_6,
  current_state,
  blur_din
);

input                 clk;
input                 rst_n;
input         [3:0]   current_state;
input       [5119:0]   buffer_data_0;
input       [5119:0]   buffer_data_1;
input       [5119:0]   buffer_data_2;
input       [5119:0]   buffer_data_3;
input       [5119:0]   buffer_data_4;
input       [5119:0]   buffer_data_5;
input       [5119:0]   buffer_data_6;
output reg  [5119:0]  blur_din;

parameter ST_IDLE        = 0,
          ST_READY       = 1,/*Idle 1 state for SRAM to get READY*/
          ST_GAUSSIAN_0  = 2,
          ST_GAUSSIAN_1  = 3,
          ST_GAUSSIAN_2  = 4,
          ST_GAUSSIAN_3  = 5,
          ST_GAUSSIAN_4  = 6,
          ST_GAUSSIAN_5  = 7,
          ST_GAUSSIAN_6  = 8,
          ST_GAUSSIAN_7  = 9,
          ST_GAUSSIAN_8  = 10,
          ST_GAUSSIAN_9  = 11;

reg       [223:0] G_Kernel_7x7  [0:3];
always @(posedge clk) begin
  if (!rst_n) begin
    G_Kernel_7x7[0][31:0]    <= 32'h03C6EBCB; //18'b000000111100011011;//'d014754;
    G_Kernel_7x7[0][63:32]   <= 32'h046AA8A8; //18'b000001000110101010;//'d017252;
    G_Kernel_7x7[0][95:64]   <= 32'h04D9ED31; //18'b000001001101100111;//'d018950;
    G_Kernel_7x7[0][127:96]   <= 32'h050165DE; //18'b000001010000000101;//'d019552;
    G_Kernel_7x7[0][159:128]   <= 32'h04D9ED31; //18'b000001001101100111;//'d018950;
    G_Kernel_7x7[0][191:160]  <= 32'h046AA8A8; //18'b000001000110101010;//'d017252;
    G_Kernel_7x7[0][223:192] <= 32'h03C6EBCB; //18'b000000111100011011;//'d014754;
    G_Kernel_7x7[1][31:0]    <= 32'h046AA8A8; //18'b000001000110101010;//'d017252;
    G_Kernel_7x7[1][63:32]   <= 32'h052A1FB1; //18'b000001010010101000;//'d020174;
    G_Kernel_7x7[1][95:64]   <= 32'h05AC3BC7; //18'b000001011010110000;//'d022159;
    G_Kernel_7x7[1][127:96]   <= 32'h05DA6392; //18'b000001011101101001;//'d022863;
    G_Kernel_7x7[1][159:128]   <= 32'h05AC3BC7; //18'b000001011010110000;//'d022159;
    G_Kernel_7x7[1][191:160]  <= 32'h052A1FB1; //18'b000001010010101000;//'d020174;
    G_Kernel_7x7[1][223:192] <= 32'h046AA8A8; //18'b000001000110101010;//'d017252;
    G_Kernel_7x7[2][31:0]    <= 32'h04D9ED31; //18'b000001001101100111;//'d018950;
    G_Kernel_7x7[2][63:32]   <= 32'h05AC3BC7; //18'b000001011010110000;//'d022159;
    G_Kernel_7x7[2][95:64]   <= 32'h063B25B2; //18'b000001100011101100;//'d024340;
    G_Kernel_7x7[2][127:96]   <= 32'h066DD847; //18'b000001100110110111;//'d025113;
    G_Kernel_7x7[2][159:128]   <= 32'h063B25B2; //18'b000001100011101100;//'d024340;
    G_Kernel_7x7[2][191:160]  <= 32'h05AC3BC7; //18'b000001011010110000;//'d022159;
    G_Kernel_7x7[2][223:192] <= 32'h04D9ED31; //18'b000001001101100111;//'d018950;
    G_Kernel_7x7[3][31:0]    <= 32'h050165DE; //18'b000001010000000101;//'d019552;
    G_Kernel_7x7[3][63:32]   <= 32'h05DA6392; //18'b000001011101101001;//'d022863;
    G_Kernel_7x7[3][95:64]   <= 32'h066DD847; //18'b000001100110110111;//'d025113;
    G_Kernel_7x7[3][127:96]   <= 32'h06A2275A; //18'b000001101010001000;//'d025911;
    G_Kernel_7x7[3][159:128]   <= 32'h066DD847; //18'b000001100110110111;//'d025113;
    G_Kernel_7x7[3][191:160]  <= 32'h05DA6392; //18'b000001011101101001;//'d022863;
    G_Kernel_7x7[3][223:192] <= 32'h050165DE; //18'b000001010000000101;//'d019552;
  end
end

reg    [55:0]    layer0[0:63]; //wire
reg    [55:0]    layer1[0:63]; //wire
reg    [55:0]    layer2[0:63]; //wire
reg    [55:0]    layer3[0:63]; //wire
reg    [55:0]    layer4[0:63]; //wire
reg    [55:0]    layer5[0:63]; //wire
reg    [55:0]    layer6[0:63]; //wire
always @(*) begin
  case(current_state)
    ST_GAUSSIAN_0: begin
        layer0[0][7:0] = 0;
        layer0[0][15:8] = 0;
        layer0[0][23:16] = 0;
        layer0[0][31:24] = buffer_data_6[7:0];
        layer0[0][39:32] = buffer_data_6[15:8];
        layer0[0][47:40] = buffer_data_6[23:16];
        layer0[0][55:48] = buffer_data_6[31:24];
        layer1[0][7:0] = 0;
        layer1[0][15:8] = 0;
        layer1[0][23:16] = 0;
        layer1[0][31:24] = buffer_data_5[7:0];
        layer1[0][39:32] = buffer_data_5[15:8];
        layer1[0][47:40] = buffer_data_5[23:16];
        layer1[0][55:48] = buffer_data_5[31:24];
        layer2[0][7:0] = 0;
        layer2[0][15:8] = 0;
        layer2[0][23:16] = 0;
        layer2[0][31:24] = buffer_data_4[7:0];
        layer2[0][39:32] = buffer_data_4[15:8];
        layer2[0][47:40] = buffer_data_4[23:16];
        layer2[0][55:48] = buffer_data_4[31:24];
        layer3[0][7:0] = 0;
        layer3[0][15:8] = 0;
        layer3[0][23:16] = 0;
        layer3[0][31:24] = buffer_data_3[7:0];
        layer3[0][39:32] = buffer_data_3[15:8];
        layer3[0][47:40] = buffer_data_3[23:16];
        layer3[0][55:48] = buffer_data_3[31:24];
        layer4[0][7:0] = 0;
        layer4[0][15:8] = 0;
        layer4[0][23:16] = 0;
        layer4[0][31:24] = buffer_data_2[7:0];
        layer4[0][39:32] = buffer_data_2[15:8];
        layer4[0][47:40] = buffer_data_2[23:16];
        layer4[0][55:48] = buffer_data_2[31:24];
        layer5[0][7:0] = 0;
        layer5[0][15:8] = 0;
        layer5[0][23:16] = 0;
        layer5[0][31:24] = buffer_data_1[7:0];
        layer5[0][39:32] = buffer_data_1[15:8];
        layer5[0][47:40] = buffer_data_1[23:16];
        layer5[0][55:48] = buffer_data_1[31:24];
        layer6[0][7:0] = 0;
        layer6[0][15:8] = 0;
        layer6[0][23:16] = 0;
        layer6[0][31:24] = buffer_data_0[7:0];
        layer6[0][39:32] = buffer_data_0[15:8];
        layer6[0][47:40] = buffer_data_0[23:16];
        layer6[0][55:48] = buffer_data_0[31:24];
        layer0[1][7:0] = 0;
        layer0[1][15:8] = 0;
        layer0[1][23:16] = buffer_data_6[7:0];
        layer0[1][31:24] = buffer_data_6[15:8];
        layer0[1][39:32] = buffer_data_6[23:16];
        layer0[1][47:40] = buffer_data_6[31:24];
        layer0[1][55:48] = buffer_data_6[39:32];
        layer1[1][7:0] = 0;
        layer1[1][15:8] = 0;
        layer1[1][23:16] = buffer_data_5[7:0];
        layer1[1][31:24] = buffer_data_5[15:8];
        layer1[1][39:32] = buffer_data_5[23:16];
        layer1[1][47:40] = buffer_data_5[31:24];
        layer1[1][55:48] = buffer_data_5[39:32];
        layer2[1][7:0] = 0;
        layer2[1][15:8] = 0;
        layer2[1][23:16] = buffer_data_4[7:0];
        layer2[1][31:24] = buffer_data_4[15:8];
        layer2[1][39:32] = buffer_data_4[23:16];
        layer2[1][47:40] = buffer_data_4[31:24];
        layer2[1][55:48] = buffer_data_4[39:32];
        layer3[1][7:0] = 0;
        layer3[1][15:8] = 0;
        layer3[1][23:16] = buffer_data_3[7:0];
        layer3[1][31:24] = buffer_data_3[15:8];
        layer3[1][39:32] = buffer_data_3[23:16];
        layer3[1][47:40] = buffer_data_3[31:24];
        layer3[1][55:48] = buffer_data_3[39:32];
        layer4[1][7:0] = 0;
        layer4[1][15:8] = 0;
        layer4[1][23:16] = buffer_data_2[7:0];
        layer4[1][31:24] = buffer_data_2[15:8];
        layer4[1][39:32] = buffer_data_2[23:16];
        layer4[1][47:40] = buffer_data_2[31:24];
        layer4[1][55:48] = buffer_data_2[39:32];
        layer5[1][7:0] = 0;
        layer5[1][15:8] = 0;
        layer5[1][23:16] = buffer_data_1[7:0];
        layer5[1][31:24] = buffer_data_1[15:8];
        layer5[1][39:32] = buffer_data_1[23:16];
        layer5[1][47:40] = buffer_data_1[31:24];
        layer5[1][55:48] = buffer_data_1[39:32];
        layer6[1][7:0] = 0;
        layer6[1][15:8] = 0;
        layer6[1][23:16] = buffer_data_0[7:0];
        layer6[1][31:24] = buffer_data_0[15:8];
        layer6[1][39:32] = buffer_data_0[23:16];
        layer6[1][47:40] = buffer_data_0[31:24];
        layer6[1][55:48] = buffer_data_0[39:32];
        layer0[2][7:0] = 0;
        layer0[2][15:8] = buffer_data_6[7:0];
        layer0[2][23:16] = buffer_data_6[15:8];
        layer0[2][31:24] = buffer_data_6[23:16];
        layer0[2][39:32] = buffer_data_6[31:24];
        layer0[2][47:40] = buffer_data_6[39:32];
        layer0[2][55:48] = buffer_data_6[47:40];
        layer1[2][7:0] = 0;
        layer1[2][15:8] = buffer_data_5[7:0];
        layer1[2][23:16] = buffer_data_5[15:8];
        layer1[2][31:24] = buffer_data_5[23:16];
        layer1[2][39:32] = buffer_data_5[31:24];
        layer1[2][47:40] = buffer_data_5[39:32];
        layer1[2][55:48] = buffer_data_5[47:40];
        layer2[2][7:0] = 0;
        layer2[2][15:8] = buffer_data_4[7:0];
        layer2[2][23:16] = buffer_data_4[15:8];
        layer2[2][31:24] = buffer_data_4[23:16];
        layer2[2][39:32] = buffer_data_4[31:24];
        layer2[2][47:40] = buffer_data_4[39:32];
        layer2[2][55:48] = buffer_data_4[47:40];
        layer3[2][7:0] = 0;
        layer3[2][15:8] = buffer_data_3[7:0];
        layer3[2][23:16] = buffer_data_3[15:8];
        layer3[2][31:24] = buffer_data_3[23:16];
        layer3[2][39:32] = buffer_data_3[31:24];
        layer3[2][47:40] = buffer_data_3[39:32];
        layer3[2][55:48] = buffer_data_3[47:40];
        layer4[2][7:0] = 0;
        layer4[2][15:8] = buffer_data_2[7:0];
        layer4[2][23:16] = buffer_data_2[15:8];
        layer4[2][31:24] = buffer_data_2[23:16];
        layer4[2][39:32] = buffer_data_2[31:24];
        layer4[2][47:40] = buffer_data_2[39:32];
        layer4[2][55:48] = buffer_data_2[47:40];
        layer5[2][7:0] = 0;
        layer5[2][15:8] = buffer_data_1[7:0];
        layer5[2][23:16] = buffer_data_1[15:8];
        layer5[2][31:24] = buffer_data_1[23:16];
        layer5[2][39:32] = buffer_data_1[31:24];
        layer5[2][47:40] = buffer_data_1[39:32];
        layer5[2][55:48] = buffer_data_1[47:40];
        layer6[2][7:0] = 0;
        layer6[2][15:8] = buffer_data_0[7:0];
        layer6[2][23:16] = buffer_data_0[15:8];
        layer6[2][31:24] = buffer_data_0[23:16];
        layer6[2][39:32] = buffer_data_0[31:24];
        layer6[2][47:40] = buffer_data_0[39:32];
        layer6[2][55:48] = buffer_data_0[47:40];
        layer0[3][7:0] = buffer_data_6[7:0];
        layer0[3][15:8] = buffer_data_6[15:8];
        layer0[3][23:16] = buffer_data_6[23:16];
        layer0[3][31:24] = buffer_data_6[31:24];
        layer0[3][39:32] = buffer_data_6[39:32];
        layer0[3][47:40] = buffer_data_6[47:40];
        layer0[3][55:48] = buffer_data_6[55:48];
        layer1[3][7:0] = buffer_data_5[7:0];
        layer1[3][15:8] = buffer_data_5[15:8];
        layer1[3][23:16] = buffer_data_5[23:16];
        layer1[3][31:24] = buffer_data_5[31:24];
        layer1[3][39:32] = buffer_data_5[39:32];
        layer1[3][47:40] = buffer_data_5[47:40];
        layer1[3][55:48] = buffer_data_5[55:48];
        layer2[3][7:0] = buffer_data_4[7:0];
        layer2[3][15:8] = buffer_data_4[15:8];
        layer2[3][23:16] = buffer_data_4[23:16];
        layer2[3][31:24] = buffer_data_4[31:24];
        layer2[3][39:32] = buffer_data_4[39:32];
        layer2[3][47:40] = buffer_data_4[47:40];
        layer2[3][55:48] = buffer_data_4[55:48];
        layer3[3][7:0] = buffer_data_3[7:0];
        layer3[3][15:8] = buffer_data_3[15:8];
        layer3[3][23:16] = buffer_data_3[23:16];
        layer3[3][31:24] = buffer_data_3[31:24];
        layer3[3][39:32] = buffer_data_3[39:32];
        layer3[3][47:40] = buffer_data_3[47:40];
        layer3[3][55:48] = buffer_data_3[55:48];
        layer4[3][7:0] = buffer_data_2[7:0];
        layer4[3][15:8] = buffer_data_2[15:8];
        layer4[3][23:16] = buffer_data_2[23:16];
        layer4[3][31:24] = buffer_data_2[31:24];
        layer4[3][39:32] = buffer_data_2[39:32];
        layer4[3][47:40] = buffer_data_2[47:40];
        layer4[3][55:48] = buffer_data_2[55:48];
        layer5[3][7:0] = buffer_data_1[7:0];
        layer5[3][15:8] = buffer_data_1[15:8];
        layer5[3][23:16] = buffer_data_1[23:16];
        layer5[3][31:24] = buffer_data_1[31:24];
        layer5[3][39:32] = buffer_data_1[39:32];
        layer5[3][47:40] = buffer_data_1[47:40];
        layer5[3][55:48] = buffer_data_1[55:48];
        layer6[3][7:0] = buffer_data_0[7:0];
        layer6[3][15:8] = buffer_data_0[15:8];
        layer6[3][23:16] = buffer_data_0[23:16];
        layer6[3][31:24] = buffer_data_0[31:24];
        layer6[3][39:32] = buffer_data_0[39:32];
        layer6[3][47:40] = buffer_data_0[47:40];
        layer6[3][55:48] = buffer_data_0[55:48];
        layer0[4][7:0] = buffer_data_6[15:8];
        layer0[4][15:8] = buffer_data_6[23:16];
        layer0[4][23:16] = buffer_data_6[31:24];
        layer0[4][31:24] = buffer_data_6[39:32];
        layer0[4][39:32] = buffer_data_6[47:40];
        layer0[4][47:40] = buffer_data_6[55:48];
        layer0[4][55:48] = buffer_data_6[63:56];
        layer1[4][7:0] = buffer_data_5[15:8];
        layer1[4][15:8] = buffer_data_5[23:16];
        layer1[4][23:16] = buffer_data_5[31:24];
        layer1[4][31:24] = buffer_data_5[39:32];
        layer1[4][39:32] = buffer_data_5[47:40];
        layer1[4][47:40] = buffer_data_5[55:48];
        layer1[4][55:48] = buffer_data_5[63:56];
        layer2[4][7:0] = buffer_data_4[15:8];
        layer2[4][15:8] = buffer_data_4[23:16];
        layer2[4][23:16] = buffer_data_4[31:24];
        layer2[4][31:24] = buffer_data_4[39:32];
        layer2[4][39:32] = buffer_data_4[47:40];
        layer2[4][47:40] = buffer_data_4[55:48];
        layer2[4][55:48] = buffer_data_4[63:56];
        layer3[4][7:0] = buffer_data_3[15:8];
        layer3[4][15:8] = buffer_data_3[23:16];
        layer3[4][23:16] = buffer_data_3[31:24];
        layer3[4][31:24] = buffer_data_3[39:32];
        layer3[4][39:32] = buffer_data_3[47:40];
        layer3[4][47:40] = buffer_data_3[55:48];
        layer3[4][55:48] = buffer_data_3[63:56];
        layer4[4][7:0] = buffer_data_2[15:8];
        layer4[4][15:8] = buffer_data_2[23:16];
        layer4[4][23:16] = buffer_data_2[31:24];
        layer4[4][31:24] = buffer_data_2[39:32];
        layer4[4][39:32] = buffer_data_2[47:40];
        layer4[4][47:40] = buffer_data_2[55:48];
        layer4[4][55:48] = buffer_data_2[63:56];
        layer5[4][7:0] = buffer_data_1[15:8];
        layer5[4][15:8] = buffer_data_1[23:16];
        layer5[4][23:16] = buffer_data_1[31:24];
        layer5[4][31:24] = buffer_data_1[39:32];
        layer5[4][39:32] = buffer_data_1[47:40];
        layer5[4][47:40] = buffer_data_1[55:48];
        layer5[4][55:48] = buffer_data_1[63:56];
        layer6[4][7:0] = buffer_data_0[15:8];
        layer6[4][15:8] = buffer_data_0[23:16];
        layer6[4][23:16] = buffer_data_0[31:24];
        layer6[4][31:24] = buffer_data_0[39:32];
        layer6[4][39:32] = buffer_data_0[47:40];
        layer6[4][47:40] = buffer_data_0[55:48];
        layer6[4][55:48] = buffer_data_0[63:56];
        layer0[5][7:0] = buffer_data_6[23:16];
        layer0[5][15:8] = buffer_data_6[31:24];
        layer0[5][23:16] = buffer_data_6[39:32];
        layer0[5][31:24] = buffer_data_6[47:40];
        layer0[5][39:32] = buffer_data_6[55:48];
        layer0[5][47:40] = buffer_data_6[63:56];
        layer0[5][55:48] = buffer_data_6[71:64];
        layer1[5][7:0] = buffer_data_5[23:16];
        layer1[5][15:8] = buffer_data_5[31:24];
        layer1[5][23:16] = buffer_data_5[39:32];
        layer1[5][31:24] = buffer_data_5[47:40];
        layer1[5][39:32] = buffer_data_5[55:48];
        layer1[5][47:40] = buffer_data_5[63:56];
        layer1[5][55:48] = buffer_data_5[71:64];
        layer2[5][7:0] = buffer_data_4[23:16];
        layer2[5][15:8] = buffer_data_4[31:24];
        layer2[5][23:16] = buffer_data_4[39:32];
        layer2[5][31:24] = buffer_data_4[47:40];
        layer2[5][39:32] = buffer_data_4[55:48];
        layer2[5][47:40] = buffer_data_4[63:56];
        layer2[5][55:48] = buffer_data_4[71:64];
        layer3[5][7:0] = buffer_data_3[23:16];
        layer3[5][15:8] = buffer_data_3[31:24];
        layer3[5][23:16] = buffer_data_3[39:32];
        layer3[5][31:24] = buffer_data_3[47:40];
        layer3[5][39:32] = buffer_data_3[55:48];
        layer3[5][47:40] = buffer_data_3[63:56];
        layer3[5][55:48] = buffer_data_3[71:64];
        layer4[5][7:0] = buffer_data_2[23:16];
        layer4[5][15:8] = buffer_data_2[31:24];
        layer4[5][23:16] = buffer_data_2[39:32];
        layer4[5][31:24] = buffer_data_2[47:40];
        layer4[5][39:32] = buffer_data_2[55:48];
        layer4[5][47:40] = buffer_data_2[63:56];
        layer4[5][55:48] = buffer_data_2[71:64];
        layer5[5][7:0] = buffer_data_1[23:16];
        layer5[5][15:8] = buffer_data_1[31:24];
        layer5[5][23:16] = buffer_data_1[39:32];
        layer5[5][31:24] = buffer_data_1[47:40];
        layer5[5][39:32] = buffer_data_1[55:48];
        layer5[5][47:40] = buffer_data_1[63:56];
        layer5[5][55:48] = buffer_data_1[71:64];
        layer6[5][7:0] = buffer_data_0[23:16];
        layer6[5][15:8] = buffer_data_0[31:24];
        layer6[5][23:16] = buffer_data_0[39:32];
        layer6[5][31:24] = buffer_data_0[47:40];
        layer6[5][39:32] = buffer_data_0[55:48];
        layer6[5][47:40] = buffer_data_0[63:56];
        layer6[5][55:48] = buffer_data_0[71:64];
        layer0[6][7:0] = buffer_data_6[31:24];
        layer0[6][15:8] = buffer_data_6[39:32];
        layer0[6][23:16] = buffer_data_6[47:40];
        layer0[6][31:24] = buffer_data_6[55:48];
        layer0[6][39:32] = buffer_data_6[63:56];
        layer0[6][47:40] = buffer_data_6[71:64];
        layer0[6][55:48] = buffer_data_6[79:72];
        layer1[6][7:0] = buffer_data_5[31:24];
        layer1[6][15:8] = buffer_data_5[39:32];
        layer1[6][23:16] = buffer_data_5[47:40];
        layer1[6][31:24] = buffer_data_5[55:48];
        layer1[6][39:32] = buffer_data_5[63:56];
        layer1[6][47:40] = buffer_data_5[71:64];
        layer1[6][55:48] = buffer_data_5[79:72];
        layer2[6][7:0] = buffer_data_4[31:24];
        layer2[6][15:8] = buffer_data_4[39:32];
        layer2[6][23:16] = buffer_data_4[47:40];
        layer2[6][31:24] = buffer_data_4[55:48];
        layer2[6][39:32] = buffer_data_4[63:56];
        layer2[6][47:40] = buffer_data_4[71:64];
        layer2[6][55:48] = buffer_data_4[79:72];
        layer3[6][7:0] = buffer_data_3[31:24];
        layer3[6][15:8] = buffer_data_3[39:32];
        layer3[6][23:16] = buffer_data_3[47:40];
        layer3[6][31:24] = buffer_data_3[55:48];
        layer3[6][39:32] = buffer_data_3[63:56];
        layer3[6][47:40] = buffer_data_3[71:64];
        layer3[6][55:48] = buffer_data_3[79:72];
        layer4[6][7:0] = buffer_data_2[31:24];
        layer4[6][15:8] = buffer_data_2[39:32];
        layer4[6][23:16] = buffer_data_2[47:40];
        layer4[6][31:24] = buffer_data_2[55:48];
        layer4[6][39:32] = buffer_data_2[63:56];
        layer4[6][47:40] = buffer_data_2[71:64];
        layer4[6][55:48] = buffer_data_2[79:72];
        layer5[6][7:0] = buffer_data_1[31:24];
        layer5[6][15:8] = buffer_data_1[39:32];
        layer5[6][23:16] = buffer_data_1[47:40];
        layer5[6][31:24] = buffer_data_1[55:48];
        layer5[6][39:32] = buffer_data_1[63:56];
        layer5[6][47:40] = buffer_data_1[71:64];
        layer5[6][55:48] = buffer_data_1[79:72];
        layer6[6][7:0] = buffer_data_0[31:24];
        layer6[6][15:8] = buffer_data_0[39:32];
        layer6[6][23:16] = buffer_data_0[47:40];
        layer6[6][31:24] = buffer_data_0[55:48];
        layer6[6][39:32] = buffer_data_0[63:56];
        layer6[6][47:40] = buffer_data_0[71:64];
        layer6[6][55:48] = buffer_data_0[79:72];
        layer0[7][7:0] = buffer_data_6[39:32];
        layer0[7][15:8] = buffer_data_6[47:40];
        layer0[7][23:16] = buffer_data_6[55:48];
        layer0[7][31:24] = buffer_data_6[63:56];
        layer0[7][39:32] = buffer_data_6[71:64];
        layer0[7][47:40] = buffer_data_6[79:72];
        layer0[7][55:48] = buffer_data_6[87:80];
        layer1[7][7:0] = buffer_data_5[39:32];
        layer1[7][15:8] = buffer_data_5[47:40];
        layer1[7][23:16] = buffer_data_5[55:48];
        layer1[7][31:24] = buffer_data_5[63:56];
        layer1[7][39:32] = buffer_data_5[71:64];
        layer1[7][47:40] = buffer_data_5[79:72];
        layer1[7][55:48] = buffer_data_5[87:80];
        layer2[7][7:0] = buffer_data_4[39:32];
        layer2[7][15:8] = buffer_data_4[47:40];
        layer2[7][23:16] = buffer_data_4[55:48];
        layer2[7][31:24] = buffer_data_4[63:56];
        layer2[7][39:32] = buffer_data_4[71:64];
        layer2[7][47:40] = buffer_data_4[79:72];
        layer2[7][55:48] = buffer_data_4[87:80];
        layer3[7][7:0] = buffer_data_3[39:32];
        layer3[7][15:8] = buffer_data_3[47:40];
        layer3[7][23:16] = buffer_data_3[55:48];
        layer3[7][31:24] = buffer_data_3[63:56];
        layer3[7][39:32] = buffer_data_3[71:64];
        layer3[7][47:40] = buffer_data_3[79:72];
        layer3[7][55:48] = buffer_data_3[87:80];
        layer4[7][7:0] = buffer_data_2[39:32];
        layer4[7][15:8] = buffer_data_2[47:40];
        layer4[7][23:16] = buffer_data_2[55:48];
        layer4[7][31:24] = buffer_data_2[63:56];
        layer4[7][39:32] = buffer_data_2[71:64];
        layer4[7][47:40] = buffer_data_2[79:72];
        layer4[7][55:48] = buffer_data_2[87:80];
        layer5[7][7:0] = buffer_data_1[39:32];
        layer5[7][15:8] = buffer_data_1[47:40];
        layer5[7][23:16] = buffer_data_1[55:48];
        layer5[7][31:24] = buffer_data_1[63:56];
        layer5[7][39:32] = buffer_data_1[71:64];
        layer5[7][47:40] = buffer_data_1[79:72];
        layer5[7][55:48] = buffer_data_1[87:80];
        layer6[7][7:0] = buffer_data_0[39:32];
        layer6[7][15:8] = buffer_data_0[47:40];
        layer6[7][23:16] = buffer_data_0[55:48];
        layer6[7][31:24] = buffer_data_0[63:56];
        layer6[7][39:32] = buffer_data_0[71:64];
        layer6[7][47:40] = buffer_data_0[79:72];
        layer6[7][55:48] = buffer_data_0[87:80];
        layer0[8][7:0] = buffer_data_6[47:40];
        layer0[8][15:8] = buffer_data_6[55:48];
        layer0[8][23:16] = buffer_data_6[63:56];
        layer0[8][31:24] = buffer_data_6[71:64];
        layer0[8][39:32] = buffer_data_6[79:72];
        layer0[8][47:40] = buffer_data_6[87:80];
        layer0[8][55:48] = buffer_data_6[95:88];
        layer1[8][7:0] = buffer_data_5[47:40];
        layer1[8][15:8] = buffer_data_5[55:48];
        layer1[8][23:16] = buffer_data_5[63:56];
        layer1[8][31:24] = buffer_data_5[71:64];
        layer1[8][39:32] = buffer_data_5[79:72];
        layer1[8][47:40] = buffer_data_5[87:80];
        layer1[8][55:48] = buffer_data_5[95:88];
        layer2[8][7:0] = buffer_data_4[47:40];
        layer2[8][15:8] = buffer_data_4[55:48];
        layer2[8][23:16] = buffer_data_4[63:56];
        layer2[8][31:24] = buffer_data_4[71:64];
        layer2[8][39:32] = buffer_data_4[79:72];
        layer2[8][47:40] = buffer_data_4[87:80];
        layer2[8][55:48] = buffer_data_4[95:88];
        layer3[8][7:0] = buffer_data_3[47:40];
        layer3[8][15:8] = buffer_data_3[55:48];
        layer3[8][23:16] = buffer_data_3[63:56];
        layer3[8][31:24] = buffer_data_3[71:64];
        layer3[8][39:32] = buffer_data_3[79:72];
        layer3[8][47:40] = buffer_data_3[87:80];
        layer3[8][55:48] = buffer_data_3[95:88];
        layer4[8][7:0] = buffer_data_2[47:40];
        layer4[8][15:8] = buffer_data_2[55:48];
        layer4[8][23:16] = buffer_data_2[63:56];
        layer4[8][31:24] = buffer_data_2[71:64];
        layer4[8][39:32] = buffer_data_2[79:72];
        layer4[8][47:40] = buffer_data_2[87:80];
        layer4[8][55:48] = buffer_data_2[95:88];
        layer5[8][7:0] = buffer_data_1[47:40];
        layer5[8][15:8] = buffer_data_1[55:48];
        layer5[8][23:16] = buffer_data_1[63:56];
        layer5[8][31:24] = buffer_data_1[71:64];
        layer5[8][39:32] = buffer_data_1[79:72];
        layer5[8][47:40] = buffer_data_1[87:80];
        layer5[8][55:48] = buffer_data_1[95:88];
        layer6[8][7:0] = buffer_data_0[47:40];
        layer6[8][15:8] = buffer_data_0[55:48];
        layer6[8][23:16] = buffer_data_0[63:56];
        layer6[8][31:24] = buffer_data_0[71:64];
        layer6[8][39:32] = buffer_data_0[79:72];
        layer6[8][47:40] = buffer_data_0[87:80];
        layer6[8][55:48] = buffer_data_0[95:88];
        layer0[9][7:0] = buffer_data_6[55:48];
        layer0[9][15:8] = buffer_data_6[63:56];
        layer0[9][23:16] = buffer_data_6[71:64];
        layer0[9][31:24] = buffer_data_6[79:72];
        layer0[9][39:32] = buffer_data_6[87:80];
        layer0[9][47:40] = buffer_data_6[95:88];
        layer0[9][55:48] = buffer_data_6[103:96];
        layer1[9][7:0] = buffer_data_5[55:48];
        layer1[9][15:8] = buffer_data_5[63:56];
        layer1[9][23:16] = buffer_data_5[71:64];
        layer1[9][31:24] = buffer_data_5[79:72];
        layer1[9][39:32] = buffer_data_5[87:80];
        layer1[9][47:40] = buffer_data_5[95:88];
        layer1[9][55:48] = buffer_data_5[103:96];
        layer2[9][7:0] = buffer_data_4[55:48];
        layer2[9][15:8] = buffer_data_4[63:56];
        layer2[9][23:16] = buffer_data_4[71:64];
        layer2[9][31:24] = buffer_data_4[79:72];
        layer2[9][39:32] = buffer_data_4[87:80];
        layer2[9][47:40] = buffer_data_4[95:88];
        layer2[9][55:48] = buffer_data_4[103:96];
        layer3[9][7:0] = buffer_data_3[55:48];
        layer3[9][15:8] = buffer_data_3[63:56];
        layer3[9][23:16] = buffer_data_3[71:64];
        layer3[9][31:24] = buffer_data_3[79:72];
        layer3[9][39:32] = buffer_data_3[87:80];
        layer3[9][47:40] = buffer_data_3[95:88];
        layer3[9][55:48] = buffer_data_3[103:96];
        layer4[9][7:0] = buffer_data_2[55:48];
        layer4[9][15:8] = buffer_data_2[63:56];
        layer4[9][23:16] = buffer_data_2[71:64];
        layer4[9][31:24] = buffer_data_2[79:72];
        layer4[9][39:32] = buffer_data_2[87:80];
        layer4[9][47:40] = buffer_data_2[95:88];
        layer4[9][55:48] = buffer_data_2[103:96];
        layer5[9][7:0] = buffer_data_1[55:48];
        layer5[9][15:8] = buffer_data_1[63:56];
        layer5[9][23:16] = buffer_data_1[71:64];
        layer5[9][31:24] = buffer_data_1[79:72];
        layer5[9][39:32] = buffer_data_1[87:80];
        layer5[9][47:40] = buffer_data_1[95:88];
        layer5[9][55:48] = buffer_data_1[103:96];
        layer6[9][7:0] = buffer_data_0[55:48];
        layer6[9][15:8] = buffer_data_0[63:56];
        layer6[9][23:16] = buffer_data_0[71:64];
        layer6[9][31:24] = buffer_data_0[79:72];
        layer6[9][39:32] = buffer_data_0[87:80];
        layer6[9][47:40] = buffer_data_0[95:88];
        layer6[9][55:48] = buffer_data_0[103:96];
        layer0[10][7:0] = buffer_data_6[63:56];
        layer0[10][15:8] = buffer_data_6[71:64];
        layer0[10][23:16] = buffer_data_6[79:72];
        layer0[10][31:24] = buffer_data_6[87:80];
        layer0[10][39:32] = buffer_data_6[95:88];
        layer0[10][47:40] = buffer_data_6[103:96];
        layer0[10][55:48] = buffer_data_6[111:104];
        layer1[10][7:0] = buffer_data_5[63:56];
        layer1[10][15:8] = buffer_data_5[71:64];
        layer1[10][23:16] = buffer_data_5[79:72];
        layer1[10][31:24] = buffer_data_5[87:80];
        layer1[10][39:32] = buffer_data_5[95:88];
        layer1[10][47:40] = buffer_data_5[103:96];
        layer1[10][55:48] = buffer_data_5[111:104];
        layer2[10][7:0] = buffer_data_4[63:56];
        layer2[10][15:8] = buffer_data_4[71:64];
        layer2[10][23:16] = buffer_data_4[79:72];
        layer2[10][31:24] = buffer_data_4[87:80];
        layer2[10][39:32] = buffer_data_4[95:88];
        layer2[10][47:40] = buffer_data_4[103:96];
        layer2[10][55:48] = buffer_data_4[111:104];
        layer3[10][7:0] = buffer_data_3[63:56];
        layer3[10][15:8] = buffer_data_3[71:64];
        layer3[10][23:16] = buffer_data_3[79:72];
        layer3[10][31:24] = buffer_data_3[87:80];
        layer3[10][39:32] = buffer_data_3[95:88];
        layer3[10][47:40] = buffer_data_3[103:96];
        layer3[10][55:48] = buffer_data_3[111:104];
        layer4[10][7:0] = buffer_data_2[63:56];
        layer4[10][15:8] = buffer_data_2[71:64];
        layer4[10][23:16] = buffer_data_2[79:72];
        layer4[10][31:24] = buffer_data_2[87:80];
        layer4[10][39:32] = buffer_data_2[95:88];
        layer4[10][47:40] = buffer_data_2[103:96];
        layer4[10][55:48] = buffer_data_2[111:104];
        layer5[10][7:0] = buffer_data_1[63:56];
        layer5[10][15:8] = buffer_data_1[71:64];
        layer5[10][23:16] = buffer_data_1[79:72];
        layer5[10][31:24] = buffer_data_1[87:80];
        layer5[10][39:32] = buffer_data_1[95:88];
        layer5[10][47:40] = buffer_data_1[103:96];
        layer5[10][55:48] = buffer_data_1[111:104];
        layer6[10][7:0] = buffer_data_0[63:56];
        layer6[10][15:8] = buffer_data_0[71:64];
        layer6[10][23:16] = buffer_data_0[79:72];
        layer6[10][31:24] = buffer_data_0[87:80];
        layer6[10][39:32] = buffer_data_0[95:88];
        layer6[10][47:40] = buffer_data_0[103:96];
        layer6[10][55:48] = buffer_data_0[111:104];
        layer0[11][7:0] = buffer_data_6[71:64];
        layer0[11][15:8] = buffer_data_6[79:72];
        layer0[11][23:16] = buffer_data_6[87:80];
        layer0[11][31:24] = buffer_data_6[95:88];
        layer0[11][39:32] = buffer_data_6[103:96];
        layer0[11][47:40] = buffer_data_6[111:104];
        layer0[11][55:48] = buffer_data_6[119:112];
        layer1[11][7:0] = buffer_data_5[71:64];
        layer1[11][15:8] = buffer_data_5[79:72];
        layer1[11][23:16] = buffer_data_5[87:80];
        layer1[11][31:24] = buffer_data_5[95:88];
        layer1[11][39:32] = buffer_data_5[103:96];
        layer1[11][47:40] = buffer_data_5[111:104];
        layer1[11][55:48] = buffer_data_5[119:112];
        layer2[11][7:0] = buffer_data_4[71:64];
        layer2[11][15:8] = buffer_data_4[79:72];
        layer2[11][23:16] = buffer_data_4[87:80];
        layer2[11][31:24] = buffer_data_4[95:88];
        layer2[11][39:32] = buffer_data_4[103:96];
        layer2[11][47:40] = buffer_data_4[111:104];
        layer2[11][55:48] = buffer_data_4[119:112];
        layer3[11][7:0] = buffer_data_3[71:64];
        layer3[11][15:8] = buffer_data_3[79:72];
        layer3[11][23:16] = buffer_data_3[87:80];
        layer3[11][31:24] = buffer_data_3[95:88];
        layer3[11][39:32] = buffer_data_3[103:96];
        layer3[11][47:40] = buffer_data_3[111:104];
        layer3[11][55:48] = buffer_data_3[119:112];
        layer4[11][7:0] = buffer_data_2[71:64];
        layer4[11][15:8] = buffer_data_2[79:72];
        layer4[11][23:16] = buffer_data_2[87:80];
        layer4[11][31:24] = buffer_data_2[95:88];
        layer4[11][39:32] = buffer_data_2[103:96];
        layer4[11][47:40] = buffer_data_2[111:104];
        layer4[11][55:48] = buffer_data_2[119:112];
        layer5[11][7:0] = buffer_data_1[71:64];
        layer5[11][15:8] = buffer_data_1[79:72];
        layer5[11][23:16] = buffer_data_1[87:80];
        layer5[11][31:24] = buffer_data_1[95:88];
        layer5[11][39:32] = buffer_data_1[103:96];
        layer5[11][47:40] = buffer_data_1[111:104];
        layer5[11][55:48] = buffer_data_1[119:112];
        layer6[11][7:0] = buffer_data_0[71:64];
        layer6[11][15:8] = buffer_data_0[79:72];
        layer6[11][23:16] = buffer_data_0[87:80];
        layer6[11][31:24] = buffer_data_0[95:88];
        layer6[11][39:32] = buffer_data_0[103:96];
        layer6[11][47:40] = buffer_data_0[111:104];
        layer6[11][55:48] = buffer_data_0[119:112];
        layer0[12][7:0] = buffer_data_6[79:72];
        layer0[12][15:8] = buffer_data_6[87:80];
        layer0[12][23:16] = buffer_data_6[95:88];
        layer0[12][31:24] = buffer_data_6[103:96];
        layer0[12][39:32] = buffer_data_6[111:104];
        layer0[12][47:40] = buffer_data_6[119:112];
        layer0[12][55:48] = buffer_data_6[127:120];
        layer1[12][7:0] = buffer_data_5[79:72];
        layer1[12][15:8] = buffer_data_5[87:80];
        layer1[12][23:16] = buffer_data_5[95:88];
        layer1[12][31:24] = buffer_data_5[103:96];
        layer1[12][39:32] = buffer_data_5[111:104];
        layer1[12][47:40] = buffer_data_5[119:112];
        layer1[12][55:48] = buffer_data_5[127:120];
        layer2[12][7:0] = buffer_data_4[79:72];
        layer2[12][15:8] = buffer_data_4[87:80];
        layer2[12][23:16] = buffer_data_4[95:88];
        layer2[12][31:24] = buffer_data_4[103:96];
        layer2[12][39:32] = buffer_data_4[111:104];
        layer2[12][47:40] = buffer_data_4[119:112];
        layer2[12][55:48] = buffer_data_4[127:120];
        layer3[12][7:0] = buffer_data_3[79:72];
        layer3[12][15:8] = buffer_data_3[87:80];
        layer3[12][23:16] = buffer_data_3[95:88];
        layer3[12][31:24] = buffer_data_3[103:96];
        layer3[12][39:32] = buffer_data_3[111:104];
        layer3[12][47:40] = buffer_data_3[119:112];
        layer3[12][55:48] = buffer_data_3[127:120];
        layer4[12][7:0] = buffer_data_2[79:72];
        layer4[12][15:8] = buffer_data_2[87:80];
        layer4[12][23:16] = buffer_data_2[95:88];
        layer4[12][31:24] = buffer_data_2[103:96];
        layer4[12][39:32] = buffer_data_2[111:104];
        layer4[12][47:40] = buffer_data_2[119:112];
        layer4[12][55:48] = buffer_data_2[127:120];
        layer5[12][7:0] = buffer_data_1[79:72];
        layer5[12][15:8] = buffer_data_1[87:80];
        layer5[12][23:16] = buffer_data_1[95:88];
        layer5[12][31:24] = buffer_data_1[103:96];
        layer5[12][39:32] = buffer_data_1[111:104];
        layer5[12][47:40] = buffer_data_1[119:112];
        layer5[12][55:48] = buffer_data_1[127:120];
        layer6[12][7:0] = buffer_data_0[79:72];
        layer6[12][15:8] = buffer_data_0[87:80];
        layer6[12][23:16] = buffer_data_0[95:88];
        layer6[12][31:24] = buffer_data_0[103:96];
        layer6[12][39:32] = buffer_data_0[111:104];
        layer6[12][47:40] = buffer_data_0[119:112];
        layer6[12][55:48] = buffer_data_0[127:120];
        layer0[13][7:0] = buffer_data_6[87:80];
        layer0[13][15:8] = buffer_data_6[95:88];
        layer0[13][23:16] = buffer_data_6[103:96];
        layer0[13][31:24] = buffer_data_6[111:104];
        layer0[13][39:32] = buffer_data_6[119:112];
        layer0[13][47:40] = buffer_data_6[127:120];
        layer0[13][55:48] = buffer_data_6[135:128];
        layer1[13][7:0] = buffer_data_5[87:80];
        layer1[13][15:8] = buffer_data_5[95:88];
        layer1[13][23:16] = buffer_data_5[103:96];
        layer1[13][31:24] = buffer_data_5[111:104];
        layer1[13][39:32] = buffer_data_5[119:112];
        layer1[13][47:40] = buffer_data_5[127:120];
        layer1[13][55:48] = buffer_data_5[135:128];
        layer2[13][7:0] = buffer_data_4[87:80];
        layer2[13][15:8] = buffer_data_4[95:88];
        layer2[13][23:16] = buffer_data_4[103:96];
        layer2[13][31:24] = buffer_data_4[111:104];
        layer2[13][39:32] = buffer_data_4[119:112];
        layer2[13][47:40] = buffer_data_4[127:120];
        layer2[13][55:48] = buffer_data_4[135:128];
        layer3[13][7:0] = buffer_data_3[87:80];
        layer3[13][15:8] = buffer_data_3[95:88];
        layer3[13][23:16] = buffer_data_3[103:96];
        layer3[13][31:24] = buffer_data_3[111:104];
        layer3[13][39:32] = buffer_data_3[119:112];
        layer3[13][47:40] = buffer_data_3[127:120];
        layer3[13][55:48] = buffer_data_3[135:128];
        layer4[13][7:0] = buffer_data_2[87:80];
        layer4[13][15:8] = buffer_data_2[95:88];
        layer4[13][23:16] = buffer_data_2[103:96];
        layer4[13][31:24] = buffer_data_2[111:104];
        layer4[13][39:32] = buffer_data_2[119:112];
        layer4[13][47:40] = buffer_data_2[127:120];
        layer4[13][55:48] = buffer_data_2[135:128];
        layer5[13][7:0] = buffer_data_1[87:80];
        layer5[13][15:8] = buffer_data_1[95:88];
        layer5[13][23:16] = buffer_data_1[103:96];
        layer5[13][31:24] = buffer_data_1[111:104];
        layer5[13][39:32] = buffer_data_1[119:112];
        layer5[13][47:40] = buffer_data_1[127:120];
        layer5[13][55:48] = buffer_data_1[135:128];
        layer6[13][7:0] = buffer_data_0[87:80];
        layer6[13][15:8] = buffer_data_0[95:88];
        layer6[13][23:16] = buffer_data_0[103:96];
        layer6[13][31:24] = buffer_data_0[111:104];
        layer6[13][39:32] = buffer_data_0[119:112];
        layer6[13][47:40] = buffer_data_0[127:120];
        layer6[13][55:48] = buffer_data_0[135:128];
        layer0[14][7:0] = buffer_data_6[95:88];
        layer0[14][15:8] = buffer_data_6[103:96];
        layer0[14][23:16] = buffer_data_6[111:104];
        layer0[14][31:24] = buffer_data_6[119:112];
        layer0[14][39:32] = buffer_data_6[127:120];
        layer0[14][47:40] = buffer_data_6[135:128];
        layer0[14][55:48] = buffer_data_6[143:136];
        layer1[14][7:0] = buffer_data_5[95:88];
        layer1[14][15:8] = buffer_data_5[103:96];
        layer1[14][23:16] = buffer_data_5[111:104];
        layer1[14][31:24] = buffer_data_5[119:112];
        layer1[14][39:32] = buffer_data_5[127:120];
        layer1[14][47:40] = buffer_data_5[135:128];
        layer1[14][55:48] = buffer_data_5[143:136];
        layer2[14][7:0] = buffer_data_4[95:88];
        layer2[14][15:8] = buffer_data_4[103:96];
        layer2[14][23:16] = buffer_data_4[111:104];
        layer2[14][31:24] = buffer_data_4[119:112];
        layer2[14][39:32] = buffer_data_4[127:120];
        layer2[14][47:40] = buffer_data_4[135:128];
        layer2[14][55:48] = buffer_data_4[143:136];
        layer3[14][7:0] = buffer_data_3[95:88];
        layer3[14][15:8] = buffer_data_3[103:96];
        layer3[14][23:16] = buffer_data_3[111:104];
        layer3[14][31:24] = buffer_data_3[119:112];
        layer3[14][39:32] = buffer_data_3[127:120];
        layer3[14][47:40] = buffer_data_3[135:128];
        layer3[14][55:48] = buffer_data_3[143:136];
        layer4[14][7:0] = buffer_data_2[95:88];
        layer4[14][15:8] = buffer_data_2[103:96];
        layer4[14][23:16] = buffer_data_2[111:104];
        layer4[14][31:24] = buffer_data_2[119:112];
        layer4[14][39:32] = buffer_data_2[127:120];
        layer4[14][47:40] = buffer_data_2[135:128];
        layer4[14][55:48] = buffer_data_2[143:136];
        layer5[14][7:0] = buffer_data_1[95:88];
        layer5[14][15:8] = buffer_data_1[103:96];
        layer5[14][23:16] = buffer_data_1[111:104];
        layer5[14][31:24] = buffer_data_1[119:112];
        layer5[14][39:32] = buffer_data_1[127:120];
        layer5[14][47:40] = buffer_data_1[135:128];
        layer5[14][55:48] = buffer_data_1[143:136];
        layer6[14][7:0] = buffer_data_0[95:88];
        layer6[14][15:8] = buffer_data_0[103:96];
        layer6[14][23:16] = buffer_data_0[111:104];
        layer6[14][31:24] = buffer_data_0[119:112];
        layer6[14][39:32] = buffer_data_0[127:120];
        layer6[14][47:40] = buffer_data_0[135:128];
        layer6[14][55:48] = buffer_data_0[143:136];
        layer0[15][7:0] = buffer_data_6[103:96];
        layer0[15][15:8] = buffer_data_6[111:104];
        layer0[15][23:16] = buffer_data_6[119:112];
        layer0[15][31:24] = buffer_data_6[127:120];
        layer0[15][39:32] = buffer_data_6[135:128];
        layer0[15][47:40] = buffer_data_6[143:136];
        layer0[15][55:48] = buffer_data_6[151:144];
        layer1[15][7:0] = buffer_data_5[103:96];
        layer1[15][15:8] = buffer_data_5[111:104];
        layer1[15][23:16] = buffer_data_5[119:112];
        layer1[15][31:24] = buffer_data_5[127:120];
        layer1[15][39:32] = buffer_data_5[135:128];
        layer1[15][47:40] = buffer_data_5[143:136];
        layer1[15][55:48] = buffer_data_5[151:144];
        layer2[15][7:0] = buffer_data_4[103:96];
        layer2[15][15:8] = buffer_data_4[111:104];
        layer2[15][23:16] = buffer_data_4[119:112];
        layer2[15][31:24] = buffer_data_4[127:120];
        layer2[15][39:32] = buffer_data_4[135:128];
        layer2[15][47:40] = buffer_data_4[143:136];
        layer2[15][55:48] = buffer_data_4[151:144];
        layer3[15][7:0] = buffer_data_3[103:96];
        layer3[15][15:8] = buffer_data_3[111:104];
        layer3[15][23:16] = buffer_data_3[119:112];
        layer3[15][31:24] = buffer_data_3[127:120];
        layer3[15][39:32] = buffer_data_3[135:128];
        layer3[15][47:40] = buffer_data_3[143:136];
        layer3[15][55:48] = buffer_data_3[151:144];
        layer4[15][7:0] = buffer_data_2[103:96];
        layer4[15][15:8] = buffer_data_2[111:104];
        layer4[15][23:16] = buffer_data_2[119:112];
        layer4[15][31:24] = buffer_data_2[127:120];
        layer4[15][39:32] = buffer_data_2[135:128];
        layer4[15][47:40] = buffer_data_2[143:136];
        layer4[15][55:48] = buffer_data_2[151:144];
        layer5[15][7:0] = buffer_data_1[103:96];
        layer5[15][15:8] = buffer_data_1[111:104];
        layer5[15][23:16] = buffer_data_1[119:112];
        layer5[15][31:24] = buffer_data_1[127:120];
        layer5[15][39:32] = buffer_data_1[135:128];
        layer5[15][47:40] = buffer_data_1[143:136];
        layer5[15][55:48] = buffer_data_1[151:144];
        layer6[15][7:0] = buffer_data_0[103:96];
        layer6[15][15:8] = buffer_data_0[111:104];
        layer6[15][23:16] = buffer_data_0[119:112];
        layer6[15][31:24] = buffer_data_0[127:120];
        layer6[15][39:32] = buffer_data_0[135:128];
        layer6[15][47:40] = buffer_data_0[143:136];
        layer6[15][55:48] = buffer_data_0[151:144];
        layer0[16][7:0] = buffer_data_6[111:104];
        layer0[16][15:8] = buffer_data_6[119:112];
        layer0[16][23:16] = buffer_data_6[127:120];
        layer0[16][31:24] = buffer_data_6[135:128];
        layer0[16][39:32] = buffer_data_6[143:136];
        layer0[16][47:40] = buffer_data_6[151:144];
        layer0[16][55:48] = buffer_data_6[159:152];
        layer1[16][7:0] = buffer_data_5[111:104];
        layer1[16][15:8] = buffer_data_5[119:112];
        layer1[16][23:16] = buffer_data_5[127:120];
        layer1[16][31:24] = buffer_data_5[135:128];
        layer1[16][39:32] = buffer_data_5[143:136];
        layer1[16][47:40] = buffer_data_5[151:144];
        layer1[16][55:48] = buffer_data_5[159:152];
        layer2[16][7:0] = buffer_data_4[111:104];
        layer2[16][15:8] = buffer_data_4[119:112];
        layer2[16][23:16] = buffer_data_4[127:120];
        layer2[16][31:24] = buffer_data_4[135:128];
        layer2[16][39:32] = buffer_data_4[143:136];
        layer2[16][47:40] = buffer_data_4[151:144];
        layer2[16][55:48] = buffer_data_4[159:152];
        layer3[16][7:0] = buffer_data_3[111:104];
        layer3[16][15:8] = buffer_data_3[119:112];
        layer3[16][23:16] = buffer_data_3[127:120];
        layer3[16][31:24] = buffer_data_3[135:128];
        layer3[16][39:32] = buffer_data_3[143:136];
        layer3[16][47:40] = buffer_data_3[151:144];
        layer3[16][55:48] = buffer_data_3[159:152];
        layer4[16][7:0] = buffer_data_2[111:104];
        layer4[16][15:8] = buffer_data_2[119:112];
        layer4[16][23:16] = buffer_data_2[127:120];
        layer4[16][31:24] = buffer_data_2[135:128];
        layer4[16][39:32] = buffer_data_2[143:136];
        layer4[16][47:40] = buffer_data_2[151:144];
        layer4[16][55:48] = buffer_data_2[159:152];
        layer5[16][7:0] = buffer_data_1[111:104];
        layer5[16][15:8] = buffer_data_1[119:112];
        layer5[16][23:16] = buffer_data_1[127:120];
        layer5[16][31:24] = buffer_data_1[135:128];
        layer5[16][39:32] = buffer_data_1[143:136];
        layer5[16][47:40] = buffer_data_1[151:144];
        layer5[16][55:48] = buffer_data_1[159:152];
        layer6[16][7:0] = buffer_data_0[111:104];
        layer6[16][15:8] = buffer_data_0[119:112];
        layer6[16][23:16] = buffer_data_0[127:120];
        layer6[16][31:24] = buffer_data_0[135:128];
        layer6[16][39:32] = buffer_data_0[143:136];
        layer6[16][47:40] = buffer_data_0[151:144];
        layer6[16][55:48] = buffer_data_0[159:152];
        layer0[17][7:0] = buffer_data_6[119:112];
        layer0[17][15:8] = buffer_data_6[127:120];
        layer0[17][23:16] = buffer_data_6[135:128];
        layer0[17][31:24] = buffer_data_6[143:136];
        layer0[17][39:32] = buffer_data_6[151:144];
        layer0[17][47:40] = buffer_data_6[159:152];
        layer0[17][55:48] = buffer_data_6[167:160];
        layer1[17][7:0] = buffer_data_5[119:112];
        layer1[17][15:8] = buffer_data_5[127:120];
        layer1[17][23:16] = buffer_data_5[135:128];
        layer1[17][31:24] = buffer_data_5[143:136];
        layer1[17][39:32] = buffer_data_5[151:144];
        layer1[17][47:40] = buffer_data_5[159:152];
        layer1[17][55:48] = buffer_data_5[167:160];
        layer2[17][7:0] = buffer_data_4[119:112];
        layer2[17][15:8] = buffer_data_4[127:120];
        layer2[17][23:16] = buffer_data_4[135:128];
        layer2[17][31:24] = buffer_data_4[143:136];
        layer2[17][39:32] = buffer_data_4[151:144];
        layer2[17][47:40] = buffer_data_4[159:152];
        layer2[17][55:48] = buffer_data_4[167:160];
        layer3[17][7:0] = buffer_data_3[119:112];
        layer3[17][15:8] = buffer_data_3[127:120];
        layer3[17][23:16] = buffer_data_3[135:128];
        layer3[17][31:24] = buffer_data_3[143:136];
        layer3[17][39:32] = buffer_data_3[151:144];
        layer3[17][47:40] = buffer_data_3[159:152];
        layer3[17][55:48] = buffer_data_3[167:160];
        layer4[17][7:0] = buffer_data_2[119:112];
        layer4[17][15:8] = buffer_data_2[127:120];
        layer4[17][23:16] = buffer_data_2[135:128];
        layer4[17][31:24] = buffer_data_2[143:136];
        layer4[17][39:32] = buffer_data_2[151:144];
        layer4[17][47:40] = buffer_data_2[159:152];
        layer4[17][55:48] = buffer_data_2[167:160];
        layer5[17][7:0] = buffer_data_1[119:112];
        layer5[17][15:8] = buffer_data_1[127:120];
        layer5[17][23:16] = buffer_data_1[135:128];
        layer5[17][31:24] = buffer_data_1[143:136];
        layer5[17][39:32] = buffer_data_1[151:144];
        layer5[17][47:40] = buffer_data_1[159:152];
        layer5[17][55:48] = buffer_data_1[167:160];
        layer6[17][7:0] = buffer_data_0[119:112];
        layer6[17][15:8] = buffer_data_0[127:120];
        layer6[17][23:16] = buffer_data_0[135:128];
        layer6[17][31:24] = buffer_data_0[143:136];
        layer6[17][39:32] = buffer_data_0[151:144];
        layer6[17][47:40] = buffer_data_0[159:152];
        layer6[17][55:48] = buffer_data_0[167:160];
        layer0[18][7:0] = buffer_data_6[127:120];
        layer0[18][15:8] = buffer_data_6[135:128];
        layer0[18][23:16] = buffer_data_6[143:136];
        layer0[18][31:24] = buffer_data_6[151:144];
        layer0[18][39:32] = buffer_data_6[159:152];
        layer0[18][47:40] = buffer_data_6[167:160];
        layer0[18][55:48] = buffer_data_6[175:168];
        layer1[18][7:0] = buffer_data_5[127:120];
        layer1[18][15:8] = buffer_data_5[135:128];
        layer1[18][23:16] = buffer_data_5[143:136];
        layer1[18][31:24] = buffer_data_5[151:144];
        layer1[18][39:32] = buffer_data_5[159:152];
        layer1[18][47:40] = buffer_data_5[167:160];
        layer1[18][55:48] = buffer_data_5[175:168];
        layer2[18][7:0] = buffer_data_4[127:120];
        layer2[18][15:8] = buffer_data_4[135:128];
        layer2[18][23:16] = buffer_data_4[143:136];
        layer2[18][31:24] = buffer_data_4[151:144];
        layer2[18][39:32] = buffer_data_4[159:152];
        layer2[18][47:40] = buffer_data_4[167:160];
        layer2[18][55:48] = buffer_data_4[175:168];
        layer3[18][7:0] = buffer_data_3[127:120];
        layer3[18][15:8] = buffer_data_3[135:128];
        layer3[18][23:16] = buffer_data_3[143:136];
        layer3[18][31:24] = buffer_data_3[151:144];
        layer3[18][39:32] = buffer_data_3[159:152];
        layer3[18][47:40] = buffer_data_3[167:160];
        layer3[18][55:48] = buffer_data_3[175:168];
        layer4[18][7:0] = buffer_data_2[127:120];
        layer4[18][15:8] = buffer_data_2[135:128];
        layer4[18][23:16] = buffer_data_2[143:136];
        layer4[18][31:24] = buffer_data_2[151:144];
        layer4[18][39:32] = buffer_data_2[159:152];
        layer4[18][47:40] = buffer_data_2[167:160];
        layer4[18][55:48] = buffer_data_2[175:168];
        layer5[18][7:0] = buffer_data_1[127:120];
        layer5[18][15:8] = buffer_data_1[135:128];
        layer5[18][23:16] = buffer_data_1[143:136];
        layer5[18][31:24] = buffer_data_1[151:144];
        layer5[18][39:32] = buffer_data_1[159:152];
        layer5[18][47:40] = buffer_data_1[167:160];
        layer5[18][55:48] = buffer_data_1[175:168];
        layer6[18][7:0] = buffer_data_0[127:120];
        layer6[18][15:8] = buffer_data_0[135:128];
        layer6[18][23:16] = buffer_data_0[143:136];
        layer6[18][31:24] = buffer_data_0[151:144];
        layer6[18][39:32] = buffer_data_0[159:152];
        layer6[18][47:40] = buffer_data_0[167:160];
        layer6[18][55:48] = buffer_data_0[175:168];
        layer0[19][7:0] = buffer_data_6[135:128];
        layer0[19][15:8] = buffer_data_6[143:136];
        layer0[19][23:16] = buffer_data_6[151:144];
        layer0[19][31:24] = buffer_data_6[159:152];
        layer0[19][39:32] = buffer_data_6[167:160];
        layer0[19][47:40] = buffer_data_6[175:168];
        layer0[19][55:48] = buffer_data_6[183:176];
        layer1[19][7:0] = buffer_data_5[135:128];
        layer1[19][15:8] = buffer_data_5[143:136];
        layer1[19][23:16] = buffer_data_5[151:144];
        layer1[19][31:24] = buffer_data_5[159:152];
        layer1[19][39:32] = buffer_data_5[167:160];
        layer1[19][47:40] = buffer_data_5[175:168];
        layer1[19][55:48] = buffer_data_5[183:176];
        layer2[19][7:0] = buffer_data_4[135:128];
        layer2[19][15:8] = buffer_data_4[143:136];
        layer2[19][23:16] = buffer_data_4[151:144];
        layer2[19][31:24] = buffer_data_4[159:152];
        layer2[19][39:32] = buffer_data_4[167:160];
        layer2[19][47:40] = buffer_data_4[175:168];
        layer2[19][55:48] = buffer_data_4[183:176];
        layer3[19][7:0] = buffer_data_3[135:128];
        layer3[19][15:8] = buffer_data_3[143:136];
        layer3[19][23:16] = buffer_data_3[151:144];
        layer3[19][31:24] = buffer_data_3[159:152];
        layer3[19][39:32] = buffer_data_3[167:160];
        layer3[19][47:40] = buffer_data_3[175:168];
        layer3[19][55:48] = buffer_data_3[183:176];
        layer4[19][7:0] = buffer_data_2[135:128];
        layer4[19][15:8] = buffer_data_2[143:136];
        layer4[19][23:16] = buffer_data_2[151:144];
        layer4[19][31:24] = buffer_data_2[159:152];
        layer4[19][39:32] = buffer_data_2[167:160];
        layer4[19][47:40] = buffer_data_2[175:168];
        layer4[19][55:48] = buffer_data_2[183:176];
        layer5[19][7:0] = buffer_data_1[135:128];
        layer5[19][15:8] = buffer_data_1[143:136];
        layer5[19][23:16] = buffer_data_1[151:144];
        layer5[19][31:24] = buffer_data_1[159:152];
        layer5[19][39:32] = buffer_data_1[167:160];
        layer5[19][47:40] = buffer_data_1[175:168];
        layer5[19][55:48] = buffer_data_1[183:176];
        layer6[19][7:0] = buffer_data_0[135:128];
        layer6[19][15:8] = buffer_data_0[143:136];
        layer6[19][23:16] = buffer_data_0[151:144];
        layer6[19][31:24] = buffer_data_0[159:152];
        layer6[19][39:32] = buffer_data_0[167:160];
        layer6[19][47:40] = buffer_data_0[175:168];
        layer6[19][55:48] = buffer_data_0[183:176];
        layer0[20][7:0] = buffer_data_6[143:136];
        layer0[20][15:8] = buffer_data_6[151:144];
        layer0[20][23:16] = buffer_data_6[159:152];
        layer0[20][31:24] = buffer_data_6[167:160];
        layer0[20][39:32] = buffer_data_6[175:168];
        layer0[20][47:40] = buffer_data_6[183:176];
        layer0[20][55:48] = buffer_data_6[191:184];
        layer1[20][7:0] = buffer_data_5[143:136];
        layer1[20][15:8] = buffer_data_5[151:144];
        layer1[20][23:16] = buffer_data_5[159:152];
        layer1[20][31:24] = buffer_data_5[167:160];
        layer1[20][39:32] = buffer_data_5[175:168];
        layer1[20][47:40] = buffer_data_5[183:176];
        layer1[20][55:48] = buffer_data_5[191:184];
        layer2[20][7:0] = buffer_data_4[143:136];
        layer2[20][15:8] = buffer_data_4[151:144];
        layer2[20][23:16] = buffer_data_4[159:152];
        layer2[20][31:24] = buffer_data_4[167:160];
        layer2[20][39:32] = buffer_data_4[175:168];
        layer2[20][47:40] = buffer_data_4[183:176];
        layer2[20][55:48] = buffer_data_4[191:184];
        layer3[20][7:0] = buffer_data_3[143:136];
        layer3[20][15:8] = buffer_data_3[151:144];
        layer3[20][23:16] = buffer_data_3[159:152];
        layer3[20][31:24] = buffer_data_3[167:160];
        layer3[20][39:32] = buffer_data_3[175:168];
        layer3[20][47:40] = buffer_data_3[183:176];
        layer3[20][55:48] = buffer_data_3[191:184];
        layer4[20][7:0] = buffer_data_2[143:136];
        layer4[20][15:8] = buffer_data_2[151:144];
        layer4[20][23:16] = buffer_data_2[159:152];
        layer4[20][31:24] = buffer_data_2[167:160];
        layer4[20][39:32] = buffer_data_2[175:168];
        layer4[20][47:40] = buffer_data_2[183:176];
        layer4[20][55:48] = buffer_data_2[191:184];
        layer5[20][7:0] = buffer_data_1[143:136];
        layer5[20][15:8] = buffer_data_1[151:144];
        layer5[20][23:16] = buffer_data_1[159:152];
        layer5[20][31:24] = buffer_data_1[167:160];
        layer5[20][39:32] = buffer_data_1[175:168];
        layer5[20][47:40] = buffer_data_1[183:176];
        layer5[20][55:48] = buffer_data_1[191:184];
        layer6[20][7:0] = buffer_data_0[143:136];
        layer6[20][15:8] = buffer_data_0[151:144];
        layer6[20][23:16] = buffer_data_0[159:152];
        layer6[20][31:24] = buffer_data_0[167:160];
        layer6[20][39:32] = buffer_data_0[175:168];
        layer6[20][47:40] = buffer_data_0[183:176];
        layer6[20][55:48] = buffer_data_0[191:184];
        layer0[21][7:0] = buffer_data_6[151:144];
        layer0[21][15:8] = buffer_data_6[159:152];
        layer0[21][23:16] = buffer_data_6[167:160];
        layer0[21][31:24] = buffer_data_6[175:168];
        layer0[21][39:32] = buffer_data_6[183:176];
        layer0[21][47:40] = buffer_data_6[191:184];
        layer0[21][55:48] = buffer_data_6[199:192];
        layer1[21][7:0] = buffer_data_5[151:144];
        layer1[21][15:8] = buffer_data_5[159:152];
        layer1[21][23:16] = buffer_data_5[167:160];
        layer1[21][31:24] = buffer_data_5[175:168];
        layer1[21][39:32] = buffer_data_5[183:176];
        layer1[21][47:40] = buffer_data_5[191:184];
        layer1[21][55:48] = buffer_data_5[199:192];
        layer2[21][7:0] = buffer_data_4[151:144];
        layer2[21][15:8] = buffer_data_4[159:152];
        layer2[21][23:16] = buffer_data_4[167:160];
        layer2[21][31:24] = buffer_data_4[175:168];
        layer2[21][39:32] = buffer_data_4[183:176];
        layer2[21][47:40] = buffer_data_4[191:184];
        layer2[21][55:48] = buffer_data_4[199:192];
        layer3[21][7:0] = buffer_data_3[151:144];
        layer3[21][15:8] = buffer_data_3[159:152];
        layer3[21][23:16] = buffer_data_3[167:160];
        layer3[21][31:24] = buffer_data_3[175:168];
        layer3[21][39:32] = buffer_data_3[183:176];
        layer3[21][47:40] = buffer_data_3[191:184];
        layer3[21][55:48] = buffer_data_3[199:192];
        layer4[21][7:0] = buffer_data_2[151:144];
        layer4[21][15:8] = buffer_data_2[159:152];
        layer4[21][23:16] = buffer_data_2[167:160];
        layer4[21][31:24] = buffer_data_2[175:168];
        layer4[21][39:32] = buffer_data_2[183:176];
        layer4[21][47:40] = buffer_data_2[191:184];
        layer4[21][55:48] = buffer_data_2[199:192];
        layer5[21][7:0] = buffer_data_1[151:144];
        layer5[21][15:8] = buffer_data_1[159:152];
        layer5[21][23:16] = buffer_data_1[167:160];
        layer5[21][31:24] = buffer_data_1[175:168];
        layer5[21][39:32] = buffer_data_1[183:176];
        layer5[21][47:40] = buffer_data_1[191:184];
        layer5[21][55:48] = buffer_data_1[199:192];
        layer6[21][7:0] = buffer_data_0[151:144];
        layer6[21][15:8] = buffer_data_0[159:152];
        layer6[21][23:16] = buffer_data_0[167:160];
        layer6[21][31:24] = buffer_data_0[175:168];
        layer6[21][39:32] = buffer_data_0[183:176];
        layer6[21][47:40] = buffer_data_0[191:184];
        layer6[21][55:48] = buffer_data_0[199:192];
        layer0[22][7:0] = buffer_data_6[159:152];
        layer0[22][15:8] = buffer_data_6[167:160];
        layer0[22][23:16] = buffer_data_6[175:168];
        layer0[22][31:24] = buffer_data_6[183:176];
        layer0[22][39:32] = buffer_data_6[191:184];
        layer0[22][47:40] = buffer_data_6[199:192];
        layer0[22][55:48] = buffer_data_6[207:200];
        layer1[22][7:0] = buffer_data_5[159:152];
        layer1[22][15:8] = buffer_data_5[167:160];
        layer1[22][23:16] = buffer_data_5[175:168];
        layer1[22][31:24] = buffer_data_5[183:176];
        layer1[22][39:32] = buffer_data_5[191:184];
        layer1[22][47:40] = buffer_data_5[199:192];
        layer1[22][55:48] = buffer_data_5[207:200];
        layer2[22][7:0] = buffer_data_4[159:152];
        layer2[22][15:8] = buffer_data_4[167:160];
        layer2[22][23:16] = buffer_data_4[175:168];
        layer2[22][31:24] = buffer_data_4[183:176];
        layer2[22][39:32] = buffer_data_4[191:184];
        layer2[22][47:40] = buffer_data_4[199:192];
        layer2[22][55:48] = buffer_data_4[207:200];
        layer3[22][7:0] = buffer_data_3[159:152];
        layer3[22][15:8] = buffer_data_3[167:160];
        layer3[22][23:16] = buffer_data_3[175:168];
        layer3[22][31:24] = buffer_data_3[183:176];
        layer3[22][39:32] = buffer_data_3[191:184];
        layer3[22][47:40] = buffer_data_3[199:192];
        layer3[22][55:48] = buffer_data_3[207:200];
        layer4[22][7:0] = buffer_data_2[159:152];
        layer4[22][15:8] = buffer_data_2[167:160];
        layer4[22][23:16] = buffer_data_2[175:168];
        layer4[22][31:24] = buffer_data_2[183:176];
        layer4[22][39:32] = buffer_data_2[191:184];
        layer4[22][47:40] = buffer_data_2[199:192];
        layer4[22][55:48] = buffer_data_2[207:200];
        layer5[22][7:0] = buffer_data_1[159:152];
        layer5[22][15:8] = buffer_data_1[167:160];
        layer5[22][23:16] = buffer_data_1[175:168];
        layer5[22][31:24] = buffer_data_1[183:176];
        layer5[22][39:32] = buffer_data_1[191:184];
        layer5[22][47:40] = buffer_data_1[199:192];
        layer5[22][55:48] = buffer_data_1[207:200];
        layer6[22][7:0] = buffer_data_0[159:152];
        layer6[22][15:8] = buffer_data_0[167:160];
        layer6[22][23:16] = buffer_data_0[175:168];
        layer6[22][31:24] = buffer_data_0[183:176];
        layer6[22][39:32] = buffer_data_0[191:184];
        layer6[22][47:40] = buffer_data_0[199:192];
        layer6[22][55:48] = buffer_data_0[207:200];
        layer0[23][7:0] = buffer_data_6[167:160];
        layer0[23][15:8] = buffer_data_6[175:168];
        layer0[23][23:16] = buffer_data_6[183:176];
        layer0[23][31:24] = buffer_data_6[191:184];
        layer0[23][39:32] = buffer_data_6[199:192];
        layer0[23][47:40] = buffer_data_6[207:200];
        layer0[23][55:48] = buffer_data_6[215:208];
        layer1[23][7:0] = buffer_data_5[167:160];
        layer1[23][15:8] = buffer_data_5[175:168];
        layer1[23][23:16] = buffer_data_5[183:176];
        layer1[23][31:24] = buffer_data_5[191:184];
        layer1[23][39:32] = buffer_data_5[199:192];
        layer1[23][47:40] = buffer_data_5[207:200];
        layer1[23][55:48] = buffer_data_5[215:208];
        layer2[23][7:0] = buffer_data_4[167:160];
        layer2[23][15:8] = buffer_data_4[175:168];
        layer2[23][23:16] = buffer_data_4[183:176];
        layer2[23][31:24] = buffer_data_4[191:184];
        layer2[23][39:32] = buffer_data_4[199:192];
        layer2[23][47:40] = buffer_data_4[207:200];
        layer2[23][55:48] = buffer_data_4[215:208];
        layer3[23][7:0] = buffer_data_3[167:160];
        layer3[23][15:8] = buffer_data_3[175:168];
        layer3[23][23:16] = buffer_data_3[183:176];
        layer3[23][31:24] = buffer_data_3[191:184];
        layer3[23][39:32] = buffer_data_3[199:192];
        layer3[23][47:40] = buffer_data_3[207:200];
        layer3[23][55:48] = buffer_data_3[215:208];
        layer4[23][7:0] = buffer_data_2[167:160];
        layer4[23][15:8] = buffer_data_2[175:168];
        layer4[23][23:16] = buffer_data_2[183:176];
        layer4[23][31:24] = buffer_data_2[191:184];
        layer4[23][39:32] = buffer_data_2[199:192];
        layer4[23][47:40] = buffer_data_2[207:200];
        layer4[23][55:48] = buffer_data_2[215:208];
        layer5[23][7:0] = buffer_data_1[167:160];
        layer5[23][15:8] = buffer_data_1[175:168];
        layer5[23][23:16] = buffer_data_1[183:176];
        layer5[23][31:24] = buffer_data_1[191:184];
        layer5[23][39:32] = buffer_data_1[199:192];
        layer5[23][47:40] = buffer_data_1[207:200];
        layer5[23][55:48] = buffer_data_1[215:208];
        layer6[23][7:0] = buffer_data_0[167:160];
        layer6[23][15:8] = buffer_data_0[175:168];
        layer6[23][23:16] = buffer_data_0[183:176];
        layer6[23][31:24] = buffer_data_0[191:184];
        layer6[23][39:32] = buffer_data_0[199:192];
        layer6[23][47:40] = buffer_data_0[207:200];
        layer6[23][55:48] = buffer_data_0[215:208];
        layer0[24][7:0] = buffer_data_6[175:168];
        layer0[24][15:8] = buffer_data_6[183:176];
        layer0[24][23:16] = buffer_data_6[191:184];
        layer0[24][31:24] = buffer_data_6[199:192];
        layer0[24][39:32] = buffer_data_6[207:200];
        layer0[24][47:40] = buffer_data_6[215:208];
        layer0[24][55:48] = buffer_data_6[223:216];
        layer1[24][7:0] = buffer_data_5[175:168];
        layer1[24][15:8] = buffer_data_5[183:176];
        layer1[24][23:16] = buffer_data_5[191:184];
        layer1[24][31:24] = buffer_data_5[199:192];
        layer1[24][39:32] = buffer_data_5[207:200];
        layer1[24][47:40] = buffer_data_5[215:208];
        layer1[24][55:48] = buffer_data_5[223:216];
        layer2[24][7:0] = buffer_data_4[175:168];
        layer2[24][15:8] = buffer_data_4[183:176];
        layer2[24][23:16] = buffer_data_4[191:184];
        layer2[24][31:24] = buffer_data_4[199:192];
        layer2[24][39:32] = buffer_data_4[207:200];
        layer2[24][47:40] = buffer_data_4[215:208];
        layer2[24][55:48] = buffer_data_4[223:216];
        layer3[24][7:0] = buffer_data_3[175:168];
        layer3[24][15:8] = buffer_data_3[183:176];
        layer3[24][23:16] = buffer_data_3[191:184];
        layer3[24][31:24] = buffer_data_3[199:192];
        layer3[24][39:32] = buffer_data_3[207:200];
        layer3[24][47:40] = buffer_data_3[215:208];
        layer3[24][55:48] = buffer_data_3[223:216];
        layer4[24][7:0] = buffer_data_2[175:168];
        layer4[24][15:8] = buffer_data_2[183:176];
        layer4[24][23:16] = buffer_data_2[191:184];
        layer4[24][31:24] = buffer_data_2[199:192];
        layer4[24][39:32] = buffer_data_2[207:200];
        layer4[24][47:40] = buffer_data_2[215:208];
        layer4[24][55:48] = buffer_data_2[223:216];
        layer5[24][7:0] = buffer_data_1[175:168];
        layer5[24][15:8] = buffer_data_1[183:176];
        layer5[24][23:16] = buffer_data_1[191:184];
        layer5[24][31:24] = buffer_data_1[199:192];
        layer5[24][39:32] = buffer_data_1[207:200];
        layer5[24][47:40] = buffer_data_1[215:208];
        layer5[24][55:48] = buffer_data_1[223:216];
        layer6[24][7:0] = buffer_data_0[175:168];
        layer6[24][15:8] = buffer_data_0[183:176];
        layer6[24][23:16] = buffer_data_0[191:184];
        layer6[24][31:24] = buffer_data_0[199:192];
        layer6[24][39:32] = buffer_data_0[207:200];
        layer6[24][47:40] = buffer_data_0[215:208];
        layer6[24][55:48] = buffer_data_0[223:216];
        layer0[25][7:0] = buffer_data_6[183:176];
        layer0[25][15:8] = buffer_data_6[191:184];
        layer0[25][23:16] = buffer_data_6[199:192];
        layer0[25][31:24] = buffer_data_6[207:200];
        layer0[25][39:32] = buffer_data_6[215:208];
        layer0[25][47:40] = buffer_data_6[223:216];
        layer0[25][55:48] = buffer_data_6[231:224];
        layer1[25][7:0] = buffer_data_5[183:176];
        layer1[25][15:8] = buffer_data_5[191:184];
        layer1[25][23:16] = buffer_data_5[199:192];
        layer1[25][31:24] = buffer_data_5[207:200];
        layer1[25][39:32] = buffer_data_5[215:208];
        layer1[25][47:40] = buffer_data_5[223:216];
        layer1[25][55:48] = buffer_data_5[231:224];
        layer2[25][7:0] = buffer_data_4[183:176];
        layer2[25][15:8] = buffer_data_4[191:184];
        layer2[25][23:16] = buffer_data_4[199:192];
        layer2[25][31:24] = buffer_data_4[207:200];
        layer2[25][39:32] = buffer_data_4[215:208];
        layer2[25][47:40] = buffer_data_4[223:216];
        layer2[25][55:48] = buffer_data_4[231:224];
        layer3[25][7:0] = buffer_data_3[183:176];
        layer3[25][15:8] = buffer_data_3[191:184];
        layer3[25][23:16] = buffer_data_3[199:192];
        layer3[25][31:24] = buffer_data_3[207:200];
        layer3[25][39:32] = buffer_data_3[215:208];
        layer3[25][47:40] = buffer_data_3[223:216];
        layer3[25][55:48] = buffer_data_3[231:224];
        layer4[25][7:0] = buffer_data_2[183:176];
        layer4[25][15:8] = buffer_data_2[191:184];
        layer4[25][23:16] = buffer_data_2[199:192];
        layer4[25][31:24] = buffer_data_2[207:200];
        layer4[25][39:32] = buffer_data_2[215:208];
        layer4[25][47:40] = buffer_data_2[223:216];
        layer4[25][55:48] = buffer_data_2[231:224];
        layer5[25][7:0] = buffer_data_1[183:176];
        layer5[25][15:8] = buffer_data_1[191:184];
        layer5[25][23:16] = buffer_data_1[199:192];
        layer5[25][31:24] = buffer_data_1[207:200];
        layer5[25][39:32] = buffer_data_1[215:208];
        layer5[25][47:40] = buffer_data_1[223:216];
        layer5[25][55:48] = buffer_data_1[231:224];
        layer6[25][7:0] = buffer_data_0[183:176];
        layer6[25][15:8] = buffer_data_0[191:184];
        layer6[25][23:16] = buffer_data_0[199:192];
        layer6[25][31:24] = buffer_data_0[207:200];
        layer6[25][39:32] = buffer_data_0[215:208];
        layer6[25][47:40] = buffer_data_0[223:216];
        layer6[25][55:48] = buffer_data_0[231:224];
        layer0[26][7:0] = buffer_data_6[191:184];
        layer0[26][15:8] = buffer_data_6[199:192];
        layer0[26][23:16] = buffer_data_6[207:200];
        layer0[26][31:24] = buffer_data_6[215:208];
        layer0[26][39:32] = buffer_data_6[223:216];
        layer0[26][47:40] = buffer_data_6[231:224];
        layer0[26][55:48] = buffer_data_6[239:232];
        layer1[26][7:0] = buffer_data_5[191:184];
        layer1[26][15:8] = buffer_data_5[199:192];
        layer1[26][23:16] = buffer_data_5[207:200];
        layer1[26][31:24] = buffer_data_5[215:208];
        layer1[26][39:32] = buffer_data_5[223:216];
        layer1[26][47:40] = buffer_data_5[231:224];
        layer1[26][55:48] = buffer_data_5[239:232];
        layer2[26][7:0] = buffer_data_4[191:184];
        layer2[26][15:8] = buffer_data_4[199:192];
        layer2[26][23:16] = buffer_data_4[207:200];
        layer2[26][31:24] = buffer_data_4[215:208];
        layer2[26][39:32] = buffer_data_4[223:216];
        layer2[26][47:40] = buffer_data_4[231:224];
        layer2[26][55:48] = buffer_data_4[239:232];
        layer3[26][7:0] = buffer_data_3[191:184];
        layer3[26][15:8] = buffer_data_3[199:192];
        layer3[26][23:16] = buffer_data_3[207:200];
        layer3[26][31:24] = buffer_data_3[215:208];
        layer3[26][39:32] = buffer_data_3[223:216];
        layer3[26][47:40] = buffer_data_3[231:224];
        layer3[26][55:48] = buffer_data_3[239:232];
        layer4[26][7:0] = buffer_data_2[191:184];
        layer4[26][15:8] = buffer_data_2[199:192];
        layer4[26][23:16] = buffer_data_2[207:200];
        layer4[26][31:24] = buffer_data_2[215:208];
        layer4[26][39:32] = buffer_data_2[223:216];
        layer4[26][47:40] = buffer_data_2[231:224];
        layer4[26][55:48] = buffer_data_2[239:232];
        layer5[26][7:0] = buffer_data_1[191:184];
        layer5[26][15:8] = buffer_data_1[199:192];
        layer5[26][23:16] = buffer_data_1[207:200];
        layer5[26][31:24] = buffer_data_1[215:208];
        layer5[26][39:32] = buffer_data_1[223:216];
        layer5[26][47:40] = buffer_data_1[231:224];
        layer5[26][55:48] = buffer_data_1[239:232];
        layer6[26][7:0] = buffer_data_0[191:184];
        layer6[26][15:8] = buffer_data_0[199:192];
        layer6[26][23:16] = buffer_data_0[207:200];
        layer6[26][31:24] = buffer_data_0[215:208];
        layer6[26][39:32] = buffer_data_0[223:216];
        layer6[26][47:40] = buffer_data_0[231:224];
        layer6[26][55:48] = buffer_data_0[239:232];
        layer0[27][7:0] = buffer_data_6[199:192];
        layer0[27][15:8] = buffer_data_6[207:200];
        layer0[27][23:16] = buffer_data_6[215:208];
        layer0[27][31:24] = buffer_data_6[223:216];
        layer0[27][39:32] = buffer_data_6[231:224];
        layer0[27][47:40] = buffer_data_6[239:232];
        layer0[27][55:48] = buffer_data_6[247:240];
        layer1[27][7:0] = buffer_data_5[199:192];
        layer1[27][15:8] = buffer_data_5[207:200];
        layer1[27][23:16] = buffer_data_5[215:208];
        layer1[27][31:24] = buffer_data_5[223:216];
        layer1[27][39:32] = buffer_data_5[231:224];
        layer1[27][47:40] = buffer_data_5[239:232];
        layer1[27][55:48] = buffer_data_5[247:240];
        layer2[27][7:0] = buffer_data_4[199:192];
        layer2[27][15:8] = buffer_data_4[207:200];
        layer2[27][23:16] = buffer_data_4[215:208];
        layer2[27][31:24] = buffer_data_4[223:216];
        layer2[27][39:32] = buffer_data_4[231:224];
        layer2[27][47:40] = buffer_data_4[239:232];
        layer2[27][55:48] = buffer_data_4[247:240];
        layer3[27][7:0] = buffer_data_3[199:192];
        layer3[27][15:8] = buffer_data_3[207:200];
        layer3[27][23:16] = buffer_data_3[215:208];
        layer3[27][31:24] = buffer_data_3[223:216];
        layer3[27][39:32] = buffer_data_3[231:224];
        layer3[27][47:40] = buffer_data_3[239:232];
        layer3[27][55:48] = buffer_data_3[247:240];
        layer4[27][7:0] = buffer_data_2[199:192];
        layer4[27][15:8] = buffer_data_2[207:200];
        layer4[27][23:16] = buffer_data_2[215:208];
        layer4[27][31:24] = buffer_data_2[223:216];
        layer4[27][39:32] = buffer_data_2[231:224];
        layer4[27][47:40] = buffer_data_2[239:232];
        layer4[27][55:48] = buffer_data_2[247:240];
        layer5[27][7:0] = buffer_data_1[199:192];
        layer5[27][15:8] = buffer_data_1[207:200];
        layer5[27][23:16] = buffer_data_1[215:208];
        layer5[27][31:24] = buffer_data_1[223:216];
        layer5[27][39:32] = buffer_data_1[231:224];
        layer5[27][47:40] = buffer_data_1[239:232];
        layer5[27][55:48] = buffer_data_1[247:240];
        layer6[27][7:0] = buffer_data_0[199:192];
        layer6[27][15:8] = buffer_data_0[207:200];
        layer6[27][23:16] = buffer_data_0[215:208];
        layer6[27][31:24] = buffer_data_0[223:216];
        layer6[27][39:32] = buffer_data_0[231:224];
        layer6[27][47:40] = buffer_data_0[239:232];
        layer6[27][55:48] = buffer_data_0[247:240];
        layer0[28][7:0] = buffer_data_6[207:200];
        layer0[28][15:8] = buffer_data_6[215:208];
        layer0[28][23:16] = buffer_data_6[223:216];
        layer0[28][31:24] = buffer_data_6[231:224];
        layer0[28][39:32] = buffer_data_6[239:232];
        layer0[28][47:40] = buffer_data_6[247:240];
        layer0[28][55:48] = buffer_data_6[255:248];
        layer1[28][7:0] = buffer_data_5[207:200];
        layer1[28][15:8] = buffer_data_5[215:208];
        layer1[28][23:16] = buffer_data_5[223:216];
        layer1[28][31:24] = buffer_data_5[231:224];
        layer1[28][39:32] = buffer_data_5[239:232];
        layer1[28][47:40] = buffer_data_5[247:240];
        layer1[28][55:48] = buffer_data_5[255:248];
        layer2[28][7:0] = buffer_data_4[207:200];
        layer2[28][15:8] = buffer_data_4[215:208];
        layer2[28][23:16] = buffer_data_4[223:216];
        layer2[28][31:24] = buffer_data_4[231:224];
        layer2[28][39:32] = buffer_data_4[239:232];
        layer2[28][47:40] = buffer_data_4[247:240];
        layer2[28][55:48] = buffer_data_4[255:248];
        layer3[28][7:0] = buffer_data_3[207:200];
        layer3[28][15:8] = buffer_data_3[215:208];
        layer3[28][23:16] = buffer_data_3[223:216];
        layer3[28][31:24] = buffer_data_3[231:224];
        layer3[28][39:32] = buffer_data_3[239:232];
        layer3[28][47:40] = buffer_data_3[247:240];
        layer3[28][55:48] = buffer_data_3[255:248];
        layer4[28][7:0] = buffer_data_2[207:200];
        layer4[28][15:8] = buffer_data_2[215:208];
        layer4[28][23:16] = buffer_data_2[223:216];
        layer4[28][31:24] = buffer_data_2[231:224];
        layer4[28][39:32] = buffer_data_2[239:232];
        layer4[28][47:40] = buffer_data_2[247:240];
        layer4[28][55:48] = buffer_data_2[255:248];
        layer5[28][7:0] = buffer_data_1[207:200];
        layer5[28][15:8] = buffer_data_1[215:208];
        layer5[28][23:16] = buffer_data_1[223:216];
        layer5[28][31:24] = buffer_data_1[231:224];
        layer5[28][39:32] = buffer_data_1[239:232];
        layer5[28][47:40] = buffer_data_1[247:240];
        layer5[28][55:48] = buffer_data_1[255:248];
        layer6[28][7:0] = buffer_data_0[207:200];
        layer6[28][15:8] = buffer_data_0[215:208];
        layer6[28][23:16] = buffer_data_0[223:216];
        layer6[28][31:24] = buffer_data_0[231:224];
        layer6[28][39:32] = buffer_data_0[239:232];
        layer6[28][47:40] = buffer_data_0[247:240];
        layer6[28][55:48] = buffer_data_0[255:248];
        layer0[29][7:0] = buffer_data_6[215:208];
        layer0[29][15:8] = buffer_data_6[223:216];
        layer0[29][23:16] = buffer_data_6[231:224];
        layer0[29][31:24] = buffer_data_6[239:232];
        layer0[29][39:32] = buffer_data_6[247:240];
        layer0[29][47:40] = buffer_data_6[255:248];
        layer0[29][55:48] = buffer_data_6[263:256];
        layer1[29][7:0] = buffer_data_5[215:208];
        layer1[29][15:8] = buffer_data_5[223:216];
        layer1[29][23:16] = buffer_data_5[231:224];
        layer1[29][31:24] = buffer_data_5[239:232];
        layer1[29][39:32] = buffer_data_5[247:240];
        layer1[29][47:40] = buffer_data_5[255:248];
        layer1[29][55:48] = buffer_data_5[263:256];
        layer2[29][7:0] = buffer_data_4[215:208];
        layer2[29][15:8] = buffer_data_4[223:216];
        layer2[29][23:16] = buffer_data_4[231:224];
        layer2[29][31:24] = buffer_data_4[239:232];
        layer2[29][39:32] = buffer_data_4[247:240];
        layer2[29][47:40] = buffer_data_4[255:248];
        layer2[29][55:48] = buffer_data_4[263:256];
        layer3[29][7:0] = buffer_data_3[215:208];
        layer3[29][15:8] = buffer_data_3[223:216];
        layer3[29][23:16] = buffer_data_3[231:224];
        layer3[29][31:24] = buffer_data_3[239:232];
        layer3[29][39:32] = buffer_data_3[247:240];
        layer3[29][47:40] = buffer_data_3[255:248];
        layer3[29][55:48] = buffer_data_3[263:256];
        layer4[29][7:0] = buffer_data_2[215:208];
        layer4[29][15:8] = buffer_data_2[223:216];
        layer4[29][23:16] = buffer_data_2[231:224];
        layer4[29][31:24] = buffer_data_2[239:232];
        layer4[29][39:32] = buffer_data_2[247:240];
        layer4[29][47:40] = buffer_data_2[255:248];
        layer4[29][55:48] = buffer_data_2[263:256];
        layer5[29][7:0] = buffer_data_1[215:208];
        layer5[29][15:8] = buffer_data_1[223:216];
        layer5[29][23:16] = buffer_data_1[231:224];
        layer5[29][31:24] = buffer_data_1[239:232];
        layer5[29][39:32] = buffer_data_1[247:240];
        layer5[29][47:40] = buffer_data_1[255:248];
        layer5[29][55:48] = buffer_data_1[263:256];
        layer6[29][7:0] = buffer_data_0[215:208];
        layer6[29][15:8] = buffer_data_0[223:216];
        layer6[29][23:16] = buffer_data_0[231:224];
        layer6[29][31:24] = buffer_data_0[239:232];
        layer6[29][39:32] = buffer_data_0[247:240];
        layer6[29][47:40] = buffer_data_0[255:248];
        layer6[29][55:48] = buffer_data_0[263:256];
        layer0[30][7:0] = buffer_data_6[223:216];
        layer0[30][15:8] = buffer_data_6[231:224];
        layer0[30][23:16] = buffer_data_6[239:232];
        layer0[30][31:24] = buffer_data_6[247:240];
        layer0[30][39:32] = buffer_data_6[255:248];
        layer0[30][47:40] = buffer_data_6[263:256];
        layer0[30][55:48] = buffer_data_6[271:264];
        layer1[30][7:0] = buffer_data_5[223:216];
        layer1[30][15:8] = buffer_data_5[231:224];
        layer1[30][23:16] = buffer_data_5[239:232];
        layer1[30][31:24] = buffer_data_5[247:240];
        layer1[30][39:32] = buffer_data_5[255:248];
        layer1[30][47:40] = buffer_data_5[263:256];
        layer1[30][55:48] = buffer_data_5[271:264];
        layer2[30][7:0] = buffer_data_4[223:216];
        layer2[30][15:8] = buffer_data_4[231:224];
        layer2[30][23:16] = buffer_data_4[239:232];
        layer2[30][31:24] = buffer_data_4[247:240];
        layer2[30][39:32] = buffer_data_4[255:248];
        layer2[30][47:40] = buffer_data_4[263:256];
        layer2[30][55:48] = buffer_data_4[271:264];
        layer3[30][7:0] = buffer_data_3[223:216];
        layer3[30][15:8] = buffer_data_3[231:224];
        layer3[30][23:16] = buffer_data_3[239:232];
        layer3[30][31:24] = buffer_data_3[247:240];
        layer3[30][39:32] = buffer_data_3[255:248];
        layer3[30][47:40] = buffer_data_3[263:256];
        layer3[30][55:48] = buffer_data_3[271:264];
        layer4[30][7:0] = buffer_data_2[223:216];
        layer4[30][15:8] = buffer_data_2[231:224];
        layer4[30][23:16] = buffer_data_2[239:232];
        layer4[30][31:24] = buffer_data_2[247:240];
        layer4[30][39:32] = buffer_data_2[255:248];
        layer4[30][47:40] = buffer_data_2[263:256];
        layer4[30][55:48] = buffer_data_2[271:264];
        layer5[30][7:0] = buffer_data_1[223:216];
        layer5[30][15:8] = buffer_data_1[231:224];
        layer5[30][23:16] = buffer_data_1[239:232];
        layer5[30][31:24] = buffer_data_1[247:240];
        layer5[30][39:32] = buffer_data_1[255:248];
        layer5[30][47:40] = buffer_data_1[263:256];
        layer5[30][55:48] = buffer_data_1[271:264];
        layer6[30][7:0] = buffer_data_0[223:216];
        layer6[30][15:8] = buffer_data_0[231:224];
        layer6[30][23:16] = buffer_data_0[239:232];
        layer6[30][31:24] = buffer_data_0[247:240];
        layer6[30][39:32] = buffer_data_0[255:248];
        layer6[30][47:40] = buffer_data_0[263:256];
        layer6[30][55:48] = buffer_data_0[271:264];
        layer0[31][7:0] = buffer_data_6[231:224];
        layer0[31][15:8] = buffer_data_6[239:232];
        layer0[31][23:16] = buffer_data_6[247:240];
        layer0[31][31:24] = buffer_data_6[255:248];
        layer0[31][39:32] = buffer_data_6[263:256];
        layer0[31][47:40] = buffer_data_6[271:264];
        layer0[31][55:48] = buffer_data_6[279:272];
        layer1[31][7:0] = buffer_data_5[231:224];
        layer1[31][15:8] = buffer_data_5[239:232];
        layer1[31][23:16] = buffer_data_5[247:240];
        layer1[31][31:24] = buffer_data_5[255:248];
        layer1[31][39:32] = buffer_data_5[263:256];
        layer1[31][47:40] = buffer_data_5[271:264];
        layer1[31][55:48] = buffer_data_5[279:272];
        layer2[31][7:0] = buffer_data_4[231:224];
        layer2[31][15:8] = buffer_data_4[239:232];
        layer2[31][23:16] = buffer_data_4[247:240];
        layer2[31][31:24] = buffer_data_4[255:248];
        layer2[31][39:32] = buffer_data_4[263:256];
        layer2[31][47:40] = buffer_data_4[271:264];
        layer2[31][55:48] = buffer_data_4[279:272];
        layer3[31][7:0] = buffer_data_3[231:224];
        layer3[31][15:8] = buffer_data_3[239:232];
        layer3[31][23:16] = buffer_data_3[247:240];
        layer3[31][31:24] = buffer_data_3[255:248];
        layer3[31][39:32] = buffer_data_3[263:256];
        layer3[31][47:40] = buffer_data_3[271:264];
        layer3[31][55:48] = buffer_data_3[279:272];
        layer4[31][7:0] = buffer_data_2[231:224];
        layer4[31][15:8] = buffer_data_2[239:232];
        layer4[31][23:16] = buffer_data_2[247:240];
        layer4[31][31:24] = buffer_data_2[255:248];
        layer4[31][39:32] = buffer_data_2[263:256];
        layer4[31][47:40] = buffer_data_2[271:264];
        layer4[31][55:48] = buffer_data_2[279:272];
        layer5[31][7:0] = buffer_data_1[231:224];
        layer5[31][15:8] = buffer_data_1[239:232];
        layer5[31][23:16] = buffer_data_1[247:240];
        layer5[31][31:24] = buffer_data_1[255:248];
        layer5[31][39:32] = buffer_data_1[263:256];
        layer5[31][47:40] = buffer_data_1[271:264];
        layer5[31][55:48] = buffer_data_1[279:272];
        layer6[31][7:0] = buffer_data_0[231:224];
        layer6[31][15:8] = buffer_data_0[239:232];
        layer6[31][23:16] = buffer_data_0[247:240];
        layer6[31][31:24] = buffer_data_0[255:248];
        layer6[31][39:32] = buffer_data_0[263:256];
        layer6[31][47:40] = buffer_data_0[271:264];
        layer6[31][55:48] = buffer_data_0[279:272];
        layer0[32][7:0] = buffer_data_6[239:232];
        layer0[32][15:8] = buffer_data_6[247:240];
        layer0[32][23:16] = buffer_data_6[255:248];
        layer0[32][31:24] = buffer_data_6[263:256];
        layer0[32][39:32] = buffer_data_6[271:264];
        layer0[32][47:40] = buffer_data_6[279:272];
        layer0[32][55:48] = buffer_data_6[287:280];
        layer1[32][7:0] = buffer_data_5[239:232];
        layer1[32][15:8] = buffer_data_5[247:240];
        layer1[32][23:16] = buffer_data_5[255:248];
        layer1[32][31:24] = buffer_data_5[263:256];
        layer1[32][39:32] = buffer_data_5[271:264];
        layer1[32][47:40] = buffer_data_5[279:272];
        layer1[32][55:48] = buffer_data_5[287:280];
        layer2[32][7:0] = buffer_data_4[239:232];
        layer2[32][15:8] = buffer_data_4[247:240];
        layer2[32][23:16] = buffer_data_4[255:248];
        layer2[32][31:24] = buffer_data_4[263:256];
        layer2[32][39:32] = buffer_data_4[271:264];
        layer2[32][47:40] = buffer_data_4[279:272];
        layer2[32][55:48] = buffer_data_4[287:280];
        layer3[32][7:0] = buffer_data_3[239:232];
        layer3[32][15:8] = buffer_data_3[247:240];
        layer3[32][23:16] = buffer_data_3[255:248];
        layer3[32][31:24] = buffer_data_3[263:256];
        layer3[32][39:32] = buffer_data_3[271:264];
        layer3[32][47:40] = buffer_data_3[279:272];
        layer3[32][55:48] = buffer_data_3[287:280];
        layer4[32][7:0] = buffer_data_2[239:232];
        layer4[32][15:8] = buffer_data_2[247:240];
        layer4[32][23:16] = buffer_data_2[255:248];
        layer4[32][31:24] = buffer_data_2[263:256];
        layer4[32][39:32] = buffer_data_2[271:264];
        layer4[32][47:40] = buffer_data_2[279:272];
        layer4[32][55:48] = buffer_data_2[287:280];
        layer5[32][7:0] = buffer_data_1[239:232];
        layer5[32][15:8] = buffer_data_1[247:240];
        layer5[32][23:16] = buffer_data_1[255:248];
        layer5[32][31:24] = buffer_data_1[263:256];
        layer5[32][39:32] = buffer_data_1[271:264];
        layer5[32][47:40] = buffer_data_1[279:272];
        layer5[32][55:48] = buffer_data_1[287:280];
        layer6[32][7:0] = buffer_data_0[239:232];
        layer6[32][15:8] = buffer_data_0[247:240];
        layer6[32][23:16] = buffer_data_0[255:248];
        layer6[32][31:24] = buffer_data_0[263:256];
        layer6[32][39:32] = buffer_data_0[271:264];
        layer6[32][47:40] = buffer_data_0[279:272];
        layer6[32][55:48] = buffer_data_0[287:280];
        layer0[33][7:0] = buffer_data_6[247:240];
        layer0[33][15:8] = buffer_data_6[255:248];
        layer0[33][23:16] = buffer_data_6[263:256];
        layer0[33][31:24] = buffer_data_6[271:264];
        layer0[33][39:32] = buffer_data_6[279:272];
        layer0[33][47:40] = buffer_data_6[287:280];
        layer0[33][55:48] = buffer_data_6[295:288];
        layer1[33][7:0] = buffer_data_5[247:240];
        layer1[33][15:8] = buffer_data_5[255:248];
        layer1[33][23:16] = buffer_data_5[263:256];
        layer1[33][31:24] = buffer_data_5[271:264];
        layer1[33][39:32] = buffer_data_5[279:272];
        layer1[33][47:40] = buffer_data_5[287:280];
        layer1[33][55:48] = buffer_data_5[295:288];
        layer2[33][7:0] = buffer_data_4[247:240];
        layer2[33][15:8] = buffer_data_4[255:248];
        layer2[33][23:16] = buffer_data_4[263:256];
        layer2[33][31:24] = buffer_data_4[271:264];
        layer2[33][39:32] = buffer_data_4[279:272];
        layer2[33][47:40] = buffer_data_4[287:280];
        layer2[33][55:48] = buffer_data_4[295:288];
        layer3[33][7:0] = buffer_data_3[247:240];
        layer3[33][15:8] = buffer_data_3[255:248];
        layer3[33][23:16] = buffer_data_3[263:256];
        layer3[33][31:24] = buffer_data_3[271:264];
        layer3[33][39:32] = buffer_data_3[279:272];
        layer3[33][47:40] = buffer_data_3[287:280];
        layer3[33][55:48] = buffer_data_3[295:288];
        layer4[33][7:0] = buffer_data_2[247:240];
        layer4[33][15:8] = buffer_data_2[255:248];
        layer4[33][23:16] = buffer_data_2[263:256];
        layer4[33][31:24] = buffer_data_2[271:264];
        layer4[33][39:32] = buffer_data_2[279:272];
        layer4[33][47:40] = buffer_data_2[287:280];
        layer4[33][55:48] = buffer_data_2[295:288];
        layer5[33][7:0] = buffer_data_1[247:240];
        layer5[33][15:8] = buffer_data_1[255:248];
        layer5[33][23:16] = buffer_data_1[263:256];
        layer5[33][31:24] = buffer_data_1[271:264];
        layer5[33][39:32] = buffer_data_1[279:272];
        layer5[33][47:40] = buffer_data_1[287:280];
        layer5[33][55:48] = buffer_data_1[295:288];
        layer6[33][7:0] = buffer_data_0[247:240];
        layer6[33][15:8] = buffer_data_0[255:248];
        layer6[33][23:16] = buffer_data_0[263:256];
        layer6[33][31:24] = buffer_data_0[271:264];
        layer6[33][39:32] = buffer_data_0[279:272];
        layer6[33][47:40] = buffer_data_0[287:280];
        layer6[33][55:48] = buffer_data_0[295:288];
        layer0[34][7:0] = buffer_data_6[255:248];
        layer0[34][15:8] = buffer_data_6[263:256];
        layer0[34][23:16] = buffer_data_6[271:264];
        layer0[34][31:24] = buffer_data_6[279:272];
        layer0[34][39:32] = buffer_data_6[287:280];
        layer0[34][47:40] = buffer_data_6[295:288];
        layer0[34][55:48] = buffer_data_6[303:296];
        layer1[34][7:0] = buffer_data_5[255:248];
        layer1[34][15:8] = buffer_data_5[263:256];
        layer1[34][23:16] = buffer_data_5[271:264];
        layer1[34][31:24] = buffer_data_5[279:272];
        layer1[34][39:32] = buffer_data_5[287:280];
        layer1[34][47:40] = buffer_data_5[295:288];
        layer1[34][55:48] = buffer_data_5[303:296];
        layer2[34][7:0] = buffer_data_4[255:248];
        layer2[34][15:8] = buffer_data_4[263:256];
        layer2[34][23:16] = buffer_data_4[271:264];
        layer2[34][31:24] = buffer_data_4[279:272];
        layer2[34][39:32] = buffer_data_4[287:280];
        layer2[34][47:40] = buffer_data_4[295:288];
        layer2[34][55:48] = buffer_data_4[303:296];
        layer3[34][7:0] = buffer_data_3[255:248];
        layer3[34][15:8] = buffer_data_3[263:256];
        layer3[34][23:16] = buffer_data_3[271:264];
        layer3[34][31:24] = buffer_data_3[279:272];
        layer3[34][39:32] = buffer_data_3[287:280];
        layer3[34][47:40] = buffer_data_3[295:288];
        layer3[34][55:48] = buffer_data_3[303:296];
        layer4[34][7:0] = buffer_data_2[255:248];
        layer4[34][15:8] = buffer_data_2[263:256];
        layer4[34][23:16] = buffer_data_2[271:264];
        layer4[34][31:24] = buffer_data_2[279:272];
        layer4[34][39:32] = buffer_data_2[287:280];
        layer4[34][47:40] = buffer_data_2[295:288];
        layer4[34][55:48] = buffer_data_2[303:296];
        layer5[34][7:0] = buffer_data_1[255:248];
        layer5[34][15:8] = buffer_data_1[263:256];
        layer5[34][23:16] = buffer_data_1[271:264];
        layer5[34][31:24] = buffer_data_1[279:272];
        layer5[34][39:32] = buffer_data_1[287:280];
        layer5[34][47:40] = buffer_data_1[295:288];
        layer5[34][55:48] = buffer_data_1[303:296];
        layer6[34][7:0] = buffer_data_0[255:248];
        layer6[34][15:8] = buffer_data_0[263:256];
        layer6[34][23:16] = buffer_data_0[271:264];
        layer6[34][31:24] = buffer_data_0[279:272];
        layer6[34][39:32] = buffer_data_0[287:280];
        layer6[34][47:40] = buffer_data_0[295:288];
        layer6[34][55:48] = buffer_data_0[303:296];
        layer0[35][7:0] = buffer_data_6[263:256];
        layer0[35][15:8] = buffer_data_6[271:264];
        layer0[35][23:16] = buffer_data_6[279:272];
        layer0[35][31:24] = buffer_data_6[287:280];
        layer0[35][39:32] = buffer_data_6[295:288];
        layer0[35][47:40] = buffer_data_6[303:296];
        layer0[35][55:48] = buffer_data_6[311:304];
        layer1[35][7:0] = buffer_data_5[263:256];
        layer1[35][15:8] = buffer_data_5[271:264];
        layer1[35][23:16] = buffer_data_5[279:272];
        layer1[35][31:24] = buffer_data_5[287:280];
        layer1[35][39:32] = buffer_data_5[295:288];
        layer1[35][47:40] = buffer_data_5[303:296];
        layer1[35][55:48] = buffer_data_5[311:304];
        layer2[35][7:0] = buffer_data_4[263:256];
        layer2[35][15:8] = buffer_data_4[271:264];
        layer2[35][23:16] = buffer_data_4[279:272];
        layer2[35][31:24] = buffer_data_4[287:280];
        layer2[35][39:32] = buffer_data_4[295:288];
        layer2[35][47:40] = buffer_data_4[303:296];
        layer2[35][55:48] = buffer_data_4[311:304];
        layer3[35][7:0] = buffer_data_3[263:256];
        layer3[35][15:8] = buffer_data_3[271:264];
        layer3[35][23:16] = buffer_data_3[279:272];
        layer3[35][31:24] = buffer_data_3[287:280];
        layer3[35][39:32] = buffer_data_3[295:288];
        layer3[35][47:40] = buffer_data_3[303:296];
        layer3[35][55:48] = buffer_data_3[311:304];
        layer4[35][7:0] = buffer_data_2[263:256];
        layer4[35][15:8] = buffer_data_2[271:264];
        layer4[35][23:16] = buffer_data_2[279:272];
        layer4[35][31:24] = buffer_data_2[287:280];
        layer4[35][39:32] = buffer_data_2[295:288];
        layer4[35][47:40] = buffer_data_2[303:296];
        layer4[35][55:48] = buffer_data_2[311:304];
        layer5[35][7:0] = buffer_data_1[263:256];
        layer5[35][15:8] = buffer_data_1[271:264];
        layer5[35][23:16] = buffer_data_1[279:272];
        layer5[35][31:24] = buffer_data_1[287:280];
        layer5[35][39:32] = buffer_data_1[295:288];
        layer5[35][47:40] = buffer_data_1[303:296];
        layer5[35][55:48] = buffer_data_1[311:304];
        layer6[35][7:0] = buffer_data_0[263:256];
        layer6[35][15:8] = buffer_data_0[271:264];
        layer6[35][23:16] = buffer_data_0[279:272];
        layer6[35][31:24] = buffer_data_0[287:280];
        layer6[35][39:32] = buffer_data_0[295:288];
        layer6[35][47:40] = buffer_data_0[303:296];
        layer6[35][55:48] = buffer_data_0[311:304];
        layer0[36][7:0] = buffer_data_6[271:264];
        layer0[36][15:8] = buffer_data_6[279:272];
        layer0[36][23:16] = buffer_data_6[287:280];
        layer0[36][31:24] = buffer_data_6[295:288];
        layer0[36][39:32] = buffer_data_6[303:296];
        layer0[36][47:40] = buffer_data_6[311:304];
        layer0[36][55:48] = buffer_data_6[319:312];
        layer1[36][7:0] = buffer_data_5[271:264];
        layer1[36][15:8] = buffer_data_5[279:272];
        layer1[36][23:16] = buffer_data_5[287:280];
        layer1[36][31:24] = buffer_data_5[295:288];
        layer1[36][39:32] = buffer_data_5[303:296];
        layer1[36][47:40] = buffer_data_5[311:304];
        layer1[36][55:48] = buffer_data_5[319:312];
        layer2[36][7:0] = buffer_data_4[271:264];
        layer2[36][15:8] = buffer_data_4[279:272];
        layer2[36][23:16] = buffer_data_4[287:280];
        layer2[36][31:24] = buffer_data_4[295:288];
        layer2[36][39:32] = buffer_data_4[303:296];
        layer2[36][47:40] = buffer_data_4[311:304];
        layer2[36][55:48] = buffer_data_4[319:312];
        layer3[36][7:0] = buffer_data_3[271:264];
        layer3[36][15:8] = buffer_data_3[279:272];
        layer3[36][23:16] = buffer_data_3[287:280];
        layer3[36][31:24] = buffer_data_3[295:288];
        layer3[36][39:32] = buffer_data_3[303:296];
        layer3[36][47:40] = buffer_data_3[311:304];
        layer3[36][55:48] = buffer_data_3[319:312];
        layer4[36][7:0] = buffer_data_2[271:264];
        layer4[36][15:8] = buffer_data_2[279:272];
        layer4[36][23:16] = buffer_data_2[287:280];
        layer4[36][31:24] = buffer_data_2[295:288];
        layer4[36][39:32] = buffer_data_2[303:296];
        layer4[36][47:40] = buffer_data_2[311:304];
        layer4[36][55:48] = buffer_data_2[319:312];
        layer5[36][7:0] = buffer_data_1[271:264];
        layer5[36][15:8] = buffer_data_1[279:272];
        layer5[36][23:16] = buffer_data_1[287:280];
        layer5[36][31:24] = buffer_data_1[295:288];
        layer5[36][39:32] = buffer_data_1[303:296];
        layer5[36][47:40] = buffer_data_1[311:304];
        layer5[36][55:48] = buffer_data_1[319:312];
        layer6[36][7:0] = buffer_data_0[271:264];
        layer6[36][15:8] = buffer_data_0[279:272];
        layer6[36][23:16] = buffer_data_0[287:280];
        layer6[36][31:24] = buffer_data_0[295:288];
        layer6[36][39:32] = buffer_data_0[303:296];
        layer6[36][47:40] = buffer_data_0[311:304];
        layer6[36][55:48] = buffer_data_0[319:312];
        layer0[37][7:0] = buffer_data_6[279:272];
        layer0[37][15:8] = buffer_data_6[287:280];
        layer0[37][23:16] = buffer_data_6[295:288];
        layer0[37][31:24] = buffer_data_6[303:296];
        layer0[37][39:32] = buffer_data_6[311:304];
        layer0[37][47:40] = buffer_data_6[319:312];
        layer0[37][55:48] = buffer_data_6[327:320];
        layer1[37][7:0] = buffer_data_5[279:272];
        layer1[37][15:8] = buffer_data_5[287:280];
        layer1[37][23:16] = buffer_data_5[295:288];
        layer1[37][31:24] = buffer_data_5[303:296];
        layer1[37][39:32] = buffer_data_5[311:304];
        layer1[37][47:40] = buffer_data_5[319:312];
        layer1[37][55:48] = buffer_data_5[327:320];
        layer2[37][7:0] = buffer_data_4[279:272];
        layer2[37][15:8] = buffer_data_4[287:280];
        layer2[37][23:16] = buffer_data_4[295:288];
        layer2[37][31:24] = buffer_data_4[303:296];
        layer2[37][39:32] = buffer_data_4[311:304];
        layer2[37][47:40] = buffer_data_4[319:312];
        layer2[37][55:48] = buffer_data_4[327:320];
        layer3[37][7:0] = buffer_data_3[279:272];
        layer3[37][15:8] = buffer_data_3[287:280];
        layer3[37][23:16] = buffer_data_3[295:288];
        layer3[37][31:24] = buffer_data_3[303:296];
        layer3[37][39:32] = buffer_data_3[311:304];
        layer3[37][47:40] = buffer_data_3[319:312];
        layer3[37][55:48] = buffer_data_3[327:320];
        layer4[37][7:0] = buffer_data_2[279:272];
        layer4[37][15:8] = buffer_data_2[287:280];
        layer4[37][23:16] = buffer_data_2[295:288];
        layer4[37][31:24] = buffer_data_2[303:296];
        layer4[37][39:32] = buffer_data_2[311:304];
        layer4[37][47:40] = buffer_data_2[319:312];
        layer4[37][55:48] = buffer_data_2[327:320];
        layer5[37][7:0] = buffer_data_1[279:272];
        layer5[37][15:8] = buffer_data_1[287:280];
        layer5[37][23:16] = buffer_data_1[295:288];
        layer5[37][31:24] = buffer_data_1[303:296];
        layer5[37][39:32] = buffer_data_1[311:304];
        layer5[37][47:40] = buffer_data_1[319:312];
        layer5[37][55:48] = buffer_data_1[327:320];
        layer6[37][7:0] = buffer_data_0[279:272];
        layer6[37][15:8] = buffer_data_0[287:280];
        layer6[37][23:16] = buffer_data_0[295:288];
        layer6[37][31:24] = buffer_data_0[303:296];
        layer6[37][39:32] = buffer_data_0[311:304];
        layer6[37][47:40] = buffer_data_0[319:312];
        layer6[37][55:48] = buffer_data_0[327:320];
        layer0[38][7:0] = buffer_data_6[287:280];
        layer0[38][15:8] = buffer_data_6[295:288];
        layer0[38][23:16] = buffer_data_6[303:296];
        layer0[38][31:24] = buffer_data_6[311:304];
        layer0[38][39:32] = buffer_data_6[319:312];
        layer0[38][47:40] = buffer_data_6[327:320];
        layer0[38][55:48] = buffer_data_6[335:328];
        layer1[38][7:0] = buffer_data_5[287:280];
        layer1[38][15:8] = buffer_data_5[295:288];
        layer1[38][23:16] = buffer_data_5[303:296];
        layer1[38][31:24] = buffer_data_5[311:304];
        layer1[38][39:32] = buffer_data_5[319:312];
        layer1[38][47:40] = buffer_data_5[327:320];
        layer1[38][55:48] = buffer_data_5[335:328];
        layer2[38][7:0] = buffer_data_4[287:280];
        layer2[38][15:8] = buffer_data_4[295:288];
        layer2[38][23:16] = buffer_data_4[303:296];
        layer2[38][31:24] = buffer_data_4[311:304];
        layer2[38][39:32] = buffer_data_4[319:312];
        layer2[38][47:40] = buffer_data_4[327:320];
        layer2[38][55:48] = buffer_data_4[335:328];
        layer3[38][7:0] = buffer_data_3[287:280];
        layer3[38][15:8] = buffer_data_3[295:288];
        layer3[38][23:16] = buffer_data_3[303:296];
        layer3[38][31:24] = buffer_data_3[311:304];
        layer3[38][39:32] = buffer_data_3[319:312];
        layer3[38][47:40] = buffer_data_3[327:320];
        layer3[38][55:48] = buffer_data_3[335:328];
        layer4[38][7:0] = buffer_data_2[287:280];
        layer4[38][15:8] = buffer_data_2[295:288];
        layer4[38][23:16] = buffer_data_2[303:296];
        layer4[38][31:24] = buffer_data_2[311:304];
        layer4[38][39:32] = buffer_data_2[319:312];
        layer4[38][47:40] = buffer_data_2[327:320];
        layer4[38][55:48] = buffer_data_2[335:328];
        layer5[38][7:0] = buffer_data_1[287:280];
        layer5[38][15:8] = buffer_data_1[295:288];
        layer5[38][23:16] = buffer_data_1[303:296];
        layer5[38][31:24] = buffer_data_1[311:304];
        layer5[38][39:32] = buffer_data_1[319:312];
        layer5[38][47:40] = buffer_data_1[327:320];
        layer5[38][55:48] = buffer_data_1[335:328];
        layer6[38][7:0] = buffer_data_0[287:280];
        layer6[38][15:8] = buffer_data_0[295:288];
        layer6[38][23:16] = buffer_data_0[303:296];
        layer6[38][31:24] = buffer_data_0[311:304];
        layer6[38][39:32] = buffer_data_0[319:312];
        layer6[38][47:40] = buffer_data_0[327:320];
        layer6[38][55:48] = buffer_data_0[335:328];
        layer0[39][7:0] = buffer_data_6[295:288];
        layer0[39][15:8] = buffer_data_6[303:296];
        layer0[39][23:16] = buffer_data_6[311:304];
        layer0[39][31:24] = buffer_data_6[319:312];
        layer0[39][39:32] = buffer_data_6[327:320];
        layer0[39][47:40] = buffer_data_6[335:328];
        layer0[39][55:48] = buffer_data_6[343:336];
        layer1[39][7:0] = buffer_data_5[295:288];
        layer1[39][15:8] = buffer_data_5[303:296];
        layer1[39][23:16] = buffer_data_5[311:304];
        layer1[39][31:24] = buffer_data_5[319:312];
        layer1[39][39:32] = buffer_data_5[327:320];
        layer1[39][47:40] = buffer_data_5[335:328];
        layer1[39][55:48] = buffer_data_5[343:336];
        layer2[39][7:0] = buffer_data_4[295:288];
        layer2[39][15:8] = buffer_data_4[303:296];
        layer2[39][23:16] = buffer_data_4[311:304];
        layer2[39][31:24] = buffer_data_4[319:312];
        layer2[39][39:32] = buffer_data_4[327:320];
        layer2[39][47:40] = buffer_data_4[335:328];
        layer2[39][55:48] = buffer_data_4[343:336];
        layer3[39][7:0] = buffer_data_3[295:288];
        layer3[39][15:8] = buffer_data_3[303:296];
        layer3[39][23:16] = buffer_data_3[311:304];
        layer3[39][31:24] = buffer_data_3[319:312];
        layer3[39][39:32] = buffer_data_3[327:320];
        layer3[39][47:40] = buffer_data_3[335:328];
        layer3[39][55:48] = buffer_data_3[343:336];
        layer4[39][7:0] = buffer_data_2[295:288];
        layer4[39][15:8] = buffer_data_2[303:296];
        layer4[39][23:16] = buffer_data_2[311:304];
        layer4[39][31:24] = buffer_data_2[319:312];
        layer4[39][39:32] = buffer_data_2[327:320];
        layer4[39][47:40] = buffer_data_2[335:328];
        layer4[39][55:48] = buffer_data_2[343:336];
        layer5[39][7:0] = buffer_data_1[295:288];
        layer5[39][15:8] = buffer_data_1[303:296];
        layer5[39][23:16] = buffer_data_1[311:304];
        layer5[39][31:24] = buffer_data_1[319:312];
        layer5[39][39:32] = buffer_data_1[327:320];
        layer5[39][47:40] = buffer_data_1[335:328];
        layer5[39][55:48] = buffer_data_1[343:336];
        layer6[39][7:0] = buffer_data_0[295:288];
        layer6[39][15:8] = buffer_data_0[303:296];
        layer6[39][23:16] = buffer_data_0[311:304];
        layer6[39][31:24] = buffer_data_0[319:312];
        layer6[39][39:32] = buffer_data_0[327:320];
        layer6[39][47:40] = buffer_data_0[335:328];
        layer6[39][55:48] = buffer_data_0[343:336];
        layer0[40][7:0] = buffer_data_6[303:296];
        layer0[40][15:8] = buffer_data_6[311:304];
        layer0[40][23:16] = buffer_data_6[319:312];
        layer0[40][31:24] = buffer_data_6[327:320];
        layer0[40][39:32] = buffer_data_6[335:328];
        layer0[40][47:40] = buffer_data_6[343:336];
        layer0[40][55:48] = buffer_data_6[351:344];
        layer1[40][7:0] = buffer_data_5[303:296];
        layer1[40][15:8] = buffer_data_5[311:304];
        layer1[40][23:16] = buffer_data_5[319:312];
        layer1[40][31:24] = buffer_data_5[327:320];
        layer1[40][39:32] = buffer_data_5[335:328];
        layer1[40][47:40] = buffer_data_5[343:336];
        layer1[40][55:48] = buffer_data_5[351:344];
        layer2[40][7:0] = buffer_data_4[303:296];
        layer2[40][15:8] = buffer_data_4[311:304];
        layer2[40][23:16] = buffer_data_4[319:312];
        layer2[40][31:24] = buffer_data_4[327:320];
        layer2[40][39:32] = buffer_data_4[335:328];
        layer2[40][47:40] = buffer_data_4[343:336];
        layer2[40][55:48] = buffer_data_4[351:344];
        layer3[40][7:0] = buffer_data_3[303:296];
        layer3[40][15:8] = buffer_data_3[311:304];
        layer3[40][23:16] = buffer_data_3[319:312];
        layer3[40][31:24] = buffer_data_3[327:320];
        layer3[40][39:32] = buffer_data_3[335:328];
        layer3[40][47:40] = buffer_data_3[343:336];
        layer3[40][55:48] = buffer_data_3[351:344];
        layer4[40][7:0] = buffer_data_2[303:296];
        layer4[40][15:8] = buffer_data_2[311:304];
        layer4[40][23:16] = buffer_data_2[319:312];
        layer4[40][31:24] = buffer_data_2[327:320];
        layer4[40][39:32] = buffer_data_2[335:328];
        layer4[40][47:40] = buffer_data_2[343:336];
        layer4[40][55:48] = buffer_data_2[351:344];
        layer5[40][7:0] = buffer_data_1[303:296];
        layer5[40][15:8] = buffer_data_1[311:304];
        layer5[40][23:16] = buffer_data_1[319:312];
        layer5[40][31:24] = buffer_data_1[327:320];
        layer5[40][39:32] = buffer_data_1[335:328];
        layer5[40][47:40] = buffer_data_1[343:336];
        layer5[40][55:48] = buffer_data_1[351:344];
        layer6[40][7:0] = buffer_data_0[303:296];
        layer6[40][15:8] = buffer_data_0[311:304];
        layer6[40][23:16] = buffer_data_0[319:312];
        layer6[40][31:24] = buffer_data_0[327:320];
        layer6[40][39:32] = buffer_data_0[335:328];
        layer6[40][47:40] = buffer_data_0[343:336];
        layer6[40][55:48] = buffer_data_0[351:344];
        layer0[41][7:0] = buffer_data_6[311:304];
        layer0[41][15:8] = buffer_data_6[319:312];
        layer0[41][23:16] = buffer_data_6[327:320];
        layer0[41][31:24] = buffer_data_6[335:328];
        layer0[41][39:32] = buffer_data_6[343:336];
        layer0[41][47:40] = buffer_data_6[351:344];
        layer0[41][55:48] = buffer_data_6[359:352];
        layer1[41][7:0] = buffer_data_5[311:304];
        layer1[41][15:8] = buffer_data_5[319:312];
        layer1[41][23:16] = buffer_data_5[327:320];
        layer1[41][31:24] = buffer_data_5[335:328];
        layer1[41][39:32] = buffer_data_5[343:336];
        layer1[41][47:40] = buffer_data_5[351:344];
        layer1[41][55:48] = buffer_data_5[359:352];
        layer2[41][7:0] = buffer_data_4[311:304];
        layer2[41][15:8] = buffer_data_4[319:312];
        layer2[41][23:16] = buffer_data_4[327:320];
        layer2[41][31:24] = buffer_data_4[335:328];
        layer2[41][39:32] = buffer_data_4[343:336];
        layer2[41][47:40] = buffer_data_4[351:344];
        layer2[41][55:48] = buffer_data_4[359:352];
        layer3[41][7:0] = buffer_data_3[311:304];
        layer3[41][15:8] = buffer_data_3[319:312];
        layer3[41][23:16] = buffer_data_3[327:320];
        layer3[41][31:24] = buffer_data_3[335:328];
        layer3[41][39:32] = buffer_data_3[343:336];
        layer3[41][47:40] = buffer_data_3[351:344];
        layer3[41][55:48] = buffer_data_3[359:352];
        layer4[41][7:0] = buffer_data_2[311:304];
        layer4[41][15:8] = buffer_data_2[319:312];
        layer4[41][23:16] = buffer_data_2[327:320];
        layer4[41][31:24] = buffer_data_2[335:328];
        layer4[41][39:32] = buffer_data_2[343:336];
        layer4[41][47:40] = buffer_data_2[351:344];
        layer4[41][55:48] = buffer_data_2[359:352];
        layer5[41][7:0] = buffer_data_1[311:304];
        layer5[41][15:8] = buffer_data_1[319:312];
        layer5[41][23:16] = buffer_data_1[327:320];
        layer5[41][31:24] = buffer_data_1[335:328];
        layer5[41][39:32] = buffer_data_1[343:336];
        layer5[41][47:40] = buffer_data_1[351:344];
        layer5[41][55:48] = buffer_data_1[359:352];
        layer6[41][7:0] = buffer_data_0[311:304];
        layer6[41][15:8] = buffer_data_0[319:312];
        layer6[41][23:16] = buffer_data_0[327:320];
        layer6[41][31:24] = buffer_data_0[335:328];
        layer6[41][39:32] = buffer_data_0[343:336];
        layer6[41][47:40] = buffer_data_0[351:344];
        layer6[41][55:48] = buffer_data_0[359:352];
        layer0[42][7:0] = buffer_data_6[319:312];
        layer0[42][15:8] = buffer_data_6[327:320];
        layer0[42][23:16] = buffer_data_6[335:328];
        layer0[42][31:24] = buffer_data_6[343:336];
        layer0[42][39:32] = buffer_data_6[351:344];
        layer0[42][47:40] = buffer_data_6[359:352];
        layer0[42][55:48] = buffer_data_6[367:360];
        layer1[42][7:0] = buffer_data_5[319:312];
        layer1[42][15:8] = buffer_data_5[327:320];
        layer1[42][23:16] = buffer_data_5[335:328];
        layer1[42][31:24] = buffer_data_5[343:336];
        layer1[42][39:32] = buffer_data_5[351:344];
        layer1[42][47:40] = buffer_data_5[359:352];
        layer1[42][55:48] = buffer_data_5[367:360];
        layer2[42][7:0] = buffer_data_4[319:312];
        layer2[42][15:8] = buffer_data_4[327:320];
        layer2[42][23:16] = buffer_data_4[335:328];
        layer2[42][31:24] = buffer_data_4[343:336];
        layer2[42][39:32] = buffer_data_4[351:344];
        layer2[42][47:40] = buffer_data_4[359:352];
        layer2[42][55:48] = buffer_data_4[367:360];
        layer3[42][7:0] = buffer_data_3[319:312];
        layer3[42][15:8] = buffer_data_3[327:320];
        layer3[42][23:16] = buffer_data_3[335:328];
        layer3[42][31:24] = buffer_data_3[343:336];
        layer3[42][39:32] = buffer_data_3[351:344];
        layer3[42][47:40] = buffer_data_3[359:352];
        layer3[42][55:48] = buffer_data_3[367:360];
        layer4[42][7:0] = buffer_data_2[319:312];
        layer4[42][15:8] = buffer_data_2[327:320];
        layer4[42][23:16] = buffer_data_2[335:328];
        layer4[42][31:24] = buffer_data_2[343:336];
        layer4[42][39:32] = buffer_data_2[351:344];
        layer4[42][47:40] = buffer_data_2[359:352];
        layer4[42][55:48] = buffer_data_2[367:360];
        layer5[42][7:0] = buffer_data_1[319:312];
        layer5[42][15:8] = buffer_data_1[327:320];
        layer5[42][23:16] = buffer_data_1[335:328];
        layer5[42][31:24] = buffer_data_1[343:336];
        layer5[42][39:32] = buffer_data_1[351:344];
        layer5[42][47:40] = buffer_data_1[359:352];
        layer5[42][55:48] = buffer_data_1[367:360];
        layer6[42][7:0] = buffer_data_0[319:312];
        layer6[42][15:8] = buffer_data_0[327:320];
        layer6[42][23:16] = buffer_data_0[335:328];
        layer6[42][31:24] = buffer_data_0[343:336];
        layer6[42][39:32] = buffer_data_0[351:344];
        layer6[42][47:40] = buffer_data_0[359:352];
        layer6[42][55:48] = buffer_data_0[367:360];
        layer0[43][7:0] = buffer_data_6[327:320];
        layer0[43][15:8] = buffer_data_6[335:328];
        layer0[43][23:16] = buffer_data_6[343:336];
        layer0[43][31:24] = buffer_data_6[351:344];
        layer0[43][39:32] = buffer_data_6[359:352];
        layer0[43][47:40] = buffer_data_6[367:360];
        layer0[43][55:48] = buffer_data_6[375:368];
        layer1[43][7:0] = buffer_data_5[327:320];
        layer1[43][15:8] = buffer_data_5[335:328];
        layer1[43][23:16] = buffer_data_5[343:336];
        layer1[43][31:24] = buffer_data_5[351:344];
        layer1[43][39:32] = buffer_data_5[359:352];
        layer1[43][47:40] = buffer_data_5[367:360];
        layer1[43][55:48] = buffer_data_5[375:368];
        layer2[43][7:0] = buffer_data_4[327:320];
        layer2[43][15:8] = buffer_data_4[335:328];
        layer2[43][23:16] = buffer_data_4[343:336];
        layer2[43][31:24] = buffer_data_4[351:344];
        layer2[43][39:32] = buffer_data_4[359:352];
        layer2[43][47:40] = buffer_data_4[367:360];
        layer2[43][55:48] = buffer_data_4[375:368];
        layer3[43][7:0] = buffer_data_3[327:320];
        layer3[43][15:8] = buffer_data_3[335:328];
        layer3[43][23:16] = buffer_data_3[343:336];
        layer3[43][31:24] = buffer_data_3[351:344];
        layer3[43][39:32] = buffer_data_3[359:352];
        layer3[43][47:40] = buffer_data_3[367:360];
        layer3[43][55:48] = buffer_data_3[375:368];
        layer4[43][7:0] = buffer_data_2[327:320];
        layer4[43][15:8] = buffer_data_2[335:328];
        layer4[43][23:16] = buffer_data_2[343:336];
        layer4[43][31:24] = buffer_data_2[351:344];
        layer4[43][39:32] = buffer_data_2[359:352];
        layer4[43][47:40] = buffer_data_2[367:360];
        layer4[43][55:48] = buffer_data_2[375:368];
        layer5[43][7:0] = buffer_data_1[327:320];
        layer5[43][15:8] = buffer_data_1[335:328];
        layer5[43][23:16] = buffer_data_1[343:336];
        layer5[43][31:24] = buffer_data_1[351:344];
        layer5[43][39:32] = buffer_data_1[359:352];
        layer5[43][47:40] = buffer_data_1[367:360];
        layer5[43][55:48] = buffer_data_1[375:368];
        layer6[43][7:0] = buffer_data_0[327:320];
        layer6[43][15:8] = buffer_data_0[335:328];
        layer6[43][23:16] = buffer_data_0[343:336];
        layer6[43][31:24] = buffer_data_0[351:344];
        layer6[43][39:32] = buffer_data_0[359:352];
        layer6[43][47:40] = buffer_data_0[367:360];
        layer6[43][55:48] = buffer_data_0[375:368];
        layer0[44][7:0] = buffer_data_6[335:328];
        layer0[44][15:8] = buffer_data_6[343:336];
        layer0[44][23:16] = buffer_data_6[351:344];
        layer0[44][31:24] = buffer_data_6[359:352];
        layer0[44][39:32] = buffer_data_6[367:360];
        layer0[44][47:40] = buffer_data_6[375:368];
        layer0[44][55:48] = buffer_data_6[383:376];
        layer1[44][7:0] = buffer_data_5[335:328];
        layer1[44][15:8] = buffer_data_5[343:336];
        layer1[44][23:16] = buffer_data_5[351:344];
        layer1[44][31:24] = buffer_data_5[359:352];
        layer1[44][39:32] = buffer_data_5[367:360];
        layer1[44][47:40] = buffer_data_5[375:368];
        layer1[44][55:48] = buffer_data_5[383:376];
        layer2[44][7:0] = buffer_data_4[335:328];
        layer2[44][15:8] = buffer_data_4[343:336];
        layer2[44][23:16] = buffer_data_4[351:344];
        layer2[44][31:24] = buffer_data_4[359:352];
        layer2[44][39:32] = buffer_data_4[367:360];
        layer2[44][47:40] = buffer_data_4[375:368];
        layer2[44][55:48] = buffer_data_4[383:376];
        layer3[44][7:0] = buffer_data_3[335:328];
        layer3[44][15:8] = buffer_data_3[343:336];
        layer3[44][23:16] = buffer_data_3[351:344];
        layer3[44][31:24] = buffer_data_3[359:352];
        layer3[44][39:32] = buffer_data_3[367:360];
        layer3[44][47:40] = buffer_data_3[375:368];
        layer3[44][55:48] = buffer_data_3[383:376];
        layer4[44][7:0] = buffer_data_2[335:328];
        layer4[44][15:8] = buffer_data_2[343:336];
        layer4[44][23:16] = buffer_data_2[351:344];
        layer4[44][31:24] = buffer_data_2[359:352];
        layer4[44][39:32] = buffer_data_2[367:360];
        layer4[44][47:40] = buffer_data_2[375:368];
        layer4[44][55:48] = buffer_data_2[383:376];
        layer5[44][7:0] = buffer_data_1[335:328];
        layer5[44][15:8] = buffer_data_1[343:336];
        layer5[44][23:16] = buffer_data_1[351:344];
        layer5[44][31:24] = buffer_data_1[359:352];
        layer5[44][39:32] = buffer_data_1[367:360];
        layer5[44][47:40] = buffer_data_1[375:368];
        layer5[44][55:48] = buffer_data_1[383:376];
        layer6[44][7:0] = buffer_data_0[335:328];
        layer6[44][15:8] = buffer_data_0[343:336];
        layer6[44][23:16] = buffer_data_0[351:344];
        layer6[44][31:24] = buffer_data_0[359:352];
        layer6[44][39:32] = buffer_data_0[367:360];
        layer6[44][47:40] = buffer_data_0[375:368];
        layer6[44][55:48] = buffer_data_0[383:376];
        layer0[45][7:0] = buffer_data_6[343:336];
        layer0[45][15:8] = buffer_data_6[351:344];
        layer0[45][23:16] = buffer_data_6[359:352];
        layer0[45][31:24] = buffer_data_6[367:360];
        layer0[45][39:32] = buffer_data_6[375:368];
        layer0[45][47:40] = buffer_data_6[383:376];
        layer0[45][55:48] = buffer_data_6[391:384];
        layer1[45][7:0] = buffer_data_5[343:336];
        layer1[45][15:8] = buffer_data_5[351:344];
        layer1[45][23:16] = buffer_data_5[359:352];
        layer1[45][31:24] = buffer_data_5[367:360];
        layer1[45][39:32] = buffer_data_5[375:368];
        layer1[45][47:40] = buffer_data_5[383:376];
        layer1[45][55:48] = buffer_data_5[391:384];
        layer2[45][7:0] = buffer_data_4[343:336];
        layer2[45][15:8] = buffer_data_4[351:344];
        layer2[45][23:16] = buffer_data_4[359:352];
        layer2[45][31:24] = buffer_data_4[367:360];
        layer2[45][39:32] = buffer_data_4[375:368];
        layer2[45][47:40] = buffer_data_4[383:376];
        layer2[45][55:48] = buffer_data_4[391:384];
        layer3[45][7:0] = buffer_data_3[343:336];
        layer3[45][15:8] = buffer_data_3[351:344];
        layer3[45][23:16] = buffer_data_3[359:352];
        layer3[45][31:24] = buffer_data_3[367:360];
        layer3[45][39:32] = buffer_data_3[375:368];
        layer3[45][47:40] = buffer_data_3[383:376];
        layer3[45][55:48] = buffer_data_3[391:384];
        layer4[45][7:0] = buffer_data_2[343:336];
        layer4[45][15:8] = buffer_data_2[351:344];
        layer4[45][23:16] = buffer_data_2[359:352];
        layer4[45][31:24] = buffer_data_2[367:360];
        layer4[45][39:32] = buffer_data_2[375:368];
        layer4[45][47:40] = buffer_data_2[383:376];
        layer4[45][55:48] = buffer_data_2[391:384];
        layer5[45][7:0] = buffer_data_1[343:336];
        layer5[45][15:8] = buffer_data_1[351:344];
        layer5[45][23:16] = buffer_data_1[359:352];
        layer5[45][31:24] = buffer_data_1[367:360];
        layer5[45][39:32] = buffer_data_1[375:368];
        layer5[45][47:40] = buffer_data_1[383:376];
        layer5[45][55:48] = buffer_data_1[391:384];
        layer6[45][7:0] = buffer_data_0[343:336];
        layer6[45][15:8] = buffer_data_0[351:344];
        layer6[45][23:16] = buffer_data_0[359:352];
        layer6[45][31:24] = buffer_data_0[367:360];
        layer6[45][39:32] = buffer_data_0[375:368];
        layer6[45][47:40] = buffer_data_0[383:376];
        layer6[45][55:48] = buffer_data_0[391:384];
        layer0[46][7:0] = buffer_data_6[351:344];
        layer0[46][15:8] = buffer_data_6[359:352];
        layer0[46][23:16] = buffer_data_6[367:360];
        layer0[46][31:24] = buffer_data_6[375:368];
        layer0[46][39:32] = buffer_data_6[383:376];
        layer0[46][47:40] = buffer_data_6[391:384];
        layer0[46][55:48] = buffer_data_6[399:392];
        layer1[46][7:0] = buffer_data_5[351:344];
        layer1[46][15:8] = buffer_data_5[359:352];
        layer1[46][23:16] = buffer_data_5[367:360];
        layer1[46][31:24] = buffer_data_5[375:368];
        layer1[46][39:32] = buffer_data_5[383:376];
        layer1[46][47:40] = buffer_data_5[391:384];
        layer1[46][55:48] = buffer_data_5[399:392];
        layer2[46][7:0] = buffer_data_4[351:344];
        layer2[46][15:8] = buffer_data_4[359:352];
        layer2[46][23:16] = buffer_data_4[367:360];
        layer2[46][31:24] = buffer_data_4[375:368];
        layer2[46][39:32] = buffer_data_4[383:376];
        layer2[46][47:40] = buffer_data_4[391:384];
        layer2[46][55:48] = buffer_data_4[399:392];
        layer3[46][7:0] = buffer_data_3[351:344];
        layer3[46][15:8] = buffer_data_3[359:352];
        layer3[46][23:16] = buffer_data_3[367:360];
        layer3[46][31:24] = buffer_data_3[375:368];
        layer3[46][39:32] = buffer_data_3[383:376];
        layer3[46][47:40] = buffer_data_3[391:384];
        layer3[46][55:48] = buffer_data_3[399:392];
        layer4[46][7:0] = buffer_data_2[351:344];
        layer4[46][15:8] = buffer_data_2[359:352];
        layer4[46][23:16] = buffer_data_2[367:360];
        layer4[46][31:24] = buffer_data_2[375:368];
        layer4[46][39:32] = buffer_data_2[383:376];
        layer4[46][47:40] = buffer_data_2[391:384];
        layer4[46][55:48] = buffer_data_2[399:392];
        layer5[46][7:0] = buffer_data_1[351:344];
        layer5[46][15:8] = buffer_data_1[359:352];
        layer5[46][23:16] = buffer_data_1[367:360];
        layer5[46][31:24] = buffer_data_1[375:368];
        layer5[46][39:32] = buffer_data_1[383:376];
        layer5[46][47:40] = buffer_data_1[391:384];
        layer5[46][55:48] = buffer_data_1[399:392];
        layer6[46][7:0] = buffer_data_0[351:344];
        layer6[46][15:8] = buffer_data_0[359:352];
        layer6[46][23:16] = buffer_data_0[367:360];
        layer6[46][31:24] = buffer_data_0[375:368];
        layer6[46][39:32] = buffer_data_0[383:376];
        layer6[46][47:40] = buffer_data_0[391:384];
        layer6[46][55:48] = buffer_data_0[399:392];
        layer0[47][7:0] = buffer_data_6[359:352];
        layer0[47][15:8] = buffer_data_6[367:360];
        layer0[47][23:16] = buffer_data_6[375:368];
        layer0[47][31:24] = buffer_data_6[383:376];
        layer0[47][39:32] = buffer_data_6[391:384];
        layer0[47][47:40] = buffer_data_6[399:392];
        layer0[47][55:48] = buffer_data_6[407:400];
        layer1[47][7:0] = buffer_data_5[359:352];
        layer1[47][15:8] = buffer_data_5[367:360];
        layer1[47][23:16] = buffer_data_5[375:368];
        layer1[47][31:24] = buffer_data_5[383:376];
        layer1[47][39:32] = buffer_data_5[391:384];
        layer1[47][47:40] = buffer_data_5[399:392];
        layer1[47][55:48] = buffer_data_5[407:400];
        layer2[47][7:0] = buffer_data_4[359:352];
        layer2[47][15:8] = buffer_data_4[367:360];
        layer2[47][23:16] = buffer_data_4[375:368];
        layer2[47][31:24] = buffer_data_4[383:376];
        layer2[47][39:32] = buffer_data_4[391:384];
        layer2[47][47:40] = buffer_data_4[399:392];
        layer2[47][55:48] = buffer_data_4[407:400];
        layer3[47][7:0] = buffer_data_3[359:352];
        layer3[47][15:8] = buffer_data_3[367:360];
        layer3[47][23:16] = buffer_data_3[375:368];
        layer3[47][31:24] = buffer_data_3[383:376];
        layer3[47][39:32] = buffer_data_3[391:384];
        layer3[47][47:40] = buffer_data_3[399:392];
        layer3[47][55:48] = buffer_data_3[407:400];
        layer4[47][7:0] = buffer_data_2[359:352];
        layer4[47][15:8] = buffer_data_2[367:360];
        layer4[47][23:16] = buffer_data_2[375:368];
        layer4[47][31:24] = buffer_data_2[383:376];
        layer4[47][39:32] = buffer_data_2[391:384];
        layer4[47][47:40] = buffer_data_2[399:392];
        layer4[47][55:48] = buffer_data_2[407:400];
        layer5[47][7:0] = buffer_data_1[359:352];
        layer5[47][15:8] = buffer_data_1[367:360];
        layer5[47][23:16] = buffer_data_1[375:368];
        layer5[47][31:24] = buffer_data_1[383:376];
        layer5[47][39:32] = buffer_data_1[391:384];
        layer5[47][47:40] = buffer_data_1[399:392];
        layer5[47][55:48] = buffer_data_1[407:400];
        layer6[47][7:0] = buffer_data_0[359:352];
        layer6[47][15:8] = buffer_data_0[367:360];
        layer6[47][23:16] = buffer_data_0[375:368];
        layer6[47][31:24] = buffer_data_0[383:376];
        layer6[47][39:32] = buffer_data_0[391:384];
        layer6[47][47:40] = buffer_data_0[399:392];
        layer6[47][55:48] = buffer_data_0[407:400];
        layer0[48][7:0] = buffer_data_6[367:360];
        layer0[48][15:8] = buffer_data_6[375:368];
        layer0[48][23:16] = buffer_data_6[383:376];
        layer0[48][31:24] = buffer_data_6[391:384];
        layer0[48][39:32] = buffer_data_6[399:392];
        layer0[48][47:40] = buffer_data_6[407:400];
        layer0[48][55:48] = buffer_data_6[415:408];
        layer1[48][7:0] = buffer_data_5[367:360];
        layer1[48][15:8] = buffer_data_5[375:368];
        layer1[48][23:16] = buffer_data_5[383:376];
        layer1[48][31:24] = buffer_data_5[391:384];
        layer1[48][39:32] = buffer_data_5[399:392];
        layer1[48][47:40] = buffer_data_5[407:400];
        layer1[48][55:48] = buffer_data_5[415:408];
        layer2[48][7:0] = buffer_data_4[367:360];
        layer2[48][15:8] = buffer_data_4[375:368];
        layer2[48][23:16] = buffer_data_4[383:376];
        layer2[48][31:24] = buffer_data_4[391:384];
        layer2[48][39:32] = buffer_data_4[399:392];
        layer2[48][47:40] = buffer_data_4[407:400];
        layer2[48][55:48] = buffer_data_4[415:408];
        layer3[48][7:0] = buffer_data_3[367:360];
        layer3[48][15:8] = buffer_data_3[375:368];
        layer3[48][23:16] = buffer_data_3[383:376];
        layer3[48][31:24] = buffer_data_3[391:384];
        layer3[48][39:32] = buffer_data_3[399:392];
        layer3[48][47:40] = buffer_data_3[407:400];
        layer3[48][55:48] = buffer_data_3[415:408];
        layer4[48][7:0] = buffer_data_2[367:360];
        layer4[48][15:8] = buffer_data_2[375:368];
        layer4[48][23:16] = buffer_data_2[383:376];
        layer4[48][31:24] = buffer_data_2[391:384];
        layer4[48][39:32] = buffer_data_2[399:392];
        layer4[48][47:40] = buffer_data_2[407:400];
        layer4[48][55:48] = buffer_data_2[415:408];
        layer5[48][7:0] = buffer_data_1[367:360];
        layer5[48][15:8] = buffer_data_1[375:368];
        layer5[48][23:16] = buffer_data_1[383:376];
        layer5[48][31:24] = buffer_data_1[391:384];
        layer5[48][39:32] = buffer_data_1[399:392];
        layer5[48][47:40] = buffer_data_1[407:400];
        layer5[48][55:48] = buffer_data_1[415:408];
        layer6[48][7:0] = buffer_data_0[367:360];
        layer6[48][15:8] = buffer_data_0[375:368];
        layer6[48][23:16] = buffer_data_0[383:376];
        layer6[48][31:24] = buffer_data_0[391:384];
        layer6[48][39:32] = buffer_data_0[399:392];
        layer6[48][47:40] = buffer_data_0[407:400];
        layer6[48][55:48] = buffer_data_0[415:408];
        layer0[49][7:0] = buffer_data_6[375:368];
        layer0[49][15:8] = buffer_data_6[383:376];
        layer0[49][23:16] = buffer_data_6[391:384];
        layer0[49][31:24] = buffer_data_6[399:392];
        layer0[49][39:32] = buffer_data_6[407:400];
        layer0[49][47:40] = buffer_data_6[415:408];
        layer0[49][55:48] = buffer_data_6[423:416];
        layer1[49][7:0] = buffer_data_5[375:368];
        layer1[49][15:8] = buffer_data_5[383:376];
        layer1[49][23:16] = buffer_data_5[391:384];
        layer1[49][31:24] = buffer_data_5[399:392];
        layer1[49][39:32] = buffer_data_5[407:400];
        layer1[49][47:40] = buffer_data_5[415:408];
        layer1[49][55:48] = buffer_data_5[423:416];
        layer2[49][7:0] = buffer_data_4[375:368];
        layer2[49][15:8] = buffer_data_4[383:376];
        layer2[49][23:16] = buffer_data_4[391:384];
        layer2[49][31:24] = buffer_data_4[399:392];
        layer2[49][39:32] = buffer_data_4[407:400];
        layer2[49][47:40] = buffer_data_4[415:408];
        layer2[49][55:48] = buffer_data_4[423:416];
        layer3[49][7:0] = buffer_data_3[375:368];
        layer3[49][15:8] = buffer_data_3[383:376];
        layer3[49][23:16] = buffer_data_3[391:384];
        layer3[49][31:24] = buffer_data_3[399:392];
        layer3[49][39:32] = buffer_data_3[407:400];
        layer3[49][47:40] = buffer_data_3[415:408];
        layer3[49][55:48] = buffer_data_3[423:416];
        layer4[49][7:0] = buffer_data_2[375:368];
        layer4[49][15:8] = buffer_data_2[383:376];
        layer4[49][23:16] = buffer_data_2[391:384];
        layer4[49][31:24] = buffer_data_2[399:392];
        layer4[49][39:32] = buffer_data_2[407:400];
        layer4[49][47:40] = buffer_data_2[415:408];
        layer4[49][55:48] = buffer_data_2[423:416];
        layer5[49][7:0] = buffer_data_1[375:368];
        layer5[49][15:8] = buffer_data_1[383:376];
        layer5[49][23:16] = buffer_data_1[391:384];
        layer5[49][31:24] = buffer_data_1[399:392];
        layer5[49][39:32] = buffer_data_1[407:400];
        layer5[49][47:40] = buffer_data_1[415:408];
        layer5[49][55:48] = buffer_data_1[423:416];
        layer6[49][7:0] = buffer_data_0[375:368];
        layer6[49][15:8] = buffer_data_0[383:376];
        layer6[49][23:16] = buffer_data_0[391:384];
        layer6[49][31:24] = buffer_data_0[399:392];
        layer6[49][39:32] = buffer_data_0[407:400];
        layer6[49][47:40] = buffer_data_0[415:408];
        layer6[49][55:48] = buffer_data_0[423:416];
        layer0[50][7:0] = buffer_data_6[383:376];
        layer0[50][15:8] = buffer_data_6[391:384];
        layer0[50][23:16] = buffer_data_6[399:392];
        layer0[50][31:24] = buffer_data_6[407:400];
        layer0[50][39:32] = buffer_data_6[415:408];
        layer0[50][47:40] = buffer_data_6[423:416];
        layer0[50][55:48] = buffer_data_6[431:424];
        layer1[50][7:0] = buffer_data_5[383:376];
        layer1[50][15:8] = buffer_data_5[391:384];
        layer1[50][23:16] = buffer_data_5[399:392];
        layer1[50][31:24] = buffer_data_5[407:400];
        layer1[50][39:32] = buffer_data_5[415:408];
        layer1[50][47:40] = buffer_data_5[423:416];
        layer1[50][55:48] = buffer_data_5[431:424];
        layer2[50][7:0] = buffer_data_4[383:376];
        layer2[50][15:8] = buffer_data_4[391:384];
        layer2[50][23:16] = buffer_data_4[399:392];
        layer2[50][31:24] = buffer_data_4[407:400];
        layer2[50][39:32] = buffer_data_4[415:408];
        layer2[50][47:40] = buffer_data_4[423:416];
        layer2[50][55:48] = buffer_data_4[431:424];
        layer3[50][7:0] = buffer_data_3[383:376];
        layer3[50][15:8] = buffer_data_3[391:384];
        layer3[50][23:16] = buffer_data_3[399:392];
        layer3[50][31:24] = buffer_data_3[407:400];
        layer3[50][39:32] = buffer_data_3[415:408];
        layer3[50][47:40] = buffer_data_3[423:416];
        layer3[50][55:48] = buffer_data_3[431:424];
        layer4[50][7:0] = buffer_data_2[383:376];
        layer4[50][15:8] = buffer_data_2[391:384];
        layer4[50][23:16] = buffer_data_2[399:392];
        layer4[50][31:24] = buffer_data_2[407:400];
        layer4[50][39:32] = buffer_data_2[415:408];
        layer4[50][47:40] = buffer_data_2[423:416];
        layer4[50][55:48] = buffer_data_2[431:424];
        layer5[50][7:0] = buffer_data_1[383:376];
        layer5[50][15:8] = buffer_data_1[391:384];
        layer5[50][23:16] = buffer_data_1[399:392];
        layer5[50][31:24] = buffer_data_1[407:400];
        layer5[50][39:32] = buffer_data_1[415:408];
        layer5[50][47:40] = buffer_data_1[423:416];
        layer5[50][55:48] = buffer_data_1[431:424];
        layer6[50][7:0] = buffer_data_0[383:376];
        layer6[50][15:8] = buffer_data_0[391:384];
        layer6[50][23:16] = buffer_data_0[399:392];
        layer6[50][31:24] = buffer_data_0[407:400];
        layer6[50][39:32] = buffer_data_0[415:408];
        layer6[50][47:40] = buffer_data_0[423:416];
        layer6[50][55:48] = buffer_data_0[431:424];
        layer0[51][7:0] = buffer_data_6[391:384];
        layer0[51][15:8] = buffer_data_6[399:392];
        layer0[51][23:16] = buffer_data_6[407:400];
        layer0[51][31:24] = buffer_data_6[415:408];
        layer0[51][39:32] = buffer_data_6[423:416];
        layer0[51][47:40] = buffer_data_6[431:424];
        layer0[51][55:48] = buffer_data_6[439:432];
        layer1[51][7:0] = buffer_data_5[391:384];
        layer1[51][15:8] = buffer_data_5[399:392];
        layer1[51][23:16] = buffer_data_5[407:400];
        layer1[51][31:24] = buffer_data_5[415:408];
        layer1[51][39:32] = buffer_data_5[423:416];
        layer1[51][47:40] = buffer_data_5[431:424];
        layer1[51][55:48] = buffer_data_5[439:432];
        layer2[51][7:0] = buffer_data_4[391:384];
        layer2[51][15:8] = buffer_data_4[399:392];
        layer2[51][23:16] = buffer_data_4[407:400];
        layer2[51][31:24] = buffer_data_4[415:408];
        layer2[51][39:32] = buffer_data_4[423:416];
        layer2[51][47:40] = buffer_data_4[431:424];
        layer2[51][55:48] = buffer_data_4[439:432];
        layer3[51][7:0] = buffer_data_3[391:384];
        layer3[51][15:8] = buffer_data_3[399:392];
        layer3[51][23:16] = buffer_data_3[407:400];
        layer3[51][31:24] = buffer_data_3[415:408];
        layer3[51][39:32] = buffer_data_3[423:416];
        layer3[51][47:40] = buffer_data_3[431:424];
        layer3[51][55:48] = buffer_data_3[439:432];
        layer4[51][7:0] = buffer_data_2[391:384];
        layer4[51][15:8] = buffer_data_2[399:392];
        layer4[51][23:16] = buffer_data_2[407:400];
        layer4[51][31:24] = buffer_data_2[415:408];
        layer4[51][39:32] = buffer_data_2[423:416];
        layer4[51][47:40] = buffer_data_2[431:424];
        layer4[51][55:48] = buffer_data_2[439:432];
        layer5[51][7:0] = buffer_data_1[391:384];
        layer5[51][15:8] = buffer_data_1[399:392];
        layer5[51][23:16] = buffer_data_1[407:400];
        layer5[51][31:24] = buffer_data_1[415:408];
        layer5[51][39:32] = buffer_data_1[423:416];
        layer5[51][47:40] = buffer_data_1[431:424];
        layer5[51][55:48] = buffer_data_1[439:432];
        layer6[51][7:0] = buffer_data_0[391:384];
        layer6[51][15:8] = buffer_data_0[399:392];
        layer6[51][23:16] = buffer_data_0[407:400];
        layer6[51][31:24] = buffer_data_0[415:408];
        layer6[51][39:32] = buffer_data_0[423:416];
        layer6[51][47:40] = buffer_data_0[431:424];
        layer6[51][55:48] = buffer_data_0[439:432];
        layer0[52][7:0] = buffer_data_6[399:392];
        layer0[52][15:8] = buffer_data_6[407:400];
        layer0[52][23:16] = buffer_data_6[415:408];
        layer0[52][31:24] = buffer_data_6[423:416];
        layer0[52][39:32] = buffer_data_6[431:424];
        layer0[52][47:40] = buffer_data_6[439:432];
        layer0[52][55:48] = buffer_data_6[447:440];
        layer1[52][7:0] = buffer_data_5[399:392];
        layer1[52][15:8] = buffer_data_5[407:400];
        layer1[52][23:16] = buffer_data_5[415:408];
        layer1[52][31:24] = buffer_data_5[423:416];
        layer1[52][39:32] = buffer_data_5[431:424];
        layer1[52][47:40] = buffer_data_5[439:432];
        layer1[52][55:48] = buffer_data_5[447:440];
        layer2[52][7:0] = buffer_data_4[399:392];
        layer2[52][15:8] = buffer_data_4[407:400];
        layer2[52][23:16] = buffer_data_4[415:408];
        layer2[52][31:24] = buffer_data_4[423:416];
        layer2[52][39:32] = buffer_data_4[431:424];
        layer2[52][47:40] = buffer_data_4[439:432];
        layer2[52][55:48] = buffer_data_4[447:440];
        layer3[52][7:0] = buffer_data_3[399:392];
        layer3[52][15:8] = buffer_data_3[407:400];
        layer3[52][23:16] = buffer_data_3[415:408];
        layer3[52][31:24] = buffer_data_3[423:416];
        layer3[52][39:32] = buffer_data_3[431:424];
        layer3[52][47:40] = buffer_data_3[439:432];
        layer3[52][55:48] = buffer_data_3[447:440];
        layer4[52][7:0] = buffer_data_2[399:392];
        layer4[52][15:8] = buffer_data_2[407:400];
        layer4[52][23:16] = buffer_data_2[415:408];
        layer4[52][31:24] = buffer_data_2[423:416];
        layer4[52][39:32] = buffer_data_2[431:424];
        layer4[52][47:40] = buffer_data_2[439:432];
        layer4[52][55:48] = buffer_data_2[447:440];
        layer5[52][7:0] = buffer_data_1[399:392];
        layer5[52][15:8] = buffer_data_1[407:400];
        layer5[52][23:16] = buffer_data_1[415:408];
        layer5[52][31:24] = buffer_data_1[423:416];
        layer5[52][39:32] = buffer_data_1[431:424];
        layer5[52][47:40] = buffer_data_1[439:432];
        layer5[52][55:48] = buffer_data_1[447:440];
        layer6[52][7:0] = buffer_data_0[399:392];
        layer6[52][15:8] = buffer_data_0[407:400];
        layer6[52][23:16] = buffer_data_0[415:408];
        layer6[52][31:24] = buffer_data_0[423:416];
        layer6[52][39:32] = buffer_data_0[431:424];
        layer6[52][47:40] = buffer_data_0[439:432];
        layer6[52][55:48] = buffer_data_0[447:440];
        layer0[53][7:0] = buffer_data_6[407:400];
        layer0[53][15:8] = buffer_data_6[415:408];
        layer0[53][23:16] = buffer_data_6[423:416];
        layer0[53][31:24] = buffer_data_6[431:424];
        layer0[53][39:32] = buffer_data_6[439:432];
        layer0[53][47:40] = buffer_data_6[447:440];
        layer0[53][55:48] = buffer_data_6[455:448];
        layer1[53][7:0] = buffer_data_5[407:400];
        layer1[53][15:8] = buffer_data_5[415:408];
        layer1[53][23:16] = buffer_data_5[423:416];
        layer1[53][31:24] = buffer_data_5[431:424];
        layer1[53][39:32] = buffer_data_5[439:432];
        layer1[53][47:40] = buffer_data_5[447:440];
        layer1[53][55:48] = buffer_data_5[455:448];
        layer2[53][7:0] = buffer_data_4[407:400];
        layer2[53][15:8] = buffer_data_4[415:408];
        layer2[53][23:16] = buffer_data_4[423:416];
        layer2[53][31:24] = buffer_data_4[431:424];
        layer2[53][39:32] = buffer_data_4[439:432];
        layer2[53][47:40] = buffer_data_4[447:440];
        layer2[53][55:48] = buffer_data_4[455:448];
        layer3[53][7:0] = buffer_data_3[407:400];
        layer3[53][15:8] = buffer_data_3[415:408];
        layer3[53][23:16] = buffer_data_3[423:416];
        layer3[53][31:24] = buffer_data_3[431:424];
        layer3[53][39:32] = buffer_data_3[439:432];
        layer3[53][47:40] = buffer_data_3[447:440];
        layer3[53][55:48] = buffer_data_3[455:448];
        layer4[53][7:0] = buffer_data_2[407:400];
        layer4[53][15:8] = buffer_data_2[415:408];
        layer4[53][23:16] = buffer_data_2[423:416];
        layer4[53][31:24] = buffer_data_2[431:424];
        layer4[53][39:32] = buffer_data_2[439:432];
        layer4[53][47:40] = buffer_data_2[447:440];
        layer4[53][55:48] = buffer_data_2[455:448];
        layer5[53][7:0] = buffer_data_1[407:400];
        layer5[53][15:8] = buffer_data_1[415:408];
        layer5[53][23:16] = buffer_data_1[423:416];
        layer5[53][31:24] = buffer_data_1[431:424];
        layer5[53][39:32] = buffer_data_1[439:432];
        layer5[53][47:40] = buffer_data_1[447:440];
        layer5[53][55:48] = buffer_data_1[455:448];
        layer6[53][7:0] = buffer_data_0[407:400];
        layer6[53][15:8] = buffer_data_0[415:408];
        layer6[53][23:16] = buffer_data_0[423:416];
        layer6[53][31:24] = buffer_data_0[431:424];
        layer6[53][39:32] = buffer_data_0[439:432];
        layer6[53][47:40] = buffer_data_0[447:440];
        layer6[53][55:48] = buffer_data_0[455:448];
        layer0[54][7:0] = buffer_data_6[415:408];
        layer0[54][15:8] = buffer_data_6[423:416];
        layer0[54][23:16] = buffer_data_6[431:424];
        layer0[54][31:24] = buffer_data_6[439:432];
        layer0[54][39:32] = buffer_data_6[447:440];
        layer0[54][47:40] = buffer_data_6[455:448];
        layer0[54][55:48] = buffer_data_6[463:456];
        layer1[54][7:0] = buffer_data_5[415:408];
        layer1[54][15:8] = buffer_data_5[423:416];
        layer1[54][23:16] = buffer_data_5[431:424];
        layer1[54][31:24] = buffer_data_5[439:432];
        layer1[54][39:32] = buffer_data_5[447:440];
        layer1[54][47:40] = buffer_data_5[455:448];
        layer1[54][55:48] = buffer_data_5[463:456];
        layer2[54][7:0] = buffer_data_4[415:408];
        layer2[54][15:8] = buffer_data_4[423:416];
        layer2[54][23:16] = buffer_data_4[431:424];
        layer2[54][31:24] = buffer_data_4[439:432];
        layer2[54][39:32] = buffer_data_4[447:440];
        layer2[54][47:40] = buffer_data_4[455:448];
        layer2[54][55:48] = buffer_data_4[463:456];
        layer3[54][7:0] = buffer_data_3[415:408];
        layer3[54][15:8] = buffer_data_3[423:416];
        layer3[54][23:16] = buffer_data_3[431:424];
        layer3[54][31:24] = buffer_data_3[439:432];
        layer3[54][39:32] = buffer_data_3[447:440];
        layer3[54][47:40] = buffer_data_3[455:448];
        layer3[54][55:48] = buffer_data_3[463:456];
        layer4[54][7:0] = buffer_data_2[415:408];
        layer4[54][15:8] = buffer_data_2[423:416];
        layer4[54][23:16] = buffer_data_2[431:424];
        layer4[54][31:24] = buffer_data_2[439:432];
        layer4[54][39:32] = buffer_data_2[447:440];
        layer4[54][47:40] = buffer_data_2[455:448];
        layer4[54][55:48] = buffer_data_2[463:456];
        layer5[54][7:0] = buffer_data_1[415:408];
        layer5[54][15:8] = buffer_data_1[423:416];
        layer5[54][23:16] = buffer_data_1[431:424];
        layer5[54][31:24] = buffer_data_1[439:432];
        layer5[54][39:32] = buffer_data_1[447:440];
        layer5[54][47:40] = buffer_data_1[455:448];
        layer5[54][55:48] = buffer_data_1[463:456];
        layer6[54][7:0] = buffer_data_0[415:408];
        layer6[54][15:8] = buffer_data_0[423:416];
        layer6[54][23:16] = buffer_data_0[431:424];
        layer6[54][31:24] = buffer_data_0[439:432];
        layer6[54][39:32] = buffer_data_0[447:440];
        layer6[54][47:40] = buffer_data_0[455:448];
        layer6[54][55:48] = buffer_data_0[463:456];
        layer0[55][7:0] = buffer_data_6[423:416];
        layer0[55][15:8] = buffer_data_6[431:424];
        layer0[55][23:16] = buffer_data_6[439:432];
        layer0[55][31:24] = buffer_data_6[447:440];
        layer0[55][39:32] = buffer_data_6[455:448];
        layer0[55][47:40] = buffer_data_6[463:456];
        layer0[55][55:48] = buffer_data_6[471:464];
        layer1[55][7:0] = buffer_data_5[423:416];
        layer1[55][15:8] = buffer_data_5[431:424];
        layer1[55][23:16] = buffer_data_5[439:432];
        layer1[55][31:24] = buffer_data_5[447:440];
        layer1[55][39:32] = buffer_data_5[455:448];
        layer1[55][47:40] = buffer_data_5[463:456];
        layer1[55][55:48] = buffer_data_5[471:464];
        layer2[55][7:0] = buffer_data_4[423:416];
        layer2[55][15:8] = buffer_data_4[431:424];
        layer2[55][23:16] = buffer_data_4[439:432];
        layer2[55][31:24] = buffer_data_4[447:440];
        layer2[55][39:32] = buffer_data_4[455:448];
        layer2[55][47:40] = buffer_data_4[463:456];
        layer2[55][55:48] = buffer_data_4[471:464];
        layer3[55][7:0] = buffer_data_3[423:416];
        layer3[55][15:8] = buffer_data_3[431:424];
        layer3[55][23:16] = buffer_data_3[439:432];
        layer3[55][31:24] = buffer_data_3[447:440];
        layer3[55][39:32] = buffer_data_3[455:448];
        layer3[55][47:40] = buffer_data_3[463:456];
        layer3[55][55:48] = buffer_data_3[471:464];
        layer4[55][7:0] = buffer_data_2[423:416];
        layer4[55][15:8] = buffer_data_2[431:424];
        layer4[55][23:16] = buffer_data_2[439:432];
        layer4[55][31:24] = buffer_data_2[447:440];
        layer4[55][39:32] = buffer_data_2[455:448];
        layer4[55][47:40] = buffer_data_2[463:456];
        layer4[55][55:48] = buffer_data_2[471:464];
        layer5[55][7:0] = buffer_data_1[423:416];
        layer5[55][15:8] = buffer_data_1[431:424];
        layer5[55][23:16] = buffer_data_1[439:432];
        layer5[55][31:24] = buffer_data_1[447:440];
        layer5[55][39:32] = buffer_data_1[455:448];
        layer5[55][47:40] = buffer_data_1[463:456];
        layer5[55][55:48] = buffer_data_1[471:464];
        layer6[55][7:0] = buffer_data_0[423:416];
        layer6[55][15:8] = buffer_data_0[431:424];
        layer6[55][23:16] = buffer_data_0[439:432];
        layer6[55][31:24] = buffer_data_0[447:440];
        layer6[55][39:32] = buffer_data_0[455:448];
        layer6[55][47:40] = buffer_data_0[463:456];
        layer6[55][55:48] = buffer_data_0[471:464];
        layer0[56][7:0] = buffer_data_6[431:424];
        layer0[56][15:8] = buffer_data_6[439:432];
        layer0[56][23:16] = buffer_data_6[447:440];
        layer0[56][31:24] = buffer_data_6[455:448];
        layer0[56][39:32] = buffer_data_6[463:456];
        layer0[56][47:40] = buffer_data_6[471:464];
        layer0[56][55:48] = buffer_data_6[479:472];
        layer1[56][7:0] = buffer_data_5[431:424];
        layer1[56][15:8] = buffer_data_5[439:432];
        layer1[56][23:16] = buffer_data_5[447:440];
        layer1[56][31:24] = buffer_data_5[455:448];
        layer1[56][39:32] = buffer_data_5[463:456];
        layer1[56][47:40] = buffer_data_5[471:464];
        layer1[56][55:48] = buffer_data_5[479:472];
        layer2[56][7:0] = buffer_data_4[431:424];
        layer2[56][15:8] = buffer_data_4[439:432];
        layer2[56][23:16] = buffer_data_4[447:440];
        layer2[56][31:24] = buffer_data_4[455:448];
        layer2[56][39:32] = buffer_data_4[463:456];
        layer2[56][47:40] = buffer_data_4[471:464];
        layer2[56][55:48] = buffer_data_4[479:472];
        layer3[56][7:0] = buffer_data_3[431:424];
        layer3[56][15:8] = buffer_data_3[439:432];
        layer3[56][23:16] = buffer_data_3[447:440];
        layer3[56][31:24] = buffer_data_3[455:448];
        layer3[56][39:32] = buffer_data_3[463:456];
        layer3[56][47:40] = buffer_data_3[471:464];
        layer3[56][55:48] = buffer_data_3[479:472];
        layer4[56][7:0] = buffer_data_2[431:424];
        layer4[56][15:8] = buffer_data_2[439:432];
        layer4[56][23:16] = buffer_data_2[447:440];
        layer4[56][31:24] = buffer_data_2[455:448];
        layer4[56][39:32] = buffer_data_2[463:456];
        layer4[56][47:40] = buffer_data_2[471:464];
        layer4[56][55:48] = buffer_data_2[479:472];
        layer5[56][7:0] = buffer_data_1[431:424];
        layer5[56][15:8] = buffer_data_1[439:432];
        layer5[56][23:16] = buffer_data_1[447:440];
        layer5[56][31:24] = buffer_data_1[455:448];
        layer5[56][39:32] = buffer_data_1[463:456];
        layer5[56][47:40] = buffer_data_1[471:464];
        layer5[56][55:48] = buffer_data_1[479:472];
        layer6[56][7:0] = buffer_data_0[431:424];
        layer6[56][15:8] = buffer_data_0[439:432];
        layer6[56][23:16] = buffer_data_0[447:440];
        layer6[56][31:24] = buffer_data_0[455:448];
        layer6[56][39:32] = buffer_data_0[463:456];
        layer6[56][47:40] = buffer_data_0[471:464];
        layer6[56][55:48] = buffer_data_0[479:472];
        layer0[57][7:0] = buffer_data_6[439:432];
        layer0[57][15:8] = buffer_data_6[447:440];
        layer0[57][23:16] = buffer_data_6[455:448];
        layer0[57][31:24] = buffer_data_6[463:456];
        layer0[57][39:32] = buffer_data_6[471:464];
        layer0[57][47:40] = buffer_data_6[479:472];
        layer0[57][55:48] = buffer_data_6[487:480];
        layer1[57][7:0] = buffer_data_5[439:432];
        layer1[57][15:8] = buffer_data_5[447:440];
        layer1[57][23:16] = buffer_data_5[455:448];
        layer1[57][31:24] = buffer_data_5[463:456];
        layer1[57][39:32] = buffer_data_5[471:464];
        layer1[57][47:40] = buffer_data_5[479:472];
        layer1[57][55:48] = buffer_data_5[487:480];
        layer2[57][7:0] = buffer_data_4[439:432];
        layer2[57][15:8] = buffer_data_4[447:440];
        layer2[57][23:16] = buffer_data_4[455:448];
        layer2[57][31:24] = buffer_data_4[463:456];
        layer2[57][39:32] = buffer_data_4[471:464];
        layer2[57][47:40] = buffer_data_4[479:472];
        layer2[57][55:48] = buffer_data_4[487:480];
        layer3[57][7:0] = buffer_data_3[439:432];
        layer3[57][15:8] = buffer_data_3[447:440];
        layer3[57][23:16] = buffer_data_3[455:448];
        layer3[57][31:24] = buffer_data_3[463:456];
        layer3[57][39:32] = buffer_data_3[471:464];
        layer3[57][47:40] = buffer_data_3[479:472];
        layer3[57][55:48] = buffer_data_3[487:480];
        layer4[57][7:0] = buffer_data_2[439:432];
        layer4[57][15:8] = buffer_data_2[447:440];
        layer4[57][23:16] = buffer_data_2[455:448];
        layer4[57][31:24] = buffer_data_2[463:456];
        layer4[57][39:32] = buffer_data_2[471:464];
        layer4[57][47:40] = buffer_data_2[479:472];
        layer4[57][55:48] = buffer_data_2[487:480];
        layer5[57][7:0] = buffer_data_1[439:432];
        layer5[57][15:8] = buffer_data_1[447:440];
        layer5[57][23:16] = buffer_data_1[455:448];
        layer5[57][31:24] = buffer_data_1[463:456];
        layer5[57][39:32] = buffer_data_1[471:464];
        layer5[57][47:40] = buffer_data_1[479:472];
        layer5[57][55:48] = buffer_data_1[487:480];
        layer6[57][7:0] = buffer_data_0[439:432];
        layer6[57][15:8] = buffer_data_0[447:440];
        layer6[57][23:16] = buffer_data_0[455:448];
        layer6[57][31:24] = buffer_data_0[463:456];
        layer6[57][39:32] = buffer_data_0[471:464];
        layer6[57][47:40] = buffer_data_0[479:472];
        layer6[57][55:48] = buffer_data_0[487:480];
        layer0[58][7:0] = buffer_data_6[447:440];
        layer0[58][15:8] = buffer_data_6[455:448];
        layer0[58][23:16] = buffer_data_6[463:456];
        layer0[58][31:24] = buffer_data_6[471:464];
        layer0[58][39:32] = buffer_data_6[479:472];
        layer0[58][47:40] = buffer_data_6[487:480];
        layer0[58][55:48] = buffer_data_6[495:488];
        layer1[58][7:0] = buffer_data_5[447:440];
        layer1[58][15:8] = buffer_data_5[455:448];
        layer1[58][23:16] = buffer_data_5[463:456];
        layer1[58][31:24] = buffer_data_5[471:464];
        layer1[58][39:32] = buffer_data_5[479:472];
        layer1[58][47:40] = buffer_data_5[487:480];
        layer1[58][55:48] = buffer_data_5[495:488];
        layer2[58][7:0] = buffer_data_4[447:440];
        layer2[58][15:8] = buffer_data_4[455:448];
        layer2[58][23:16] = buffer_data_4[463:456];
        layer2[58][31:24] = buffer_data_4[471:464];
        layer2[58][39:32] = buffer_data_4[479:472];
        layer2[58][47:40] = buffer_data_4[487:480];
        layer2[58][55:48] = buffer_data_4[495:488];
        layer3[58][7:0] = buffer_data_3[447:440];
        layer3[58][15:8] = buffer_data_3[455:448];
        layer3[58][23:16] = buffer_data_3[463:456];
        layer3[58][31:24] = buffer_data_3[471:464];
        layer3[58][39:32] = buffer_data_3[479:472];
        layer3[58][47:40] = buffer_data_3[487:480];
        layer3[58][55:48] = buffer_data_3[495:488];
        layer4[58][7:0] = buffer_data_2[447:440];
        layer4[58][15:8] = buffer_data_2[455:448];
        layer4[58][23:16] = buffer_data_2[463:456];
        layer4[58][31:24] = buffer_data_2[471:464];
        layer4[58][39:32] = buffer_data_2[479:472];
        layer4[58][47:40] = buffer_data_2[487:480];
        layer4[58][55:48] = buffer_data_2[495:488];
        layer5[58][7:0] = buffer_data_1[447:440];
        layer5[58][15:8] = buffer_data_1[455:448];
        layer5[58][23:16] = buffer_data_1[463:456];
        layer5[58][31:24] = buffer_data_1[471:464];
        layer5[58][39:32] = buffer_data_1[479:472];
        layer5[58][47:40] = buffer_data_1[487:480];
        layer5[58][55:48] = buffer_data_1[495:488];
        layer6[58][7:0] = buffer_data_0[447:440];
        layer6[58][15:8] = buffer_data_0[455:448];
        layer6[58][23:16] = buffer_data_0[463:456];
        layer6[58][31:24] = buffer_data_0[471:464];
        layer6[58][39:32] = buffer_data_0[479:472];
        layer6[58][47:40] = buffer_data_0[487:480];
        layer6[58][55:48] = buffer_data_0[495:488];
        layer0[59][7:0] = buffer_data_6[455:448];
        layer0[59][15:8] = buffer_data_6[463:456];
        layer0[59][23:16] = buffer_data_6[471:464];
        layer0[59][31:24] = buffer_data_6[479:472];
        layer0[59][39:32] = buffer_data_6[487:480];
        layer0[59][47:40] = buffer_data_6[495:488];
        layer0[59][55:48] = buffer_data_6[503:496];
        layer1[59][7:0] = buffer_data_5[455:448];
        layer1[59][15:8] = buffer_data_5[463:456];
        layer1[59][23:16] = buffer_data_5[471:464];
        layer1[59][31:24] = buffer_data_5[479:472];
        layer1[59][39:32] = buffer_data_5[487:480];
        layer1[59][47:40] = buffer_data_5[495:488];
        layer1[59][55:48] = buffer_data_5[503:496];
        layer2[59][7:0] = buffer_data_4[455:448];
        layer2[59][15:8] = buffer_data_4[463:456];
        layer2[59][23:16] = buffer_data_4[471:464];
        layer2[59][31:24] = buffer_data_4[479:472];
        layer2[59][39:32] = buffer_data_4[487:480];
        layer2[59][47:40] = buffer_data_4[495:488];
        layer2[59][55:48] = buffer_data_4[503:496];
        layer3[59][7:0] = buffer_data_3[455:448];
        layer3[59][15:8] = buffer_data_3[463:456];
        layer3[59][23:16] = buffer_data_3[471:464];
        layer3[59][31:24] = buffer_data_3[479:472];
        layer3[59][39:32] = buffer_data_3[487:480];
        layer3[59][47:40] = buffer_data_3[495:488];
        layer3[59][55:48] = buffer_data_3[503:496];
        layer4[59][7:0] = buffer_data_2[455:448];
        layer4[59][15:8] = buffer_data_2[463:456];
        layer4[59][23:16] = buffer_data_2[471:464];
        layer4[59][31:24] = buffer_data_2[479:472];
        layer4[59][39:32] = buffer_data_2[487:480];
        layer4[59][47:40] = buffer_data_2[495:488];
        layer4[59][55:48] = buffer_data_2[503:496];
        layer5[59][7:0] = buffer_data_1[455:448];
        layer5[59][15:8] = buffer_data_1[463:456];
        layer5[59][23:16] = buffer_data_1[471:464];
        layer5[59][31:24] = buffer_data_1[479:472];
        layer5[59][39:32] = buffer_data_1[487:480];
        layer5[59][47:40] = buffer_data_1[495:488];
        layer5[59][55:48] = buffer_data_1[503:496];
        layer6[59][7:0] = buffer_data_0[455:448];
        layer6[59][15:8] = buffer_data_0[463:456];
        layer6[59][23:16] = buffer_data_0[471:464];
        layer6[59][31:24] = buffer_data_0[479:472];
        layer6[59][39:32] = buffer_data_0[487:480];
        layer6[59][47:40] = buffer_data_0[495:488];
        layer6[59][55:48] = buffer_data_0[503:496];
        layer0[60][7:0] = buffer_data_6[463:456];
        layer0[60][15:8] = buffer_data_6[471:464];
        layer0[60][23:16] = buffer_data_6[479:472];
        layer0[60][31:24] = buffer_data_6[487:480];
        layer0[60][39:32] = buffer_data_6[495:488];
        layer0[60][47:40] = buffer_data_6[503:496];
        layer0[60][55:48] = buffer_data_6[511:504];
        layer1[60][7:0] = buffer_data_5[463:456];
        layer1[60][15:8] = buffer_data_5[471:464];
        layer1[60][23:16] = buffer_data_5[479:472];
        layer1[60][31:24] = buffer_data_5[487:480];
        layer1[60][39:32] = buffer_data_5[495:488];
        layer1[60][47:40] = buffer_data_5[503:496];
        layer1[60][55:48] = buffer_data_5[511:504];
        layer2[60][7:0] = buffer_data_4[463:456];
        layer2[60][15:8] = buffer_data_4[471:464];
        layer2[60][23:16] = buffer_data_4[479:472];
        layer2[60][31:24] = buffer_data_4[487:480];
        layer2[60][39:32] = buffer_data_4[495:488];
        layer2[60][47:40] = buffer_data_4[503:496];
        layer2[60][55:48] = buffer_data_4[511:504];
        layer3[60][7:0] = buffer_data_3[463:456];
        layer3[60][15:8] = buffer_data_3[471:464];
        layer3[60][23:16] = buffer_data_3[479:472];
        layer3[60][31:24] = buffer_data_3[487:480];
        layer3[60][39:32] = buffer_data_3[495:488];
        layer3[60][47:40] = buffer_data_3[503:496];
        layer3[60][55:48] = buffer_data_3[511:504];
        layer4[60][7:0] = buffer_data_2[463:456];
        layer4[60][15:8] = buffer_data_2[471:464];
        layer4[60][23:16] = buffer_data_2[479:472];
        layer4[60][31:24] = buffer_data_2[487:480];
        layer4[60][39:32] = buffer_data_2[495:488];
        layer4[60][47:40] = buffer_data_2[503:496];
        layer4[60][55:48] = buffer_data_2[511:504];
        layer5[60][7:0] = buffer_data_1[463:456];
        layer5[60][15:8] = buffer_data_1[471:464];
        layer5[60][23:16] = buffer_data_1[479:472];
        layer5[60][31:24] = buffer_data_1[487:480];
        layer5[60][39:32] = buffer_data_1[495:488];
        layer5[60][47:40] = buffer_data_1[503:496];
        layer5[60][55:48] = buffer_data_1[511:504];
        layer6[60][7:0] = buffer_data_0[463:456];
        layer6[60][15:8] = buffer_data_0[471:464];
        layer6[60][23:16] = buffer_data_0[479:472];
        layer6[60][31:24] = buffer_data_0[487:480];
        layer6[60][39:32] = buffer_data_0[495:488];
        layer6[60][47:40] = buffer_data_0[503:496];
        layer6[60][55:48] = buffer_data_0[511:504];
        layer0[61][7:0] = buffer_data_6[471:464];
        layer0[61][15:8] = buffer_data_6[479:472];
        layer0[61][23:16] = buffer_data_6[487:480];
        layer0[61][31:24] = buffer_data_6[495:488];
        layer0[61][39:32] = buffer_data_6[503:496];
        layer0[61][47:40] = buffer_data_6[511:504];
        layer0[61][55:48] = buffer_data_6[519:512];
        layer1[61][7:0] = buffer_data_5[471:464];
        layer1[61][15:8] = buffer_data_5[479:472];
        layer1[61][23:16] = buffer_data_5[487:480];
        layer1[61][31:24] = buffer_data_5[495:488];
        layer1[61][39:32] = buffer_data_5[503:496];
        layer1[61][47:40] = buffer_data_5[511:504];
        layer1[61][55:48] = buffer_data_5[519:512];
        layer2[61][7:0] = buffer_data_4[471:464];
        layer2[61][15:8] = buffer_data_4[479:472];
        layer2[61][23:16] = buffer_data_4[487:480];
        layer2[61][31:24] = buffer_data_4[495:488];
        layer2[61][39:32] = buffer_data_4[503:496];
        layer2[61][47:40] = buffer_data_4[511:504];
        layer2[61][55:48] = buffer_data_4[519:512];
        layer3[61][7:0] = buffer_data_3[471:464];
        layer3[61][15:8] = buffer_data_3[479:472];
        layer3[61][23:16] = buffer_data_3[487:480];
        layer3[61][31:24] = buffer_data_3[495:488];
        layer3[61][39:32] = buffer_data_3[503:496];
        layer3[61][47:40] = buffer_data_3[511:504];
        layer3[61][55:48] = buffer_data_3[519:512];
        layer4[61][7:0] = buffer_data_2[471:464];
        layer4[61][15:8] = buffer_data_2[479:472];
        layer4[61][23:16] = buffer_data_2[487:480];
        layer4[61][31:24] = buffer_data_2[495:488];
        layer4[61][39:32] = buffer_data_2[503:496];
        layer4[61][47:40] = buffer_data_2[511:504];
        layer4[61][55:48] = buffer_data_2[519:512];
        layer5[61][7:0] = buffer_data_1[471:464];
        layer5[61][15:8] = buffer_data_1[479:472];
        layer5[61][23:16] = buffer_data_1[487:480];
        layer5[61][31:24] = buffer_data_1[495:488];
        layer5[61][39:32] = buffer_data_1[503:496];
        layer5[61][47:40] = buffer_data_1[511:504];
        layer5[61][55:48] = buffer_data_1[519:512];
        layer6[61][7:0] = buffer_data_0[471:464];
        layer6[61][15:8] = buffer_data_0[479:472];
        layer6[61][23:16] = buffer_data_0[487:480];
        layer6[61][31:24] = buffer_data_0[495:488];
        layer6[61][39:32] = buffer_data_0[503:496];
        layer6[61][47:40] = buffer_data_0[511:504];
        layer6[61][55:48] = buffer_data_0[519:512];
        layer0[62][7:0] = buffer_data_6[479:472];
        layer0[62][15:8] = buffer_data_6[487:480];
        layer0[62][23:16] = buffer_data_6[495:488];
        layer0[62][31:24] = buffer_data_6[503:496];
        layer0[62][39:32] = buffer_data_6[511:504];
        layer0[62][47:40] = buffer_data_6[519:512];
        layer0[62][55:48] = buffer_data_6[527:520];
        layer1[62][7:0] = buffer_data_5[479:472];
        layer1[62][15:8] = buffer_data_5[487:480];
        layer1[62][23:16] = buffer_data_5[495:488];
        layer1[62][31:24] = buffer_data_5[503:496];
        layer1[62][39:32] = buffer_data_5[511:504];
        layer1[62][47:40] = buffer_data_5[519:512];
        layer1[62][55:48] = buffer_data_5[527:520];
        layer2[62][7:0] = buffer_data_4[479:472];
        layer2[62][15:8] = buffer_data_4[487:480];
        layer2[62][23:16] = buffer_data_4[495:488];
        layer2[62][31:24] = buffer_data_4[503:496];
        layer2[62][39:32] = buffer_data_4[511:504];
        layer2[62][47:40] = buffer_data_4[519:512];
        layer2[62][55:48] = buffer_data_4[527:520];
        layer3[62][7:0] = buffer_data_3[479:472];
        layer3[62][15:8] = buffer_data_3[487:480];
        layer3[62][23:16] = buffer_data_3[495:488];
        layer3[62][31:24] = buffer_data_3[503:496];
        layer3[62][39:32] = buffer_data_3[511:504];
        layer3[62][47:40] = buffer_data_3[519:512];
        layer3[62][55:48] = buffer_data_3[527:520];
        layer4[62][7:0] = buffer_data_2[479:472];
        layer4[62][15:8] = buffer_data_2[487:480];
        layer4[62][23:16] = buffer_data_2[495:488];
        layer4[62][31:24] = buffer_data_2[503:496];
        layer4[62][39:32] = buffer_data_2[511:504];
        layer4[62][47:40] = buffer_data_2[519:512];
        layer4[62][55:48] = buffer_data_2[527:520];
        layer5[62][7:0] = buffer_data_1[479:472];
        layer5[62][15:8] = buffer_data_1[487:480];
        layer5[62][23:16] = buffer_data_1[495:488];
        layer5[62][31:24] = buffer_data_1[503:496];
        layer5[62][39:32] = buffer_data_1[511:504];
        layer5[62][47:40] = buffer_data_1[519:512];
        layer5[62][55:48] = buffer_data_1[527:520];
        layer6[62][7:0] = buffer_data_0[479:472];
        layer6[62][15:8] = buffer_data_0[487:480];
        layer6[62][23:16] = buffer_data_0[495:488];
        layer6[62][31:24] = buffer_data_0[503:496];
        layer6[62][39:32] = buffer_data_0[511:504];
        layer6[62][47:40] = buffer_data_0[519:512];
        layer6[62][55:48] = buffer_data_0[527:520];
        layer0[63][7:0] = buffer_data_6[487:480];
        layer0[63][15:8] = buffer_data_6[495:488];
        layer0[63][23:16] = buffer_data_6[503:496];
        layer0[63][31:24] = buffer_data_6[511:504];
        layer0[63][39:32] = buffer_data_6[519:512];
        layer0[63][47:40] = buffer_data_6[527:520];
        layer0[63][55:48] = buffer_data_6[535:528];
        layer1[63][7:0] = buffer_data_5[487:480];
        layer1[63][15:8] = buffer_data_5[495:488];
        layer1[63][23:16] = buffer_data_5[503:496];
        layer1[63][31:24] = buffer_data_5[511:504];
        layer1[63][39:32] = buffer_data_5[519:512];
        layer1[63][47:40] = buffer_data_5[527:520];
        layer1[63][55:48] = buffer_data_5[535:528];
        layer2[63][7:0] = buffer_data_4[487:480];
        layer2[63][15:8] = buffer_data_4[495:488];
        layer2[63][23:16] = buffer_data_4[503:496];
        layer2[63][31:24] = buffer_data_4[511:504];
        layer2[63][39:32] = buffer_data_4[519:512];
        layer2[63][47:40] = buffer_data_4[527:520];
        layer2[63][55:48] = buffer_data_4[535:528];
        layer3[63][7:0] = buffer_data_3[487:480];
        layer3[63][15:8] = buffer_data_3[495:488];
        layer3[63][23:16] = buffer_data_3[503:496];
        layer3[63][31:24] = buffer_data_3[511:504];
        layer3[63][39:32] = buffer_data_3[519:512];
        layer3[63][47:40] = buffer_data_3[527:520];
        layer3[63][55:48] = buffer_data_3[535:528];
        layer4[63][7:0] = buffer_data_2[487:480];
        layer4[63][15:8] = buffer_data_2[495:488];
        layer4[63][23:16] = buffer_data_2[503:496];
        layer4[63][31:24] = buffer_data_2[511:504];
        layer4[63][39:32] = buffer_data_2[519:512];
        layer4[63][47:40] = buffer_data_2[527:520];
        layer4[63][55:48] = buffer_data_2[535:528];
        layer5[63][7:0] = buffer_data_1[487:480];
        layer5[63][15:8] = buffer_data_1[495:488];
        layer5[63][23:16] = buffer_data_1[503:496];
        layer5[63][31:24] = buffer_data_1[511:504];
        layer5[63][39:32] = buffer_data_1[519:512];
        layer5[63][47:40] = buffer_data_1[527:520];
        layer5[63][55:48] = buffer_data_1[535:528];
        layer6[63][7:0] = buffer_data_0[487:480];
        layer6[63][15:8] = buffer_data_0[495:488];
        layer6[63][23:16] = buffer_data_0[503:496];
        layer6[63][31:24] = buffer_data_0[511:504];
        layer6[63][39:32] = buffer_data_0[519:512];
        layer6[63][47:40] = buffer_data_0[527:520];
        layer6[63][55:48] = buffer_data_0[535:528];
    end
    ST_GAUSSIAN_1: begin
        layer0[0][7:0] = buffer_data_6[495:488];
        layer0[0][15:8] = buffer_data_6[503:496];
        layer0[0][23:16] = buffer_data_6[511:504];
        layer0[0][31:24] = buffer_data_6[519:512];
        layer0[0][39:32] = buffer_data_6[527:520];
        layer0[0][47:40] = buffer_data_6[535:528];
        layer0[0][55:48] = buffer_data_6[543:536];
        layer1[0][7:0] = buffer_data_5[495:488];
        layer1[0][15:8] = buffer_data_5[503:496];
        layer1[0][23:16] = buffer_data_5[511:504];
        layer1[0][31:24] = buffer_data_5[519:512];
        layer1[0][39:32] = buffer_data_5[527:520];
        layer1[0][47:40] = buffer_data_5[535:528];
        layer1[0][55:48] = buffer_data_5[543:536];
        layer2[0][7:0] = buffer_data_4[495:488];
        layer2[0][15:8] = buffer_data_4[503:496];
        layer2[0][23:16] = buffer_data_4[511:504];
        layer2[0][31:24] = buffer_data_4[519:512];
        layer2[0][39:32] = buffer_data_4[527:520];
        layer2[0][47:40] = buffer_data_4[535:528];
        layer2[0][55:48] = buffer_data_4[543:536];
        layer3[0][7:0] = buffer_data_3[495:488];
        layer3[0][15:8] = buffer_data_3[503:496];
        layer3[0][23:16] = buffer_data_3[511:504];
        layer3[0][31:24] = buffer_data_3[519:512];
        layer3[0][39:32] = buffer_data_3[527:520];
        layer3[0][47:40] = buffer_data_3[535:528];
        layer3[0][55:48] = buffer_data_3[543:536];
        layer4[0][7:0] = buffer_data_2[495:488];
        layer4[0][15:8] = buffer_data_2[503:496];
        layer4[0][23:16] = buffer_data_2[511:504];
        layer4[0][31:24] = buffer_data_2[519:512];
        layer4[0][39:32] = buffer_data_2[527:520];
        layer4[0][47:40] = buffer_data_2[535:528];
        layer4[0][55:48] = buffer_data_2[543:536];
        layer5[0][7:0] = buffer_data_1[495:488];
        layer5[0][15:8] = buffer_data_1[503:496];
        layer5[0][23:16] = buffer_data_1[511:504];
        layer5[0][31:24] = buffer_data_1[519:512];
        layer5[0][39:32] = buffer_data_1[527:520];
        layer5[0][47:40] = buffer_data_1[535:528];
        layer5[0][55:48] = buffer_data_1[543:536];
        layer6[0][7:0] = buffer_data_0[495:488];
        layer6[0][15:8] = buffer_data_0[503:496];
        layer6[0][23:16] = buffer_data_0[511:504];
        layer6[0][31:24] = buffer_data_0[519:512];
        layer6[0][39:32] = buffer_data_0[527:520];
        layer6[0][47:40] = buffer_data_0[535:528];
        layer6[0][55:48] = buffer_data_0[543:536];
        layer0[1][7:0] = buffer_data_6[503:496];
        layer0[1][15:8] = buffer_data_6[511:504];
        layer0[1][23:16] = buffer_data_6[519:512];
        layer0[1][31:24] = buffer_data_6[527:520];
        layer0[1][39:32] = buffer_data_6[535:528];
        layer0[1][47:40] = buffer_data_6[543:536];
        layer0[1][55:48] = buffer_data_6[551:544];
        layer1[1][7:0] = buffer_data_5[503:496];
        layer1[1][15:8] = buffer_data_5[511:504];
        layer1[1][23:16] = buffer_data_5[519:512];
        layer1[1][31:24] = buffer_data_5[527:520];
        layer1[1][39:32] = buffer_data_5[535:528];
        layer1[1][47:40] = buffer_data_5[543:536];
        layer1[1][55:48] = buffer_data_5[551:544];
        layer2[1][7:0] = buffer_data_4[503:496];
        layer2[1][15:8] = buffer_data_4[511:504];
        layer2[1][23:16] = buffer_data_4[519:512];
        layer2[1][31:24] = buffer_data_4[527:520];
        layer2[1][39:32] = buffer_data_4[535:528];
        layer2[1][47:40] = buffer_data_4[543:536];
        layer2[1][55:48] = buffer_data_4[551:544];
        layer3[1][7:0] = buffer_data_3[503:496];
        layer3[1][15:8] = buffer_data_3[511:504];
        layer3[1][23:16] = buffer_data_3[519:512];
        layer3[1][31:24] = buffer_data_3[527:520];
        layer3[1][39:32] = buffer_data_3[535:528];
        layer3[1][47:40] = buffer_data_3[543:536];
        layer3[1][55:48] = buffer_data_3[551:544];
        layer4[1][7:0] = buffer_data_2[503:496];
        layer4[1][15:8] = buffer_data_2[511:504];
        layer4[1][23:16] = buffer_data_2[519:512];
        layer4[1][31:24] = buffer_data_2[527:520];
        layer4[1][39:32] = buffer_data_2[535:528];
        layer4[1][47:40] = buffer_data_2[543:536];
        layer4[1][55:48] = buffer_data_2[551:544];
        layer5[1][7:0] = buffer_data_1[503:496];
        layer5[1][15:8] = buffer_data_1[511:504];
        layer5[1][23:16] = buffer_data_1[519:512];
        layer5[1][31:24] = buffer_data_1[527:520];
        layer5[1][39:32] = buffer_data_1[535:528];
        layer5[1][47:40] = buffer_data_1[543:536];
        layer5[1][55:48] = buffer_data_1[551:544];
        layer6[1][7:0] = buffer_data_0[503:496];
        layer6[1][15:8] = buffer_data_0[511:504];
        layer6[1][23:16] = buffer_data_0[519:512];
        layer6[1][31:24] = buffer_data_0[527:520];
        layer6[1][39:32] = buffer_data_0[535:528];
        layer6[1][47:40] = buffer_data_0[543:536];
        layer6[1][55:48] = buffer_data_0[551:544];
        layer0[2][7:0] = buffer_data_6[511:504];
        layer0[2][15:8] = buffer_data_6[519:512];
        layer0[2][23:16] = buffer_data_6[527:520];
        layer0[2][31:24] = buffer_data_6[535:528];
        layer0[2][39:32] = buffer_data_6[543:536];
        layer0[2][47:40] = buffer_data_6[551:544];
        layer0[2][55:48] = buffer_data_6[559:552];
        layer1[2][7:0] = buffer_data_5[511:504];
        layer1[2][15:8] = buffer_data_5[519:512];
        layer1[2][23:16] = buffer_data_5[527:520];
        layer1[2][31:24] = buffer_data_5[535:528];
        layer1[2][39:32] = buffer_data_5[543:536];
        layer1[2][47:40] = buffer_data_5[551:544];
        layer1[2][55:48] = buffer_data_5[559:552];
        layer2[2][7:0] = buffer_data_4[511:504];
        layer2[2][15:8] = buffer_data_4[519:512];
        layer2[2][23:16] = buffer_data_4[527:520];
        layer2[2][31:24] = buffer_data_4[535:528];
        layer2[2][39:32] = buffer_data_4[543:536];
        layer2[2][47:40] = buffer_data_4[551:544];
        layer2[2][55:48] = buffer_data_4[559:552];
        layer3[2][7:0] = buffer_data_3[511:504];
        layer3[2][15:8] = buffer_data_3[519:512];
        layer3[2][23:16] = buffer_data_3[527:520];
        layer3[2][31:24] = buffer_data_3[535:528];
        layer3[2][39:32] = buffer_data_3[543:536];
        layer3[2][47:40] = buffer_data_3[551:544];
        layer3[2][55:48] = buffer_data_3[559:552];
        layer4[2][7:0] = buffer_data_2[511:504];
        layer4[2][15:8] = buffer_data_2[519:512];
        layer4[2][23:16] = buffer_data_2[527:520];
        layer4[2][31:24] = buffer_data_2[535:528];
        layer4[2][39:32] = buffer_data_2[543:536];
        layer4[2][47:40] = buffer_data_2[551:544];
        layer4[2][55:48] = buffer_data_2[559:552];
        layer5[2][7:0] = buffer_data_1[511:504];
        layer5[2][15:8] = buffer_data_1[519:512];
        layer5[2][23:16] = buffer_data_1[527:520];
        layer5[2][31:24] = buffer_data_1[535:528];
        layer5[2][39:32] = buffer_data_1[543:536];
        layer5[2][47:40] = buffer_data_1[551:544];
        layer5[2][55:48] = buffer_data_1[559:552];
        layer6[2][7:0] = buffer_data_0[511:504];
        layer6[2][15:8] = buffer_data_0[519:512];
        layer6[2][23:16] = buffer_data_0[527:520];
        layer6[2][31:24] = buffer_data_0[535:528];
        layer6[2][39:32] = buffer_data_0[543:536];
        layer6[2][47:40] = buffer_data_0[551:544];
        layer6[2][55:48] = buffer_data_0[559:552];
        layer0[3][7:0] = buffer_data_6[519:512];
        layer0[3][15:8] = buffer_data_6[527:520];
        layer0[3][23:16] = buffer_data_6[535:528];
        layer0[3][31:24] = buffer_data_6[543:536];
        layer0[3][39:32] = buffer_data_6[551:544];
        layer0[3][47:40] = buffer_data_6[559:552];
        layer0[3][55:48] = buffer_data_6[567:560];
        layer1[3][7:0] = buffer_data_5[519:512];
        layer1[3][15:8] = buffer_data_5[527:520];
        layer1[3][23:16] = buffer_data_5[535:528];
        layer1[3][31:24] = buffer_data_5[543:536];
        layer1[3][39:32] = buffer_data_5[551:544];
        layer1[3][47:40] = buffer_data_5[559:552];
        layer1[3][55:48] = buffer_data_5[567:560];
        layer2[3][7:0] = buffer_data_4[519:512];
        layer2[3][15:8] = buffer_data_4[527:520];
        layer2[3][23:16] = buffer_data_4[535:528];
        layer2[3][31:24] = buffer_data_4[543:536];
        layer2[3][39:32] = buffer_data_4[551:544];
        layer2[3][47:40] = buffer_data_4[559:552];
        layer2[3][55:48] = buffer_data_4[567:560];
        layer3[3][7:0] = buffer_data_3[519:512];
        layer3[3][15:8] = buffer_data_3[527:520];
        layer3[3][23:16] = buffer_data_3[535:528];
        layer3[3][31:24] = buffer_data_3[543:536];
        layer3[3][39:32] = buffer_data_3[551:544];
        layer3[3][47:40] = buffer_data_3[559:552];
        layer3[3][55:48] = buffer_data_3[567:560];
        layer4[3][7:0] = buffer_data_2[519:512];
        layer4[3][15:8] = buffer_data_2[527:520];
        layer4[3][23:16] = buffer_data_2[535:528];
        layer4[3][31:24] = buffer_data_2[543:536];
        layer4[3][39:32] = buffer_data_2[551:544];
        layer4[3][47:40] = buffer_data_2[559:552];
        layer4[3][55:48] = buffer_data_2[567:560];
        layer5[3][7:0] = buffer_data_1[519:512];
        layer5[3][15:8] = buffer_data_1[527:520];
        layer5[3][23:16] = buffer_data_1[535:528];
        layer5[3][31:24] = buffer_data_1[543:536];
        layer5[3][39:32] = buffer_data_1[551:544];
        layer5[3][47:40] = buffer_data_1[559:552];
        layer5[3][55:48] = buffer_data_1[567:560];
        layer6[3][7:0] = buffer_data_0[519:512];
        layer6[3][15:8] = buffer_data_0[527:520];
        layer6[3][23:16] = buffer_data_0[535:528];
        layer6[3][31:24] = buffer_data_0[543:536];
        layer6[3][39:32] = buffer_data_0[551:544];
        layer6[3][47:40] = buffer_data_0[559:552];
        layer6[3][55:48] = buffer_data_0[567:560];
        layer0[4][7:0] = buffer_data_6[527:520];
        layer0[4][15:8] = buffer_data_6[535:528];
        layer0[4][23:16] = buffer_data_6[543:536];
        layer0[4][31:24] = buffer_data_6[551:544];
        layer0[4][39:32] = buffer_data_6[559:552];
        layer0[4][47:40] = buffer_data_6[567:560];
        layer0[4][55:48] = buffer_data_6[575:568];
        layer1[4][7:0] = buffer_data_5[527:520];
        layer1[4][15:8] = buffer_data_5[535:528];
        layer1[4][23:16] = buffer_data_5[543:536];
        layer1[4][31:24] = buffer_data_5[551:544];
        layer1[4][39:32] = buffer_data_5[559:552];
        layer1[4][47:40] = buffer_data_5[567:560];
        layer1[4][55:48] = buffer_data_5[575:568];
        layer2[4][7:0] = buffer_data_4[527:520];
        layer2[4][15:8] = buffer_data_4[535:528];
        layer2[4][23:16] = buffer_data_4[543:536];
        layer2[4][31:24] = buffer_data_4[551:544];
        layer2[4][39:32] = buffer_data_4[559:552];
        layer2[4][47:40] = buffer_data_4[567:560];
        layer2[4][55:48] = buffer_data_4[575:568];
        layer3[4][7:0] = buffer_data_3[527:520];
        layer3[4][15:8] = buffer_data_3[535:528];
        layer3[4][23:16] = buffer_data_3[543:536];
        layer3[4][31:24] = buffer_data_3[551:544];
        layer3[4][39:32] = buffer_data_3[559:552];
        layer3[4][47:40] = buffer_data_3[567:560];
        layer3[4][55:48] = buffer_data_3[575:568];
        layer4[4][7:0] = buffer_data_2[527:520];
        layer4[4][15:8] = buffer_data_2[535:528];
        layer4[4][23:16] = buffer_data_2[543:536];
        layer4[4][31:24] = buffer_data_2[551:544];
        layer4[4][39:32] = buffer_data_2[559:552];
        layer4[4][47:40] = buffer_data_2[567:560];
        layer4[4][55:48] = buffer_data_2[575:568];
        layer5[4][7:0] = buffer_data_1[527:520];
        layer5[4][15:8] = buffer_data_1[535:528];
        layer5[4][23:16] = buffer_data_1[543:536];
        layer5[4][31:24] = buffer_data_1[551:544];
        layer5[4][39:32] = buffer_data_1[559:552];
        layer5[4][47:40] = buffer_data_1[567:560];
        layer5[4][55:48] = buffer_data_1[575:568];
        layer6[4][7:0] = buffer_data_0[527:520];
        layer6[4][15:8] = buffer_data_0[535:528];
        layer6[4][23:16] = buffer_data_0[543:536];
        layer6[4][31:24] = buffer_data_0[551:544];
        layer6[4][39:32] = buffer_data_0[559:552];
        layer6[4][47:40] = buffer_data_0[567:560];
        layer6[4][55:48] = buffer_data_0[575:568];
        layer0[5][7:0] = buffer_data_6[535:528];
        layer0[5][15:8] = buffer_data_6[543:536];
        layer0[5][23:16] = buffer_data_6[551:544];
        layer0[5][31:24] = buffer_data_6[559:552];
        layer0[5][39:32] = buffer_data_6[567:560];
        layer0[5][47:40] = buffer_data_6[575:568];
        layer0[5][55:48] = buffer_data_6[583:576];
        layer1[5][7:0] = buffer_data_5[535:528];
        layer1[5][15:8] = buffer_data_5[543:536];
        layer1[5][23:16] = buffer_data_5[551:544];
        layer1[5][31:24] = buffer_data_5[559:552];
        layer1[5][39:32] = buffer_data_5[567:560];
        layer1[5][47:40] = buffer_data_5[575:568];
        layer1[5][55:48] = buffer_data_5[583:576];
        layer2[5][7:0] = buffer_data_4[535:528];
        layer2[5][15:8] = buffer_data_4[543:536];
        layer2[5][23:16] = buffer_data_4[551:544];
        layer2[5][31:24] = buffer_data_4[559:552];
        layer2[5][39:32] = buffer_data_4[567:560];
        layer2[5][47:40] = buffer_data_4[575:568];
        layer2[5][55:48] = buffer_data_4[583:576];
        layer3[5][7:0] = buffer_data_3[535:528];
        layer3[5][15:8] = buffer_data_3[543:536];
        layer3[5][23:16] = buffer_data_3[551:544];
        layer3[5][31:24] = buffer_data_3[559:552];
        layer3[5][39:32] = buffer_data_3[567:560];
        layer3[5][47:40] = buffer_data_3[575:568];
        layer3[5][55:48] = buffer_data_3[583:576];
        layer4[5][7:0] = buffer_data_2[535:528];
        layer4[5][15:8] = buffer_data_2[543:536];
        layer4[5][23:16] = buffer_data_2[551:544];
        layer4[5][31:24] = buffer_data_2[559:552];
        layer4[5][39:32] = buffer_data_2[567:560];
        layer4[5][47:40] = buffer_data_2[575:568];
        layer4[5][55:48] = buffer_data_2[583:576];
        layer5[5][7:0] = buffer_data_1[535:528];
        layer5[5][15:8] = buffer_data_1[543:536];
        layer5[5][23:16] = buffer_data_1[551:544];
        layer5[5][31:24] = buffer_data_1[559:552];
        layer5[5][39:32] = buffer_data_1[567:560];
        layer5[5][47:40] = buffer_data_1[575:568];
        layer5[5][55:48] = buffer_data_1[583:576];
        layer6[5][7:0] = buffer_data_0[535:528];
        layer6[5][15:8] = buffer_data_0[543:536];
        layer6[5][23:16] = buffer_data_0[551:544];
        layer6[5][31:24] = buffer_data_0[559:552];
        layer6[5][39:32] = buffer_data_0[567:560];
        layer6[5][47:40] = buffer_data_0[575:568];
        layer6[5][55:48] = buffer_data_0[583:576];
        layer0[6][7:0] = buffer_data_6[543:536];
        layer0[6][15:8] = buffer_data_6[551:544];
        layer0[6][23:16] = buffer_data_6[559:552];
        layer0[6][31:24] = buffer_data_6[567:560];
        layer0[6][39:32] = buffer_data_6[575:568];
        layer0[6][47:40] = buffer_data_6[583:576];
        layer0[6][55:48] = buffer_data_6[591:584];
        layer1[6][7:0] = buffer_data_5[543:536];
        layer1[6][15:8] = buffer_data_5[551:544];
        layer1[6][23:16] = buffer_data_5[559:552];
        layer1[6][31:24] = buffer_data_5[567:560];
        layer1[6][39:32] = buffer_data_5[575:568];
        layer1[6][47:40] = buffer_data_5[583:576];
        layer1[6][55:48] = buffer_data_5[591:584];
        layer2[6][7:0] = buffer_data_4[543:536];
        layer2[6][15:8] = buffer_data_4[551:544];
        layer2[6][23:16] = buffer_data_4[559:552];
        layer2[6][31:24] = buffer_data_4[567:560];
        layer2[6][39:32] = buffer_data_4[575:568];
        layer2[6][47:40] = buffer_data_4[583:576];
        layer2[6][55:48] = buffer_data_4[591:584];
        layer3[6][7:0] = buffer_data_3[543:536];
        layer3[6][15:8] = buffer_data_3[551:544];
        layer3[6][23:16] = buffer_data_3[559:552];
        layer3[6][31:24] = buffer_data_3[567:560];
        layer3[6][39:32] = buffer_data_3[575:568];
        layer3[6][47:40] = buffer_data_3[583:576];
        layer3[6][55:48] = buffer_data_3[591:584];
        layer4[6][7:0] = buffer_data_2[543:536];
        layer4[6][15:8] = buffer_data_2[551:544];
        layer4[6][23:16] = buffer_data_2[559:552];
        layer4[6][31:24] = buffer_data_2[567:560];
        layer4[6][39:32] = buffer_data_2[575:568];
        layer4[6][47:40] = buffer_data_2[583:576];
        layer4[6][55:48] = buffer_data_2[591:584];
        layer5[6][7:0] = buffer_data_1[543:536];
        layer5[6][15:8] = buffer_data_1[551:544];
        layer5[6][23:16] = buffer_data_1[559:552];
        layer5[6][31:24] = buffer_data_1[567:560];
        layer5[6][39:32] = buffer_data_1[575:568];
        layer5[6][47:40] = buffer_data_1[583:576];
        layer5[6][55:48] = buffer_data_1[591:584];
        layer6[6][7:0] = buffer_data_0[543:536];
        layer6[6][15:8] = buffer_data_0[551:544];
        layer6[6][23:16] = buffer_data_0[559:552];
        layer6[6][31:24] = buffer_data_0[567:560];
        layer6[6][39:32] = buffer_data_0[575:568];
        layer6[6][47:40] = buffer_data_0[583:576];
        layer6[6][55:48] = buffer_data_0[591:584];
        layer0[7][7:0] = buffer_data_6[551:544];
        layer0[7][15:8] = buffer_data_6[559:552];
        layer0[7][23:16] = buffer_data_6[567:560];
        layer0[7][31:24] = buffer_data_6[575:568];
        layer0[7][39:32] = buffer_data_6[583:576];
        layer0[7][47:40] = buffer_data_6[591:584];
        layer0[7][55:48] = buffer_data_6[599:592];
        layer1[7][7:0] = buffer_data_5[551:544];
        layer1[7][15:8] = buffer_data_5[559:552];
        layer1[7][23:16] = buffer_data_5[567:560];
        layer1[7][31:24] = buffer_data_5[575:568];
        layer1[7][39:32] = buffer_data_5[583:576];
        layer1[7][47:40] = buffer_data_5[591:584];
        layer1[7][55:48] = buffer_data_5[599:592];
        layer2[7][7:0] = buffer_data_4[551:544];
        layer2[7][15:8] = buffer_data_4[559:552];
        layer2[7][23:16] = buffer_data_4[567:560];
        layer2[7][31:24] = buffer_data_4[575:568];
        layer2[7][39:32] = buffer_data_4[583:576];
        layer2[7][47:40] = buffer_data_4[591:584];
        layer2[7][55:48] = buffer_data_4[599:592];
        layer3[7][7:0] = buffer_data_3[551:544];
        layer3[7][15:8] = buffer_data_3[559:552];
        layer3[7][23:16] = buffer_data_3[567:560];
        layer3[7][31:24] = buffer_data_3[575:568];
        layer3[7][39:32] = buffer_data_3[583:576];
        layer3[7][47:40] = buffer_data_3[591:584];
        layer3[7][55:48] = buffer_data_3[599:592];
        layer4[7][7:0] = buffer_data_2[551:544];
        layer4[7][15:8] = buffer_data_2[559:552];
        layer4[7][23:16] = buffer_data_2[567:560];
        layer4[7][31:24] = buffer_data_2[575:568];
        layer4[7][39:32] = buffer_data_2[583:576];
        layer4[7][47:40] = buffer_data_2[591:584];
        layer4[7][55:48] = buffer_data_2[599:592];
        layer5[7][7:0] = buffer_data_1[551:544];
        layer5[7][15:8] = buffer_data_1[559:552];
        layer5[7][23:16] = buffer_data_1[567:560];
        layer5[7][31:24] = buffer_data_1[575:568];
        layer5[7][39:32] = buffer_data_1[583:576];
        layer5[7][47:40] = buffer_data_1[591:584];
        layer5[7][55:48] = buffer_data_1[599:592];
        layer6[7][7:0] = buffer_data_0[551:544];
        layer6[7][15:8] = buffer_data_0[559:552];
        layer6[7][23:16] = buffer_data_0[567:560];
        layer6[7][31:24] = buffer_data_0[575:568];
        layer6[7][39:32] = buffer_data_0[583:576];
        layer6[7][47:40] = buffer_data_0[591:584];
        layer6[7][55:48] = buffer_data_0[599:592];
        layer0[8][7:0] = buffer_data_6[559:552];
        layer0[8][15:8] = buffer_data_6[567:560];
        layer0[8][23:16] = buffer_data_6[575:568];
        layer0[8][31:24] = buffer_data_6[583:576];
        layer0[8][39:32] = buffer_data_6[591:584];
        layer0[8][47:40] = buffer_data_6[599:592];
        layer0[8][55:48] = buffer_data_6[607:600];
        layer1[8][7:0] = buffer_data_5[559:552];
        layer1[8][15:8] = buffer_data_5[567:560];
        layer1[8][23:16] = buffer_data_5[575:568];
        layer1[8][31:24] = buffer_data_5[583:576];
        layer1[8][39:32] = buffer_data_5[591:584];
        layer1[8][47:40] = buffer_data_5[599:592];
        layer1[8][55:48] = buffer_data_5[607:600];
        layer2[8][7:0] = buffer_data_4[559:552];
        layer2[8][15:8] = buffer_data_4[567:560];
        layer2[8][23:16] = buffer_data_4[575:568];
        layer2[8][31:24] = buffer_data_4[583:576];
        layer2[8][39:32] = buffer_data_4[591:584];
        layer2[8][47:40] = buffer_data_4[599:592];
        layer2[8][55:48] = buffer_data_4[607:600];
        layer3[8][7:0] = buffer_data_3[559:552];
        layer3[8][15:8] = buffer_data_3[567:560];
        layer3[8][23:16] = buffer_data_3[575:568];
        layer3[8][31:24] = buffer_data_3[583:576];
        layer3[8][39:32] = buffer_data_3[591:584];
        layer3[8][47:40] = buffer_data_3[599:592];
        layer3[8][55:48] = buffer_data_3[607:600];
        layer4[8][7:0] = buffer_data_2[559:552];
        layer4[8][15:8] = buffer_data_2[567:560];
        layer4[8][23:16] = buffer_data_2[575:568];
        layer4[8][31:24] = buffer_data_2[583:576];
        layer4[8][39:32] = buffer_data_2[591:584];
        layer4[8][47:40] = buffer_data_2[599:592];
        layer4[8][55:48] = buffer_data_2[607:600];
        layer5[8][7:0] = buffer_data_1[559:552];
        layer5[8][15:8] = buffer_data_1[567:560];
        layer5[8][23:16] = buffer_data_1[575:568];
        layer5[8][31:24] = buffer_data_1[583:576];
        layer5[8][39:32] = buffer_data_1[591:584];
        layer5[8][47:40] = buffer_data_1[599:592];
        layer5[8][55:48] = buffer_data_1[607:600];
        layer6[8][7:0] = buffer_data_0[559:552];
        layer6[8][15:8] = buffer_data_0[567:560];
        layer6[8][23:16] = buffer_data_0[575:568];
        layer6[8][31:24] = buffer_data_0[583:576];
        layer6[8][39:32] = buffer_data_0[591:584];
        layer6[8][47:40] = buffer_data_0[599:592];
        layer6[8][55:48] = buffer_data_0[607:600];
        layer0[9][7:0] = buffer_data_6[567:560];
        layer0[9][15:8] = buffer_data_6[575:568];
        layer0[9][23:16] = buffer_data_6[583:576];
        layer0[9][31:24] = buffer_data_6[591:584];
        layer0[9][39:32] = buffer_data_6[599:592];
        layer0[9][47:40] = buffer_data_6[607:600];
        layer0[9][55:48] = buffer_data_6[615:608];
        layer1[9][7:0] = buffer_data_5[567:560];
        layer1[9][15:8] = buffer_data_5[575:568];
        layer1[9][23:16] = buffer_data_5[583:576];
        layer1[9][31:24] = buffer_data_5[591:584];
        layer1[9][39:32] = buffer_data_5[599:592];
        layer1[9][47:40] = buffer_data_5[607:600];
        layer1[9][55:48] = buffer_data_5[615:608];
        layer2[9][7:0] = buffer_data_4[567:560];
        layer2[9][15:8] = buffer_data_4[575:568];
        layer2[9][23:16] = buffer_data_4[583:576];
        layer2[9][31:24] = buffer_data_4[591:584];
        layer2[9][39:32] = buffer_data_4[599:592];
        layer2[9][47:40] = buffer_data_4[607:600];
        layer2[9][55:48] = buffer_data_4[615:608];
        layer3[9][7:0] = buffer_data_3[567:560];
        layer3[9][15:8] = buffer_data_3[575:568];
        layer3[9][23:16] = buffer_data_3[583:576];
        layer3[9][31:24] = buffer_data_3[591:584];
        layer3[9][39:32] = buffer_data_3[599:592];
        layer3[9][47:40] = buffer_data_3[607:600];
        layer3[9][55:48] = buffer_data_3[615:608];
        layer4[9][7:0] = buffer_data_2[567:560];
        layer4[9][15:8] = buffer_data_2[575:568];
        layer4[9][23:16] = buffer_data_2[583:576];
        layer4[9][31:24] = buffer_data_2[591:584];
        layer4[9][39:32] = buffer_data_2[599:592];
        layer4[9][47:40] = buffer_data_2[607:600];
        layer4[9][55:48] = buffer_data_2[615:608];
        layer5[9][7:0] = buffer_data_1[567:560];
        layer5[9][15:8] = buffer_data_1[575:568];
        layer5[9][23:16] = buffer_data_1[583:576];
        layer5[9][31:24] = buffer_data_1[591:584];
        layer5[9][39:32] = buffer_data_1[599:592];
        layer5[9][47:40] = buffer_data_1[607:600];
        layer5[9][55:48] = buffer_data_1[615:608];
        layer6[9][7:0] = buffer_data_0[567:560];
        layer6[9][15:8] = buffer_data_0[575:568];
        layer6[9][23:16] = buffer_data_0[583:576];
        layer6[9][31:24] = buffer_data_0[591:584];
        layer6[9][39:32] = buffer_data_0[599:592];
        layer6[9][47:40] = buffer_data_0[607:600];
        layer6[9][55:48] = buffer_data_0[615:608];
        layer0[10][7:0] = buffer_data_6[575:568];
        layer0[10][15:8] = buffer_data_6[583:576];
        layer0[10][23:16] = buffer_data_6[591:584];
        layer0[10][31:24] = buffer_data_6[599:592];
        layer0[10][39:32] = buffer_data_6[607:600];
        layer0[10][47:40] = buffer_data_6[615:608];
        layer0[10][55:48] = buffer_data_6[623:616];
        layer1[10][7:0] = buffer_data_5[575:568];
        layer1[10][15:8] = buffer_data_5[583:576];
        layer1[10][23:16] = buffer_data_5[591:584];
        layer1[10][31:24] = buffer_data_5[599:592];
        layer1[10][39:32] = buffer_data_5[607:600];
        layer1[10][47:40] = buffer_data_5[615:608];
        layer1[10][55:48] = buffer_data_5[623:616];
        layer2[10][7:0] = buffer_data_4[575:568];
        layer2[10][15:8] = buffer_data_4[583:576];
        layer2[10][23:16] = buffer_data_4[591:584];
        layer2[10][31:24] = buffer_data_4[599:592];
        layer2[10][39:32] = buffer_data_4[607:600];
        layer2[10][47:40] = buffer_data_4[615:608];
        layer2[10][55:48] = buffer_data_4[623:616];
        layer3[10][7:0] = buffer_data_3[575:568];
        layer3[10][15:8] = buffer_data_3[583:576];
        layer3[10][23:16] = buffer_data_3[591:584];
        layer3[10][31:24] = buffer_data_3[599:592];
        layer3[10][39:32] = buffer_data_3[607:600];
        layer3[10][47:40] = buffer_data_3[615:608];
        layer3[10][55:48] = buffer_data_3[623:616];
        layer4[10][7:0] = buffer_data_2[575:568];
        layer4[10][15:8] = buffer_data_2[583:576];
        layer4[10][23:16] = buffer_data_2[591:584];
        layer4[10][31:24] = buffer_data_2[599:592];
        layer4[10][39:32] = buffer_data_2[607:600];
        layer4[10][47:40] = buffer_data_2[615:608];
        layer4[10][55:48] = buffer_data_2[623:616];
        layer5[10][7:0] = buffer_data_1[575:568];
        layer5[10][15:8] = buffer_data_1[583:576];
        layer5[10][23:16] = buffer_data_1[591:584];
        layer5[10][31:24] = buffer_data_1[599:592];
        layer5[10][39:32] = buffer_data_1[607:600];
        layer5[10][47:40] = buffer_data_1[615:608];
        layer5[10][55:48] = buffer_data_1[623:616];
        layer6[10][7:0] = buffer_data_0[575:568];
        layer6[10][15:8] = buffer_data_0[583:576];
        layer6[10][23:16] = buffer_data_0[591:584];
        layer6[10][31:24] = buffer_data_0[599:592];
        layer6[10][39:32] = buffer_data_0[607:600];
        layer6[10][47:40] = buffer_data_0[615:608];
        layer6[10][55:48] = buffer_data_0[623:616];
        layer0[11][7:0] = buffer_data_6[583:576];
        layer0[11][15:8] = buffer_data_6[591:584];
        layer0[11][23:16] = buffer_data_6[599:592];
        layer0[11][31:24] = buffer_data_6[607:600];
        layer0[11][39:32] = buffer_data_6[615:608];
        layer0[11][47:40] = buffer_data_6[623:616];
        layer0[11][55:48] = buffer_data_6[631:624];
        layer1[11][7:0] = buffer_data_5[583:576];
        layer1[11][15:8] = buffer_data_5[591:584];
        layer1[11][23:16] = buffer_data_5[599:592];
        layer1[11][31:24] = buffer_data_5[607:600];
        layer1[11][39:32] = buffer_data_5[615:608];
        layer1[11][47:40] = buffer_data_5[623:616];
        layer1[11][55:48] = buffer_data_5[631:624];
        layer2[11][7:0] = buffer_data_4[583:576];
        layer2[11][15:8] = buffer_data_4[591:584];
        layer2[11][23:16] = buffer_data_4[599:592];
        layer2[11][31:24] = buffer_data_4[607:600];
        layer2[11][39:32] = buffer_data_4[615:608];
        layer2[11][47:40] = buffer_data_4[623:616];
        layer2[11][55:48] = buffer_data_4[631:624];
        layer3[11][7:0] = buffer_data_3[583:576];
        layer3[11][15:8] = buffer_data_3[591:584];
        layer3[11][23:16] = buffer_data_3[599:592];
        layer3[11][31:24] = buffer_data_3[607:600];
        layer3[11][39:32] = buffer_data_3[615:608];
        layer3[11][47:40] = buffer_data_3[623:616];
        layer3[11][55:48] = buffer_data_3[631:624];
        layer4[11][7:0] = buffer_data_2[583:576];
        layer4[11][15:8] = buffer_data_2[591:584];
        layer4[11][23:16] = buffer_data_2[599:592];
        layer4[11][31:24] = buffer_data_2[607:600];
        layer4[11][39:32] = buffer_data_2[615:608];
        layer4[11][47:40] = buffer_data_2[623:616];
        layer4[11][55:48] = buffer_data_2[631:624];
        layer5[11][7:0] = buffer_data_1[583:576];
        layer5[11][15:8] = buffer_data_1[591:584];
        layer5[11][23:16] = buffer_data_1[599:592];
        layer5[11][31:24] = buffer_data_1[607:600];
        layer5[11][39:32] = buffer_data_1[615:608];
        layer5[11][47:40] = buffer_data_1[623:616];
        layer5[11][55:48] = buffer_data_1[631:624];
        layer6[11][7:0] = buffer_data_0[583:576];
        layer6[11][15:8] = buffer_data_0[591:584];
        layer6[11][23:16] = buffer_data_0[599:592];
        layer6[11][31:24] = buffer_data_0[607:600];
        layer6[11][39:32] = buffer_data_0[615:608];
        layer6[11][47:40] = buffer_data_0[623:616];
        layer6[11][55:48] = buffer_data_0[631:624];
        layer0[12][7:0] = buffer_data_6[591:584];
        layer0[12][15:8] = buffer_data_6[599:592];
        layer0[12][23:16] = buffer_data_6[607:600];
        layer0[12][31:24] = buffer_data_6[615:608];
        layer0[12][39:32] = buffer_data_6[623:616];
        layer0[12][47:40] = buffer_data_6[631:624];
        layer0[12][55:48] = buffer_data_6[639:632];
        layer1[12][7:0] = buffer_data_5[591:584];
        layer1[12][15:8] = buffer_data_5[599:592];
        layer1[12][23:16] = buffer_data_5[607:600];
        layer1[12][31:24] = buffer_data_5[615:608];
        layer1[12][39:32] = buffer_data_5[623:616];
        layer1[12][47:40] = buffer_data_5[631:624];
        layer1[12][55:48] = buffer_data_5[639:632];
        layer2[12][7:0] = buffer_data_4[591:584];
        layer2[12][15:8] = buffer_data_4[599:592];
        layer2[12][23:16] = buffer_data_4[607:600];
        layer2[12][31:24] = buffer_data_4[615:608];
        layer2[12][39:32] = buffer_data_4[623:616];
        layer2[12][47:40] = buffer_data_4[631:624];
        layer2[12][55:48] = buffer_data_4[639:632];
        layer3[12][7:0] = buffer_data_3[591:584];
        layer3[12][15:8] = buffer_data_3[599:592];
        layer3[12][23:16] = buffer_data_3[607:600];
        layer3[12][31:24] = buffer_data_3[615:608];
        layer3[12][39:32] = buffer_data_3[623:616];
        layer3[12][47:40] = buffer_data_3[631:624];
        layer3[12][55:48] = buffer_data_3[639:632];
        layer4[12][7:0] = buffer_data_2[591:584];
        layer4[12][15:8] = buffer_data_2[599:592];
        layer4[12][23:16] = buffer_data_2[607:600];
        layer4[12][31:24] = buffer_data_2[615:608];
        layer4[12][39:32] = buffer_data_2[623:616];
        layer4[12][47:40] = buffer_data_2[631:624];
        layer4[12][55:48] = buffer_data_2[639:632];
        layer5[12][7:0] = buffer_data_1[591:584];
        layer5[12][15:8] = buffer_data_1[599:592];
        layer5[12][23:16] = buffer_data_1[607:600];
        layer5[12][31:24] = buffer_data_1[615:608];
        layer5[12][39:32] = buffer_data_1[623:616];
        layer5[12][47:40] = buffer_data_1[631:624];
        layer5[12][55:48] = buffer_data_1[639:632];
        layer6[12][7:0] = buffer_data_0[591:584];
        layer6[12][15:8] = buffer_data_0[599:592];
        layer6[12][23:16] = buffer_data_0[607:600];
        layer6[12][31:24] = buffer_data_0[615:608];
        layer6[12][39:32] = buffer_data_0[623:616];
        layer6[12][47:40] = buffer_data_0[631:624];
        layer6[12][55:48] = buffer_data_0[639:632];
        layer0[13][7:0] = buffer_data_6[599:592];
        layer0[13][15:8] = buffer_data_6[607:600];
        layer0[13][23:16] = buffer_data_6[615:608];
        layer0[13][31:24] = buffer_data_6[623:616];
        layer0[13][39:32] = buffer_data_6[631:624];
        layer0[13][47:40] = buffer_data_6[639:632];
        layer0[13][55:48] = buffer_data_6[647:640];
        layer1[13][7:0] = buffer_data_5[599:592];
        layer1[13][15:8] = buffer_data_5[607:600];
        layer1[13][23:16] = buffer_data_5[615:608];
        layer1[13][31:24] = buffer_data_5[623:616];
        layer1[13][39:32] = buffer_data_5[631:624];
        layer1[13][47:40] = buffer_data_5[639:632];
        layer1[13][55:48] = buffer_data_5[647:640];
        layer2[13][7:0] = buffer_data_4[599:592];
        layer2[13][15:8] = buffer_data_4[607:600];
        layer2[13][23:16] = buffer_data_4[615:608];
        layer2[13][31:24] = buffer_data_4[623:616];
        layer2[13][39:32] = buffer_data_4[631:624];
        layer2[13][47:40] = buffer_data_4[639:632];
        layer2[13][55:48] = buffer_data_4[647:640];
        layer3[13][7:0] = buffer_data_3[599:592];
        layer3[13][15:8] = buffer_data_3[607:600];
        layer3[13][23:16] = buffer_data_3[615:608];
        layer3[13][31:24] = buffer_data_3[623:616];
        layer3[13][39:32] = buffer_data_3[631:624];
        layer3[13][47:40] = buffer_data_3[639:632];
        layer3[13][55:48] = buffer_data_3[647:640];
        layer4[13][7:0] = buffer_data_2[599:592];
        layer4[13][15:8] = buffer_data_2[607:600];
        layer4[13][23:16] = buffer_data_2[615:608];
        layer4[13][31:24] = buffer_data_2[623:616];
        layer4[13][39:32] = buffer_data_2[631:624];
        layer4[13][47:40] = buffer_data_2[639:632];
        layer4[13][55:48] = buffer_data_2[647:640];
        layer5[13][7:0] = buffer_data_1[599:592];
        layer5[13][15:8] = buffer_data_1[607:600];
        layer5[13][23:16] = buffer_data_1[615:608];
        layer5[13][31:24] = buffer_data_1[623:616];
        layer5[13][39:32] = buffer_data_1[631:624];
        layer5[13][47:40] = buffer_data_1[639:632];
        layer5[13][55:48] = buffer_data_1[647:640];
        layer6[13][7:0] = buffer_data_0[599:592];
        layer6[13][15:8] = buffer_data_0[607:600];
        layer6[13][23:16] = buffer_data_0[615:608];
        layer6[13][31:24] = buffer_data_0[623:616];
        layer6[13][39:32] = buffer_data_0[631:624];
        layer6[13][47:40] = buffer_data_0[639:632];
        layer6[13][55:48] = buffer_data_0[647:640];
        layer0[14][7:0] = buffer_data_6[607:600];
        layer0[14][15:8] = buffer_data_6[615:608];
        layer0[14][23:16] = buffer_data_6[623:616];
        layer0[14][31:24] = buffer_data_6[631:624];
        layer0[14][39:32] = buffer_data_6[639:632];
        layer0[14][47:40] = buffer_data_6[647:640];
        layer0[14][55:48] = buffer_data_6[655:648];
        layer1[14][7:0] = buffer_data_5[607:600];
        layer1[14][15:8] = buffer_data_5[615:608];
        layer1[14][23:16] = buffer_data_5[623:616];
        layer1[14][31:24] = buffer_data_5[631:624];
        layer1[14][39:32] = buffer_data_5[639:632];
        layer1[14][47:40] = buffer_data_5[647:640];
        layer1[14][55:48] = buffer_data_5[655:648];
        layer2[14][7:0] = buffer_data_4[607:600];
        layer2[14][15:8] = buffer_data_4[615:608];
        layer2[14][23:16] = buffer_data_4[623:616];
        layer2[14][31:24] = buffer_data_4[631:624];
        layer2[14][39:32] = buffer_data_4[639:632];
        layer2[14][47:40] = buffer_data_4[647:640];
        layer2[14][55:48] = buffer_data_4[655:648];
        layer3[14][7:0] = buffer_data_3[607:600];
        layer3[14][15:8] = buffer_data_3[615:608];
        layer3[14][23:16] = buffer_data_3[623:616];
        layer3[14][31:24] = buffer_data_3[631:624];
        layer3[14][39:32] = buffer_data_3[639:632];
        layer3[14][47:40] = buffer_data_3[647:640];
        layer3[14][55:48] = buffer_data_3[655:648];
        layer4[14][7:0] = buffer_data_2[607:600];
        layer4[14][15:8] = buffer_data_2[615:608];
        layer4[14][23:16] = buffer_data_2[623:616];
        layer4[14][31:24] = buffer_data_2[631:624];
        layer4[14][39:32] = buffer_data_2[639:632];
        layer4[14][47:40] = buffer_data_2[647:640];
        layer4[14][55:48] = buffer_data_2[655:648];
        layer5[14][7:0] = buffer_data_1[607:600];
        layer5[14][15:8] = buffer_data_1[615:608];
        layer5[14][23:16] = buffer_data_1[623:616];
        layer5[14][31:24] = buffer_data_1[631:624];
        layer5[14][39:32] = buffer_data_1[639:632];
        layer5[14][47:40] = buffer_data_1[647:640];
        layer5[14][55:48] = buffer_data_1[655:648];
        layer6[14][7:0] = buffer_data_0[607:600];
        layer6[14][15:8] = buffer_data_0[615:608];
        layer6[14][23:16] = buffer_data_0[623:616];
        layer6[14][31:24] = buffer_data_0[631:624];
        layer6[14][39:32] = buffer_data_0[639:632];
        layer6[14][47:40] = buffer_data_0[647:640];
        layer6[14][55:48] = buffer_data_0[655:648];
        layer0[15][7:0] = buffer_data_6[615:608];
        layer0[15][15:8] = buffer_data_6[623:616];
        layer0[15][23:16] = buffer_data_6[631:624];
        layer0[15][31:24] = buffer_data_6[639:632];
        layer0[15][39:32] = buffer_data_6[647:640];
        layer0[15][47:40] = buffer_data_6[655:648];
        layer0[15][55:48] = buffer_data_6[663:656];
        layer1[15][7:0] = buffer_data_5[615:608];
        layer1[15][15:8] = buffer_data_5[623:616];
        layer1[15][23:16] = buffer_data_5[631:624];
        layer1[15][31:24] = buffer_data_5[639:632];
        layer1[15][39:32] = buffer_data_5[647:640];
        layer1[15][47:40] = buffer_data_5[655:648];
        layer1[15][55:48] = buffer_data_5[663:656];
        layer2[15][7:0] = buffer_data_4[615:608];
        layer2[15][15:8] = buffer_data_4[623:616];
        layer2[15][23:16] = buffer_data_4[631:624];
        layer2[15][31:24] = buffer_data_4[639:632];
        layer2[15][39:32] = buffer_data_4[647:640];
        layer2[15][47:40] = buffer_data_4[655:648];
        layer2[15][55:48] = buffer_data_4[663:656];
        layer3[15][7:0] = buffer_data_3[615:608];
        layer3[15][15:8] = buffer_data_3[623:616];
        layer3[15][23:16] = buffer_data_3[631:624];
        layer3[15][31:24] = buffer_data_3[639:632];
        layer3[15][39:32] = buffer_data_3[647:640];
        layer3[15][47:40] = buffer_data_3[655:648];
        layer3[15][55:48] = buffer_data_3[663:656];
        layer4[15][7:0] = buffer_data_2[615:608];
        layer4[15][15:8] = buffer_data_2[623:616];
        layer4[15][23:16] = buffer_data_2[631:624];
        layer4[15][31:24] = buffer_data_2[639:632];
        layer4[15][39:32] = buffer_data_2[647:640];
        layer4[15][47:40] = buffer_data_2[655:648];
        layer4[15][55:48] = buffer_data_2[663:656];
        layer5[15][7:0] = buffer_data_1[615:608];
        layer5[15][15:8] = buffer_data_1[623:616];
        layer5[15][23:16] = buffer_data_1[631:624];
        layer5[15][31:24] = buffer_data_1[639:632];
        layer5[15][39:32] = buffer_data_1[647:640];
        layer5[15][47:40] = buffer_data_1[655:648];
        layer5[15][55:48] = buffer_data_1[663:656];
        layer6[15][7:0] = buffer_data_0[615:608];
        layer6[15][15:8] = buffer_data_0[623:616];
        layer6[15][23:16] = buffer_data_0[631:624];
        layer6[15][31:24] = buffer_data_0[639:632];
        layer6[15][39:32] = buffer_data_0[647:640];
        layer6[15][47:40] = buffer_data_0[655:648];
        layer6[15][55:48] = buffer_data_0[663:656];
        layer0[16][7:0] = buffer_data_6[623:616];
        layer0[16][15:8] = buffer_data_6[631:624];
        layer0[16][23:16] = buffer_data_6[639:632];
        layer0[16][31:24] = buffer_data_6[647:640];
        layer0[16][39:32] = buffer_data_6[655:648];
        layer0[16][47:40] = buffer_data_6[663:656];
        layer0[16][55:48] = buffer_data_6[671:664];
        layer1[16][7:0] = buffer_data_5[623:616];
        layer1[16][15:8] = buffer_data_5[631:624];
        layer1[16][23:16] = buffer_data_5[639:632];
        layer1[16][31:24] = buffer_data_5[647:640];
        layer1[16][39:32] = buffer_data_5[655:648];
        layer1[16][47:40] = buffer_data_5[663:656];
        layer1[16][55:48] = buffer_data_5[671:664];
        layer2[16][7:0] = buffer_data_4[623:616];
        layer2[16][15:8] = buffer_data_4[631:624];
        layer2[16][23:16] = buffer_data_4[639:632];
        layer2[16][31:24] = buffer_data_4[647:640];
        layer2[16][39:32] = buffer_data_4[655:648];
        layer2[16][47:40] = buffer_data_4[663:656];
        layer2[16][55:48] = buffer_data_4[671:664];
        layer3[16][7:0] = buffer_data_3[623:616];
        layer3[16][15:8] = buffer_data_3[631:624];
        layer3[16][23:16] = buffer_data_3[639:632];
        layer3[16][31:24] = buffer_data_3[647:640];
        layer3[16][39:32] = buffer_data_3[655:648];
        layer3[16][47:40] = buffer_data_3[663:656];
        layer3[16][55:48] = buffer_data_3[671:664];
        layer4[16][7:0] = buffer_data_2[623:616];
        layer4[16][15:8] = buffer_data_2[631:624];
        layer4[16][23:16] = buffer_data_2[639:632];
        layer4[16][31:24] = buffer_data_2[647:640];
        layer4[16][39:32] = buffer_data_2[655:648];
        layer4[16][47:40] = buffer_data_2[663:656];
        layer4[16][55:48] = buffer_data_2[671:664];
        layer5[16][7:0] = buffer_data_1[623:616];
        layer5[16][15:8] = buffer_data_1[631:624];
        layer5[16][23:16] = buffer_data_1[639:632];
        layer5[16][31:24] = buffer_data_1[647:640];
        layer5[16][39:32] = buffer_data_1[655:648];
        layer5[16][47:40] = buffer_data_1[663:656];
        layer5[16][55:48] = buffer_data_1[671:664];
        layer6[16][7:0] = buffer_data_0[623:616];
        layer6[16][15:8] = buffer_data_0[631:624];
        layer6[16][23:16] = buffer_data_0[639:632];
        layer6[16][31:24] = buffer_data_0[647:640];
        layer6[16][39:32] = buffer_data_0[655:648];
        layer6[16][47:40] = buffer_data_0[663:656];
        layer6[16][55:48] = buffer_data_0[671:664];
        layer0[17][7:0] = buffer_data_6[631:624];
        layer0[17][15:8] = buffer_data_6[639:632];
        layer0[17][23:16] = buffer_data_6[647:640];
        layer0[17][31:24] = buffer_data_6[655:648];
        layer0[17][39:32] = buffer_data_6[663:656];
        layer0[17][47:40] = buffer_data_6[671:664];
        layer0[17][55:48] = buffer_data_6[679:672];
        layer1[17][7:0] = buffer_data_5[631:624];
        layer1[17][15:8] = buffer_data_5[639:632];
        layer1[17][23:16] = buffer_data_5[647:640];
        layer1[17][31:24] = buffer_data_5[655:648];
        layer1[17][39:32] = buffer_data_5[663:656];
        layer1[17][47:40] = buffer_data_5[671:664];
        layer1[17][55:48] = buffer_data_5[679:672];
        layer2[17][7:0] = buffer_data_4[631:624];
        layer2[17][15:8] = buffer_data_4[639:632];
        layer2[17][23:16] = buffer_data_4[647:640];
        layer2[17][31:24] = buffer_data_4[655:648];
        layer2[17][39:32] = buffer_data_4[663:656];
        layer2[17][47:40] = buffer_data_4[671:664];
        layer2[17][55:48] = buffer_data_4[679:672];
        layer3[17][7:0] = buffer_data_3[631:624];
        layer3[17][15:8] = buffer_data_3[639:632];
        layer3[17][23:16] = buffer_data_3[647:640];
        layer3[17][31:24] = buffer_data_3[655:648];
        layer3[17][39:32] = buffer_data_3[663:656];
        layer3[17][47:40] = buffer_data_3[671:664];
        layer3[17][55:48] = buffer_data_3[679:672];
        layer4[17][7:0] = buffer_data_2[631:624];
        layer4[17][15:8] = buffer_data_2[639:632];
        layer4[17][23:16] = buffer_data_2[647:640];
        layer4[17][31:24] = buffer_data_2[655:648];
        layer4[17][39:32] = buffer_data_2[663:656];
        layer4[17][47:40] = buffer_data_2[671:664];
        layer4[17][55:48] = buffer_data_2[679:672];
        layer5[17][7:0] = buffer_data_1[631:624];
        layer5[17][15:8] = buffer_data_1[639:632];
        layer5[17][23:16] = buffer_data_1[647:640];
        layer5[17][31:24] = buffer_data_1[655:648];
        layer5[17][39:32] = buffer_data_1[663:656];
        layer5[17][47:40] = buffer_data_1[671:664];
        layer5[17][55:48] = buffer_data_1[679:672];
        layer6[17][7:0] = buffer_data_0[631:624];
        layer6[17][15:8] = buffer_data_0[639:632];
        layer6[17][23:16] = buffer_data_0[647:640];
        layer6[17][31:24] = buffer_data_0[655:648];
        layer6[17][39:32] = buffer_data_0[663:656];
        layer6[17][47:40] = buffer_data_0[671:664];
        layer6[17][55:48] = buffer_data_0[679:672];
        layer0[18][7:0] = buffer_data_6[639:632];
        layer0[18][15:8] = buffer_data_6[647:640];
        layer0[18][23:16] = buffer_data_6[655:648];
        layer0[18][31:24] = buffer_data_6[663:656];
        layer0[18][39:32] = buffer_data_6[671:664];
        layer0[18][47:40] = buffer_data_6[679:672];
        layer0[18][55:48] = buffer_data_6[687:680];
        layer1[18][7:0] = buffer_data_5[639:632];
        layer1[18][15:8] = buffer_data_5[647:640];
        layer1[18][23:16] = buffer_data_5[655:648];
        layer1[18][31:24] = buffer_data_5[663:656];
        layer1[18][39:32] = buffer_data_5[671:664];
        layer1[18][47:40] = buffer_data_5[679:672];
        layer1[18][55:48] = buffer_data_5[687:680];
        layer2[18][7:0] = buffer_data_4[639:632];
        layer2[18][15:8] = buffer_data_4[647:640];
        layer2[18][23:16] = buffer_data_4[655:648];
        layer2[18][31:24] = buffer_data_4[663:656];
        layer2[18][39:32] = buffer_data_4[671:664];
        layer2[18][47:40] = buffer_data_4[679:672];
        layer2[18][55:48] = buffer_data_4[687:680];
        layer3[18][7:0] = buffer_data_3[639:632];
        layer3[18][15:8] = buffer_data_3[647:640];
        layer3[18][23:16] = buffer_data_3[655:648];
        layer3[18][31:24] = buffer_data_3[663:656];
        layer3[18][39:32] = buffer_data_3[671:664];
        layer3[18][47:40] = buffer_data_3[679:672];
        layer3[18][55:48] = buffer_data_3[687:680];
        layer4[18][7:0] = buffer_data_2[639:632];
        layer4[18][15:8] = buffer_data_2[647:640];
        layer4[18][23:16] = buffer_data_2[655:648];
        layer4[18][31:24] = buffer_data_2[663:656];
        layer4[18][39:32] = buffer_data_2[671:664];
        layer4[18][47:40] = buffer_data_2[679:672];
        layer4[18][55:48] = buffer_data_2[687:680];
        layer5[18][7:0] = buffer_data_1[639:632];
        layer5[18][15:8] = buffer_data_1[647:640];
        layer5[18][23:16] = buffer_data_1[655:648];
        layer5[18][31:24] = buffer_data_1[663:656];
        layer5[18][39:32] = buffer_data_1[671:664];
        layer5[18][47:40] = buffer_data_1[679:672];
        layer5[18][55:48] = buffer_data_1[687:680];
        layer6[18][7:0] = buffer_data_0[639:632];
        layer6[18][15:8] = buffer_data_0[647:640];
        layer6[18][23:16] = buffer_data_0[655:648];
        layer6[18][31:24] = buffer_data_0[663:656];
        layer6[18][39:32] = buffer_data_0[671:664];
        layer6[18][47:40] = buffer_data_0[679:672];
        layer6[18][55:48] = buffer_data_0[687:680];
        layer0[19][7:0] = buffer_data_6[647:640];
        layer0[19][15:8] = buffer_data_6[655:648];
        layer0[19][23:16] = buffer_data_6[663:656];
        layer0[19][31:24] = buffer_data_6[671:664];
        layer0[19][39:32] = buffer_data_6[679:672];
        layer0[19][47:40] = buffer_data_6[687:680];
        layer0[19][55:48] = buffer_data_6[695:688];
        layer1[19][7:0] = buffer_data_5[647:640];
        layer1[19][15:8] = buffer_data_5[655:648];
        layer1[19][23:16] = buffer_data_5[663:656];
        layer1[19][31:24] = buffer_data_5[671:664];
        layer1[19][39:32] = buffer_data_5[679:672];
        layer1[19][47:40] = buffer_data_5[687:680];
        layer1[19][55:48] = buffer_data_5[695:688];
        layer2[19][7:0] = buffer_data_4[647:640];
        layer2[19][15:8] = buffer_data_4[655:648];
        layer2[19][23:16] = buffer_data_4[663:656];
        layer2[19][31:24] = buffer_data_4[671:664];
        layer2[19][39:32] = buffer_data_4[679:672];
        layer2[19][47:40] = buffer_data_4[687:680];
        layer2[19][55:48] = buffer_data_4[695:688];
        layer3[19][7:0] = buffer_data_3[647:640];
        layer3[19][15:8] = buffer_data_3[655:648];
        layer3[19][23:16] = buffer_data_3[663:656];
        layer3[19][31:24] = buffer_data_3[671:664];
        layer3[19][39:32] = buffer_data_3[679:672];
        layer3[19][47:40] = buffer_data_3[687:680];
        layer3[19][55:48] = buffer_data_3[695:688];
        layer4[19][7:0] = buffer_data_2[647:640];
        layer4[19][15:8] = buffer_data_2[655:648];
        layer4[19][23:16] = buffer_data_2[663:656];
        layer4[19][31:24] = buffer_data_2[671:664];
        layer4[19][39:32] = buffer_data_2[679:672];
        layer4[19][47:40] = buffer_data_2[687:680];
        layer4[19][55:48] = buffer_data_2[695:688];
        layer5[19][7:0] = buffer_data_1[647:640];
        layer5[19][15:8] = buffer_data_1[655:648];
        layer5[19][23:16] = buffer_data_1[663:656];
        layer5[19][31:24] = buffer_data_1[671:664];
        layer5[19][39:32] = buffer_data_1[679:672];
        layer5[19][47:40] = buffer_data_1[687:680];
        layer5[19][55:48] = buffer_data_1[695:688];
        layer6[19][7:0] = buffer_data_0[647:640];
        layer6[19][15:8] = buffer_data_0[655:648];
        layer6[19][23:16] = buffer_data_0[663:656];
        layer6[19][31:24] = buffer_data_0[671:664];
        layer6[19][39:32] = buffer_data_0[679:672];
        layer6[19][47:40] = buffer_data_0[687:680];
        layer6[19][55:48] = buffer_data_0[695:688];
        layer0[20][7:0] = buffer_data_6[655:648];
        layer0[20][15:8] = buffer_data_6[663:656];
        layer0[20][23:16] = buffer_data_6[671:664];
        layer0[20][31:24] = buffer_data_6[679:672];
        layer0[20][39:32] = buffer_data_6[687:680];
        layer0[20][47:40] = buffer_data_6[695:688];
        layer0[20][55:48] = buffer_data_6[703:696];
        layer1[20][7:0] = buffer_data_5[655:648];
        layer1[20][15:8] = buffer_data_5[663:656];
        layer1[20][23:16] = buffer_data_5[671:664];
        layer1[20][31:24] = buffer_data_5[679:672];
        layer1[20][39:32] = buffer_data_5[687:680];
        layer1[20][47:40] = buffer_data_5[695:688];
        layer1[20][55:48] = buffer_data_5[703:696];
        layer2[20][7:0] = buffer_data_4[655:648];
        layer2[20][15:8] = buffer_data_4[663:656];
        layer2[20][23:16] = buffer_data_4[671:664];
        layer2[20][31:24] = buffer_data_4[679:672];
        layer2[20][39:32] = buffer_data_4[687:680];
        layer2[20][47:40] = buffer_data_4[695:688];
        layer2[20][55:48] = buffer_data_4[703:696];
        layer3[20][7:0] = buffer_data_3[655:648];
        layer3[20][15:8] = buffer_data_3[663:656];
        layer3[20][23:16] = buffer_data_3[671:664];
        layer3[20][31:24] = buffer_data_3[679:672];
        layer3[20][39:32] = buffer_data_3[687:680];
        layer3[20][47:40] = buffer_data_3[695:688];
        layer3[20][55:48] = buffer_data_3[703:696];
        layer4[20][7:0] = buffer_data_2[655:648];
        layer4[20][15:8] = buffer_data_2[663:656];
        layer4[20][23:16] = buffer_data_2[671:664];
        layer4[20][31:24] = buffer_data_2[679:672];
        layer4[20][39:32] = buffer_data_2[687:680];
        layer4[20][47:40] = buffer_data_2[695:688];
        layer4[20][55:48] = buffer_data_2[703:696];
        layer5[20][7:0] = buffer_data_1[655:648];
        layer5[20][15:8] = buffer_data_1[663:656];
        layer5[20][23:16] = buffer_data_1[671:664];
        layer5[20][31:24] = buffer_data_1[679:672];
        layer5[20][39:32] = buffer_data_1[687:680];
        layer5[20][47:40] = buffer_data_1[695:688];
        layer5[20][55:48] = buffer_data_1[703:696];
        layer6[20][7:0] = buffer_data_0[655:648];
        layer6[20][15:8] = buffer_data_0[663:656];
        layer6[20][23:16] = buffer_data_0[671:664];
        layer6[20][31:24] = buffer_data_0[679:672];
        layer6[20][39:32] = buffer_data_0[687:680];
        layer6[20][47:40] = buffer_data_0[695:688];
        layer6[20][55:48] = buffer_data_0[703:696];
        layer0[21][7:0] = buffer_data_6[663:656];
        layer0[21][15:8] = buffer_data_6[671:664];
        layer0[21][23:16] = buffer_data_6[679:672];
        layer0[21][31:24] = buffer_data_6[687:680];
        layer0[21][39:32] = buffer_data_6[695:688];
        layer0[21][47:40] = buffer_data_6[703:696];
        layer0[21][55:48] = buffer_data_6[711:704];
        layer1[21][7:0] = buffer_data_5[663:656];
        layer1[21][15:8] = buffer_data_5[671:664];
        layer1[21][23:16] = buffer_data_5[679:672];
        layer1[21][31:24] = buffer_data_5[687:680];
        layer1[21][39:32] = buffer_data_5[695:688];
        layer1[21][47:40] = buffer_data_5[703:696];
        layer1[21][55:48] = buffer_data_5[711:704];
        layer2[21][7:0] = buffer_data_4[663:656];
        layer2[21][15:8] = buffer_data_4[671:664];
        layer2[21][23:16] = buffer_data_4[679:672];
        layer2[21][31:24] = buffer_data_4[687:680];
        layer2[21][39:32] = buffer_data_4[695:688];
        layer2[21][47:40] = buffer_data_4[703:696];
        layer2[21][55:48] = buffer_data_4[711:704];
        layer3[21][7:0] = buffer_data_3[663:656];
        layer3[21][15:8] = buffer_data_3[671:664];
        layer3[21][23:16] = buffer_data_3[679:672];
        layer3[21][31:24] = buffer_data_3[687:680];
        layer3[21][39:32] = buffer_data_3[695:688];
        layer3[21][47:40] = buffer_data_3[703:696];
        layer3[21][55:48] = buffer_data_3[711:704];
        layer4[21][7:0] = buffer_data_2[663:656];
        layer4[21][15:8] = buffer_data_2[671:664];
        layer4[21][23:16] = buffer_data_2[679:672];
        layer4[21][31:24] = buffer_data_2[687:680];
        layer4[21][39:32] = buffer_data_2[695:688];
        layer4[21][47:40] = buffer_data_2[703:696];
        layer4[21][55:48] = buffer_data_2[711:704];
        layer5[21][7:0] = buffer_data_1[663:656];
        layer5[21][15:8] = buffer_data_1[671:664];
        layer5[21][23:16] = buffer_data_1[679:672];
        layer5[21][31:24] = buffer_data_1[687:680];
        layer5[21][39:32] = buffer_data_1[695:688];
        layer5[21][47:40] = buffer_data_1[703:696];
        layer5[21][55:48] = buffer_data_1[711:704];
        layer6[21][7:0] = buffer_data_0[663:656];
        layer6[21][15:8] = buffer_data_0[671:664];
        layer6[21][23:16] = buffer_data_0[679:672];
        layer6[21][31:24] = buffer_data_0[687:680];
        layer6[21][39:32] = buffer_data_0[695:688];
        layer6[21][47:40] = buffer_data_0[703:696];
        layer6[21][55:48] = buffer_data_0[711:704];
        layer0[22][7:0] = buffer_data_6[671:664];
        layer0[22][15:8] = buffer_data_6[679:672];
        layer0[22][23:16] = buffer_data_6[687:680];
        layer0[22][31:24] = buffer_data_6[695:688];
        layer0[22][39:32] = buffer_data_6[703:696];
        layer0[22][47:40] = buffer_data_6[711:704];
        layer0[22][55:48] = buffer_data_6[719:712];
        layer1[22][7:0] = buffer_data_5[671:664];
        layer1[22][15:8] = buffer_data_5[679:672];
        layer1[22][23:16] = buffer_data_5[687:680];
        layer1[22][31:24] = buffer_data_5[695:688];
        layer1[22][39:32] = buffer_data_5[703:696];
        layer1[22][47:40] = buffer_data_5[711:704];
        layer1[22][55:48] = buffer_data_5[719:712];
        layer2[22][7:0] = buffer_data_4[671:664];
        layer2[22][15:8] = buffer_data_4[679:672];
        layer2[22][23:16] = buffer_data_4[687:680];
        layer2[22][31:24] = buffer_data_4[695:688];
        layer2[22][39:32] = buffer_data_4[703:696];
        layer2[22][47:40] = buffer_data_4[711:704];
        layer2[22][55:48] = buffer_data_4[719:712];
        layer3[22][7:0] = buffer_data_3[671:664];
        layer3[22][15:8] = buffer_data_3[679:672];
        layer3[22][23:16] = buffer_data_3[687:680];
        layer3[22][31:24] = buffer_data_3[695:688];
        layer3[22][39:32] = buffer_data_3[703:696];
        layer3[22][47:40] = buffer_data_3[711:704];
        layer3[22][55:48] = buffer_data_3[719:712];
        layer4[22][7:0] = buffer_data_2[671:664];
        layer4[22][15:8] = buffer_data_2[679:672];
        layer4[22][23:16] = buffer_data_2[687:680];
        layer4[22][31:24] = buffer_data_2[695:688];
        layer4[22][39:32] = buffer_data_2[703:696];
        layer4[22][47:40] = buffer_data_2[711:704];
        layer4[22][55:48] = buffer_data_2[719:712];
        layer5[22][7:0] = buffer_data_1[671:664];
        layer5[22][15:8] = buffer_data_1[679:672];
        layer5[22][23:16] = buffer_data_1[687:680];
        layer5[22][31:24] = buffer_data_1[695:688];
        layer5[22][39:32] = buffer_data_1[703:696];
        layer5[22][47:40] = buffer_data_1[711:704];
        layer5[22][55:48] = buffer_data_1[719:712];
        layer6[22][7:0] = buffer_data_0[671:664];
        layer6[22][15:8] = buffer_data_0[679:672];
        layer6[22][23:16] = buffer_data_0[687:680];
        layer6[22][31:24] = buffer_data_0[695:688];
        layer6[22][39:32] = buffer_data_0[703:696];
        layer6[22][47:40] = buffer_data_0[711:704];
        layer6[22][55:48] = buffer_data_0[719:712];
        layer0[23][7:0] = buffer_data_6[679:672];
        layer0[23][15:8] = buffer_data_6[687:680];
        layer0[23][23:16] = buffer_data_6[695:688];
        layer0[23][31:24] = buffer_data_6[703:696];
        layer0[23][39:32] = buffer_data_6[711:704];
        layer0[23][47:40] = buffer_data_6[719:712];
        layer0[23][55:48] = buffer_data_6[727:720];
        layer1[23][7:0] = buffer_data_5[679:672];
        layer1[23][15:8] = buffer_data_5[687:680];
        layer1[23][23:16] = buffer_data_5[695:688];
        layer1[23][31:24] = buffer_data_5[703:696];
        layer1[23][39:32] = buffer_data_5[711:704];
        layer1[23][47:40] = buffer_data_5[719:712];
        layer1[23][55:48] = buffer_data_5[727:720];
        layer2[23][7:0] = buffer_data_4[679:672];
        layer2[23][15:8] = buffer_data_4[687:680];
        layer2[23][23:16] = buffer_data_4[695:688];
        layer2[23][31:24] = buffer_data_4[703:696];
        layer2[23][39:32] = buffer_data_4[711:704];
        layer2[23][47:40] = buffer_data_4[719:712];
        layer2[23][55:48] = buffer_data_4[727:720];
        layer3[23][7:0] = buffer_data_3[679:672];
        layer3[23][15:8] = buffer_data_3[687:680];
        layer3[23][23:16] = buffer_data_3[695:688];
        layer3[23][31:24] = buffer_data_3[703:696];
        layer3[23][39:32] = buffer_data_3[711:704];
        layer3[23][47:40] = buffer_data_3[719:712];
        layer3[23][55:48] = buffer_data_3[727:720];
        layer4[23][7:0] = buffer_data_2[679:672];
        layer4[23][15:8] = buffer_data_2[687:680];
        layer4[23][23:16] = buffer_data_2[695:688];
        layer4[23][31:24] = buffer_data_2[703:696];
        layer4[23][39:32] = buffer_data_2[711:704];
        layer4[23][47:40] = buffer_data_2[719:712];
        layer4[23][55:48] = buffer_data_2[727:720];
        layer5[23][7:0] = buffer_data_1[679:672];
        layer5[23][15:8] = buffer_data_1[687:680];
        layer5[23][23:16] = buffer_data_1[695:688];
        layer5[23][31:24] = buffer_data_1[703:696];
        layer5[23][39:32] = buffer_data_1[711:704];
        layer5[23][47:40] = buffer_data_1[719:712];
        layer5[23][55:48] = buffer_data_1[727:720];
        layer6[23][7:0] = buffer_data_0[679:672];
        layer6[23][15:8] = buffer_data_0[687:680];
        layer6[23][23:16] = buffer_data_0[695:688];
        layer6[23][31:24] = buffer_data_0[703:696];
        layer6[23][39:32] = buffer_data_0[711:704];
        layer6[23][47:40] = buffer_data_0[719:712];
        layer6[23][55:48] = buffer_data_0[727:720];
        layer0[24][7:0] = buffer_data_6[687:680];
        layer0[24][15:8] = buffer_data_6[695:688];
        layer0[24][23:16] = buffer_data_6[703:696];
        layer0[24][31:24] = buffer_data_6[711:704];
        layer0[24][39:32] = buffer_data_6[719:712];
        layer0[24][47:40] = buffer_data_6[727:720];
        layer0[24][55:48] = buffer_data_6[735:728];
        layer1[24][7:0] = buffer_data_5[687:680];
        layer1[24][15:8] = buffer_data_5[695:688];
        layer1[24][23:16] = buffer_data_5[703:696];
        layer1[24][31:24] = buffer_data_5[711:704];
        layer1[24][39:32] = buffer_data_5[719:712];
        layer1[24][47:40] = buffer_data_5[727:720];
        layer1[24][55:48] = buffer_data_5[735:728];
        layer2[24][7:0] = buffer_data_4[687:680];
        layer2[24][15:8] = buffer_data_4[695:688];
        layer2[24][23:16] = buffer_data_4[703:696];
        layer2[24][31:24] = buffer_data_4[711:704];
        layer2[24][39:32] = buffer_data_4[719:712];
        layer2[24][47:40] = buffer_data_4[727:720];
        layer2[24][55:48] = buffer_data_4[735:728];
        layer3[24][7:0] = buffer_data_3[687:680];
        layer3[24][15:8] = buffer_data_3[695:688];
        layer3[24][23:16] = buffer_data_3[703:696];
        layer3[24][31:24] = buffer_data_3[711:704];
        layer3[24][39:32] = buffer_data_3[719:712];
        layer3[24][47:40] = buffer_data_3[727:720];
        layer3[24][55:48] = buffer_data_3[735:728];
        layer4[24][7:0] = buffer_data_2[687:680];
        layer4[24][15:8] = buffer_data_2[695:688];
        layer4[24][23:16] = buffer_data_2[703:696];
        layer4[24][31:24] = buffer_data_2[711:704];
        layer4[24][39:32] = buffer_data_2[719:712];
        layer4[24][47:40] = buffer_data_2[727:720];
        layer4[24][55:48] = buffer_data_2[735:728];
        layer5[24][7:0] = buffer_data_1[687:680];
        layer5[24][15:8] = buffer_data_1[695:688];
        layer5[24][23:16] = buffer_data_1[703:696];
        layer5[24][31:24] = buffer_data_1[711:704];
        layer5[24][39:32] = buffer_data_1[719:712];
        layer5[24][47:40] = buffer_data_1[727:720];
        layer5[24][55:48] = buffer_data_1[735:728];
        layer6[24][7:0] = buffer_data_0[687:680];
        layer6[24][15:8] = buffer_data_0[695:688];
        layer6[24][23:16] = buffer_data_0[703:696];
        layer6[24][31:24] = buffer_data_0[711:704];
        layer6[24][39:32] = buffer_data_0[719:712];
        layer6[24][47:40] = buffer_data_0[727:720];
        layer6[24][55:48] = buffer_data_0[735:728];
        layer0[25][7:0] = buffer_data_6[695:688];
        layer0[25][15:8] = buffer_data_6[703:696];
        layer0[25][23:16] = buffer_data_6[711:704];
        layer0[25][31:24] = buffer_data_6[719:712];
        layer0[25][39:32] = buffer_data_6[727:720];
        layer0[25][47:40] = buffer_data_6[735:728];
        layer0[25][55:48] = buffer_data_6[743:736];
        layer1[25][7:0] = buffer_data_5[695:688];
        layer1[25][15:8] = buffer_data_5[703:696];
        layer1[25][23:16] = buffer_data_5[711:704];
        layer1[25][31:24] = buffer_data_5[719:712];
        layer1[25][39:32] = buffer_data_5[727:720];
        layer1[25][47:40] = buffer_data_5[735:728];
        layer1[25][55:48] = buffer_data_5[743:736];
        layer2[25][7:0] = buffer_data_4[695:688];
        layer2[25][15:8] = buffer_data_4[703:696];
        layer2[25][23:16] = buffer_data_4[711:704];
        layer2[25][31:24] = buffer_data_4[719:712];
        layer2[25][39:32] = buffer_data_4[727:720];
        layer2[25][47:40] = buffer_data_4[735:728];
        layer2[25][55:48] = buffer_data_4[743:736];
        layer3[25][7:0] = buffer_data_3[695:688];
        layer3[25][15:8] = buffer_data_3[703:696];
        layer3[25][23:16] = buffer_data_3[711:704];
        layer3[25][31:24] = buffer_data_3[719:712];
        layer3[25][39:32] = buffer_data_3[727:720];
        layer3[25][47:40] = buffer_data_3[735:728];
        layer3[25][55:48] = buffer_data_3[743:736];
        layer4[25][7:0] = buffer_data_2[695:688];
        layer4[25][15:8] = buffer_data_2[703:696];
        layer4[25][23:16] = buffer_data_2[711:704];
        layer4[25][31:24] = buffer_data_2[719:712];
        layer4[25][39:32] = buffer_data_2[727:720];
        layer4[25][47:40] = buffer_data_2[735:728];
        layer4[25][55:48] = buffer_data_2[743:736];
        layer5[25][7:0] = buffer_data_1[695:688];
        layer5[25][15:8] = buffer_data_1[703:696];
        layer5[25][23:16] = buffer_data_1[711:704];
        layer5[25][31:24] = buffer_data_1[719:712];
        layer5[25][39:32] = buffer_data_1[727:720];
        layer5[25][47:40] = buffer_data_1[735:728];
        layer5[25][55:48] = buffer_data_1[743:736];
        layer6[25][7:0] = buffer_data_0[695:688];
        layer6[25][15:8] = buffer_data_0[703:696];
        layer6[25][23:16] = buffer_data_0[711:704];
        layer6[25][31:24] = buffer_data_0[719:712];
        layer6[25][39:32] = buffer_data_0[727:720];
        layer6[25][47:40] = buffer_data_0[735:728];
        layer6[25][55:48] = buffer_data_0[743:736];
        layer0[26][7:0] = buffer_data_6[703:696];
        layer0[26][15:8] = buffer_data_6[711:704];
        layer0[26][23:16] = buffer_data_6[719:712];
        layer0[26][31:24] = buffer_data_6[727:720];
        layer0[26][39:32] = buffer_data_6[735:728];
        layer0[26][47:40] = buffer_data_6[743:736];
        layer0[26][55:48] = buffer_data_6[751:744];
        layer1[26][7:0] = buffer_data_5[703:696];
        layer1[26][15:8] = buffer_data_5[711:704];
        layer1[26][23:16] = buffer_data_5[719:712];
        layer1[26][31:24] = buffer_data_5[727:720];
        layer1[26][39:32] = buffer_data_5[735:728];
        layer1[26][47:40] = buffer_data_5[743:736];
        layer1[26][55:48] = buffer_data_5[751:744];
        layer2[26][7:0] = buffer_data_4[703:696];
        layer2[26][15:8] = buffer_data_4[711:704];
        layer2[26][23:16] = buffer_data_4[719:712];
        layer2[26][31:24] = buffer_data_4[727:720];
        layer2[26][39:32] = buffer_data_4[735:728];
        layer2[26][47:40] = buffer_data_4[743:736];
        layer2[26][55:48] = buffer_data_4[751:744];
        layer3[26][7:0] = buffer_data_3[703:696];
        layer3[26][15:8] = buffer_data_3[711:704];
        layer3[26][23:16] = buffer_data_3[719:712];
        layer3[26][31:24] = buffer_data_3[727:720];
        layer3[26][39:32] = buffer_data_3[735:728];
        layer3[26][47:40] = buffer_data_3[743:736];
        layer3[26][55:48] = buffer_data_3[751:744];
        layer4[26][7:0] = buffer_data_2[703:696];
        layer4[26][15:8] = buffer_data_2[711:704];
        layer4[26][23:16] = buffer_data_2[719:712];
        layer4[26][31:24] = buffer_data_2[727:720];
        layer4[26][39:32] = buffer_data_2[735:728];
        layer4[26][47:40] = buffer_data_2[743:736];
        layer4[26][55:48] = buffer_data_2[751:744];
        layer5[26][7:0] = buffer_data_1[703:696];
        layer5[26][15:8] = buffer_data_1[711:704];
        layer5[26][23:16] = buffer_data_1[719:712];
        layer5[26][31:24] = buffer_data_1[727:720];
        layer5[26][39:32] = buffer_data_1[735:728];
        layer5[26][47:40] = buffer_data_1[743:736];
        layer5[26][55:48] = buffer_data_1[751:744];
        layer6[26][7:0] = buffer_data_0[703:696];
        layer6[26][15:8] = buffer_data_0[711:704];
        layer6[26][23:16] = buffer_data_0[719:712];
        layer6[26][31:24] = buffer_data_0[727:720];
        layer6[26][39:32] = buffer_data_0[735:728];
        layer6[26][47:40] = buffer_data_0[743:736];
        layer6[26][55:48] = buffer_data_0[751:744];
        layer0[27][7:0] = buffer_data_6[711:704];
        layer0[27][15:8] = buffer_data_6[719:712];
        layer0[27][23:16] = buffer_data_6[727:720];
        layer0[27][31:24] = buffer_data_6[735:728];
        layer0[27][39:32] = buffer_data_6[743:736];
        layer0[27][47:40] = buffer_data_6[751:744];
        layer0[27][55:48] = buffer_data_6[759:752];
        layer1[27][7:0] = buffer_data_5[711:704];
        layer1[27][15:8] = buffer_data_5[719:712];
        layer1[27][23:16] = buffer_data_5[727:720];
        layer1[27][31:24] = buffer_data_5[735:728];
        layer1[27][39:32] = buffer_data_5[743:736];
        layer1[27][47:40] = buffer_data_5[751:744];
        layer1[27][55:48] = buffer_data_5[759:752];
        layer2[27][7:0] = buffer_data_4[711:704];
        layer2[27][15:8] = buffer_data_4[719:712];
        layer2[27][23:16] = buffer_data_4[727:720];
        layer2[27][31:24] = buffer_data_4[735:728];
        layer2[27][39:32] = buffer_data_4[743:736];
        layer2[27][47:40] = buffer_data_4[751:744];
        layer2[27][55:48] = buffer_data_4[759:752];
        layer3[27][7:0] = buffer_data_3[711:704];
        layer3[27][15:8] = buffer_data_3[719:712];
        layer3[27][23:16] = buffer_data_3[727:720];
        layer3[27][31:24] = buffer_data_3[735:728];
        layer3[27][39:32] = buffer_data_3[743:736];
        layer3[27][47:40] = buffer_data_3[751:744];
        layer3[27][55:48] = buffer_data_3[759:752];
        layer4[27][7:0] = buffer_data_2[711:704];
        layer4[27][15:8] = buffer_data_2[719:712];
        layer4[27][23:16] = buffer_data_2[727:720];
        layer4[27][31:24] = buffer_data_2[735:728];
        layer4[27][39:32] = buffer_data_2[743:736];
        layer4[27][47:40] = buffer_data_2[751:744];
        layer4[27][55:48] = buffer_data_2[759:752];
        layer5[27][7:0] = buffer_data_1[711:704];
        layer5[27][15:8] = buffer_data_1[719:712];
        layer5[27][23:16] = buffer_data_1[727:720];
        layer5[27][31:24] = buffer_data_1[735:728];
        layer5[27][39:32] = buffer_data_1[743:736];
        layer5[27][47:40] = buffer_data_1[751:744];
        layer5[27][55:48] = buffer_data_1[759:752];
        layer6[27][7:0] = buffer_data_0[711:704];
        layer6[27][15:8] = buffer_data_0[719:712];
        layer6[27][23:16] = buffer_data_0[727:720];
        layer6[27][31:24] = buffer_data_0[735:728];
        layer6[27][39:32] = buffer_data_0[743:736];
        layer6[27][47:40] = buffer_data_0[751:744];
        layer6[27][55:48] = buffer_data_0[759:752];
        layer0[28][7:0] = buffer_data_6[719:712];
        layer0[28][15:8] = buffer_data_6[727:720];
        layer0[28][23:16] = buffer_data_6[735:728];
        layer0[28][31:24] = buffer_data_6[743:736];
        layer0[28][39:32] = buffer_data_6[751:744];
        layer0[28][47:40] = buffer_data_6[759:752];
        layer0[28][55:48] = buffer_data_6[767:760];
        layer1[28][7:0] = buffer_data_5[719:712];
        layer1[28][15:8] = buffer_data_5[727:720];
        layer1[28][23:16] = buffer_data_5[735:728];
        layer1[28][31:24] = buffer_data_5[743:736];
        layer1[28][39:32] = buffer_data_5[751:744];
        layer1[28][47:40] = buffer_data_5[759:752];
        layer1[28][55:48] = buffer_data_5[767:760];
        layer2[28][7:0] = buffer_data_4[719:712];
        layer2[28][15:8] = buffer_data_4[727:720];
        layer2[28][23:16] = buffer_data_4[735:728];
        layer2[28][31:24] = buffer_data_4[743:736];
        layer2[28][39:32] = buffer_data_4[751:744];
        layer2[28][47:40] = buffer_data_4[759:752];
        layer2[28][55:48] = buffer_data_4[767:760];
        layer3[28][7:0] = buffer_data_3[719:712];
        layer3[28][15:8] = buffer_data_3[727:720];
        layer3[28][23:16] = buffer_data_3[735:728];
        layer3[28][31:24] = buffer_data_3[743:736];
        layer3[28][39:32] = buffer_data_3[751:744];
        layer3[28][47:40] = buffer_data_3[759:752];
        layer3[28][55:48] = buffer_data_3[767:760];
        layer4[28][7:0] = buffer_data_2[719:712];
        layer4[28][15:8] = buffer_data_2[727:720];
        layer4[28][23:16] = buffer_data_2[735:728];
        layer4[28][31:24] = buffer_data_2[743:736];
        layer4[28][39:32] = buffer_data_2[751:744];
        layer4[28][47:40] = buffer_data_2[759:752];
        layer4[28][55:48] = buffer_data_2[767:760];
        layer5[28][7:0] = buffer_data_1[719:712];
        layer5[28][15:8] = buffer_data_1[727:720];
        layer5[28][23:16] = buffer_data_1[735:728];
        layer5[28][31:24] = buffer_data_1[743:736];
        layer5[28][39:32] = buffer_data_1[751:744];
        layer5[28][47:40] = buffer_data_1[759:752];
        layer5[28][55:48] = buffer_data_1[767:760];
        layer6[28][7:0] = buffer_data_0[719:712];
        layer6[28][15:8] = buffer_data_0[727:720];
        layer6[28][23:16] = buffer_data_0[735:728];
        layer6[28][31:24] = buffer_data_0[743:736];
        layer6[28][39:32] = buffer_data_0[751:744];
        layer6[28][47:40] = buffer_data_0[759:752];
        layer6[28][55:48] = buffer_data_0[767:760];
        layer0[29][7:0] = buffer_data_6[727:720];
        layer0[29][15:8] = buffer_data_6[735:728];
        layer0[29][23:16] = buffer_data_6[743:736];
        layer0[29][31:24] = buffer_data_6[751:744];
        layer0[29][39:32] = buffer_data_6[759:752];
        layer0[29][47:40] = buffer_data_6[767:760];
        layer0[29][55:48] = buffer_data_6[775:768];
        layer1[29][7:0] = buffer_data_5[727:720];
        layer1[29][15:8] = buffer_data_5[735:728];
        layer1[29][23:16] = buffer_data_5[743:736];
        layer1[29][31:24] = buffer_data_5[751:744];
        layer1[29][39:32] = buffer_data_5[759:752];
        layer1[29][47:40] = buffer_data_5[767:760];
        layer1[29][55:48] = buffer_data_5[775:768];
        layer2[29][7:0] = buffer_data_4[727:720];
        layer2[29][15:8] = buffer_data_4[735:728];
        layer2[29][23:16] = buffer_data_4[743:736];
        layer2[29][31:24] = buffer_data_4[751:744];
        layer2[29][39:32] = buffer_data_4[759:752];
        layer2[29][47:40] = buffer_data_4[767:760];
        layer2[29][55:48] = buffer_data_4[775:768];
        layer3[29][7:0] = buffer_data_3[727:720];
        layer3[29][15:8] = buffer_data_3[735:728];
        layer3[29][23:16] = buffer_data_3[743:736];
        layer3[29][31:24] = buffer_data_3[751:744];
        layer3[29][39:32] = buffer_data_3[759:752];
        layer3[29][47:40] = buffer_data_3[767:760];
        layer3[29][55:48] = buffer_data_3[775:768];
        layer4[29][7:0] = buffer_data_2[727:720];
        layer4[29][15:8] = buffer_data_2[735:728];
        layer4[29][23:16] = buffer_data_2[743:736];
        layer4[29][31:24] = buffer_data_2[751:744];
        layer4[29][39:32] = buffer_data_2[759:752];
        layer4[29][47:40] = buffer_data_2[767:760];
        layer4[29][55:48] = buffer_data_2[775:768];
        layer5[29][7:0] = buffer_data_1[727:720];
        layer5[29][15:8] = buffer_data_1[735:728];
        layer5[29][23:16] = buffer_data_1[743:736];
        layer5[29][31:24] = buffer_data_1[751:744];
        layer5[29][39:32] = buffer_data_1[759:752];
        layer5[29][47:40] = buffer_data_1[767:760];
        layer5[29][55:48] = buffer_data_1[775:768];
        layer6[29][7:0] = buffer_data_0[727:720];
        layer6[29][15:8] = buffer_data_0[735:728];
        layer6[29][23:16] = buffer_data_0[743:736];
        layer6[29][31:24] = buffer_data_0[751:744];
        layer6[29][39:32] = buffer_data_0[759:752];
        layer6[29][47:40] = buffer_data_0[767:760];
        layer6[29][55:48] = buffer_data_0[775:768];
        layer0[30][7:0] = buffer_data_6[735:728];
        layer0[30][15:8] = buffer_data_6[743:736];
        layer0[30][23:16] = buffer_data_6[751:744];
        layer0[30][31:24] = buffer_data_6[759:752];
        layer0[30][39:32] = buffer_data_6[767:760];
        layer0[30][47:40] = buffer_data_6[775:768];
        layer0[30][55:48] = buffer_data_6[783:776];
        layer1[30][7:0] = buffer_data_5[735:728];
        layer1[30][15:8] = buffer_data_5[743:736];
        layer1[30][23:16] = buffer_data_5[751:744];
        layer1[30][31:24] = buffer_data_5[759:752];
        layer1[30][39:32] = buffer_data_5[767:760];
        layer1[30][47:40] = buffer_data_5[775:768];
        layer1[30][55:48] = buffer_data_5[783:776];
        layer2[30][7:0] = buffer_data_4[735:728];
        layer2[30][15:8] = buffer_data_4[743:736];
        layer2[30][23:16] = buffer_data_4[751:744];
        layer2[30][31:24] = buffer_data_4[759:752];
        layer2[30][39:32] = buffer_data_4[767:760];
        layer2[30][47:40] = buffer_data_4[775:768];
        layer2[30][55:48] = buffer_data_4[783:776];
        layer3[30][7:0] = buffer_data_3[735:728];
        layer3[30][15:8] = buffer_data_3[743:736];
        layer3[30][23:16] = buffer_data_3[751:744];
        layer3[30][31:24] = buffer_data_3[759:752];
        layer3[30][39:32] = buffer_data_3[767:760];
        layer3[30][47:40] = buffer_data_3[775:768];
        layer3[30][55:48] = buffer_data_3[783:776];
        layer4[30][7:0] = buffer_data_2[735:728];
        layer4[30][15:8] = buffer_data_2[743:736];
        layer4[30][23:16] = buffer_data_2[751:744];
        layer4[30][31:24] = buffer_data_2[759:752];
        layer4[30][39:32] = buffer_data_2[767:760];
        layer4[30][47:40] = buffer_data_2[775:768];
        layer4[30][55:48] = buffer_data_2[783:776];
        layer5[30][7:0] = buffer_data_1[735:728];
        layer5[30][15:8] = buffer_data_1[743:736];
        layer5[30][23:16] = buffer_data_1[751:744];
        layer5[30][31:24] = buffer_data_1[759:752];
        layer5[30][39:32] = buffer_data_1[767:760];
        layer5[30][47:40] = buffer_data_1[775:768];
        layer5[30][55:48] = buffer_data_1[783:776];
        layer6[30][7:0] = buffer_data_0[735:728];
        layer6[30][15:8] = buffer_data_0[743:736];
        layer6[30][23:16] = buffer_data_0[751:744];
        layer6[30][31:24] = buffer_data_0[759:752];
        layer6[30][39:32] = buffer_data_0[767:760];
        layer6[30][47:40] = buffer_data_0[775:768];
        layer6[30][55:48] = buffer_data_0[783:776];
        layer0[31][7:0] = buffer_data_6[743:736];
        layer0[31][15:8] = buffer_data_6[751:744];
        layer0[31][23:16] = buffer_data_6[759:752];
        layer0[31][31:24] = buffer_data_6[767:760];
        layer0[31][39:32] = buffer_data_6[775:768];
        layer0[31][47:40] = buffer_data_6[783:776];
        layer0[31][55:48] = buffer_data_6[791:784];
        layer1[31][7:0] = buffer_data_5[743:736];
        layer1[31][15:8] = buffer_data_5[751:744];
        layer1[31][23:16] = buffer_data_5[759:752];
        layer1[31][31:24] = buffer_data_5[767:760];
        layer1[31][39:32] = buffer_data_5[775:768];
        layer1[31][47:40] = buffer_data_5[783:776];
        layer1[31][55:48] = buffer_data_5[791:784];
        layer2[31][7:0] = buffer_data_4[743:736];
        layer2[31][15:8] = buffer_data_4[751:744];
        layer2[31][23:16] = buffer_data_4[759:752];
        layer2[31][31:24] = buffer_data_4[767:760];
        layer2[31][39:32] = buffer_data_4[775:768];
        layer2[31][47:40] = buffer_data_4[783:776];
        layer2[31][55:48] = buffer_data_4[791:784];
        layer3[31][7:0] = buffer_data_3[743:736];
        layer3[31][15:8] = buffer_data_3[751:744];
        layer3[31][23:16] = buffer_data_3[759:752];
        layer3[31][31:24] = buffer_data_3[767:760];
        layer3[31][39:32] = buffer_data_3[775:768];
        layer3[31][47:40] = buffer_data_3[783:776];
        layer3[31][55:48] = buffer_data_3[791:784];
        layer4[31][7:0] = buffer_data_2[743:736];
        layer4[31][15:8] = buffer_data_2[751:744];
        layer4[31][23:16] = buffer_data_2[759:752];
        layer4[31][31:24] = buffer_data_2[767:760];
        layer4[31][39:32] = buffer_data_2[775:768];
        layer4[31][47:40] = buffer_data_2[783:776];
        layer4[31][55:48] = buffer_data_2[791:784];
        layer5[31][7:0] = buffer_data_1[743:736];
        layer5[31][15:8] = buffer_data_1[751:744];
        layer5[31][23:16] = buffer_data_1[759:752];
        layer5[31][31:24] = buffer_data_1[767:760];
        layer5[31][39:32] = buffer_data_1[775:768];
        layer5[31][47:40] = buffer_data_1[783:776];
        layer5[31][55:48] = buffer_data_1[791:784];
        layer6[31][7:0] = buffer_data_0[743:736];
        layer6[31][15:8] = buffer_data_0[751:744];
        layer6[31][23:16] = buffer_data_0[759:752];
        layer6[31][31:24] = buffer_data_0[767:760];
        layer6[31][39:32] = buffer_data_0[775:768];
        layer6[31][47:40] = buffer_data_0[783:776];
        layer6[31][55:48] = buffer_data_0[791:784];
        layer0[32][7:0] = buffer_data_6[751:744];
        layer0[32][15:8] = buffer_data_6[759:752];
        layer0[32][23:16] = buffer_data_6[767:760];
        layer0[32][31:24] = buffer_data_6[775:768];
        layer0[32][39:32] = buffer_data_6[783:776];
        layer0[32][47:40] = buffer_data_6[791:784];
        layer0[32][55:48] = buffer_data_6[799:792];
        layer1[32][7:0] = buffer_data_5[751:744];
        layer1[32][15:8] = buffer_data_5[759:752];
        layer1[32][23:16] = buffer_data_5[767:760];
        layer1[32][31:24] = buffer_data_5[775:768];
        layer1[32][39:32] = buffer_data_5[783:776];
        layer1[32][47:40] = buffer_data_5[791:784];
        layer1[32][55:48] = buffer_data_5[799:792];
        layer2[32][7:0] = buffer_data_4[751:744];
        layer2[32][15:8] = buffer_data_4[759:752];
        layer2[32][23:16] = buffer_data_4[767:760];
        layer2[32][31:24] = buffer_data_4[775:768];
        layer2[32][39:32] = buffer_data_4[783:776];
        layer2[32][47:40] = buffer_data_4[791:784];
        layer2[32][55:48] = buffer_data_4[799:792];
        layer3[32][7:0] = buffer_data_3[751:744];
        layer3[32][15:8] = buffer_data_3[759:752];
        layer3[32][23:16] = buffer_data_3[767:760];
        layer3[32][31:24] = buffer_data_3[775:768];
        layer3[32][39:32] = buffer_data_3[783:776];
        layer3[32][47:40] = buffer_data_3[791:784];
        layer3[32][55:48] = buffer_data_3[799:792];
        layer4[32][7:0] = buffer_data_2[751:744];
        layer4[32][15:8] = buffer_data_2[759:752];
        layer4[32][23:16] = buffer_data_2[767:760];
        layer4[32][31:24] = buffer_data_2[775:768];
        layer4[32][39:32] = buffer_data_2[783:776];
        layer4[32][47:40] = buffer_data_2[791:784];
        layer4[32][55:48] = buffer_data_2[799:792];
        layer5[32][7:0] = buffer_data_1[751:744];
        layer5[32][15:8] = buffer_data_1[759:752];
        layer5[32][23:16] = buffer_data_1[767:760];
        layer5[32][31:24] = buffer_data_1[775:768];
        layer5[32][39:32] = buffer_data_1[783:776];
        layer5[32][47:40] = buffer_data_1[791:784];
        layer5[32][55:48] = buffer_data_1[799:792];
        layer6[32][7:0] = buffer_data_0[751:744];
        layer6[32][15:8] = buffer_data_0[759:752];
        layer6[32][23:16] = buffer_data_0[767:760];
        layer6[32][31:24] = buffer_data_0[775:768];
        layer6[32][39:32] = buffer_data_0[783:776];
        layer6[32][47:40] = buffer_data_0[791:784];
        layer6[32][55:48] = buffer_data_0[799:792];
        layer0[33][7:0] = buffer_data_6[759:752];
        layer0[33][15:8] = buffer_data_6[767:760];
        layer0[33][23:16] = buffer_data_6[775:768];
        layer0[33][31:24] = buffer_data_6[783:776];
        layer0[33][39:32] = buffer_data_6[791:784];
        layer0[33][47:40] = buffer_data_6[799:792];
        layer0[33][55:48] = buffer_data_6[807:800];
        layer1[33][7:0] = buffer_data_5[759:752];
        layer1[33][15:8] = buffer_data_5[767:760];
        layer1[33][23:16] = buffer_data_5[775:768];
        layer1[33][31:24] = buffer_data_5[783:776];
        layer1[33][39:32] = buffer_data_5[791:784];
        layer1[33][47:40] = buffer_data_5[799:792];
        layer1[33][55:48] = buffer_data_5[807:800];
        layer2[33][7:0] = buffer_data_4[759:752];
        layer2[33][15:8] = buffer_data_4[767:760];
        layer2[33][23:16] = buffer_data_4[775:768];
        layer2[33][31:24] = buffer_data_4[783:776];
        layer2[33][39:32] = buffer_data_4[791:784];
        layer2[33][47:40] = buffer_data_4[799:792];
        layer2[33][55:48] = buffer_data_4[807:800];
        layer3[33][7:0] = buffer_data_3[759:752];
        layer3[33][15:8] = buffer_data_3[767:760];
        layer3[33][23:16] = buffer_data_3[775:768];
        layer3[33][31:24] = buffer_data_3[783:776];
        layer3[33][39:32] = buffer_data_3[791:784];
        layer3[33][47:40] = buffer_data_3[799:792];
        layer3[33][55:48] = buffer_data_3[807:800];
        layer4[33][7:0] = buffer_data_2[759:752];
        layer4[33][15:8] = buffer_data_2[767:760];
        layer4[33][23:16] = buffer_data_2[775:768];
        layer4[33][31:24] = buffer_data_2[783:776];
        layer4[33][39:32] = buffer_data_2[791:784];
        layer4[33][47:40] = buffer_data_2[799:792];
        layer4[33][55:48] = buffer_data_2[807:800];
        layer5[33][7:0] = buffer_data_1[759:752];
        layer5[33][15:8] = buffer_data_1[767:760];
        layer5[33][23:16] = buffer_data_1[775:768];
        layer5[33][31:24] = buffer_data_1[783:776];
        layer5[33][39:32] = buffer_data_1[791:784];
        layer5[33][47:40] = buffer_data_1[799:792];
        layer5[33][55:48] = buffer_data_1[807:800];
        layer6[33][7:0] = buffer_data_0[759:752];
        layer6[33][15:8] = buffer_data_0[767:760];
        layer6[33][23:16] = buffer_data_0[775:768];
        layer6[33][31:24] = buffer_data_0[783:776];
        layer6[33][39:32] = buffer_data_0[791:784];
        layer6[33][47:40] = buffer_data_0[799:792];
        layer6[33][55:48] = buffer_data_0[807:800];
        layer0[34][7:0] = buffer_data_6[767:760];
        layer0[34][15:8] = buffer_data_6[775:768];
        layer0[34][23:16] = buffer_data_6[783:776];
        layer0[34][31:24] = buffer_data_6[791:784];
        layer0[34][39:32] = buffer_data_6[799:792];
        layer0[34][47:40] = buffer_data_6[807:800];
        layer0[34][55:48] = buffer_data_6[815:808];
        layer1[34][7:0] = buffer_data_5[767:760];
        layer1[34][15:8] = buffer_data_5[775:768];
        layer1[34][23:16] = buffer_data_5[783:776];
        layer1[34][31:24] = buffer_data_5[791:784];
        layer1[34][39:32] = buffer_data_5[799:792];
        layer1[34][47:40] = buffer_data_5[807:800];
        layer1[34][55:48] = buffer_data_5[815:808];
        layer2[34][7:0] = buffer_data_4[767:760];
        layer2[34][15:8] = buffer_data_4[775:768];
        layer2[34][23:16] = buffer_data_4[783:776];
        layer2[34][31:24] = buffer_data_4[791:784];
        layer2[34][39:32] = buffer_data_4[799:792];
        layer2[34][47:40] = buffer_data_4[807:800];
        layer2[34][55:48] = buffer_data_4[815:808];
        layer3[34][7:0] = buffer_data_3[767:760];
        layer3[34][15:8] = buffer_data_3[775:768];
        layer3[34][23:16] = buffer_data_3[783:776];
        layer3[34][31:24] = buffer_data_3[791:784];
        layer3[34][39:32] = buffer_data_3[799:792];
        layer3[34][47:40] = buffer_data_3[807:800];
        layer3[34][55:48] = buffer_data_3[815:808];
        layer4[34][7:0] = buffer_data_2[767:760];
        layer4[34][15:8] = buffer_data_2[775:768];
        layer4[34][23:16] = buffer_data_2[783:776];
        layer4[34][31:24] = buffer_data_2[791:784];
        layer4[34][39:32] = buffer_data_2[799:792];
        layer4[34][47:40] = buffer_data_2[807:800];
        layer4[34][55:48] = buffer_data_2[815:808];
        layer5[34][7:0] = buffer_data_1[767:760];
        layer5[34][15:8] = buffer_data_1[775:768];
        layer5[34][23:16] = buffer_data_1[783:776];
        layer5[34][31:24] = buffer_data_1[791:784];
        layer5[34][39:32] = buffer_data_1[799:792];
        layer5[34][47:40] = buffer_data_1[807:800];
        layer5[34][55:48] = buffer_data_1[815:808];
        layer6[34][7:0] = buffer_data_0[767:760];
        layer6[34][15:8] = buffer_data_0[775:768];
        layer6[34][23:16] = buffer_data_0[783:776];
        layer6[34][31:24] = buffer_data_0[791:784];
        layer6[34][39:32] = buffer_data_0[799:792];
        layer6[34][47:40] = buffer_data_0[807:800];
        layer6[34][55:48] = buffer_data_0[815:808];
        layer0[35][7:0] = buffer_data_6[775:768];
        layer0[35][15:8] = buffer_data_6[783:776];
        layer0[35][23:16] = buffer_data_6[791:784];
        layer0[35][31:24] = buffer_data_6[799:792];
        layer0[35][39:32] = buffer_data_6[807:800];
        layer0[35][47:40] = buffer_data_6[815:808];
        layer0[35][55:48] = buffer_data_6[823:816];
        layer1[35][7:0] = buffer_data_5[775:768];
        layer1[35][15:8] = buffer_data_5[783:776];
        layer1[35][23:16] = buffer_data_5[791:784];
        layer1[35][31:24] = buffer_data_5[799:792];
        layer1[35][39:32] = buffer_data_5[807:800];
        layer1[35][47:40] = buffer_data_5[815:808];
        layer1[35][55:48] = buffer_data_5[823:816];
        layer2[35][7:0] = buffer_data_4[775:768];
        layer2[35][15:8] = buffer_data_4[783:776];
        layer2[35][23:16] = buffer_data_4[791:784];
        layer2[35][31:24] = buffer_data_4[799:792];
        layer2[35][39:32] = buffer_data_4[807:800];
        layer2[35][47:40] = buffer_data_4[815:808];
        layer2[35][55:48] = buffer_data_4[823:816];
        layer3[35][7:0] = buffer_data_3[775:768];
        layer3[35][15:8] = buffer_data_3[783:776];
        layer3[35][23:16] = buffer_data_3[791:784];
        layer3[35][31:24] = buffer_data_3[799:792];
        layer3[35][39:32] = buffer_data_3[807:800];
        layer3[35][47:40] = buffer_data_3[815:808];
        layer3[35][55:48] = buffer_data_3[823:816];
        layer4[35][7:0] = buffer_data_2[775:768];
        layer4[35][15:8] = buffer_data_2[783:776];
        layer4[35][23:16] = buffer_data_2[791:784];
        layer4[35][31:24] = buffer_data_2[799:792];
        layer4[35][39:32] = buffer_data_2[807:800];
        layer4[35][47:40] = buffer_data_2[815:808];
        layer4[35][55:48] = buffer_data_2[823:816];
        layer5[35][7:0] = buffer_data_1[775:768];
        layer5[35][15:8] = buffer_data_1[783:776];
        layer5[35][23:16] = buffer_data_1[791:784];
        layer5[35][31:24] = buffer_data_1[799:792];
        layer5[35][39:32] = buffer_data_1[807:800];
        layer5[35][47:40] = buffer_data_1[815:808];
        layer5[35][55:48] = buffer_data_1[823:816];
        layer6[35][7:0] = buffer_data_0[775:768];
        layer6[35][15:8] = buffer_data_0[783:776];
        layer6[35][23:16] = buffer_data_0[791:784];
        layer6[35][31:24] = buffer_data_0[799:792];
        layer6[35][39:32] = buffer_data_0[807:800];
        layer6[35][47:40] = buffer_data_0[815:808];
        layer6[35][55:48] = buffer_data_0[823:816];
        layer0[36][7:0] = buffer_data_6[783:776];
        layer0[36][15:8] = buffer_data_6[791:784];
        layer0[36][23:16] = buffer_data_6[799:792];
        layer0[36][31:24] = buffer_data_6[807:800];
        layer0[36][39:32] = buffer_data_6[815:808];
        layer0[36][47:40] = buffer_data_6[823:816];
        layer0[36][55:48] = buffer_data_6[831:824];
        layer1[36][7:0] = buffer_data_5[783:776];
        layer1[36][15:8] = buffer_data_5[791:784];
        layer1[36][23:16] = buffer_data_5[799:792];
        layer1[36][31:24] = buffer_data_5[807:800];
        layer1[36][39:32] = buffer_data_5[815:808];
        layer1[36][47:40] = buffer_data_5[823:816];
        layer1[36][55:48] = buffer_data_5[831:824];
        layer2[36][7:0] = buffer_data_4[783:776];
        layer2[36][15:8] = buffer_data_4[791:784];
        layer2[36][23:16] = buffer_data_4[799:792];
        layer2[36][31:24] = buffer_data_4[807:800];
        layer2[36][39:32] = buffer_data_4[815:808];
        layer2[36][47:40] = buffer_data_4[823:816];
        layer2[36][55:48] = buffer_data_4[831:824];
        layer3[36][7:0] = buffer_data_3[783:776];
        layer3[36][15:8] = buffer_data_3[791:784];
        layer3[36][23:16] = buffer_data_3[799:792];
        layer3[36][31:24] = buffer_data_3[807:800];
        layer3[36][39:32] = buffer_data_3[815:808];
        layer3[36][47:40] = buffer_data_3[823:816];
        layer3[36][55:48] = buffer_data_3[831:824];
        layer4[36][7:0] = buffer_data_2[783:776];
        layer4[36][15:8] = buffer_data_2[791:784];
        layer4[36][23:16] = buffer_data_2[799:792];
        layer4[36][31:24] = buffer_data_2[807:800];
        layer4[36][39:32] = buffer_data_2[815:808];
        layer4[36][47:40] = buffer_data_2[823:816];
        layer4[36][55:48] = buffer_data_2[831:824];
        layer5[36][7:0] = buffer_data_1[783:776];
        layer5[36][15:8] = buffer_data_1[791:784];
        layer5[36][23:16] = buffer_data_1[799:792];
        layer5[36][31:24] = buffer_data_1[807:800];
        layer5[36][39:32] = buffer_data_1[815:808];
        layer5[36][47:40] = buffer_data_1[823:816];
        layer5[36][55:48] = buffer_data_1[831:824];
        layer6[36][7:0] = buffer_data_0[783:776];
        layer6[36][15:8] = buffer_data_0[791:784];
        layer6[36][23:16] = buffer_data_0[799:792];
        layer6[36][31:24] = buffer_data_0[807:800];
        layer6[36][39:32] = buffer_data_0[815:808];
        layer6[36][47:40] = buffer_data_0[823:816];
        layer6[36][55:48] = buffer_data_0[831:824];
        layer0[37][7:0] = buffer_data_6[791:784];
        layer0[37][15:8] = buffer_data_6[799:792];
        layer0[37][23:16] = buffer_data_6[807:800];
        layer0[37][31:24] = buffer_data_6[815:808];
        layer0[37][39:32] = buffer_data_6[823:816];
        layer0[37][47:40] = buffer_data_6[831:824];
        layer0[37][55:48] = buffer_data_6[839:832];
        layer1[37][7:0] = buffer_data_5[791:784];
        layer1[37][15:8] = buffer_data_5[799:792];
        layer1[37][23:16] = buffer_data_5[807:800];
        layer1[37][31:24] = buffer_data_5[815:808];
        layer1[37][39:32] = buffer_data_5[823:816];
        layer1[37][47:40] = buffer_data_5[831:824];
        layer1[37][55:48] = buffer_data_5[839:832];
        layer2[37][7:0] = buffer_data_4[791:784];
        layer2[37][15:8] = buffer_data_4[799:792];
        layer2[37][23:16] = buffer_data_4[807:800];
        layer2[37][31:24] = buffer_data_4[815:808];
        layer2[37][39:32] = buffer_data_4[823:816];
        layer2[37][47:40] = buffer_data_4[831:824];
        layer2[37][55:48] = buffer_data_4[839:832];
        layer3[37][7:0] = buffer_data_3[791:784];
        layer3[37][15:8] = buffer_data_3[799:792];
        layer3[37][23:16] = buffer_data_3[807:800];
        layer3[37][31:24] = buffer_data_3[815:808];
        layer3[37][39:32] = buffer_data_3[823:816];
        layer3[37][47:40] = buffer_data_3[831:824];
        layer3[37][55:48] = buffer_data_3[839:832];
        layer4[37][7:0] = buffer_data_2[791:784];
        layer4[37][15:8] = buffer_data_2[799:792];
        layer4[37][23:16] = buffer_data_2[807:800];
        layer4[37][31:24] = buffer_data_2[815:808];
        layer4[37][39:32] = buffer_data_2[823:816];
        layer4[37][47:40] = buffer_data_2[831:824];
        layer4[37][55:48] = buffer_data_2[839:832];
        layer5[37][7:0] = buffer_data_1[791:784];
        layer5[37][15:8] = buffer_data_1[799:792];
        layer5[37][23:16] = buffer_data_1[807:800];
        layer5[37][31:24] = buffer_data_1[815:808];
        layer5[37][39:32] = buffer_data_1[823:816];
        layer5[37][47:40] = buffer_data_1[831:824];
        layer5[37][55:48] = buffer_data_1[839:832];
        layer6[37][7:0] = buffer_data_0[791:784];
        layer6[37][15:8] = buffer_data_0[799:792];
        layer6[37][23:16] = buffer_data_0[807:800];
        layer6[37][31:24] = buffer_data_0[815:808];
        layer6[37][39:32] = buffer_data_0[823:816];
        layer6[37][47:40] = buffer_data_0[831:824];
        layer6[37][55:48] = buffer_data_0[839:832];
        layer0[38][7:0] = buffer_data_6[799:792];
        layer0[38][15:8] = buffer_data_6[807:800];
        layer0[38][23:16] = buffer_data_6[815:808];
        layer0[38][31:24] = buffer_data_6[823:816];
        layer0[38][39:32] = buffer_data_6[831:824];
        layer0[38][47:40] = buffer_data_6[839:832];
        layer0[38][55:48] = buffer_data_6[847:840];
        layer1[38][7:0] = buffer_data_5[799:792];
        layer1[38][15:8] = buffer_data_5[807:800];
        layer1[38][23:16] = buffer_data_5[815:808];
        layer1[38][31:24] = buffer_data_5[823:816];
        layer1[38][39:32] = buffer_data_5[831:824];
        layer1[38][47:40] = buffer_data_5[839:832];
        layer1[38][55:48] = buffer_data_5[847:840];
        layer2[38][7:0] = buffer_data_4[799:792];
        layer2[38][15:8] = buffer_data_4[807:800];
        layer2[38][23:16] = buffer_data_4[815:808];
        layer2[38][31:24] = buffer_data_4[823:816];
        layer2[38][39:32] = buffer_data_4[831:824];
        layer2[38][47:40] = buffer_data_4[839:832];
        layer2[38][55:48] = buffer_data_4[847:840];
        layer3[38][7:0] = buffer_data_3[799:792];
        layer3[38][15:8] = buffer_data_3[807:800];
        layer3[38][23:16] = buffer_data_3[815:808];
        layer3[38][31:24] = buffer_data_3[823:816];
        layer3[38][39:32] = buffer_data_3[831:824];
        layer3[38][47:40] = buffer_data_3[839:832];
        layer3[38][55:48] = buffer_data_3[847:840];
        layer4[38][7:0] = buffer_data_2[799:792];
        layer4[38][15:8] = buffer_data_2[807:800];
        layer4[38][23:16] = buffer_data_2[815:808];
        layer4[38][31:24] = buffer_data_2[823:816];
        layer4[38][39:32] = buffer_data_2[831:824];
        layer4[38][47:40] = buffer_data_2[839:832];
        layer4[38][55:48] = buffer_data_2[847:840];
        layer5[38][7:0] = buffer_data_1[799:792];
        layer5[38][15:8] = buffer_data_1[807:800];
        layer5[38][23:16] = buffer_data_1[815:808];
        layer5[38][31:24] = buffer_data_1[823:816];
        layer5[38][39:32] = buffer_data_1[831:824];
        layer5[38][47:40] = buffer_data_1[839:832];
        layer5[38][55:48] = buffer_data_1[847:840];
        layer6[38][7:0] = buffer_data_0[799:792];
        layer6[38][15:8] = buffer_data_0[807:800];
        layer6[38][23:16] = buffer_data_0[815:808];
        layer6[38][31:24] = buffer_data_0[823:816];
        layer6[38][39:32] = buffer_data_0[831:824];
        layer6[38][47:40] = buffer_data_0[839:832];
        layer6[38][55:48] = buffer_data_0[847:840];
        layer0[39][7:0] = buffer_data_6[807:800];
        layer0[39][15:8] = buffer_data_6[815:808];
        layer0[39][23:16] = buffer_data_6[823:816];
        layer0[39][31:24] = buffer_data_6[831:824];
        layer0[39][39:32] = buffer_data_6[839:832];
        layer0[39][47:40] = buffer_data_6[847:840];
        layer0[39][55:48] = buffer_data_6[855:848];
        layer1[39][7:0] = buffer_data_5[807:800];
        layer1[39][15:8] = buffer_data_5[815:808];
        layer1[39][23:16] = buffer_data_5[823:816];
        layer1[39][31:24] = buffer_data_5[831:824];
        layer1[39][39:32] = buffer_data_5[839:832];
        layer1[39][47:40] = buffer_data_5[847:840];
        layer1[39][55:48] = buffer_data_5[855:848];
        layer2[39][7:0] = buffer_data_4[807:800];
        layer2[39][15:8] = buffer_data_4[815:808];
        layer2[39][23:16] = buffer_data_4[823:816];
        layer2[39][31:24] = buffer_data_4[831:824];
        layer2[39][39:32] = buffer_data_4[839:832];
        layer2[39][47:40] = buffer_data_4[847:840];
        layer2[39][55:48] = buffer_data_4[855:848];
        layer3[39][7:0] = buffer_data_3[807:800];
        layer3[39][15:8] = buffer_data_3[815:808];
        layer3[39][23:16] = buffer_data_3[823:816];
        layer3[39][31:24] = buffer_data_3[831:824];
        layer3[39][39:32] = buffer_data_3[839:832];
        layer3[39][47:40] = buffer_data_3[847:840];
        layer3[39][55:48] = buffer_data_3[855:848];
        layer4[39][7:0] = buffer_data_2[807:800];
        layer4[39][15:8] = buffer_data_2[815:808];
        layer4[39][23:16] = buffer_data_2[823:816];
        layer4[39][31:24] = buffer_data_2[831:824];
        layer4[39][39:32] = buffer_data_2[839:832];
        layer4[39][47:40] = buffer_data_2[847:840];
        layer4[39][55:48] = buffer_data_2[855:848];
        layer5[39][7:0] = buffer_data_1[807:800];
        layer5[39][15:8] = buffer_data_1[815:808];
        layer5[39][23:16] = buffer_data_1[823:816];
        layer5[39][31:24] = buffer_data_1[831:824];
        layer5[39][39:32] = buffer_data_1[839:832];
        layer5[39][47:40] = buffer_data_1[847:840];
        layer5[39][55:48] = buffer_data_1[855:848];
        layer6[39][7:0] = buffer_data_0[807:800];
        layer6[39][15:8] = buffer_data_0[815:808];
        layer6[39][23:16] = buffer_data_0[823:816];
        layer6[39][31:24] = buffer_data_0[831:824];
        layer6[39][39:32] = buffer_data_0[839:832];
        layer6[39][47:40] = buffer_data_0[847:840];
        layer6[39][55:48] = buffer_data_0[855:848];
        layer0[40][7:0] = buffer_data_6[815:808];
        layer0[40][15:8] = buffer_data_6[823:816];
        layer0[40][23:16] = buffer_data_6[831:824];
        layer0[40][31:24] = buffer_data_6[839:832];
        layer0[40][39:32] = buffer_data_6[847:840];
        layer0[40][47:40] = buffer_data_6[855:848];
        layer0[40][55:48] = buffer_data_6[863:856];
        layer1[40][7:0] = buffer_data_5[815:808];
        layer1[40][15:8] = buffer_data_5[823:816];
        layer1[40][23:16] = buffer_data_5[831:824];
        layer1[40][31:24] = buffer_data_5[839:832];
        layer1[40][39:32] = buffer_data_5[847:840];
        layer1[40][47:40] = buffer_data_5[855:848];
        layer1[40][55:48] = buffer_data_5[863:856];
        layer2[40][7:0] = buffer_data_4[815:808];
        layer2[40][15:8] = buffer_data_4[823:816];
        layer2[40][23:16] = buffer_data_4[831:824];
        layer2[40][31:24] = buffer_data_4[839:832];
        layer2[40][39:32] = buffer_data_4[847:840];
        layer2[40][47:40] = buffer_data_4[855:848];
        layer2[40][55:48] = buffer_data_4[863:856];
        layer3[40][7:0] = buffer_data_3[815:808];
        layer3[40][15:8] = buffer_data_3[823:816];
        layer3[40][23:16] = buffer_data_3[831:824];
        layer3[40][31:24] = buffer_data_3[839:832];
        layer3[40][39:32] = buffer_data_3[847:840];
        layer3[40][47:40] = buffer_data_3[855:848];
        layer3[40][55:48] = buffer_data_3[863:856];
        layer4[40][7:0] = buffer_data_2[815:808];
        layer4[40][15:8] = buffer_data_2[823:816];
        layer4[40][23:16] = buffer_data_2[831:824];
        layer4[40][31:24] = buffer_data_2[839:832];
        layer4[40][39:32] = buffer_data_2[847:840];
        layer4[40][47:40] = buffer_data_2[855:848];
        layer4[40][55:48] = buffer_data_2[863:856];
        layer5[40][7:0] = buffer_data_1[815:808];
        layer5[40][15:8] = buffer_data_1[823:816];
        layer5[40][23:16] = buffer_data_1[831:824];
        layer5[40][31:24] = buffer_data_1[839:832];
        layer5[40][39:32] = buffer_data_1[847:840];
        layer5[40][47:40] = buffer_data_1[855:848];
        layer5[40][55:48] = buffer_data_1[863:856];
        layer6[40][7:0] = buffer_data_0[815:808];
        layer6[40][15:8] = buffer_data_0[823:816];
        layer6[40][23:16] = buffer_data_0[831:824];
        layer6[40][31:24] = buffer_data_0[839:832];
        layer6[40][39:32] = buffer_data_0[847:840];
        layer6[40][47:40] = buffer_data_0[855:848];
        layer6[40][55:48] = buffer_data_0[863:856];
        layer0[41][7:0] = buffer_data_6[823:816];
        layer0[41][15:8] = buffer_data_6[831:824];
        layer0[41][23:16] = buffer_data_6[839:832];
        layer0[41][31:24] = buffer_data_6[847:840];
        layer0[41][39:32] = buffer_data_6[855:848];
        layer0[41][47:40] = buffer_data_6[863:856];
        layer0[41][55:48] = buffer_data_6[871:864];
        layer1[41][7:0] = buffer_data_5[823:816];
        layer1[41][15:8] = buffer_data_5[831:824];
        layer1[41][23:16] = buffer_data_5[839:832];
        layer1[41][31:24] = buffer_data_5[847:840];
        layer1[41][39:32] = buffer_data_5[855:848];
        layer1[41][47:40] = buffer_data_5[863:856];
        layer1[41][55:48] = buffer_data_5[871:864];
        layer2[41][7:0] = buffer_data_4[823:816];
        layer2[41][15:8] = buffer_data_4[831:824];
        layer2[41][23:16] = buffer_data_4[839:832];
        layer2[41][31:24] = buffer_data_4[847:840];
        layer2[41][39:32] = buffer_data_4[855:848];
        layer2[41][47:40] = buffer_data_4[863:856];
        layer2[41][55:48] = buffer_data_4[871:864];
        layer3[41][7:0] = buffer_data_3[823:816];
        layer3[41][15:8] = buffer_data_3[831:824];
        layer3[41][23:16] = buffer_data_3[839:832];
        layer3[41][31:24] = buffer_data_3[847:840];
        layer3[41][39:32] = buffer_data_3[855:848];
        layer3[41][47:40] = buffer_data_3[863:856];
        layer3[41][55:48] = buffer_data_3[871:864];
        layer4[41][7:0] = buffer_data_2[823:816];
        layer4[41][15:8] = buffer_data_2[831:824];
        layer4[41][23:16] = buffer_data_2[839:832];
        layer4[41][31:24] = buffer_data_2[847:840];
        layer4[41][39:32] = buffer_data_2[855:848];
        layer4[41][47:40] = buffer_data_2[863:856];
        layer4[41][55:48] = buffer_data_2[871:864];
        layer5[41][7:0] = buffer_data_1[823:816];
        layer5[41][15:8] = buffer_data_1[831:824];
        layer5[41][23:16] = buffer_data_1[839:832];
        layer5[41][31:24] = buffer_data_1[847:840];
        layer5[41][39:32] = buffer_data_1[855:848];
        layer5[41][47:40] = buffer_data_1[863:856];
        layer5[41][55:48] = buffer_data_1[871:864];
        layer6[41][7:0] = buffer_data_0[823:816];
        layer6[41][15:8] = buffer_data_0[831:824];
        layer6[41][23:16] = buffer_data_0[839:832];
        layer6[41][31:24] = buffer_data_0[847:840];
        layer6[41][39:32] = buffer_data_0[855:848];
        layer6[41][47:40] = buffer_data_0[863:856];
        layer6[41][55:48] = buffer_data_0[871:864];
        layer0[42][7:0] = buffer_data_6[831:824];
        layer0[42][15:8] = buffer_data_6[839:832];
        layer0[42][23:16] = buffer_data_6[847:840];
        layer0[42][31:24] = buffer_data_6[855:848];
        layer0[42][39:32] = buffer_data_6[863:856];
        layer0[42][47:40] = buffer_data_6[871:864];
        layer0[42][55:48] = buffer_data_6[879:872];
        layer1[42][7:0] = buffer_data_5[831:824];
        layer1[42][15:8] = buffer_data_5[839:832];
        layer1[42][23:16] = buffer_data_5[847:840];
        layer1[42][31:24] = buffer_data_5[855:848];
        layer1[42][39:32] = buffer_data_5[863:856];
        layer1[42][47:40] = buffer_data_5[871:864];
        layer1[42][55:48] = buffer_data_5[879:872];
        layer2[42][7:0] = buffer_data_4[831:824];
        layer2[42][15:8] = buffer_data_4[839:832];
        layer2[42][23:16] = buffer_data_4[847:840];
        layer2[42][31:24] = buffer_data_4[855:848];
        layer2[42][39:32] = buffer_data_4[863:856];
        layer2[42][47:40] = buffer_data_4[871:864];
        layer2[42][55:48] = buffer_data_4[879:872];
        layer3[42][7:0] = buffer_data_3[831:824];
        layer3[42][15:8] = buffer_data_3[839:832];
        layer3[42][23:16] = buffer_data_3[847:840];
        layer3[42][31:24] = buffer_data_3[855:848];
        layer3[42][39:32] = buffer_data_3[863:856];
        layer3[42][47:40] = buffer_data_3[871:864];
        layer3[42][55:48] = buffer_data_3[879:872];
        layer4[42][7:0] = buffer_data_2[831:824];
        layer4[42][15:8] = buffer_data_2[839:832];
        layer4[42][23:16] = buffer_data_2[847:840];
        layer4[42][31:24] = buffer_data_2[855:848];
        layer4[42][39:32] = buffer_data_2[863:856];
        layer4[42][47:40] = buffer_data_2[871:864];
        layer4[42][55:48] = buffer_data_2[879:872];
        layer5[42][7:0] = buffer_data_1[831:824];
        layer5[42][15:8] = buffer_data_1[839:832];
        layer5[42][23:16] = buffer_data_1[847:840];
        layer5[42][31:24] = buffer_data_1[855:848];
        layer5[42][39:32] = buffer_data_1[863:856];
        layer5[42][47:40] = buffer_data_1[871:864];
        layer5[42][55:48] = buffer_data_1[879:872];
        layer6[42][7:0] = buffer_data_0[831:824];
        layer6[42][15:8] = buffer_data_0[839:832];
        layer6[42][23:16] = buffer_data_0[847:840];
        layer6[42][31:24] = buffer_data_0[855:848];
        layer6[42][39:32] = buffer_data_0[863:856];
        layer6[42][47:40] = buffer_data_0[871:864];
        layer6[42][55:48] = buffer_data_0[879:872];
        layer0[43][7:0] = buffer_data_6[839:832];
        layer0[43][15:8] = buffer_data_6[847:840];
        layer0[43][23:16] = buffer_data_6[855:848];
        layer0[43][31:24] = buffer_data_6[863:856];
        layer0[43][39:32] = buffer_data_6[871:864];
        layer0[43][47:40] = buffer_data_6[879:872];
        layer0[43][55:48] = buffer_data_6[887:880];
        layer1[43][7:0] = buffer_data_5[839:832];
        layer1[43][15:8] = buffer_data_5[847:840];
        layer1[43][23:16] = buffer_data_5[855:848];
        layer1[43][31:24] = buffer_data_5[863:856];
        layer1[43][39:32] = buffer_data_5[871:864];
        layer1[43][47:40] = buffer_data_5[879:872];
        layer1[43][55:48] = buffer_data_5[887:880];
        layer2[43][7:0] = buffer_data_4[839:832];
        layer2[43][15:8] = buffer_data_4[847:840];
        layer2[43][23:16] = buffer_data_4[855:848];
        layer2[43][31:24] = buffer_data_4[863:856];
        layer2[43][39:32] = buffer_data_4[871:864];
        layer2[43][47:40] = buffer_data_4[879:872];
        layer2[43][55:48] = buffer_data_4[887:880];
        layer3[43][7:0] = buffer_data_3[839:832];
        layer3[43][15:8] = buffer_data_3[847:840];
        layer3[43][23:16] = buffer_data_3[855:848];
        layer3[43][31:24] = buffer_data_3[863:856];
        layer3[43][39:32] = buffer_data_3[871:864];
        layer3[43][47:40] = buffer_data_3[879:872];
        layer3[43][55:48] = buffer_data_3[887:880];
        layer4[43][7:0] = buffer_data_2[839:832];
        layer4[43][15:8] = buffer_data_2[847:840];
        layer4[43][23:16] = buffer_data_2[855:848];
        layer4[43][31:24] = buffer_data_2[863:856];
        layer4[43][39:32] = buffer_data_2[871:864];
        layer4[43][47:40] = buffer_data_2[879:872];
        layer4[43][55:48] = buffer_data_2[887:880];
        layer5[43][7:0] = buffer_data_1[839:832];
        layer5[43][15:8] = buffer_data_1[847:840];
        layer5[43][23:16] = buffer_data_1[855:848];
        layer5[43][31:24] = buffer_data_1[863:856];
        layer5[43][39:32] = buffer_data_1[871:864];
        layer5[43][47:40] = buffer_data_1[879:872];
        layer5[43][55:48] = buffer_data_1[887:880];
        layer6[43][7:0] = buffer_data_0[839:832];
        layer6[43][15:8] = buffer_data_0[847:840];
        layer6[43][23:16] = buffer_data_0[855:848];
        layer6[43][31:24] = buffer_data_0[863:856];
        layer6[43][39:32] = buffer_data_0[871:864];
        layer6[43][47:40] = buffer_data_0[879:872];
        layer6[43][55:48] = buffer_data_0[887:880];
        layer0[44][7:0] = buffer_data_6[847:840];
        layer0[44][15:8] = buffer_data_6[855:848];
        layer0[44][23:16] = buffer_data_6[863:856];
        layer0[44][31:24] = buffer_data_6[871:864];
        layer0[44][39:32] = buffer_data_6[879:872];
        layer0[44][47:40] = buffer_data_6[887:880];
        layer0[44][55:48] = buffer_data_6[895:888];
        layer1[44][7:0] = buffer_data_5[847:840];
        layer1[44][15:8] = buffer_data_5[855:848];
        layer1[44][23:16] = buffer_data_5[863:856];
        layer1[44][31:24] = buffer_data_5[871:864];
        layer1[44][39:32] = buffer_data_5[879:872];
        layer1[44][47:40] = buffer_data_5[887:880];
        layer1[44][55:48] = buffer_data_5[895:888];
        layer2[44][7:0] = buffer_data_4[847:840];
        layer2[44][15:8] = buffer_data_4[855:848];
        layer2[44][23:16] = buffer_data_4[863:856];
        layer2[44][31:24] = buffer_data_4[871:864];
        layer2[44][39:32] = buffer_data_4[879:872];
        layer2[44][47:40] = buffer_data_4[887:880];
        layer2[44][55:48] = buffer_data_4[895:888];
        layer3[44][7:0] = buffer_data_3[847:840];
        layer3[44][15:8] = buffer_data_3[855:848];
        layer3[44][23:16] = buffer_data_3[863:856];
        layer3[44][31:24] = buffer_data_3[871:864];
        layer3[44][39:32] = buffer_data_3[879:872];
        layer3[44][47:40] = buffer_data_3[887:880];
        layer3[44][55:48] = buffer_data_3[895:888];
        layer4[44][7:0] = buffer_data_2[847:840];
        layer4[44][15:8] = buffer_data_2[855:848];
        layer4[44][23:16] = buffer_data_2[863:856];
        layer4[44][31:24] = buffer_data_2[871:864];
        layer4[44][39:32] = buffer_data_2[879:872];
        layer4[44][47:40] = buffer_data_2[887:880];
        layer4[44][55:48] = buffer_data_2[895:888];
        layer5[44][7:0] = buffer_data_1[847:840];
        layer5[44][15:8] = buffer_data_1[855:848];
        layer5[44][23:16] = buffer_data_1[863:856];
        layer5[44][31:24] = buffer_data_1[871:864];
        layer5[44][39:32] = buffer_data_1[879:872];
        layer5[44][47:40] = buffer_data_1[887:880];
        layer5[44][55:48] = buffer_data_1[895:888];
        layer6[44][7:0] = buffer_data_0[847:840];
        layer6[44][15:8] = buffer_data_0[855:848];
        layer6[44][23:16] = buffer_data_0[863:856];
        layer6[44][31:24] = buffer_data_0[871:864];
        layer6[44][39:32] = buffer_data_0[879:872];
        layer6[44][47:40] = buffer_data_0[887:880];
        layer6[44][55:48] = buffer_data_0[895:888];
        layer0[45][7:0] = buffer_data_6[855:848];
        layer0[45][15:8] = buffer_data_6[863:856];
        layer0[45][23:16] = buffer_data_6[871:864];
        layer0[45][31:24] = buffer_data_6[879:872];
        layer0[45][39:32] = buffer_data_6[887:880];
        layer0[45][47:40] = buffer_data_6[895:888];
        layer0[45][55:48] = buffer_data_6[903:896];
        layer1[45][7:0] = buffer_data_5[855:848];
        layer1[45][15:8] = buffer_data_5[863:856];
        layer1[45][23:16] = buffer_data_5[871:864];
        layer1[45][31:24] = buffer_data_5[879:872];
        layer1[45][39:32] = buffer_data_5[887:880];
        layer1[45][47:40] = buffer_data_5[895:888];
        layer1[45][55:48] = buffer_data_5[903:896];
        layer2[45][7:0] = buffer_data_4[855:848];
        layer2[45][15:8] = buffer_data_4[863:856];
        layer2[45][23:16] = buffer_data_4[871:864];
        layer2[45][31:24] = buffer_data_4[879:872];
        layer2[45][39:32] = buffer_data_4[887:880];
        layer2[45][47:40] = buffer_data_4[895:888];
        layer2[45][55:48] = buffer_data_4[903:896];
        layer3[45][7:0] = buffer_data_3[855:848];
        layer3[45][15:8] = buffer_data_3[863:856];
        layer3[45][23:16] = buffer_data_3[871:864];
        layer3[45][31:24] = buffer_data_3[879:872];
        layer3[45][39:32] = buffer_data_3[887:880];
        layer3[45][47:40] = buffer_data_3[895:888];
        layer3[45][55:48] = buffer_data_3[903:896];
        layer4[45][7:0] = buffer_data_2[855:848];
        layer4[45][15:8] = buffer_data_2[863:856];
        layer4[45][23:16] = buffer_data_2[871:864];
        layer4[45][31:24] = buffer_data_2[879:872];
        layer4[45][39:32] = buffer_data_2[887:880];
        layer4[45][47:40] = buffer_data_2[895:888];
        layer4[45][55:48] = buffer_data_2[903:896];
        layer5[45][7:0] = buffer_data_1[855:848];
        layer5[45][15:8] = buffer_data_1[863:856];
        layer5[45][23:16] = buffer_data_1[871:864];
        layer5[45][31:24] = buffer_data_1[879:872];
        layer5[45][39:32] = buffer_data_1[887:880];
        layer5[45][47:40] = buffer_data_1[895:888];
        layer5[45][55:48] = buffer_data_1[903:896];
        layer6[45][7:0] = buffer_data_0[855:848];
        layer6[45][15:8] = buffer_data_0[863:856];
        layer6[45][23:16] = buffer_data_0[871:864];
        layer6[45][31:24] = buffer_data_0[879:872];
        layer6[45][39:32] = buffer_data_0[887:880];
        layer6[45][47:40] = buffer_data_0[895:888];
        layer6[45][55:48] = buffer_data_0[903:896];
        layer0[46][7:0] = buffer_data_6[863:856];
        layer0[46][15:8] = buffer_data_6[871:864];
        layer0[46][23:16] = buffer_data_6[879:872];
        layer0[46][31:24] = buffer_data_6[887:880];
        layer0[46][39:32] = buffer_data_6[895:888];
        layer0[46][47:40] = buffer_data_6[903:896];
        layer0[46][55:48] = buffer_data_6[911:904];
        layer1[46][7:0] = buffer_data_5[863:856];
        layer1[46][15:8] = buffer_data_5[871:864];
        layer1[46][23:16] = buffer_data_5[879:872];
        layer1[46][31:24] = buffer_data_5[887:880];
        layer1[46][39:32] = buffer_data_5[895:888];
        layer1[46][47:40] = buffer_data_5[903:896];
        layer1[46][55:48] = buffer_data_5[911:904];
        layer2[46][7:0] = buffer_data_4[863:856];
        layer2[46][15:8] = buffer_data_4[871:864];
        layer2[46][23:16] = buffer_data_4[879:872];
        layer2[46][31:24] = buffer_data_4[887:880];
        layer2[46][39:32] = buffer_data_4[895:888];
        layer2[46][47:40] = buffer_data_4[903:896];
        layer2[46][55:48] = buffer_data_4[911:904];
        layer3[46][7:0] = buffer_data_3[863:856];
        layer3[46][15:8] = buffer_data_3[871:864];
        layer3[46][23:16] = buffer_data_3[879:872];
        layer3[46][31:24] = buffer_data_3[887:880];
        layer3[46][39:32] = buffer_data_3[895:888];
        layer3[46][47:40] = buffer_data_3[903:896];
        layer3[46][55:48] = buffer_data_3[911:904];
        layer4[46][7:0] = buffer_data_2[863:856];
        layer4[46][15:8] = buffer_data_2[871:864];
        layer4[46][23:16] = buffer_data_2[879:872];
        layer4[46][31:24] = buffer_data_2[887:880];
        layer4[46][39:32] = buffer_data_2[895:888];
        layer4[46][47:40] = buffer_data_2[903:896];
        layer4[46][55:48] = buffer_data_2[911:904];
        layer5[46][7:0] = buffer_data_1[863:856];
        layer5[46][15:8] = buffer_data_1[871:864];
        layer5[46][23:16] = buffer_data_1[879:872];
        layer5[46][31:24] = buffer_data_1[887:880];
        layer5[46][39:32] = buffer_data_1[895:888];
        layer5[46][47:40] = buffer_data_1[903:896];
        layer5[46][55:48] = buffer_data_1[911:904];
        layer6[46][7:0] = buffer_data_0[863:856];
        layer6[46][15:8] = buffer_data_0[871:864];
        layer6[46][23:16] = buffer_data_0[879:872];
        layer6[46][31:24] = buffer_data_0[887:880];
        layer6[46][39:32] = buffer_data_0[895:888];
        layer6[46][47:40] = buffer_data_0[903:896];
        layer6[46][55:48] = buffer_data_0[911:904];
        layer0[47][7:0] = buffer_data_6[871:864];
        layer0[47][15:8] = buffer_data_6[879:872];
        layer0[47][23:16] = buffer_data_6[887:880];
        layer0[47][31:24] = buffer_data_6[895:888];
        layer0[47][39:32] = buffer_data_6[903:896];
        layer0[47][47:40] = buffer_data_6[911:904];
        layer0[47][55:48] = buffer_data_6[919:912];
        layer1[47][7:0] = buffer_data_5[871:864];
        layer1[47][15:8] = buffer_data_5[879:872];
        layer1[47][23:16] = buffer_data_5[887:880];
        layer1[47][31:24] = buffer_data_5[895:888];
        layer1[47][39:32] = buffer_data_5[903:896];
        layer1[47][47:40] = buffer_data_5[911:904];
        layer1[47][55:48] = buffer_data_5[919:912];
        layer2[47][7:0] = buffer_data_4[871:864];
        layer2[47][15:8] = buffer_data_4[879:872];
        layer2[47][23:16] = buffer_data_4[887:880];
        layer2[47][31:24] = buffer_data_4[895:888];
        layer2[47][39:32] = buffer_data_4[903:896];
        layer2[47][47:40] = buffer_data_4[911:904];
        layer2[47][55:48] = buffer_data_4[919:912];
        layer3[47][7:0] = buffer_data_3[871:864];
        layer3[47][15:8] = buffer_data_3[879:872];
        layer3[47][23:16] = buffer_data_3[887:880];
        layer3[47][31:24] = buffer_data_3[895:888];
        layer3[47][39:32] = buffer_data_3[903:896];
        layer3[47][47:40] = buffer_data_3[911:904];
        layer3[47][55:48] = buffer_data_3[919:912];
        layer4[47][7:0] = buffer_data_2[871:864];
        layer4[47][15:8] = buffer_data_2[879:872];
        layer4[47][23:16] = buffer_data_2[887:880];
        layer4[47][31:24] = buffer_data_2[895:888];
        layer4[47][39:32] = buffer_data_2[903:896];
        layer4[47][47:40] = buffer_data_2[911:904];
        layer4[47][55:48] = buffer_data_2[919:912];
        layer5[47][7:0] = buffer_data_1[871:864];
        layer5[47][15:8] = buffer_data_1[879:872];
        layer5[47][23:16] = buffer_data_1[887:880];
        layer5[47][31:24] = buffer_data_1[895:888];
        layer5[47][39:32] = buffer_data_1[903:896];
        layer5[47][47:40] = buffer_data_1[911:904];
        layer5[47][55:48] = buffer_data_1[919:912];
        layer6[47][7:0] = buffer_data_0[871:864];
        layer6[47][15:8] = buffer_data_0[879:872];
        layer6[47][23:16] = buffer_data_0[887:880];
        layer6[47][31:24] = buffer_data_0[895:888];
        layer6[47][39:32] = buffer_data_0[903:896];
        layer6[47][47:40] = buffer_data_0[911:904];
        layer6[47][55:48] = buffer_data_0[919:912];
        layer0[48][7:0] = buffer_data_6[879:872];
        layer0[48][15:8] = buffer_data_6[887:880];
        layer0[48][23:16] = buffer_data_6[895:888];
        layer0[48][31:24] = buffer_data_6[903:896];
        layer0[48][39:32] = buffer_data_6[911:904];
        layer0[48][47:40] = buffer_data_6[919:912];
        layer0[48][55:48] = buffer_data_6[927:920];
        layer1[48][7:0] = buffer_data_5[879:872];
        layer1[48][15:8] = buffer_data_5[887:880];
        layer1[48][23:16] = buffer_data_5[895:888];
        layer1[48][31:24] = buffer_data_5[903:896];
        layer1[48][39:32] = buffer_data_5[911:904];
        layer1[48][47:40] = buffer_data_5[919:912];
        layer1[48][55:48] = buffer_data_5[927:920];
        layer2[48][7:0] = buffer_data_4[879:872];
        layer2[48][15:8] = buffer_data_4[887:880];
        layer2[48][23:16] = buffer_data_4[895:888];
        layer2[48][31:24] = buffer_data_4[903:896];
        layer2[48][39:32] = buffer_data_4[911:904];
        layer2[48][47:40] = buffer_data_4[919:912];
        layer2[48][55:48] = buffer_data_4[927:920];
        layer3[48][7:0] = buffer_data_3[879:872];
        layer3[48][15:8] = buffer_data_3[887:880];
        layer3[48][23:16] = buffer_data_3[895:888];
        layer3[48][31:24] = buffer_data_3[903:896];
        layer3[48][39:32] = buffer_data_3[911:904];
        layer3[48][47:40] = buffer_data_3[919:912];
        layer3[48][55:48] = buffer_data_3[927:920];
        layer4[48][7:0] = buffer_data_2[879:872];
        layer4[48][15:8] = buffer_data_2[887:880];
        layer4[48][23:16] = buffer_data_2[895:888];
        layer4[48][31:24] = buffer_data_2[903:896];
        layer4[48][39:32] = buffer_data_2[911:904];
        layer4[48][47:40] = buffer_data_2[919:912];
        layer4[48][55:48] = buffer_data_2[927:920];
        layer5[48][7:0] = buffer_data_1[879:872];
        layer5[48][15:8] = buffer_data_1[887:880];
        layer5[48][23:16] = buffer_data_1[895:888];
        layer5[48][31:24] = buffer_data_1[903:896];
        layer5[48][39:32] = buffer_data_1[911:904];
        layer5[48][47:40] = buffer_data_1[919:912];
        layer5[48][55:48] = buffer_data_1[927:920];
        layer6[48][7:0] = buffer_data_0[879:872];
        layer6[48][15:8] = buffer_data_0[887:880];
        layer6[48][23:16] = buffer_data_0[895:888];
        layer6[48][31:24] = buffer_data_0[903:896];
        layer6[48][39:32] = buffer_data_0[911:904];
        layer6[48][47:40] = buffer_data_0[919:912];
        layer6[48][55:48] = buffer_data_0[927:920];
        layer0[49][7:0] = buffer_data_6[887:880];
        layer0[49][15:8] = buffer_data_6[895:888];
        layer0[49][23:16] = buffer_data_6[903:896];
        layer0[49][31:24] = buffer_data_6[911:904];
        layer0[49][39:32] = buffer_data_6[919:912];
        layer0[49][47:40] = buffer_data_6[927:920];
        layer0[49][55:48] = buffer_data_6[935:928];
        layer1[49][7:0] = buffer_data_5[887:880];
        layer1[49][15:8] = buffer_data_5[895:888];
        layer1[49][23:16] = buffer_data_5[903:896];
        layer1[49][31:24] = buffer_data_5[911:904];
        layer1[49][39:32] = buffer_data_5[919:912];
        layer1[49][47:40] = buffer_data_5[927:920];
        layer1[49][55:48] = buffer_data_5[935:928];
        layer2[49][7:0] = buffer_data_4[887:880];
        layer2[49][15:8] = buffer_data_4[895:888];
        layer2[49][23:16] = buffer_data_4[903:896];
        layer2[49][31:24] = buffer_data_4[911:904];
        layer2[49][39:32] = buffer_data_4[919:912];
        layer2[49][47:40] = buffer_data_4[927:920];
        layer2[49][55:48] = buffer_data_4[935:928];
        layer3[49][7:0] = buffer_data_3[887:880];
        layer3[49][15:8] = buffer_data_3[895:888];
        layer3[49][23:16] = buffer_data_3[903:896];
        layer3[49][31:24] = buffer_data_3[911:904];
        layer3[49][39:32] = buffer_data_3[919:912];
        layer3[49][47:40] = buffer_data_3[927:920];
        layer3[49][55:48] = buffer_data_3[935:928];
        layer4[49][7:0] = buffer_data_2[887:880];
        layer4[49][15:8] = buffer_data_2[895:888];
        layer4[49][23:16] = buffer_data_2[903:896];
        layer4[49][31:24] = buffer_data_2[911:904];
        layer4[49][39:32] = buffer_data_2[919:912];
        layer4[49][47:40] = buffer_data_2[927:920];
        layer4[49][55:48] = buffer_data_2[935:928];
        layer5[49][7:0] = buffer_data_1[887:880];
        layer5[49][15:8] = buffer_data_1[895:888];
        layer5[49][23:16] = buffer_data_1[903:896];
        layer5[49][31:24] = buffer_data_1[911:904];
        layer5[49][39:32] = buffer_data_1[919:912];
        layer5[49][47:40] = buffer_data_1[927:920];
        layer5[49][55:48] = buffer_data_1[935:928];
        layer6[49][7:0] = buffer_data_0[887:880];
        layer6[49][15:8] = buffer_data_0[895:888];
        layer6[49][23:16] = buffer_data_0[903:896];
        layer6[49][31:24] = buffer_data_0[911:904];
        layer6[49][39:32] = buffer_data_0[919:912];
        layer6[49][47:40] = buffer_data_0[927:920];
        layer6[49][55:48] = buffer_data_0[935:928];
        layer0[50][7:0] = buffer_data_6[895:888];
        layer0[50][15:8] = buffer_data_6[903:896];
        layer0[50][23:16] = buffer_data_6[911:904];
        layer0[50][31:24] = buffer_data_6[919:912];
        layer0[50][39:32] = buffer_data_6[927:920];
        layer0[50][47:40] = buffer_data_6[935:928];
        layer0[50][55:48] = buffer_data_6[943:936];
        layer1[50][7:0] = buffer_data_5[895:888];
        layer1[50][15:8] = buffer_data_5[903:896];
        layer1[50][23:16] = buffer_data_5[911:904];
        layer1[50][31:24] = buffer_data_5[919:912];
        layer1[50][39:32] = buffer_data_5[927:920];
        layer1[50][47:40] = buffer_data_5[935:928];
        layer1[50][55:48] = buffer_data_5[943:936];
        layer2[50][7:0] = buffer_data_4[895:888];
        layer2[50][15:8] = buffer_data_4[903:896];
        layer2[50][23:16] = buffer_data_4[911:904];
        layer2[50][31:24] = buffer_data_4[919:912];
        layer2[50][39:32] = buffer_data_4[927:920];
        layer2[50][47:40] = buffer_data_4[935:928];
        layer2[50][55:48] = buffer_data_4[943:936];
        layer3[50][7:0] = buffer_data_3[895:888];
        layer3[50][15:8] = buffer_data_3[903:896];
        layer3[50][23:16] = buffer_data_3[911:904];
        layer3[50][31:24] = buffer_data_3[919:912];
        layer3[50][39:32] = buffer_data_3[927:920];
        layer3[50][47:40] = buffer_data_3[935:928];
        layer3[50][55:48] = buffer_data_3[943:936];
        layer4[50][7:0] = buffer_data_2[895:888];
        layer4[50][15:8] = buffer_data_2[903:896];
        layer4[50][23:16] = buffer_data_2[911:904];
        layer4[50][31:24] = buffer_data_2[919:912];
        layer4[50][39:32] = buffer_data_2[927:920];
        layer4[50][47:40] = buffer_data_2[935:928];
        layer4[50][55:48] = buffer_data_2[943:936];
        layer5[50][7:0] = buffer_data_1[895:888];
        layer5[50][15:8] = buffer_data_1[903:896];
        layer5[50][23:16] = buffer_data_1[911:904];
        layer5[50][31:24] = buffer_data_1[919:912];
        layer5[50][39:32] = buffer_data_1[927:920];
        layer5[50][47:40] = buffer_data_1[935:928];
        layer5[50][55:48] = buffer_data_1[943:936];
        layer6[50][7:0] = buffer_data_0[895:888];
        layer6[50][15:8] = buffer_data_0[903:896];
        layer6[50][23:16] = buffer_data_0[911:904];
        layer6[50][31:24] = buffer_data_0[919:912];
        layer6[50][39:32] = buffer_data_0[927:920];
        layer6[50][47:40] = buffer_data_0[935:928];
        layer6[50][55:48] = buffer_data_0[943:936];
        layer0[51][7:0] = buffer_data_6[903:896];
        layer0[51][15:8] = buffer_data_6[911:904];
        layer0[51][23:16] = buffer_data_6[919:912];
        layer0[51][31:24] = buffer_data_6[927:920];
        layer0[51][39:32] = buffer_data_6[935:928];
        layer0[51][47:40] = buffer_data_6[943:936];
        layer0[51][55:48] = buffer_data_6[951:944];
        layer1[51][7:0] = buffer_data_5[903:896];
        layer1[51][15:8] = buffer_data_5[911:904];
        layer1[51][23:16] = buffer_data_5[919:912];
        layer1[51][31:24] = buffer_data_5[927:920];
        layer1[51][39:32] = buffer_data_5[935:928];
        layer1[51][47:40] = buffer_data_5[943:936];
        layer1[51][55:48] = buffer_data_5[951:944];
        layer2[51][7:0] = buffer_data_4[903:896];
        layer2[51][15:8] = buffer_data_4[911:904];
        layer2[51][23:16] = buffer_data_4[919:912];
        layer2[51][31:24] = buffer_data_4[927:920];
        layer2[51][39:32] = buffer_data_4[935:928];
        layer2[51][47:40] = buffer_data_4[943:936];
        layer2[51][55:48] = buffer_data_4[951:944];
        layer3[51][7:0] = buffer_data_3[903:896];
        layer3[51][15:8] = buffer_data_3[911:904];
        layer3[51][23:16] = buffer_data_3[919:912];
        layer3[51][31:24] = buffer_data_3[927:920];
        layer3[51][39:32] = buffer_data_3[935:928];
        layer3[51][47:40] = buffer_data_3[943:936];
        layer3[51][55:48] = buffer_data_3[951:944];
        layer4[51][7:0] = buffer_data_2[903:896];
        layer4[51][15:8] = buffer_data_2[911:904];
        layer4[51][23:16] = buffer_data_2[919:912];
        layer4[51][31:24] = buffer_data_2[927:920];
        layer4[51][39:32] = buffer_data_2[935:928];
        layer4[51][47:40] = buffer_data_2[943:936];
        layer4[51][55:48] = buffer_data_2[951:944];
        layer5[51][7:0] = buffer_data_1[903:896];
        layer5[51][15:8] = buffer_data_1[911:904];
        layer5[51][23:16] = buffer_data_1[919:912];
        layer5[51][31:24] = buffer_data_1[927:920];
        layer5[51][39:32] = buffer_data_1[935:928];
        layer5[51][47:40] = buffer_data_1[943:936];
        layer5[51][55:48] = buffer_data_1[951:944];
        layer6[51][7:0] = buffer_data_0[903:896];
        layer6[51][15:8] = buffer_data_0[911:904];
        layer6[51][23:16] = buffer_data_0[919:912];
        layer6[51][31:24] = buffer_data_0[927:920];
        layer6[51][39:32] = buffer_data_0[935:928];
        layer6[51][47:40] = buffer_data_0[943:936];
        layer6[51][55:48] = buffer_data_0[951:944];
        layer0[52][7:0] = buffer_data_6[911:904];
        layer0[52][15:8] = buffer_data_6[919:912];
        layer0[52][23:16] = buffer_data_6[927:920];
        layer0[52][31:24] = buffer_data_6[935:928];
        layer0[52][39:32] = buffer_data_6[943:936];
        layer0[52][47:40] = buffer_data_6[951:944];
        layer0[52][55:48] = buffer_data_6[959:952];
        layer1[52][7:0] = buffer_data_5[911:904];
        layer1[52][15:8] = buffer_data_5[919:912];
        layer1[52][23:16] = buffer_data_5[927:920];
        layer1[52][31:24] = buffer_data_5[935:928];
        layer1[52][39:32] = buffer_data_5[943:936];
        layer1[52][47:40] = buffer_data_5[951:944];
        layer1[52][55:48] = buffer_data_5[959:952];
        layer2[52][7:0] = buffer_data_4[911:904];
        layer2[52][15:8] = buffer_data_4[919:912];
        layer2[52][23:16] = buffer_data_4[927:920];
        layer2[52][31:24] = buffer_data_4[935:928];
        layer2[52][39:32] = buffer_data_4[943:936];
        layer2[52][47:40] = buffer_data_4[951:944];
        layer2[52][55:48] = buffer_data_4[959:952];
        layer3[52][7:0] = buffer_data_3[911:904];
        layer3[52][15:8] = buffer_data_3[919:912];
        layer3[52][23:16] = buffer_data_3[927:920];
        layer3[52][31:24] = buffer_data_3[935:928];
        layer3[52][39:32] = buffer_data_3[943:936];
        layer3[52][47:40] = buffer_data_3[951:944];
        layer3[52][55:48] = buffer_data_3[959:952];
        layer4[52][7:0] = buffer_data_2[911:904];
        layer4[52][15:8] = buffer_data_2[919:912];
        layer4[52][23:16] = buffer_data_2[927:920];
        layer4[52][31:24] = buffer_data_2[935:928];
        layer4[52][39:32] = buffer_data_2[943:936];
        layer4[52][47:40] = buffer_data_2[951:944];
        layer4[52][55:48] = buffer_data_2[959:952];
        layer5[52][7:0] = buffer_data_1[911:904];
        layer5[52][15:8] = buffer_data_1[919:912];
        layer5[52][23:16] = buffer_data_1[927:920];
        layer5[52][31:24] = buffer_data_1[935:928];
        layer5[52][39:32] = buffer_data_1[943:936];
        layer5[52][47:40] = buffer_data_1[951:944];
        layer5[52][55:48] = buffer_data_1[959:952];
        layer6[52][7:0] = buffer_data_0[911:904];
        layer6[52][15:8] = buffer_data_0[919:912];
        layer6[52][23:16] = buffer_data_0[927:920];
        layer6[52][31:24] = buffer_data_0[935:928];
        layer6[52][39:32] = buffer_data_0[943:936];
        layer6[52][47:40] = buffer_data_0[951:944];
        layer6[52][55:48] = buffer_data_0[959:952];
        layer0[53][7:0] = buffer_data_6[919:912];
        layer0[53][15:8] = buffer_data_6[927:920];
        layer0[53][23:16] = buffer_data_6[935:928];
        layer0[53][31:24] = buffer_data_6[943:936];
        layer0[53][39:32] = buffer_data_6[951:944];
        layer0[53][47:40] = buffer_data_6[959:952];
        layer0[53][55:48] = buffer_data_6[967:960];
        layer1[53][7:0] = buffer_data_5[919:912];
        layer1[53][15:8] = buffer_data_5[927:920];
        layer1[53][23:16] = buffer_data_5[935:928];
        layer1[53][31:24] = buffer_data_5[943:936];
        layer1[53][39:32] = buffer_data_5[951:944];
        layer1[53][47:40] = buffer_data_5[959:952];
        layer1[53][55:48] = buffer_data_5[967:960];
        layer2[53][7:0] = buffer_data_4[919:912];
        layer2[53][15:8] = buffer_data_4[927:920];
        layer2[53][23:16] = buffer_data_4[935:928];
        layer2[53][31:24] = buffer_data_4[943:936];
        layer2[53][39:32] = buffer_data_4[951:944];
        layer2[53][47:40] = buffer_data_4[959:952];
        layer2[53][55:48] = buffer_data_4[967:960];
        layer3[53][7:0] = buffer_data_3[919:912];
        layer3[53][15:8] = buffer_data_3[927:920];
        layer3[53][23:16] = buffer_data_3[935:928];
        layer3[53][31:24] = buffer_data_3[943:936];
        layer3[53][39:32] = buffer_data_3[951:944];
        layer3[53][47:40] = buffer_data_3[959:952];
        layer3[53][55:48] = buffer_data_3[967:960];
        layer4[53][7:0] = buffer_data_2[919:912];
        layer4[53][15:8] = buffer_data_2[927:920];
        layer4[53][23:16] = buffer_data_2[935:928];
        layer4[53][31:24] = buffer_data_2[943:936];
        layer4[53][39:32] = buffer_data_2[951:944];
        layer4[53][47:40] = buffer_data_2[959:952];
        layer4[53][55:48] = buffer_data_2[967:960];
        layer5[53][7:0] = buffer_data_1[919:912];
        layer5[53][15:8] = buffer_data_1[927:920];
        layer5[53][23:16] = buffer_data_1[935:928];
        layer5[53][31:24] = buffer_data_1[943:936];
        layer5[53][39:32] = buffer_data_1[951:944];
        layer5[53][47:40] = buffer_data_1[959:952];
        layer5[53][55:48] = buffer_data_1[967:960];
        layer6[53][7:0] = buffer_data_0[919:912];
        layer6[53][15:8] = buffer_data_0[927:920];
        layer6[53][23:16] = buffer_data_0[935:928];
        layer6[53][31:24] = buffer_data_0[943:936];
        layer6[53][39:32] = buffer_data_0[951:944];
        layer6[53][47:40] = buffer_data_0[959:952];
        layer6[53][55:48] = buffer_data_0[967:960];
        layer0[54][7:0] = buffer_data_6[927:920];
        layer0[54][15:8] = buffer_data_6[935:928];
        layer0[54][23:16] = buffer_data_6[943:936];
        layer0[54][31:24] = buffer_data_6[951:944];
        layer0[54][39:32] = buffer_data_6[959:952];
        layer0[54][47:40] = buffer_data_6[967:960];
        layer0[54][55:48] = buffer_data_6[975:968];
        layer1[54][7:0] = buffer_data_5[927:920];
        layer1[54][15:8] = buffer_data_5[935:928];
        layer1[54][23:16] = buffer_data_5[943:936];
        layer1[54][31:24] = buffer_data_5[951:944];
        layer1[54][39:32] = buffer_data_5[959:952];
        layer1[54][47:40] = buffer_data_5[967:960];
        layer1[54][55:48] = buffer_data_5[975:968];
        layer2[54][7:0] = buffer_data_4[927:920];
        layer2[54][15:8] = buffer_data_4[935:928];
        layer2[54][23:16] = buffer_data_4[943:936];
        layer2[54][31:24] = buffer_data_4[951:944];
        layer2[54][39:32] = buffer_data_4[959:952];
        layer2[54][47:40] = buffer_data_4[967:960];
        layer2[54][55:48] = buffer_data_4[975:968];
        layer3[54][7:0] = buffer_data_3[927:920];
        layer3[54][15:8] = buffer_data_3[935:928];
        layer3[54][23:16] = buffer_data_3[943:936];
        layer3[54][31:24] = buffer_data_3[951:944];
        layer3[54][39:32] = buffer_data_3[959:952];
        layer3[54][47:40] = buffer_data_3[967:960];
        layer3[54][55:48] = buffer_data_3[975:968];
        layer4[54][7:0] = buffer_data_2[927:920];
        layer4[54][15:8] = buffer_data_2[935:928];
        layer4[54][23:16] = buffer_data_2[943:936];
        layer4[54][31:24] = buffer_data_2[951:944];
        layer4[54][39:32] = buffer_data_2[959:952];
        layer4[54][47:40] = buffer_data_2[967:960];
        layer4[54][55:48] = buffer_data_2[975:968];
        layer5[54][7:0] = buffer_data_1[927:920];
        layer5[54][15:8] = buffer_data_1[935:928];
        layer5[54][23:16] = buffer_data_1[943:936];
        layer5[54][31:24] = buffer_data_1[951:944];
        layer5[54][39:32] = buffer_data_1[959:952];
        layer5[54][47:40] = buffer_data_1[967:960];
        layer5[54][55:48] = buffer_data_1[975:968];
        layer6[54][7:0] = buffer_data_0[927:920];
        layer6[54][15:8] = buffer_data_0[935:928];
        layer6[54][23:16] = buffer_data_0[943:936];
        layer6[54][31:24] = buffer_data_0[951:944];
        layer6[54][39:32] = buffer_data_0[959:952];
        layer6[54][47:40] = buffer_data_0[967:960];
        layer6[54][55:48] = buffer_data_0[975:968];
        layer0[55][7:0] = buffer_data_6[935:928];
        layer0[55][15:8] = buffer_data_6[943:936];
        layer0[55][23:16] = buffer_data_6[951:944];
        layer0[55][31:24] = buffer_data_6[959:952];
        layer0[55][39:32] = buffer_data_6[967:960];
        layer0[55][47:40] = buffer_data_6[975:968];
        layer0[55][55:48] = buffer_data_6[983:976];
        layer1[55][7:0] = buffer_data_5[935:928];
        layer1[55][15:8] = buffer_data_5[943:936];
        layer1[55][23:16] = buffer_data_5[951:944];
        layer1[55][31:24] = buffer_data_5[959:952];
        layer1[55][39:32] = buffer_data_5[967:960];
        layer1[55][47:40] = buffer_data_5[975:968];
        layer1[55][55:48] = buffer_data_5[983:976];
        layer2[55][7:0] = buffer_data_4[935:928];
        layer2[55][15:8] = buffer_data_4[943:936];
        layer2[55][23:16] = buffer_data_4[951:944];
        layer2[55][31:24] = buffer_data_4[959:952];
        layer2[55][39:32] = buffer_data_4[967:960];
        layer2[55][47:40] = buffer_data_4[975:968];
        layer2[55][55:48] = buffer_data_4[983:976];
        layer3[55][7:0] = buffer_data_3[935:928];
        layer3[55][15:8] = buffer_data_3[943:936];
        layer3[55][23:16] = buffer_data_3[951:944];
        layer3[55][31:24] = buffer_data_3[959:952];
        layer3[55][39:32] = buffer_data_3[967:960];
        layer3[55][47:40] = buffer_data_3[975:968];
        layer3[55][55:48] = buffer_data_3[983:976];
        layer4[55][7:0] = buffer_data_2[935:928];
        layer4[55][15:8] = buffer_data_2[943:936];
        layer4[55][23:16] = buffer_data_2[951:944];
        layer4[55][31:24] = buffer_data_2[959:952];
        layer4[55][39:32] = buffer_data_2[967:960];
        layer4[55][47:40] = buffer_data_2[975:968];
        layer4[55][55:48] = buffer_data_2[983:976];
        layer5[55][7:0] = buffer_data_1[935:928];
        layer5[55][15:8] = buffer_data_1[943:936];
        layer5[55][23:16] = buffer_data_1[951:944];
        layer5[55][31:24] = buffer_data_1[959:952];
        layer5[55][39:32] = buffer_data_1[967:960];
        layer5[55][47:40] = buffer_data_1[975:968];
        layer5[55][55:48] = buffer_data_1[983:976];
        layer6[55][7:0] = buffer_data_0[935:928];
        layer6[55][15:8] = buffer_data_0[943:936];
        layer6[55][23:16] = buffer_data_0[951:944];
        layer6[55][31:24] = buffer_data_0[959:952];
        layer6[55][39:32] = buffer_data_0[967:960];
        layer6[55][47:40] = buffer_data_0[975:968];
        layer6[55][55:48] = buffer_data_0[983:976];
        layer0[56][7:0] = buffer_data_6[943:936];
        layer0[56][15:8] = buffer_data_6[951:944];
        layer0[56][23:16] = buffer_data_6[959:952];
        layer0[56][31:24] = buffer_data_6[967:960];
        layer0[56][39:32] = buffer_data_6[975:968];
        layer0[56][47:40] = buffer_data_6[983:976];
        layer0[56][55:48] = buffer_data_6[991:984];
        layer1[56][7:0] = buffer_data_5[943:936];
        layer1[56][15:8] = buffer_data_5[951:944];
        layer1[56][23:16] = buffer_data_5[959:952];
        layer1[56][31:24] = buffer_data_5[967:960];
        layer1[56][39:32] = buffer_data_5[975:968];
        layer1[56][47:40] = buffer_data_5[983:976];
        layer1[56][55:48] = buffer_data_5[991:984];
        layer2[56][7:0] = buffer_data_4[943:936];
        layer2[56][15:8] = buffer_data_4[951:944];
        layer2[56][23:16] = buffer_data_4[959:952];
        layer2[56][31:24] = buffer_data_4[967:960];
        layer2[56][39:32] = buffer_data_4[975:968];
        layer2[56][47:40] = buffer_data_4[983:976];
        layer2[56][55:48] = buffer_data_4[991:984];
        layer3[56][7:0] = buffer_data_3[943:936];
        layer3[56][15:8] = buffer_data_3[951:944];
        layer3[56][23:16] = buffer_data_3[959:952];
        layer3[56][31:24] = buffer_data_3[967:960];
        layer3[56][39:32] = buffer_data_3[975:968];
        layer3[56][47:40] = buffer_data_3[983:976];
        layer3[56][55:48] = buffer_data_3[991:984];
        layer4[56][7:0] = buffer_data_2[943:936];
        layer4[56][15:8] = buffer_data_2[951:944];
        layer4[56][23:16] = buffer_data_2[959:952];
        layer4[56][31:24] = buffer_data_2[967:960];
        layer4[56][39:32] = buffer_data_2[975:968];
        layer4[56][47:40] = buffer_data_2[983:976];
        layer4[56][55:48] = buffer_data_2[991:984];
        layer5[56][7:0] = buffer_data_1[943:936];
        layer5[56][15:8] = buffer_data_1[951:944];
        layer5[56][23:16] = buffer_data_1[959:952];
        layer5[56][31:24] = buffer_data_1[967:960];
        layer5[56][39:32] = buffer_data_1[975:968];
        layer5[56][47:40] = buffer_data_1[983:976];
        layer5[56][55:48] = buffer_data_1[991:984];
        layer6[56][7:0] = buffer_data_0[943:936];
        layer6[56][15:8] = buffer_data_0[951:944];
        layer6[56][23:16] = buffer_data_0[959:952];
        layer6[56][31:24] = buffer_data_0[967:960];
        layer6[56][39:32] = buffer_data_0[975:968];
        layer6[56][47:40] = buffer_data_0[983:976];
        layer6[56][55:48] = buffer_data_0[991:984];
        layer0[57][7:0] = buffer_data_6[951:944];
        layer0[57][15:8] = buffer_data_6[959:952];
        layer0[57][23:16] = buffer_data_6[967:960];
        layer0[57][31:24] = buffer_data_6[975:968];
        layer0[57][39:32] = buffer_data_6[983:976];
        layer0[57][47:40] = buffer_data_6[991:984];
        layer0[57][55:48] = buffer_data_6[999:992];
        layer1[57][7:0] = buffer_data_5[951:944];
        layer1[57][15:8] = buffer_data_5[959:952];
        layer1[57][23:16] = buffer_data_5[967:960];
        layer1[57][31:24] = buffer_data_5[975:968];
        layer1[57][39:32] = buffer_data_5[983:976];
        layer1[57][47:40] = buffer_data_5[991:984];
        layer1[57][55:48] = buffer_data_5[999:992];
        layer2[57][7:0] = buffer_data_4[951:944];
        layer2[57][15:8] = buffer_data_4[959:952];
        layer2[57][23:16] = buffer_data_4[967:960];
        layer2[57][31:24] = buffer_data_4[975:968];
        layer2[57][39:32] = buffer_data_4[983:976];
        layer2[57][47:40] = buffer_data_4[991:984];
        layer2[57][55:48] = buffer_data_4[999:992];
        layer3[57][7:0] = buffer_data_3[951:944];
        layer3[57][15:8] = buffer_data_3[959:952];
        layer3[57][23:16] = buffer_data_3[967:960];
        layer3[57][31:24] = buffer_data_3[975:968];
        layer3[57][39:32] = buffer_data_3[983:976];
        layer3[57][47:40] = buffer_data_3[991:984];
        layer3[57][55:48] = buffer_data_3[999:992];
        layer4[57][7:0] = buffer_data_2[951:944];
        layer4[57][15:8] = buffer_data_2[959:952];
        layer4[57][23:16] = buffer_data_2[967:960];
        layer4[57][31:24] = buffer_data_2[975:968];
        layer4[57][39:32] = buffer_data_2[983:976];
        layer4[57][47:40] = buffer_data_2[991:984];
        layer4[57][55:48] = buffer_data_2[999:992];
        layer5[57][7:0] = buffer_data_1[951:944];
        layer5[57][15:8] = buffer_data_1[959:952];
        layer5[57][23:16] = buffer_data_1[967:960];
        layer5[57][31:24] = buffer_data_1[975:968];
        layer5[57][39:32] = buffer_data_1[983:976];
        layer5[57][47:40] = buffer_data_1[991:984];
        layer5[57][55:48] = buffer_data_1[999:992];
        layer6[57][7:0] = buffer_data_0[951:944];
        layer6[57][15:8] = buffer_data_0[959:952];
        layer6[57][23:16] = buffer_data_0[967:960];
        layer6[57][31:24] = buffer_data_0[975:968];
        layer6[57][39:32] = buffer_data_0[983:976];
        layer6[57][47:40] = buffer_data_0[991:984];
        layer6[57][55:48] = buffer_data_0[999:992];
        layer0[58][7:0] = buffer_data_6[959:952];
        layer0[58][15:8] = buffer_data_6[967:960];
        layer0[58][23:16] = buffer_data_6[975:968];
        layer0[58][31:24] = buffer_data_6[983:976];
        layer0[58][39:32] = buffer_data_6[991:984];
        layer0[58][47:40] = buffer_data_6[999:992];
        layer0[58][55:48] = buffer_data_6[1007:1000];
        layer1[58][7:0] = buffer_data_5[959:952];
        layer1[58][15:8] = buffer_data_5[967:960];
        layer1[58][23:16] = buffer_data_5[975:968];
        layer1[58][31:24] = buffer_data_5[983:976];
        layer1[58][39:32] = buffer_data_5[991:984];
        layer1[58][47:40] = buffer_data_5[999:992];
        layer1[58][55:48] = buffer_data_5[1007:1000];
        layer2[58][7:0] = buffer_data_4[959:952];
        layer2[58][15:8] = buffer_data_4[967:960];
        layer2[58][23:16] = buffer_data_4[975:968];
        layer2[58][31:24] = buffer_data_4[983:976];
        layer2[58][39:32] = buffer_data_4[991:984];
        layer2[58][47:40] = buffer_data_4[999:992];
        layer2[58][55:48] = buffer_data_4[1007:1000];
        layer3[58][7:0] = buffer_data_3[959:952];
        layer3[58][15:8] = buffer_data_3[967:960];
        layer3[58][23:16] = buffer_data_3[975:968];
        layer3[58][31:24] = buffer_data_3[983:976];
        layer3[58][39:32] = buffer_data_3[991:984];
        layer3[58][47:40] = buffer_data_3[999:992];
        layer3[58][55:48] = buffer_data_3[1007:1000];
        layer4[58][7:0] = buffer_data_2[959:952];
        layer4[58][15:8] = buffer_data_2[967:960];
        layer4[58][23:16] = buffer_data_2[975:968];
        layer4[58][31:24] = buffer_data_2[983:976];
        layer4[58][39:32] = buffer_data_2[991:984];
        layer4[58][47:40] = buffer_data_2[999:992];
        layer4[58][55:48] = buffer_data_2[1007:1000];
        layer5[58][7:0] = buffer_data_1[959:952];
        layer5[58][15:8] = buffer_data_1[967:960];
        layer5[58][23:16] = buffer_data_1[975:968];
        layer5[58][31:24] = buffer_data_1[983:976];
        layer5[58][39:32] = buffer_data_1[991:984];
        layer5[58][47:40] = buffer_data_1[999:992];
        layer5[58][55:48] = buffer_data_1[1007:1000];
        layer6[58][7:0] = buffer_data_0[959:952];
        layer6[58][15:8] = buffer_data_0[967:960];
        layer6[58][23:16] = buffer_data_0[975:968];
        layer6[58][31:24] = buffer_data_0[983:976];
        layer6[58][39:32] = buffer_data_0[991:984];
        layer6[58][47:40] = buffer_data_0[999:992];
        layer6[58][55:48] = buffer_data_0[1007:1000];
        layer0[59][7:0] = buffer_data_6[967:960];
        layer0[59][15:8] = buffer_data_6[975:968];
        layer0[59][23:16] = buffer_data_6[983:976];
        layer0[59][31:24] = buffer_data_6[991:984];
        layer0[59][39:32] = buffer_data_6[999:992];
        layer0[59][47:40] = buffer_data_6[1007:1000];
        layer0[59][55:48] = buffer_data_6[1015:1008];
        layer1[59][7:0] = buffer_data_5[967:960];
        layer1[59][15:8] = buffer_data_5[975:968];
        layer1[59][23:16] = buffer_data_5[983:976];
        layer1[59][31:24] = buffer_data_5[991:984];
        layer1[59][39:32] = buffer_data_5[999:992];
        layer1[59][47:40] = buffer_data_5[1007:1000];
        layer1[59][55:48] = buffer_data_5[1015:1008];
        layer2[59][7:0] = buffer_data_4[967:960];
        layer2[59][15:8] = buffer_data_4[975:968];
        layer2[59][23:16] = buffer_data_4[983:976];
        layer2[59][31:24] = buffer_data_4[991:984];
        layer2[59][39:32] = buffer_data_4[999:992];
        layer2[59][47:40] = buffer_data_4[1007:1000];
        layer2[59][55:48] = buffer_data_4[1015:1008];
        layer3[59][7:0] = buffer_data_3[967:960];
        layer3[59][15:8] = buffer_data_3[975:968];
        layer3[59][23:16] = buffer_data_3[983:976];
        layer3[59][31:24] = buffer_data_3[991:984];
        layer3[59][39:32] = buffer_data_3[999:992];
        layer3[59][47:40] = buffer_data_3[1007:1000];
        layer3[59][55:48] = buffer_data_3[1015:1008];
        layer4[59][7:0] = buffer_data_2[967:960];
        layer4[59][15:8] = buffer_data_2[975:968];
        layer4[59][23:16] = buffer_data_2[983:976];
        layer4[59][31:24] = buffer_data_2[991:984];
        layer4[59][39:32] = buffer_data_2[999:992];
        layer4[59][47:40] = buffer_data_2[1007:1000];
        layer4[59][55:48] = buffer_data_2[1015:1008];
        layer5[59][7:0] = buffer_data_1[967:960];
        layer5[59][15:8] = buffer_data_1[975:968];
        layer5[59][23:16] = buffer_data_1[983:976];
        layer5[59][31:24] = buffer_data_1[991:984];
        layer5[59][39:32] = buffer_data_1[999:992];
        layer5[59][47:40] = buffer_data_1[1007:1000];
        layer5[59][55:48] = buffer_data_1[1015:1008];
        layer6[59][7:0] = buffer_data_0[967:960];
        layer6[59][15:8] = buffer_data_0[975:968];
        layer6[59][23:16] = buffer_data_0[983:976];
        layer6[59][31:24] = buffer_data_0[991:984];
        layer6[59][39:32] = buffer_data_0[999:992];
        layer6[59][47:40] = buffer_data_0[1007:1000];
        layer6[59][55:48] = buffer_data_0[1015:1008];
        layer0[60][7:0] = buffer_data_6[975:968];
        layer0[60][15:8] = buffer_data_6[983:976];
        layer0[60][23:16] = buffer_data_6[991:984];
        layer0[60][31:24] = buffer_data_6[999:992];
        layer0[60][39:32] = buffer_data_6[1007:1000];
        layer0[60][47:40] = buffer_data_6[1015:1008];
        layer0[60][55:48] = buffer_data_6[1023:1016];
        layer1[60][7:0] = buffer_data_5[975:968];
        layer1[60][15:8] = buffer_data_5[983:976];
        layer1[60][23:16] = buffer_data_5[991:984];
        layer1[60][31:24] = buffer_data_5[999:992];
        layer1[60][39:32] = buffer_data_5[1007:1000];
        layer1[60][47:40] = buffer_data_5[1015:1008];
        layer1[60][55:48] = buffer_data_5[1023:1016];
        layer2[60][7:0] = buffer_data_4[975:968];
        layer2[60][15:8] = buffer_data_4[983:976];
        layer2[60][23:16] = buffer_data_4[991:984];
        layer2[60][31:24] = buffer_data_4[999:992];
        layer2[60][39:32] = buffer_data_4[1007:1000];
        layer2[60][47:40] = buffer_data_4[1015:1008];
        layer2[60][55:48] = buffer_data_4[1023:1016];
        layer3[60][7:0] = buffer_data_3[975:968];
        layer3[60][15:8] = buffer_data_3[983:976];
        layer3[60][23:16] = buffer_data_3[991:984];
        layer3[60][31:24] = buffer_data_3[999:992];
        layer3[60][39:32] = buffer_data_3[1007:1000];
        layer3[60][47:40] = buffer_data_3[1015:1008];
        layer3[60][55:48] = buffer_data_3[1023:1016];
        layer4[60][7:0] = buffer_data_2[975:968];
        layer4[60][15:8] = buffer_data_2[983:976];
        layer4[60][23:16] = buffer_data_2[991:984];
        layer4[60][31:24] = buffer_data_2[999:992];
        layer4[60][39:32] = buffer_data_2[1007:1000];
        layer4[60][47:40] = buffer_data_2[1015:1008];
        layer4[60][55:48] = buffer_data_2[1023:1016];
        layer5[60][7:0] = buffer_data_1[975:968];
        layer5[60][15:8] = buffer_data_1[983:976];
        layer5[60][23:16] = buffer_data_1[991:984];
        layer5[60][31:24] = buffer_data_1[999:992];
        layer5[60][39:32] = buffer_data_1[1007:1000];
        layer5[60][47:40] = buffer_data_1[1015:1008];
        layer5[60][55:48] = buffer_data_1[1023:1016];
        layer6[60][7:0] = buffer_data_0[975:968];
        layer6[60][15:8] = buffer_data_0[983:976];
        layer6[60][23:16] = buffer_data_0[991:984];
        layer6[60][31:24] = buffer_data_0[999:992];
        layer6[60][39:32] = buffer_data_0[1007:1000];
        layer6[60][47:40] = buffer_data_0[1015:1008];
        layer6[60][55:48] = buffer_data_0[1023:1016];
        layer0[61][7:0] = buffer_data_6[983:976];
        layer0[61][15:8] = buffer_data_6[991:984];
        layer0[61][23:16] = buffer_data_6[999:992];
        layer0[61][31:24] = buffer_data_6[1007:1000];
        layer0[61][39:32] = buffer_data_6[1015:1008];
        layer0[61][47:40] = buffer_data_6[1023:1016];
        layer0[61][55:48] = buffer_data_6[1031:1024];
        layer1[61][7:0] = buffer_data_5[983:976];
        layer1[61][15:8] = buffer_data_5[991:984];
        layer1[61][23:16] = buffer_data_5[999:992];
        layer1[61][31:24] = buffer_data_5[1007:1000];
        layer1[61][39:32] = buffer_data_5[1015:1008];
        layer1[61][47:40] = buffer_data_5[1023:1016];
        layer1[61][55:48] = buffer_data_5[1031:1024];
        layer2[61][7:0] = buffer_data_4[983:976];
        layer2[61][15:8] = buffer_data_4[991:984];
        layer2[61][23:16] = buffer_data_4[999:992];
        layer2[61][31:24] = buffer_data_4[1007:1000];
        layer2[61][39:32] = buffer_data_4[1015:1008];
        layer2[61][47:40] = buffer_data_4[1023:1016];
        layer2[61][55:48] = buffer_data_4[1031:1024];
        layer3[61][7:0] = buffer_data_3[983:976];
        layer3[61][15:8] = buffer_data_3[991:984];
        layer3[61][23:16] = buffer_data_3[999:992];
        layer3[61][31:24] = buffer_data_3[1007:1000];
        layer3[61][39:32] = buffer_data_3[1015:1008];
        layer3[61][47:40] = buffer_data_3[1023:1016];
        layer3[61][55:48] = buffer_data_3[1031:1024];
        layer4[61][7:0] = buffer_data_2[983:976];
        layer4[61][15:8] = buffer_data_2[991:984];
        layer4[61][23:16] = buffer_data_2[999:992];
        layer4[61][31:24] = buffer_data_2[1007:1000];
        layer4[61][39:32] = buffer_data_2[1015:1008];
        layer4[61][47:40] = buffer_data_2[1023:1016];
        layer4[61][55:48] = buffer_data_2[1031:1024];
        layer5[61][7:0] = buffer_data_1[983:976];
        layer5[61][15:8] = buffer_data_1[991:984];
        layer5[61][23:16] = buffer_data_1[999:992];
        layer5[61][31:24] = buffer_data_1[1007:1000];
        layer5[61][39:32] = buffer_data_1[1015:1008];
        layer5[61][47:40] = buffer_data_1[1023:1016];
        layer5[61][55:48] = buffer_data_1[1031:1024];
        layer6[61][7:0] = buffer_data_0[983:976];
        layer6[61][15:8] = buffer_data_0[991:984];
        layer6[61][23:16] = buffer_data_0[999:992];
        layer6[61][31:24] = buffer_data_0[1007:1000];
        layer6[61][39:32] = buffer_data_0[1015:1008];
        layer6[61][47:40] = buffer_data_0[1023:1016];
        layer6[61][55:48] = buffer_data_0[1031:1024];
        layer0[62][7:0] = buffer_data_6[991:984];
        layer0[62][15:8] = buffer_data_6[999:992];
        layer0[62][23:16] = buffer_data_6[1007:1000];
        layer0[62][31:24] = buffer_data_6[1015:1008];
        layer0[62][39:32] = buffer_data_6[1023:1016];
        layer0[62][47:40] = buffer_data_6[1031:1024];
        layer0[62][55:48] = buffer_data_6[1039:1032];
        layer1[62][7:0] = buffer_data_5[991:984];
        layer1[62][15:8] = buffer_data_5[999:992];
        layer1[62][23:16] = buffer_data_5[1007:1000];
        layer1[62][31:24] = buffer_data_5[1015:1008];
        layer1[62][39:32] = buffer_data_5[1023:1016];
        layer1[62][47:40] = buffer_data_5[1031:1024];
        layer1[62][55:48] = buffer_data_5[1039:1032];
        layer2[62][7:0] = buffer_data_4[991:984];
        layer2[62][15:8] = buffer_data_4[999:992];
        layer2[62][23:16] = buffer_data_4[1007:1000];
        layer2[62][31:24] = buffer_data_4[1015:1008];
        layer2[62][39:32] = buffer_data_4[1023:1016];
        layer2[62][47:40] = buffer_data_4[1031:1024];
        layer2[62][55:48] = buffer_data_4[1039:1032];
        layer3[62][7:0] = buffer_data_3[991:984];
        layer3[62][15:8] = buffer_data_3[999:992];
        layer3[62][23:16] = buffer_data_3[1007:1000];
        layer3[62][31:24] = buffer_data_3[1015:1008];
        layer3[62][39:32] = buffer_data_3[1023:1016];
        layer3[62][47:40] = buffer_data_3[1031:1024];
        layer3[62][55:48] = buffer_data_3[1039:1032];
        layer4[62][7:0] = buffer_data_2[991:984];
        layer4[62][15:8] = buffer_data_2[999:992];
        layer4[62][23:16] = buffer_data_2[1007:1000];
        layer4[62][31:24] = buffer_data_2[1015:1008];
        layer4[62][39:32] = buffer_data_2[1023:1016];
        layer4[62][47:40] = buffer_data_2[1031:1024];
        layer4[62][55:48] = buffer_data_2[1039:1032];
        layer5[62][7:0] = buffer_data_1[991:984];
        layer5[62][15:8] = buffer_data_1[999:992];
        layer5[62][23:16] = buffer_data_1[1007:1000];
        layer5[62][31:24] = buffer_data_1[1015:1008];
        layer5[62][39:32] = buffer_data_1[1023:1016];
        layer5[62][47:40] = buffer_data_1[1031:1024];
        layer5[62][55:48] = buffer_data_1[1039:1032];
        layer6[62][7:0] = buffer_data_0[991:984];
        layer6[62][15:8] = buffer_data_0[999:992];
        layer6[62][23:16] = buffer_data_0[1007:1000];
        layer6[62][31:24] = buffer_data_0[1015:1008];
        layer6[62][39:32] = buffer_data_0[1023:1016];
        layer6[62][47:40] = buffer_data_0[1031:1024];
        layer6[62][55:48] = buffer_data_0[1039:1032];
        layer0[63][7:0] = buffer_data_6[999:992];
        layer0[63][15:8] = buffer_data_6[1007:1000];
        layer0[63][23:16] = buffer_data_6[1015:1008];
        layer0[63][31:24] = buffer_data_6[1023:1016];
        layer0[63][39:32] = buffer_data_6[1031:1024];
        layer0[63][47:40] = buffer_data_6[1039:1032];
        layer0[63][55:48] = buffer_data_6[1047:1040];
        layer1[63][7:0] = buffer_data_5[999:992];
        layer1[63][15:8] = buffer_data_5[1007:1000];
        layer1[63][23:16] = buffer_data_5[1015:1008];
        layer1[63][31:24] = buffer_data_5[1023:1016];
        layer1[63][39:32] = buffer_data_5[1031:1024];
        layer1[63][47:40] = buffer_data_5[1039:1032];
        layer1[63][55:48] = buffer_data_5[1047:1040];
        layer2[63][7:0] = buffer_data_4[999:992];
        layer2[63][15:8] = buffer_data_4[1007:1000];
        layer2[63][23:16] = buffer_data_4[1015:1008];
        layer2[63][31:24] = buffer_data_4[1023:1016];
        layer2[63][39:32] = buffer_data_4[1031:1024];
        layer2[63][47:40] = buffer_data_4[1039:1032];
        layer2[63][55:48] = buffer_data_4[1047:1040];
        layer3[63][7:0] = buffer_data_3[999:992];
        layer3[63][15:8] = buffer_data_3[1007:1000];
        layer3[63][23:16] = buffer_data_3[1015:1008];
        layer3[63][31:24] = buffer_data_3[1023:1016];
        layer3[63][39:32] = buffer_data_3[1031:1024];
        layer3[63][47:40] = buffer_data_3[1039:1032];
        layer3[63][55:48] = buffer_data_3[1047:1040];
        layer4[63][7:0] = buffer_data_2[999:992];
        layer4[63][15:8] = buffer_data_2[1007:1000];
        layer4[63][23:16] = buffer_data_2[1015:1008];
        layer4[63][31:24] = buffer_data_2[1023:1016];
        layer4[63][39:32] = buffer_data_2[1031:1024];
        layer4[63][47:40] = buffer_data_2[1039:1032];
        layer4[63][55:48] = buffer_data_2[1047:1040];
        layer5[63][7:0] = buffer_data_1[999:992];
        layer5[63][15:8] = buffer_data_1[1007:1000];
        layer5[63][23:16] = buffer_data_1[1015:1008];
        layer5[63][31:24] = buffer_data_1[1023:1016];
        layer5[63][39:32] = buffer_data_1[1031:1024];
        layer5[63][47:40] = buffer_data_1[1039:1032];
        layer5[63][55:48] = buffer_data_1[1047:1040];
        layer6[63][7:0] = buffer_data_0[999:992];
        layer6[63][15:8] = buffer_data_0[1007:1000];
        layer6[63][23:16] = buffer_data_0[1015:1008];
        layer6[63][31:24] = buffer_data_0[1023:1016];
        layer6[63][39:32] = buffer_data_0[1031:1024];
        layer6[63][47:40] = buffer_data_0[1039:1032];
        layer6[63][55:48] = buffer_data_0[1047:1040];
    end
    ST_GAUSSIAN_2: begin
        layer0[0][7:0] = buffer_data_6[1007:1000];
        layer0[0][15:8] = buffer_data_6[1015:1008];
        layer0[0][23:16] = buffer_data_6[1023:1016];
        layer0[0][31:24] = buffer_data_6[1031:1024];
        layer0[0][39:32] = buffer_data_6[1039:1032];
        layer0[0][47:40] = buffer_data_6[1047:1040];
        layer0[0][55:48] = buffer_data_6[1055:1048];
        layer1[0][7:0] = buffer_data_5[1007:1000];
        layer1[0][15:8] = buffer_data_5[1015:1008];
        layer1[0][23:16] = buffer_data_5[1023:1016];
        layer1[0][31:24] = buffer_data_5[1031:1024];
        layer1[0][39:32] = buffer_data_5[1039:1032];
        layer1[0][47:40] = buffer_data_5[1047:1040];
        layer1[0][55:48] = buffer_data_5[1055:1048];
        layer2[0][7:0] = buffer_data_4[1007:1000];
        layer2[0][15:8] = buffer_data_4[1015:1008];
        layer2[0][23:16] = buffer_data_4[1023:1016];
        layer2[0][31:24] = buffer_data_4[1031:1024];
        layer2[0][39:32] = buffer_data_4[1039:1032];
        layer2[0][47:40] = buffer_data_4[1047:1040];
        layer2[0][55:48] = buffer_data_4[1055:1048];
        layer3[0][7:0] = buffer_data_3[1007:1000];
        layer3[0][15:8] = buffer_data_3[1015:1008];
        layer3[0][23:16] = buffer_data_3[1023:1016];
        layer3[0][31:24] = buffer_data_3[1031:1024];
        layer3[0][39:32] = buffer_data_3[1039:1032];
        layer3[0][47:40] = buffer_data_3[1047:1040];
        layer3[0][55:48] = buffer_data_3[1055:1048];
        layer4[0][7:0] = buffer_data_2[1007:1000];
        layer4[0][15:8] = buffer_data_2[1015:1008];
        layer4[0][23:16] = buffer_data_2[1023:1016];
        layer4[0][31:24] = buffer_data_2[1031:1024];
        layer4[0][39:32] = buffer_data_2[1039:1032];
        layer4[0][47:40] = buffer_data_2[1047:1040];
        layer4[0][55:48] = buffer_data_2[1055:1048];
        layer5[0][7:0] = buffer_data_1[1007:1000];
        layer5[0][15:8] = buffer_data_1[1015:1008];
        layer5[0][23:16] = buffer_data_1[1023:1016];
        layer5[0][31:24] = buffer_data_1[1031:1024];
        layer5[0][39:32] = buffer_data_1[1039:1032];
        layer5[0][47:40] = buffer_data_1[1047:1040];
        layer5[0][55:48] = buffer_data_1[1055:1048];
        layer6[0][7:0] = buffer_data_0[1007:1000];
        layer6[0][15:8] = buffer_data_0[1015:1008];
        layer6[0][23:16] = buffer_data_0[1023:1016];
        layer6[0][31:24] = buffer_data_0[1031:1024];
        layer6[0][39:32] = buffer_data_0[1039:1032];
        layer6[0][47:40] = buffer_data_0[1047:1040];
        layer6[0][55:48] = buffer_data_0[1055:1048];
        layer0[1][7:0] = buffer_data_6[1015:1008];
        layer0[1][15:8] = buffer_data_6[1023:1016];
        layer0[1][23:16] = buffer_data_6[1031:1024];
        layer0[1][31:24] = buffer_data_6[1039:1032];
        layer0[1][39:32] = buffer_data_6[1047:1040];
        layer0[1][47:40] = buffer_data_6[1055:1048];
        layer0[1][55:48] = buffer_data_6[1063:1056];
        layer1[1][7:0] = buffer_data_5[1015:1008];
        layer1[1][15:8] = buffer_data_5[1023:1016];
        layer1[1][23:16] = buffer_data_5[1031:1024];
        layer1[1][31:24] = buffer_data_5[1039:1032];
        layer1[1][39:32] = buffer_data_5[1047:1040];
        layer1[1][47:40] = buffer_data_5[1055:1048];
        layer1[1][55:48] = buffer_data_5[1063:1056];
        layer2[1][7:0] = buffer_data_4[1015:1008];
        layer2[1][15:8] = buffer_data_4[1023:1016];
        layer2[1][23:16] = buffer_data_4[1031:1024];
        layer2[1][31:24] = buffer_data_4[1039:1032];
        layer2[1][39:32] = buffer_data_4[1047:1040];
        layer2[1][47:40] = buffer_data_4[1055:1048];
        layer2[1][55:48] = buffer_data_4[1063:1056];
        layer3[1][7:0] = buffer_data_3[1015:1008];
        layer3[1][15:8] = buffer_data_3[1023:1016];
        layer3[1][23:16] = buffer_data_3[1031:1024];
        layer3[1][31:24] = buffer_data_3[1039:1032];
        layer3[1][39:32] = buffer_data_3[1047:1040];
        layer3[1][47:40] = buffer_data_3[1055:1048];
        layer3[1][55:48] = buffer_data_3[1063:1056];
        layer4[1][7:0] = buffer_data_2[1015:1008];
        layer4[1][15:8] = buffer_data_2[1023:1016];
        layer4[1][23:16] = buffer_data_2[1031:1024];
        layer4[1][31:24] = buffer_data_2[1039:1032];
        layer4[1][39:32] = buffer_data_2[1047:1040];
        layer4[1][47:40] = buffer_data_2[1055:1048];
        layer4[1][55:48] = buffer_data_2[1063:1056];
        layer5[1][7:0] = buffer_data_1[1015:1008];
        layer5[1][15:8] = buffer_data_1[1023:1016];
        layer5[1][23:16] = buffer_data_1[1031:1024];
        layer5[1][31:24] = buffer_data_1[1039:1032];
        layer5[1][39:32] = buffer_data_1[1047:1040];
        layer5[1][47:40] = buffer_data_1[1055:1048];
        layer5[1][55:48] = buffer_data_1[1063:1056];
        layer6[1][7:0] = buffer_data_0[1015:1008];
        layer6[1][15:8] = buffer_data_0[1023:1016];
        layer6[1][23:16] = buffer_data_0[1031:1024];
        layer6[1][31:24] = buffer_data_0[1039:1032];
        layer6[1][39:32] = buffer_data_0[1047:1040];
        layer6[1][47:40] = buffer_data_0[1055:1048];
        layer6[1][55:48] = buffer_data_0[1063:1056];
        layer0[2][7:0] = buffer_data_6[1023:1016];
        layer0[2][15:8] = buffer_data_6[1031:1024];
        layer0[2][23:16] = buffer_data_6[1039:1032];
        layer0[2][31:24] = buffer_data_6[1047:1040];
        layer0[2][39:32] = buffer_data_6[1055:1048];
        layer0[2][47:40] = buffer_data_6[1063:1056];
        layer0[2][55:48] = buffer_data_6[1071:1064];
        layer1[2][7:0] = buffer_data_5[1023:1016];
        layer1[2][15:8] = buffer_data_5[1031:1024];
        layer1[2][23:16] = buffer_data_5[1039:1032];
        layer1[2][31:24] = buffer_data_5[1047:1040];
        layer1[2][39:32] = buffer_data_5[1055:1048];
        layer1[2][47:40] = buffer_data_5[1063:1056];
        layer1[2][55:48] = buffer_data_5[1071:1064];
        layer2[2][7:0] = buffer_data_4[1023:1016];
        layer2[2][15:8] = buffer_data_4[1031:1024];
        layer2[2][23:16] = buffer_data_4[1039:1032];
        layer2[2][31:24] = buffer_data_4[1047:1040];
        layer2[2][39:32] = buffer_data_4[1055:1048];
        layer2[2][47:40] = buffer_data_4[1063:1056];
        layer2[2][55:48] = buffer_data_4[1071:1064];
        layer3[2][7:0] = buffer_data_3[1023:1016];
        layer3[2][15:8] = buffer_data_3[1031:1024];
        layer3[2][23:16] = buffer_data_3[1039:1032];
        layer3[2][31:24] = buffer_data_3[1047:1040];
        layer3[2][39:32] = buffer_data_3[1055:1048];
        layer3[2][47:40] = buffer_data_3[1063:1056];
        layer3[2][55:48] = buffer_data_3[1071:1064];
        layer4[2][7:0] = buffer_data_2[1023:1016];
        layer4[2][15:8] = buffer_data_2[1031:1024];
        layer4[2][23:16] = buffer_data_2[1039:1032];
        layer4[2][31:24] = buffer_data_2[1047:1040];
        layer4[2][39:32] = buffer_data_2[1055:1048];
        layer4[2][47:40] = buffer_data_2[1063:1056];
        layer4[2][55:48] = buffer_data_2[1071:1064];
        layer5[2][7:0] = buffer_data_1[1023:1016];
        layer5[2][15:8] = buffer_data_1[1031:1024];
        layer5[2][23:16] = buffer_data_1[1039:1032];
        layer5[2][31:24] = buffer_data_1[1047:1040];
        layer5[2][39:32] = buffer_data_1[1055:1048];
        layer5[2][47:40] = buffer_data_1[1063:1056];
        layer5[2][55:48] = buffer_data_1[1071:1064];
        layer6[2][7:0] = buffer_data_0[1023:1016];
        layer6[2][15:8] = buffer_data_0[1031:1024];
        layer6[2][23:16] = buffer_data_0[1039:1032];
        layer6[2][31:24] = buffer_data_0[1047:1040];
        layer6[2][39:32] = buffer_data_0[1055:1048];
        layer6[2][47:40] = buffer_data_0[1063:1056];
        layer6[2][55:48] = buffer_data_0[1071:1064];
        layer0[3][7:0] = buffer_data_6[1031:1024];
        layer0[3][15:8] = buffer_data_6[1039:1032];
        layer0[3][23:16] = buffer_data_6[1047:1040];
        layer0[3][31:24] = buffer_data_6[1055:1048];
        layer0[3][39:32] = buffer_data_6[1063:1056];
        layer0[3][47:40] = buffer_data_6[1071:1064];
        layer0[3][55:48] = buffer_data_6[1079:1072];
        layer1[3][7:0] = buffer_data_5[1031:1024];
        layer1[3][15:8] = buffer_data_5[1039:1032];
        layer1[3][23:16] = buffer_data_5[1047:1040];
        layer1[3][31:24] = buffer_data_5[1055:1048];
        layer1[3][39:32] = buffer_data_5[1063:1056];
        layer1[3][47:40] = buffer_data_5[1071:1064];
        layer1[3][55:48] = buffer_data_5[1079:1072];
        layer2[3][7:0] = buffer_data_4[1031:1024];
        layer2[3][15:8] = buffer_data_4[1039:1032];
        layer2[3][23:16] = buffer_data_4[1047:1040];
        layer2[3][31:24] = buffer_data_4[1055:1048];
        layer2[3][39:32] = buffer_data_4[1063:1056];
        layer2[3][47:40] = buffer_data_4[1071:1064];
        layer2[3][55:48] = buffer_data_4[1079:1072];
        layer3[3][7:0] = buffer_data_3[1031:1024];
        layer3[3][15:8] = buffer_data_3[1039:1032];
        layer3[3][23:16] = buffer_data_3[1047:1040];
        layer3[3][31:24] = buffer_data_3[1055:1048];
        layer3[3][39:32] = buffer_data_3[1063:1056];
        layer3[3][47:40] = buffer_data_3[1071:1064];
        layer3[3][55:48] = buffer_data_3[1079:1072];
        layer4[3][7:0] = buffer_data_2[1031:1024];
        layer4[3][15:8] = buffer_data_2[1039:1032];
        layer4[3][23:16] = buffer_data_2[1047:1040];
        layer4[3][31:24] = buffer_data_2[1055:1048];
        layer4[3][39:32] = buffer_data_2[1063:1056];
        layer4[3][47:40] = buffer_data_2[1071:1064];
        layer4[3][55:48] = buffer_data_2[1079:1072];
        layer5[3][7:0] = buffer_data_1[1031:1024];
        layer5[3][15:8] = buffer_data_1[1039:1032];
        layer5[3][23:16] = buffer_data_1[1047:1040];
        layer5[3][31:24] = buffer_data_1[1055:1048];
        layer5[3][39:32] = buffer_data_1[1063:1056];
        layer5[3][47:40] = buffer_data_1[1071:1064];
        layer5[3][55:48] = buffer_data_1[1079:1072];
        layer6[3][7:0] = buffer_data_0[1031:1024];
        layer6[3][15:8] = buffer_data_0[1039:1032];
        layer6[3][23:16] = buffer_data_0[1047:1040];
        layer6[3][31:24] = buffer_data_0[1055:1048];
        layer6[3][39:32] = buffer_data_0[1063:1056];
        layer6[3][47:40] = buffer_data_0[1071:1064];
        layer6[3][55:48] = buffer_data_0[1079:1072];
        layer0[4][7:0] = buffer_data_6[1039:1032];
        layer0[4][15:8] = buffer_data_6[1047:1040];
        layer0[4][23:16] = buffer_data_6[1055:1048];
        layer0[4][31:24] = buffer_data_6[1063:1056];
        layer0[4][39:32] = buffer_data_6[1071:1064];
        layer0[4][47:40] = buffer_data_6[1079:1072];
        layer0[4][55:48] = buffer_data_6[1087:1080];
        layer1[4][7:0] = buffer_data_5[1039:1032];
        layer1[4][15:8] = buffer_data_5[1047:1040];
        layer1[4][23:16] = buffer_data_5[1055:1048];
        layer1[4][31:24] = buffer_data_5[1063:1056];
        layer1[4][39:32] = buffer_data_5[1071:1064];
        layer1[4][47:40] = buffer_data_5[1079:1072];
        layer1[4][55:48] = buffer_data_5[1087:1080];
        layer2[4][7:0] = buffer_data_4[1039:1032];
        layer2[4][15:8] = buffer_data_4[1047:1040];
        layer2[4][23:16] = buffer_data_4[1055:1048];
        layer2[4][31:24] = buffer_data_4[1063:1056];
        layer2[4][39:32] = buffer_data_4[1071:1064];
        layer2[4][47:40] = buffer_data_4[1079:1072];
        layer2[4][55:48] = buffer_data_4[1087:1080];
        layer3[4][7:0] = buffer_data_3[1039:1032];
        layer3[4][15:8] = buffer_data_3[1047:1040];
        layer3[4][23:16] = buffer_data_3[1055:1048];
        layer3[4][31:24] = buffer_data_3[1063:1056];
        layer3[4][39:32] = buffer_data_3[1071:1064];
        layer3[4][47:40] = buffer_data_3[1079:1072];
        layer3[4][55:48] = buffer_data_3[1087:1080];
        layer4[4][7:0] = buffer_data_2[1039:1032];
        layer4[4][15:8] = buffer_data_2[1047:1040];
        layer4[4][23:16] = buffer_data_2[1055:1048];
        layer4[4][31:24] = buffer_data_2[1063:1056];
        layer4[4][39:32] = buffer_data_2[1071:1064];
        layer4[4][47:40] = buffer_data_2[1079:1072];
        layer4[4][55:48] = buffer_data_2[1087:1080];
        layer5[4][7:0] = buffer_data_1[1039:1032];
        layer5[4][15:8] = buffer_data_1[1047:1040];
        layer5[4][23:16] = buffer_data_1[1055:1048];
        layer5[4][31:24] = buffer_data_1[1063:1056];
        layer5[4][39:32] = buffer_data_1[1071:1064];
        layer5[4][47:40] = buffer_data_1[1079:1072];
        layer5[4][55:48] = buffer_data_1[1087:1080];
        layer6[4][7:0] = buffer_data_0[1039:1032];
        layer6[4][15:8] = buffer_data_0[1047:1040];
        layer6[4][23:16] = buffer_data_0[1055:1048];
        layer6[4][31:24] = buffer_data_0[1063:1056];
        layer6[4][39:32] = buffer_data_0[1071:1064];
        layer6[4][47:40] = buffer_data_0[1079:1072];
        layer6[4][55:48] = buffer_data_0[1087:1080];
        layer0[5][7:0] = buffer_data_6[1047:1040];
        layer0[5][15:8] = buffer_data_6[1055:1048];
        layer0[5][23:16] = buffer_data_6[1063:1056];
        layer0[5][31:24] = buffer_data_6[1071:1064];
        layer0[5][39:32] = buffer_data_6[1079:1072];
        layer0[5][47:40] = buffer_data_6[1087:1080];
        layer0[5][55:48] = buffer_data_6[1095:1088];
        layer1[5][7:0] = buffer_data_5[1047:1040];
        layer1[5][15:8] = buffer_data_5[1055:1048];
        layer1[5][23:16] = buffer_data_5[1063:1056];
        layer1[5][31:24] = buffer_data_5[1071:1064];
        layer1[5][39:32] = buffer_data_5[1079:1072];
        layer1[5][47:40] = buffer_data_5[1087:1080];
        layer1[5][55:48] = buffer_data_5[1095:1088];
        layer2[5][7:0] = buffer_data_4[1047:1040];
        layer2[5][15:8] = buffer_data_4[1055:1048];
        layer2[5][23:16] = buffer_data_4[1063:1056];
        layer2[5][31:24] = buffer_data_4[1071:1064];
        layer2[5][39:32] = buffer_data_4[1079:1072];
        layer2[5][47:40] = buffer_data_4[1087:1080];
        layer2[5][55:48] = buffer_data_4[1095:1088];
        layer3[5][7:0] = buffer_data_3[1047:1040];
        layer3[5][15:8] = buffer_data_3[1055:1048];
        layer3[5][23:16] = buffer_data_3[1063:1056];
        layer3[5][31:24] = buffer_data_3[1071:1064];
        layer3[5][39:32] = buffer_data_3[1079:1072];
        layer3[5][47:40] = buffer_data_3[1087:1080];
        layer3[5][55:48] = buffer_data_3[1095:1088];
        layer4[5][7:0] = buffer_data_2[1047:1040];
        layer4[5][15:8] = buffer_data_2[1055:1048];
        layer4[5][23:16] = buffer_data_2[1063:1056];
        layer4[5][31:24] = buffer_data_2[1071:1064];
        layer4[5][39:32] = buffer_data_2[1079:1072];
        layer4[5][47:40] = buffer_data_2[1087:1080];
        layer4[5][55:48] = buffer_data_2[1095:1088];
        layer5[5][7:0] = buffer_data_1[1047:1040];
        layer5[5][15:8] = buffer_data_1[1055:1048];
        layer5[5][23:16] = buffer_data_1[1063:1056];
        layer5[5][31:24] = buffer_data_1[1071:1064];
        layer5[5][39:32] = buffer_data_1[1079:1072];
        layer5[5][47:40] = buffer_data_1[1087:1080];
        layer5[5][55:48] = buffer_data_1[1095:1088];
        layer6[5][7:0] = buffer_data_0[1047:1040];
        layer6[5][15:8] = buffer_data_0[1055:1048];
        layer6[5][23:16] = buffer_data_0[1063:1056];
        layer6[5][31:24] = buffer_data_0[1071:1064];
        layer6[5][39:32] = buffer_data_0[1079:1072];
        layer6[5][47:40] = buffer_data_0[1087:1080];
        layer6[5][55:48] = buffer_data_0[1095:1088];
        layer0[6][7:0] = buffer_data_6[1055:1048];
        layer0[6][15:8] = buffer_data_6[1063:1056];
        layer0[6][23:16] = buffer_data_6[1071:1064];
        layer0[6][31:24] = buffer_data_6[1079:1072];
        layer0[6][39:32] = buffer_data_6[1087:1080];
        layer0[6][47:40] = buffer_data_6[1095:1088];
        layer0[6][55:48] = buffer_data_6[1103:1096];
        layer1[6][7:0] = buffer_data_5[1055:1048];
        layer1[6][15:8] = buffer_data_5[1063:1056];
        layer1[6][23:16] = buffer_data_5[1071:1064];
        layer1[6][31:24] = buffer_data_5[1079:1072];
        layer1[6][39:32] = buffer_data_5[1087:1080];
        layer1[6][47:40] = buffer_data_5[1095:1088];
        layer1[6][55:48] = buffer_data_5[1103:1096];
        layer2[6][7:0] = buffer_data_4[1055:1048];
        layer2[6][15:8] = buffer_data_4[1063:1056];
        layer2[6][23:16] = buffer_data_4[1071:1064];
        layer2[6][31:24] = buffer_data_4[1079:1072];
        layer2[6][39:32] = buffer_data_4[1087:1080];
        layer2[6][47:40] = buffer_data_4[1095:1088];
        layer2[6][55:48] = buffer_data_4[1103:1096];
        layer3[6][7:0] = buffer_data_3[1055:1048];
        layer3[6][15:8] = buffer_data_3[1063:1056];
        layer3[6][23:16] = buffer_data_3[1071:1064];
        layer3[6][31:24] = buffer_data_3[1079:1072];
        layer3[6][39:32] = buffer_data_3[1087:1080];
        layer3[6][47:40] = buffer_data_3[1095:1088];
        layer3[6][55:48] = buffer_data_3[1103:1096];
        layer4[6][7:0] = buffer_data_2[1055:1048];
        layer4[6][15:8] = buffer_data_2[1063:1056];
        layer4[6][23:16] = buffer_data_2[1071:1064];
        layer4[6][31:24] = buffer_data_2[1079:1072];
        layer4[6][39:32] = buffer_data_2[1087:1080];
        layer4[6][47:40] = buffer_data_2[1095:1088];
        layer4[6][55:48] = buffer_data_2[1103:1096];
        layer5[6][7:0] = buffer_data_1[1055:1048];
        layer5[6][15:8] = buffer_data_1[1063:1056];
        layer5[6][23:16] = buffer_data_1[1071:1064];
        layer5[6][31:24] = buffer_data_1[1079:1072];
        layer5[6][39:32] = buffer_data_1[1087:1080];
        layer5[6][47:40] = buffer_data_1[1095:1088];
        layer5[6][55:48] = buffer_data_1[1103:1096];
        layer6[6][7:0] = buffer_data_0[1055:1048];
        layer6[6][15:8] = buffer_data_0[1063:1056];
        layer6[6][23:16] = buffer_data_0[1071:1064];
        layer6[6][31:24] = buffer_data_0[1079:1072];
        layer6[6][39:32] = buffer_data_0[1087:1080];
        layer6[6][47:40] = buffer_data_0[1095:1088];
        layer6[6][55:48] = buffer_data_0[1103:1096];
        layer0[7][7:0] = buffer_data_6[1063:1056];
        layer0[7][15:8] = buffer_data_6[1071:1064];
        layer0[7][23:16] = buffer_data_6[1079:1072];
        layer0[7][31:24] = buffer_data_6[1087:1080];
        layer0[7][39:32] = buffer_data_6[1095:1088];
        layer0[7][47:40] = buffer_data_6[1103:1096];
        layer0[7][55:48] = buffer_data_6[1111:1104];
        layer1[7][7:0] = buffer_data_5[1063:1056];
        layer1[7][15:8] = buffer_data_5[1071:1064];
        layer1[7][23:16] = buffer_data_5[1079:1072];
        layer1[7][31:24] = buffer_data_5[1087:1080];
        layer1[7][39:32] = buffer_data_5[1095:1088];
        layer1[7][47:40] = buffer_data_5[1103:1096];
        layer1[7][55:48] = buffer_data_5[1111:1104];
        layer2[7][7:0] = buffer_data_4[1063:1056];
        layer2[7][15:8] = buffer_data_4[1071:1064];
        layer2[7][23:16] = buffer_data_4[1079:1072];
        layer2[7][31:24] = buffer_data_4[1087:1080];
        layer2[7][39:32] = buffer_data_4[1095:1088];
        layer2[7][47:40] = buffer_data_4[1103:1096];
        layer2[7][55:48] = buffer_data_4[1111:1104];
        layer3[7][7:0] = buffer_data_3[1063:1056];
        layer3[7][15:8] = buffer_data_3[1071:1064];
        layer3[7][23:16] = buffer_data_3[1079:1072];
        layer3[7][31:24] = buffer_data_3[1087:1080];
        layer3[7][39:32] = buffer_data_3[1095:1088];
        layer3[7][47:40] = buffer_data_3[1103:1096];
        layer3[7][55:48] = buffer_data_3[1111:1104];
        layer4[7][7:0] = buffer_data_2[1063:1056];
        layer4[7][15:8] = buffer_data_2[1071:1064];
        layer4[7][23:16] = buffer_data_2[1079:1072];
        layer4[7][31:24] = buffer_data_2[1087:1080];
        layer4[7][39:32] = buffer_data_2[1095:1088];
        layer4[7][47:40] = buffer_data_2[1103:1096];
        layer4[7][55:48] = buffer_data_2[1111:1104];
        layer5[7][7:0] = buffer_data_1[1063:1056];
        layer5[7][15:8] = buffer_data_1[1071:1064];
        layer5[7][23:16] = buffer_data_1[1079:1072];
        layer5[7][31:24] = buffer_data_1[1087:1080];
        layer5[7][39:32] = buffer_data_1[1095:1088];
        layer5[7][47:40] = buffer_data_1[1103:1096];
        layer5[7][55:48] = buffer_data_1[1111:1104];
        layer6[7][7:0] = buffer_data_0[1063:1056];
        layer6[7][15:8] = buffer_data_0[1071:1064];
        layer6[7][23:16] = buffer_data_0[1079:1072];
        layer6[7][31:24] = buffer_data_0[1087:1080];
        layer6[7][39:32] = buffer_data_0[1095:1088];
        layer6[7][47:40] = buffer_data_0[1103:1096];
        layer6[7][55:48] = buffer_data_0[1111:1104];
        layer0[8][7:0] = buffer_data_6[1071:1064];
        layer0[8][15:8] = buffer_data_6[1079:1072];
        layer0[8][23:16] = buffer_data_6[1087:1080];
        layer0[8][31:24] = buffer_data_6[1095:1088];
        layer0[8][39:32] = buffer_data_6[1103:1096];
        layer0[8][47:40] = buffer_data_6[1111:1104];
        layer0[8][55:48] = buffer_data_6[1119:1112];
        layer1[8][7:0] = buffer_data_5[1071:1064];
        layer1[8][15:8] = buffer_data_5[1079:1072];
        layer1[8][23:16] = buffer_data_5[1087:1080];
        layer1[8][31:24] = buffer_data_5[1095:1088];
        layer1[8][39:32] = buffer_data_5[1103:1096];
        layer1[8][47:40] = buffer_data_5[1111:1104];
        layer1[8][55:48] = buffer_data_5[1119:1112];
        layer2[8][7:0] = buffer_data_4[1071:1064];
        layer2[8][15:8] = buffer_data_4[1079:1072];
        layer2[8][23:16] = buffer_data_4[1087:1080];
        layer2[8][31:24] = buffer_data_4[1095:1088];
        layer2[8][39:32] = buffer_data_4[1103:1096];
        layer2[8][47:40] = buffer_data_4[1111:1104];
        layer2[8][55:48] = buffer_data_4[1119:1112];
        layer3[8][7:0] = buffer_data_3[1071:1064];
        layer3[8][15:8] = buffer_data_3[1079:1072];
        layer3[8][23:16] = buffer_data_3[1087:1080];
        layer3[8][31:24] = buffer_data_3[1095:1088];
        layer3[8][39:32] = buffer_data_3[1103:1096];
        layer3[8][47:40] = buffer_data_3[1111:1104];
        layer3[8][55:48] = buffer_data_3[1119:1112];
        layer4[8][7:0] = buffer_data_2[1071:1064];
        layer4[8][15:8] = buffer_data_2[1079:1072];
        layer4[8][23:16] = buffer_data_2[1087:1080];
        layer4[8][31:24] = buffer_data_2[1095:1088];
        layer4[8][39:32] = buffer_data_2[1103:1096];
        layer4[8][47:40] = buffer_data_2[1111:1104];
        layer4[8][55:48] = buffer_data_2[1119:1112];
        layer5[8][7:0] = buffer_data_1[1071:1064];
        layer5[8][15:8] = buffer_data_1[1079:1072];
        layer5[8][23:16] = buffer_data_1[1087:1080];
        layer5[8][31:24] = buffer_data_1[1095:1088];
        layer5[8][39:32] = buffer_data_1[1103:1096];
        layer5[8][47:40] = buffer_data_1[1111:1104];
        layer5[8][55:48] = buffer_data_1[1119:1112];
        layer6[8][7:0] = buffer_data_0[1071:1064];
        layer6[8][15:8] = buffer_data_0[1079:1072];
        layer6[8][23:16] = buffer_data_0[1087:1080];
        layer6[8][31:24] = buffer_data_0[1095:1088];
        layer6[8][39:32] = buffer_data_0[1103:1096];
        layer6[8][47:40] = buffer_data_0[1111:1104];
        layer6[8][55:48] = buffer_data_0[1119:1112];
        layer0[9][7:0] = buffer_data_6[1079:1072];
        layer0[9][15:8] = buffer_data_6[1087:1080];
        layer0[9][23:16] = buffer_data_6[1095:1088];
        layer0[9][31:24] = buffer_data_6[1103:1096];
        layer0[9][39:32] = buffer_data_6[1111:1104];
        layer0[9][47:40] = buffer_data_6[1119:1112];
        layer0[9][55:48] = buffer_data_6[1127:1120];
        layer1[9][7:0] = buffer_data_5[1079:1072];
        layer1[9][15:8] = buffer_data_5[1087:1080];
        layer1[9][23:16] = buffer_data_5[1095:1088];
        layer1[9][31:24] = buffer_data_5[1103:1096];
        layer1[9][39:32] = buffer_data_5[1111:1104];
        layer1[9][47:40] = buffer_data_5[1119:1112];
        layer1[9][55:48] = buffer_data_5[1127:1120];
        layer2[9][7:0] = buffer_data_4[1079:1072];
        layer2[9][15:8] = buffer_data_4[1087:1080];
        layer2[9][23:16] = buffer_data_4[1095:1088];
        layer2[9][31:24] = buffer_data_4[1103:1096];
        layer2[9][39:32] = buffer_data_4[1111:1104];
        layer2[9][47:40] = buffer_data_4[1119:1112];
        layer2[9][55:48] = buffer_data_4[1127:1120];
        layer3[9][7:0] = buffer_data_3[1079:1072];
        layer3[9][15:8] = buffer_data_3[1087:1080];
        layer3[9][23:16] = buffer_data_3[1095:1088];
        layer3[9][31:24] = buffer_data_3[1103:1096];
        layer3[9][39:32] = buffer_data_3[1111:1104];
        layer3[9][47:40] = buffer_data_3[1119:1112];
        layer3[9][55:48] = buffer_data_3[1127:1120];
        layer4[9][7:0] = buffer_data_2[1079:1072];
        layer4[9][15:8] = buffer_data_2[1087:1080];
        layer4[9][23:16] = buffer_data_2[1095:1088];
        layer4[9][31:24] = buffer_data_2[1103:1096];
        layer4[9][39:32] = buffer_data_2[1111:1104];
        layer4[9][47:40] = buffer_data_2[1119:1112];
        layer4[9][55:48] = buffer_data_2[1127:1120];
        layer5[9][7:0] = buffer_data_1[1079:1072];
        layer5[9][15:8] = buffer_data_1[1087:1080];
        layer5[9][23:16] = buffer_data_1[1095:1088];
        layer5[9][31:24] = buffer_data_1[1103:1096];
        layer5[9][39:32] = buffer_data_1[1111:1104];
        layer5[9][47:40] = buffer_data_1[1119:1112];
        layer5[9][55:48] = buffer_data_1[1127:1120];
        layer6[9][7:0] = buffer_data_0[1079:1072];
        layer6[9][15:8] = buffer_data_0[1087:1080];
        layer6[9][23:16] = buffer_data_0[1095:1088];
        layer6[9][31:24] = buffer_data_0[1103:1096];
        layer6[9][39:32] = buffer_data_0[1111:1104];
        layer6[9][47:40] = buffer_data_0[1119:1112];
        layer6[9][55:48] = buffer_data_0[1127:1120];
        layer0[10][7:0] = buffer_data_6[1087:1080];
        layer0[10][15:8] = buffer_data_6[1095:1088];
        layer0[10][23:16] = buffer_data_6[1103:1096];
        layer0[10][31:24] = buffer_data_6[1111:1104];
        layer0[10][39:32] = buffer_data_6[1119:1112];
        layer0[10][47:40] = buffer_data_6[1127:1120];
        layer0[10][55:48] = buffer_data_6[1135:1128];
        layer1[10][7:0] = buffer_data_5[1087:1080];
        layer1[10][15:8] = buffer_data_5[1095:1088];
        layer1[10][23:16] = buffer_data_5[1103:1096];
        layer1[10][31:24] = buffer_data_5[1111:1104];
        layer1[10][39:32] = buffer_data_5[1119:1112];
        layer1[10][47:40] = buffer_data_5[1127:1120];
        layer1[10][55:48] = buffer_data_5[1135:1128];
        layer2[10][7:0] = buffer_data_4[1087:1080];
        layer2[10][15:8] = buffer_data_4[1095:1088];
        layer2[10][23:16] = buffer_data_4[1103:1096];
        layer2[10][31:24] = buffer_data_4[1111:1104];
        layer2[10][39:32] = buffer_data_4[1119:1112];
        layer2[10][47:40] = buffer_data_4[1127:1120];
        layer2[10][55:48] = buffer_data_4[1135:1128];
        layer3[10][7:0] = buffer_data_3[1087:1080];
        layer3[10][15:8] = buffer_data_3[1095:1088];
        layer3[10][23:16] = buffer_data_3[1103:1096];
        layer3[10][31:24] = buffer_data_3[1111:1104];
        layer3[10][39:32] = buffer_data_3[1119:1112];
        layer3[10][47:40] = buffer_data_3[1127:1120];
        layer3[10][55:48] = buffer_data_3[1135:1128];
        layer4[10][7:0] = buffer_data_2[1087:1080];
        layer4[10][15:8] = buffer_data_2[1095:1088];
        layer4[10][23:16] = buffer_data_2[1103:1096];
        layer4[10][31:24] = buffer_data_2[1111:1104];
        layer4[10][39:32] = buffer_data_2[1119:1112];
        layer4[10][47:40] = buffer_data_2[1127:1120];
        layer4[10][55:48] = buffer_data_2[1135:1128];
        layer5[10][7:0] = buffer_data_1[1087:1080];
        layer5[10][15:8] = buffer_data_1[1095:1088];
        layer5[10][23:16] = buffer_data_1[1103:1096];
        layer5[10][31:24] = buffer_data_1[1111:1104];
        layer5[10][39:32] = buffer_data_1[1119:1112];
        layer5[10][47:40] = buffer_data_1[1127:1120];
        layer5[10][55:48] = buffer_data_1[1135:1128];
        layer6[10][7:0] = buffer_data_0[1087:1080];
        layer6[10][15:8] = buffer_data_0[1095:1088];
        layer6[10][23:16] = buffer_data_0[1103:1096];
        layer6[10][31:24] = buffer_data_0[1111:1104];
        layer6[10][39:32] = buffer_data_0[1119:1112];
        layer6[10][47:40] = buffer_data_0[1127:1120];
        layer6[10][55:48] = buffer_data_0[1135:1128];
        layer0[11][7:0] = buffer_data_6[1095:1088];
        layer0[11][15:8] = buffer_data_6[1103:1096];
        layer0[11][23:16] = buffer_data_6[1111:1104];
        layer0[11][31:24] = buffer_data_6[1119:1112];
        layer0[11][39:32] = buffer_data_6[1127:1120];
        layer0[11][47:40] = buffer_data_6[1135:1128];
        layer0[11][55:48] = buffer_data_6[1143:1136];
        layer1[11][7:0] = buffer_data_5[1095:1088];
        layer1[11][15:8] = buffer_data_5[1103:1096];
        layer1[11][23:16] = buffer_data_5[1111:1104];
        layer1[11][31:24] = buffer_data_5[1119:1112];
        layer1[11][39:32] = buffer_data_5[1127:1120];
        layer1[11][47:40] = buffer_data_5[1135:1128];
        layer1[11][55:48] = buffer_data_5[1143:1136];
        layer2[11][7:0] = buffer_data_4[1095:1088];
        layer2[11][15:8] = buffer_data_4[1103:1096];
        layer2[11][23:16] = buffer_data_4[1111:1104];
        layer2[11][31:24] = buffer_data_4[1119:1112];
        layer2[11][39:32] = buffer_data_4[1127:1120];
        layer2[11][47:40] = buffer_data_4[1135:1128];
        layer2[11][55:48] = buffer_data_4[1143:1136];
        layer3[11][7:0] = buffer_data_3[1095:1088];
        layer3[11][15:8] = buffer_data_3[1103:1096];
        layer3[11][23:16] = buffer_data_3[1111:1104];
        layer3[11][31:24] = buffer_data_3[1119:1112];
        layer3[11][39:32] = buffer_data_3[1127:1120];
        layer3[11][47:40] = buffer_data_3[1135:1128];
        layer3[11][55:48] = buffer_data_3[1143:1136];
        layer4[11][7:0] = buffer_data_2[1095:1088];
        layer4[11][15:8] = buffer_data_2[1103:1096];
        layer4[11][23:16] = buffer_data_2[1111:1104];
        layer4[11][31:24] = buffer_data_2[1119:1112];
        layer4[11][39:32] = buffer_data_2[1127:1120];
        layer4[11][47:40] = buffer_data_2[1135:1128];
        layer4[11][55:48] = buffer_data_2[1143:1136];
        layer5[11][7:0] = buffer_data_1[1095:1088];
        layer5[11][15:8] = buffer_data_1[1103:1096];
        layer5[11][23:16] = buffer_data_1[1111:1104];
        layer5[11][31:24] = buffer_data_1[1119:1112];
        layer5[11][39:32] = buffer_data_1[1127:1120];
        layer5[11][47:40] = buffer_data_1[1135:1128];
        layer5[11][55:48] = buffer_data_1[1143:1136];
        layer6[11][7:0] = buffer_data_0[1095:1088];
        layer6[11][15:8] = buffer_data_0[1103:1096];
        layer6[11][23:16] = buffer_data_0[1111:1104];
        layer6[11][31:24] = buffer_data_0[1119:1112];
        layer6[11][39:32] = buffer_data_0[1127:1120];
        layer6[11][47:40] = buffer_data_0[1135:1128];
        layer6[11][55:48] = buffer_data_0[1143:1136];
        layer0[12][7:0] = buffer_data_6[1103:1096];
        layer0[12][15:8] = buffer_data_6[1111:1104];
        layer0[12][23:16] = buffer_data_6[1119:1112];
        layer0[12][31:24] = buffer_data_6[1127:1120];
        layer0[12][39:32] = buffer_data_6[1135:1128];
        layer0[12][47:40] = buffer_data_6[1143:1136];
        layer0[12][55:48] = buffer_data_6[1151:1144];
        layer1[12][7:0] = buffer_data_5[1103:1096];
        layer1[12][15:8] = buffer_data_5[1111:1104];
        layer1[12][23:16] = buffer_data_5[1119:1112];
        layer1[12][31:24] = buffer_data_5[1127:1120];
        layer1[12][39:32] = buffer_data_5[1135:1128];
        layer1[12][47:40] = buffer_data_5[1143:1136];
        layer1[12][55:48] = buffer_data_5[1151:1144];
        layer2[12][7:0] = buffer_data_4[1103:1096];
        layer2[12][15:8] = buffer_data_4[1111:1104];
        layer2[12][23:16] = buffer_data_4[1119:1112];
        layer2[12][31:24] = buffer_data_4[1127:1120];
        layer2[12][39:32] = buffer_data_4[1135:1128];
        layer2[12][47:40] = buffer_data_4[1143:1136];
        layer2[12][55:48] = buffer_data_4[1151:1144];
        layer3[12][7:0] = buffer_data_3[1103:1096];
        layer3[12][15:8] = buffer_data_3[1111:1104];
        layer3[12][23:16] = buffer_data_3[1119:1112];
        layer3[12][31:24] = buffer_data_3[1127:1120];
        layer3[12][39:32] = buffer_data_3[1135:1128];
        layer3[12][47:40] = buffer_data_3[1143:1136];
        layer3[12][55:48] = buffer_data_3[1151:1144];
        layer4[12][7:0] = buffer_data_2[1103:1096];
        layer4[12][15:8] = buffer_data_2[1111:1104];
        layer4[12][23:16] = buffer_data_2[1119:1112];
        layer4[12][31:24] = buffer_data_2[1127:1120];
        layer4[12][39:32] = buffer_data_2[1135:1128];
        layer4[12][47:40] = buffer_data_2[1143:1136];
        layer4[12][55:48] = buffer_data_2[1151:1144];
        layer5[12][7:0] = buffer_data_1[1103:1096];
        layer5[12][15:8] = buffer_data_1[1111:1104];
        layer5[12][23:16] = buffer_data_1[1119:1112];
        layer5[12][31:24] = buffer_data_1[1127:1120];
        layer5[12][39:32] = buffer_data_1[1135:1128];
        layer5[12][47:40] = buffer_data_1[1143:1136];
        layer5[12][55:48] = buffer_data_1[1151:1144];
        layer6[12][7:0] = buffer_data_0[1103:1096];
        layer6[12][15:8] = buffer_data_0[1111:1104];
        layer6[12][23:16] = buffer_data_0[1119:1112];
        layer6[12][31:24] = buffer_data_0[1127:1120];
        layer6[12][39:32] = buffer_data_0[1135:1128];
        layer6[12][47:40] = buffer_data_0[1143:1136];
        layer6[12][55:48] = buffer_data_0[1151:1144];
        layer0[13][7:0] = buffer_data_6[1111:1104];
        layer0[13][15:8] = buffer_data_6[1119:1112];
        layer0[13][23:16] = buffer_data_6[1127:1120];
        layer0[13][31:24] = buffer_data_6[1135:1128];
        layer0[13][39:32] = buffer_data_6[1143:1136];
        layer0[13][47:40] = buffer_data_6[1151:1144];
        layer0[13][55:48] = buffer_data_6[1159:1152];
        layer1[13][7:0] = buffer_data_5[1111:1104];
        layer1[13][15:8] = buffer_data_5[1119:1112];
        layer1[13][23:16] = buffer_data_5[1127:1120];
        layer1[13][31:24] = buffer_data_5[1135:1128];
        layer1[13][39:32] = buffer_data_5[1143:1136];
        layer1[13][47:40] = buffer_data_5[1151:1144];
        layer1[13][55:48] = buffer_data_5[1159:1152];
        layer2[13][7:0] = buffer_data_4[1111:1104];
        layer2[13][15:8] = buffer_data_4[1119:1112];
        layer2[13][23:16] = buffer_data_4[1127:1120];
        layer2[13][31:24] = buffer_data_4[1135:1128];
        layer2[13][39:32] = buffer_data_4[1143:1136];
        layer2[13][47:40] = buffer_data_4[1151:1144];
        layer2[13][55:48] = buffer_data_4[1159:1152];
        layer3[13][7:0] = buffer_data_3[1111:1104];
        layer3[13][15:8] = buffer_data_3[1119:1112];
        layer3[13][23:16] = buffer_data_3[1127:1120];
        layer3[13][31:24] = buffer_data_3[1135:1128];
        layer3[13][39:32] = buffer_data_3[1143:1136];
        layer3[13][47:40] = buffer_data_3[1151:1144];
        layer3[13][55:48] = buffer_data_3[1159:1152];
        layer4[13][7:0] = buffer_data_2[1111:1104];
        layer4[13][15:8] = buffer_data_2[1119:1112];
        layer4[13][23:16] = buffer_data_2[1127:1120];
        layer4[13][31:24] = buffer_data_2[1135:1128];
        layer4[13][39:32] = buffer_data_2[1143:1136];
        layer4[13][47:40] = buffer_data_2[1151:1144];
        layer4[13][55:48] = buffer_data_2[1159:1152];
        layer5[13][7:0] = buffer_data_1[1111:1104];
        layer5[13][15:8] = buffer_data_1[1119:1112];
        layer5[13][23:16] = buffer_data_1[1127:1120];
        layer5[13][31:24] = buffer_data_1[1135:1128];
        layer5[13][39:32] = buffer_data_1[1143:1136];
        layer5[13][47:40] = buffer_data_1[1151:1144];
        layer5[13][55:48] = buffer_data_1[1159:1152];
        layer6[13][7:0] = buffer_data_0[1111:1104];
        layer6[13][15:8] = buffer_data_0[1119:1112];
        layer6[13][23:16] = buffer_data_0[1127:1120];
        layer6[13][31:24] = buffer_data_0[1135:1128];
        layer6[13][39:32] = buffer_data_0[1143:1136];
        layer6[13][47:40] = buffer_data_0[1151:1144];
        layer6[13][55:48] = buffer_data_0[1159:1152];
        layer0[14][7:0] = buffer_data_6[1119:1112];
        layer0[14][15:8] = buffer_data_6[1127:1120];
        layer0[14][23:16] = buffer_data_6[1135:1128];
        layer0[14][31:24] = buffer_data_6[1143:1136];
        layer0[14][39:32] = buffer_data_6[1151:1144];
        layer0[14][47:40] = buffer_data_6[1159:1152];
        layer0[14][55:48] = buffer_data_6[1167:1160];
        layer1[14][7:0] = buffer_data_5[1119:1112];
        layer1[14][15:8] = buffer_data_5[1127:1120];
        layer1[14][23:16] = buffer_data_5[1135:1128];
        layer1[14][31:24] = buffer_data_5[1143:1136];
        layer1[14][39:32] = buffer_data_5[1151:1144];
        layer1[14][47:40] = buffer_data_5[1159:1152];
        layer1[14][55:48] = buffer_data_5[1167:1160];
        layer2[14][7:0] = buffer_data_4[1119:1112];
        layer2[14][15:8] = buffer_data_4[1127:1120];
        layer2[14][23:16] = buffer_data_4[1135:1128];
        layer2[14][31:24] = buffer_data_4[1143:1136];
        layer2[14][39:32] = buffer_data_4[1151:1144];
        layer2[14][47:40] = buffer_data_4[1159:1152];
        layer2[14][55:48] = buffer_data_4[1167:1160];
        layer3[14][7:0] = buffer_data_3[1119:1112];
        layer3[14][15:8] = buffer_data_3[1127:1120];
        layer3[14][23:16] = buffer_data_3[1135:1128];
        layer3[14][31:24] = buffer_data_3[1143:1136];
        layer3[14][39:32] = buffer_data_3[1151:1144];
        layer3[14][47:40] = buffer_data_3[1159:1152];
        layer3[14][55:48] = buffer_data_3[1167:1160];
        layer4[14][7:0] = buffer_data_2[1119:1112];
        layer4[14][15:8] = buffer_data_2[1127:1120];
        layer4[14][23:16] = buffer_data_2[1135:1128];
        layer4[14][31:24] = buffer_data_2[1143:1136];
        layer4[14][39:32] = buffer_data_2[1151:1144];
        layer4[14][47:40] = buffer_data_2[1159:1152];
        layer4[14][55:48] = buffer_data_2[1167:1160];
        layer5[14][7:0] = buffer_data_1[1119:1112];
        layer5[14][15:8] = buffer_data_1[1127:1120];
        layer5[14][23:16] = buffer_data_1[1135:1128];
        layer5[14][31:24] = buffer_data_1[1143:1136];
        layer5[14][39:32] = buffer_data_1[1151:1144];
        layer5[14][47:40] = buffer_data_1[1159:1152];
        layer5[14][55:48] = buffer_data_1[1167:1160];
        layer6[14][7:0] = buffer_data_0[1119:1112];
        layer6[14][15:8] = buffer_data_0[1127:1120];
        layer6[14][23:16] = buffer_data_0[1135:1128];
        layer6[14][31:24] = buffer_data_0[1143:1136];
        layer6[14][39:32] = buffer_data_0[1151:1144];
        layer6[14][47:40] = buffer_data_0[1159:1152];
        layer6[14][55:48] = buffer_data_0[1167:1160];
        layer0[15][7:0] = buffer_data_6[1127:1120];
        layer0[15][15:8] = buffer_data_6[1135:1128];
        layer0[15][23:16] = buffer_data_6[1143:1136];
        layer0[15][31:24] = buffer_data_6[1151:1144];
        layer0[15][39:32] = buffer_data_6[1159:1152];
        layer0[15][47:40] = buffer_data_6[1167:1160];
        layer0[15][55:48] = buffer_data_6[1175:1168];
        layer1[15][7:0] = buffer_data_5[1127:1120];
        layer1[15][15:8] = buffer_data_5[1135:1128];
        layer1[15][23:16] = buffer_data_5[1143:1136];
        layer1[15][31:24] = buffer_data_5[1151:1144];
        layer1[15][39:32] = buffer_data_5[1159:1152];
        layer1[15][47:40] = buffer_data_5[1167:1160];
        layer1[15][55:48] = buffer_data_5[1175:1168];
        layer2[15][7:0] = buffer_data_4[1127:1120];
        layer2[15][15:8] = buffer_data_4[1135:1128];
        layer2[15][23:16] = buffer_data_4[1143:1136];
        layer2[15][31:24] = buffer_data_4[1151:1144];
        layer2[15][39:32] = buffer_data_4[1159:1152];
        layer2[15][47:40] = buffer_data_4[1167:1160];
        layer2[15][55:48] = buffer_data_4[1175:1168];
        layer3[15][7:0] = buffer_data_3[1127:1120];
        layer3[15][15:8] = buffer_data_3[1135:1128];
        layer3[15][23:16] = buffer_data_3[1143:1136];
        layer3[15][31:24] = buffer_data_3[1151:1144];
        layer3[15][39:32] = buffer_data_3[1159:1152];
        layer3[15][47:40] = buffer_data_3[1167:1160];
        layer3[15][55:48] = buffer_data_3[1175:1168];
        layer4[15][7:0] = buffer_data_2[1127:1120];
        layer4[15][15:8] = buffer_data_2[1135:1128];
        layer4[15][23:16] = buffer_data_2[1143:1136];
        layer4[15][31:24] = buffer_data_2[1151:1144];
        layer4[15][39:32] = buffer_data_2[1159:1152];
        layer4[15][47:40] = buffer_data_2[1167:1160];
        layer4[15][55:48] = buffer_data_2[1175:1168];
        layer5[15][7:0] = buffer_data_1[1127:1120];
        layer5[15][15:8] = buffer_data_1[1135:1128];
        layer5[15][23:16] = buffer_data_1[1143:1136];
        layer5[15][31:24] = buffer_data_1[1151:1144];
        layer5[15][39:32] = buffer_data_1[1159:1152];
        layer5[15][47:40] = buffer_data_1[1167:1160];
        layer5[15][55:48] = buffer_data_1[1175:1168];
        layer6[15][7:0] = buffer_data_0[1127:1120];
        layer6[15][15:8] = buffer_data_0[1135:1128];
        layer6[15][23:16] = buffer_data_0[1143:1136];
        layer6[15][31:24] = buffer_data_0[1151:1144];
        layer6[15][39:32] = buffer_data_0[1159:1152];
        layer6[15][47:40] = buffer_data_0[1167:1160];
        layer6[15][55:48] = buffer_data_0[1175:1168];
        layer0[16][7:0] = buffer_data_6[1135:1128];
        layer0[16][15:8] = buffer_data_6[1143:1136];
        layer0[16][23:16] = buffer_data_6[1151:1144];
        layer0[16][31:24] = buffer_data_6[1159:1152];
        layer0[16][39:32] = buffer_data_6[1167:1160];
        layer0[16][47:40] = buffer_data_6[1175:1168];
        layer0[16][55:48] = buffer_data_6[1183:1176];
        layer1[16][7:0] = buffer_data_5[1135:1128];
        layer1[16][15:8] = buffer_data_5[1143:1136];
        layer1[16][23:16] = buffer_data_5[1151:1144];
        layer1[16][31:24] = buffer_data_5[1159:1152];
        layer1[16][39:32] = buffer_data_5[1167:1160];
        layer1[16][47:40] = buffer_data_5[1175:1168];
        layer1[16][55:48] = buffer_data_5[1183:1176];
        layer2[16][7:0] = buffer_data_4[1135:1128];
        layer2[16][15:8] = buffer_data_4[1143:1136];
        layer2[16][23:16] = buffer_data_4[1151:1144];
        layer2[16][31:24] = buffer_data_4[1159:1152];
        layer2[16][39:32] = buffer_data_4[1167:1160];
        layer2[16][47:40] = buffer_data_4[1175:1168];
        layer2[16][55:48] = buffer_data_4[1183:1176];
        layer3[16][7:0] = buffer_data_3[1135:1128];
        layer3[16][15:8] = buffer_data_3[1143:1136];
        layer3[16][23:16] = buffer_data_3[1151:1144];
        layer3[16][31:24] = buffer_data_3[1159:1152];
        layer3[16][39:32] = buffer_data_3[1167:1160];
        layer3[16][47:40] = buffer_data_3[1175:1168];
        layer3[16][55:48] = buffer_data_3[1183:1176];
        layer4[16][7:0] = buffer_data_2[1135:1128];
        layer4[16][15:8] = buffer_data_2[1143:1136];
        layer4[16][23:16] = buffer_data_2[1151:1144];
        layer4[16][31:24] = buffer_data_2[1159:1152];
        layer4[16][39:32] = buffer_data_2[1167:1160];
        layer4[16][47:40] = buffer_data_2[1175:1168];
        layer4[16][55:48] = buffer_data_2[1183:1176];
        layer5[16][7:0] = buffer_data_1[1135:1128];
        layer5[16][15:8] = buffer_data_1[1143:1136];
        layer5[16][23:16] = buffer_data_1[1151:1144];
        layer5[16][31:24] = buffer_data_1[1159:1152];
        layer5[16][39:32] = buffer_data_1[1167:1160];
        layer5[16][47:40] = buffer_data_1[1175:1168];
        layer5[16][55:48] = buffer_data_1[1183:1176];
        layer6[16][7:0] = buffer_data_0[1135:1128];
        layer6[16][15:8] = buffer_data_0[1143:1136];
        layer6[16][23:16] = buffer_data_0[1151:1144];
        layer6[16][31:24] = buffer_data_0[1159:1152];
        layer6[16][39:32] = buffer_data_0[1167:1160];
        layer6[16][47:40] = buffer_data_0[1175:1168];
        layer6[16][55:48] = buffer_data_0[1183:1176];
        layer0[17][7:0] = buffer_data_6[1143:1136];
        layer0[17][15:8] = buffer_data_6[1151:1144];
        layer0[17][23:16] = buffer_data_6[1159:1152];
        layer0[17][31:24] = buffer_data_6[1167:1160];
        layer0[17][39:32] = buffer_data_6[1175:1168];
        layer0[17][47:40] = buffer_data_6[1183:1176];
        layer0[17][55:48] = buffer_data_6[1191:1184];
        layer1[17][7:0] = buffer_data_5[1143:1136];
        layer1[17][15:8] = buffer_data_5[1151:1144];
        layer1[17][23:16] = buffer_data_5[1159:1152];
        layer1[17][31:24] = buffer_data_5[1167:1160];
        layer1[17][39:32] = buffer_data_5[1175:1168];
        layer1[17][47:40] = buffer_data_5[1183:1176];
        layer1[17][55:48] = buffer_data_5[1191:1184];
        layer2[17][7:0] = buffer_data_4[1143:1136];
        layer2[17][15:8] = buffer_data_4[1151:1144];
        layer2[17][23:16] = buffer_data_4[1159:1152];
        layer2[17][31:24] = buffer_data_4[1167:1160];
        layer2[17][39:32] = buffer_data_4[1175:1168];
        layer2[17][47:40] = buffer_data_4[1183:1176];
        layer2[17][55:48] = buffer_data_4[1191:1184];
        layer3[17][7:0] = buffer_data_3[1143:1136];
        layer3[17][15:8] = buffer_data_3[1151:1144];
        layer3[17][23:16] = buffer_data_3[1159:1152];
        layer3[17][31:24] = buffer_data_3[1167:1160];
        layer3[17][39:32] = buffer_data_3[1175:1168];
        layer3[17][47:40] = buffer_data_3[1183:1176];
        layer3[17][55:48] = buffer_data_3[1191:1184];
        layer4[17][7:0] = buffer_data_2[1143:1136];
        layer4[17][15:8] = buffer_data_2[1151:1144];
        layer4[17][23:16] = buffer_data_2[1159:1152];
        layer4[17][31:24] = buffer_data_2[1167:1160];
        layer4[17][39:32] = buffer_data_2[1175:1168];
        layer4[17][47:40] = buffer_data_2[1183:1176];
        layer4[17][55:48] = buffer_data_2[1191:1184];
        layer5[17][7:0] = buffer_data_1[1143:1136];
        layer5[17][15:8] = buffer_data_1[1151:1144];
        layer5[17][23:16] = buffer_data_1[1159:1152];
        layer5[17][31:24] = buffer_data_1[1167:1160];
        layer5[17][39:32] = buffer_data_1[1175:1168];
        layer5[17][47:40] = buffer_data_1[1183:1176];
        layer5[17][55:48] = buffer_data_1[1191:1184];
        layer6[17][7:0] = buffer_data_0[1143:1136];
        layer6[17][15:8] = buffer_data_0[1151:1144];
        layer6[17][23:16] = buffer_data_0[1159:1152];
        layer6[17][31:24] = buffer_data_0[1167:1160];
        layer6[17][39:32] = buffer_data_0[1175:1168];
        layer6[17][47:40] = buffer_data_0[1183:1176];
        layer6[17][55:48] = buffer_data_0[1191:1184];
        layer0[18][7:0] = buffer_data_6[1151:1144];
        layer0[18][15:8] = buffer_data_6[1159:1152];
        layer0[18][23:16] = buffer_data_6[1167:1160];
        layer0[18][31:24] = buffer_data_6[1175:1168];
        layer0[18][39:32] = buffer_data_6[1183:1176];
        layer0[18][47:40] = buffer_data_6[1191:1184];
        layer0[18][55:48] = buffer_data_6[1199:1192];
        layer1[18][7:0] = buffer_data_5[1151:1144];
        layer1[18][15:8] = buffer_data_5[1159:1152];
        layer1[18][23:16] = buffer_data_5[1167:1160];
        layer1[18][31:24] = buffer_data_5[1175:1168];
        layer1[18][39:32] = buffer_data_5[1183:1176];
        layer1[18][47:40] = buffer_data_5[1191:1184];
        layer1[18][55:48] = buffer_data_5[1199:1192];
        layer2[18][7:0] = buffer_data_4[1151:1144];
        layer2[18][15:8] = buffer_data_4[1159:1152];
        layer2[18][23:16] = buffer_data_4[1167:1160];
        layer2[18][31:24] = buffer_data_4[1175:1168];
        layer2[18][39:32] = buffer_data_4[1183:1176];
        layer2[18][47:40] = buffer_data_4[1191:1184];
        layer2[18][55:48] = buffer_data_4[1199:1192];
        layer3[18][7:0] = buffer_data_3[1151:1144];
        layer3[18][15:8] = buffer_data_3[1159:1152];
        layer3[18][23:16] = buffer_data_3[1167:1160];
        layer3[18][31:24] = buffer_data_3[1175:1168];
        layer3[18][39:32] = buffer_data_3[1183:1176];
        layer3[18][47:40] = buffer_data_3[1191:1184];
        layer3[18][55:48] = buffer_data_3[1199:1192];
        layer4[18][7:0] = buffer_data_2[1151:1144];
        layer4[18][15:8] = buffer_data_2[1159:1152];
        layer4[18][23:16] = buffer_data_2[1167:1160];
        layer4[18][31:24] = buffer_data_2[1175:1168];
        layer4[18][39:32] = buffer_data_2[1183:1176];
        layer4[18][47:40] = buffer_data_2[1191:1184];
        layer4[18][55:48] = buffer_data_2[1199:1192];
        layer5[18][7:0] = buffer_data_1[1151:1144];
        layer5[18][15:8] = buffer_data_1[1159:1152];
        layer5[18][23:16] = buffer_data_1[1167:1160];
        layer5[18][31:24] = buffer_data_1[1175:1168];
        layer5[18][39:32] = buffer_data_1[1183:1176];
        layer5[18][47:40] = buffer_data_1[1191:1184];
        layer5[18][55:48] = buffer_data_1[1199:1192];
        layer6[18][7:0] = buffer_data_0[1151:1144];
        layer6[18][15:8] = buffer_data_0[1159:1152];
        layer6[18][23:16] = buffer_data_0[1167:1160];
        layer6[18][31:24] = buffer_data_0[1175:1168];
        layer6[18][39:32] = buffer_data_0[1183:1176];
        layer6[18][47:40] = buffer_data_0[1191:1184];
        layer6[18][55:48] = buffer_data_0[1199:1192];
        layer0[19][7:0] = buffer_data_6[1159:1152];
        layer0[19][15:8] = buffer_data_6[1167:1160];
        layer0[19][23:16] = buffer_data_6[1175:1168];
        layer0[19][31:24] = buffer_data_6[1183:1176];
        layer0[19][39:32] = buffer_data_6[1191:1184];
        layer0[19][47:40] = buffer_data_6[1199:1192];
        layer0[19][55:48] = buffer_data_6[1207:1200];
        layer1[19][7:0] = buffer_data_5[1159:1152];
        layer1[19][15:8] = buffer_data_5[1167:1160];
        layer1[19][23:16] = buffer_data_5[1175:1168];
        layer1[19][31:24] = buffer_data_5[1183:1176];
        layer1[19][39:32] = buffer_data_5[1191:1184];
        layer1[19][47:40] = buffer_data_5[1199:1192];
        layer1[19][55:48] = buffer_data_5[1207:1200];
        layer2[19][7:0] = buffer_data_4[1159:1152];
        layer2[19][15:8] = buffer_data_4[1167:1160];
        layer2[19][23:16] = buffer_data_4[1175:1168];
        layer2[19][31:24] = buffer_data_4[1183:1176];
        layer2[19][39:32] = buffer_data_4[1191:1184];
        layer2[19][47:40] = buffer_data_4[1199:1192];
        layer2[19][55:48] = buffer_data_4[1207:1200];
        layer3[19][7:0] = buffer_data_3[1159:1152];
        layer3[19][15:8] = buffer_data_3[1167:1160];
        layer3[19][23:16] = buffer_data_3[1175:1168];
        layer3[19][31:24] = buffer_data_3[1183:1176];
        layer3[19][39:32] = buffer_data_3[1191:1184];
        layer3[19][47:40] = buffer_data_3[1199:1192];
        layer3[19][55:48] = buffer_data_3[1207:1200];
        layer4[19][7:0] = buffer_data_2[1159:1152];
        layer4[19][15:8] = buffer_data_2[1167:1160];
        layer4[19][23:16] = buffer_data_2[1175:1168];
        layer4[19][31:24] = buffer_data_2[1183:1176];
        layer4[19][39:32] = buffer_data_2[1191:1184];
        layer4[19][47:40] = buffer_data_2[1199:1192];
        layer4[19][55:48] = buffer_data_2[1207:1200];
        layer5[19][7:0] = buffer_data_1[1159:1152];
        layer5[19][15:8] = buffer_data_1[1167:1160];
        layer5[19][23:16] = buffer_data_1[1175:1168];
        layer5[19][31:24] = buffer_data_1[1183:1176];
        layer5[19][39:32] = buffer_data_1[1191:1184];
        layer5[19][47:40] = buffer_data_1[1199:1192];
        layer5[19][55:48] = buffer_data_1[1207:1200];
        layer6[19][7:0] = buffer_data_0[1159:1152];
        layer6[19][15:8] = buffer_data_0[1167:1160];
        layer6[19][23:16] = buffer_data_0[1175:1168];
        layer6[19][31:24] = buffer_data_0[1183:1176];
        layer6[19][39:32] = buffer_data_0[1191:1184];
        layer6[19][47:40] = buffer_data_0[1199:1192];
        layer6[19][55:48] = buffer_data_0[1207:1200];
        layer0[20][7:0] = buffer_data_6[1167:1160];
        layer0[20][15:8] = buffer_data_6[1175:1168];
        layer0[20][23:16] = buffer_data_6[1183:1176];
        layer0[20][31:24] = buffer_data_6[1191:1184];
        layer0[20][39:32] = buffer_data_6[1199:1192];
        layer0[20][47:40] = buffer_data_6[1207:1200];
        layer0[20][55:48] = buffer_data_6[1215:1208];
        layer1[20][7:0] = buffer_data_5[1167:1160];
        layer1[20][15:8] = buffer_data_5[1175:1168];
        layer1[20][23:16] = buffer_data_5[1183:1176];
        layer1[20][31:24] = buffer_data_5[1191:1184];
        layer1[20][39:32] = buffer_data_5[1199:1192];
        layer1[20][47:40] = buffer_data_5[1207:1200];
        layer1[20][55:48] = buffer_data_5[1215:1208];
        layer2[20][7:0] = buffer_data_4[1167:1160];
        layer2[20][15:8] = buffer_data_4[1175:1168];
        layer2[20][23:16] = buffer_data_4[1183:1176];
        layer2[20][31:24] = buffer_data_4[1191:1184];
        layer2[20][39:32] = buffer_data_4[1199:1192];
        layer2[20][47:40] = buffer_data_4[1207:1200];
        layer2[20][55:48] = buffer_data_4[1215:1208];
        layer3[20][7:0] = buffer_data_3[1167:1160];
        layer3[20][15:8] = buffer_data_3[1175:1168];
        layer3[20][23:16] = buffer_data_3[1183:1176];
        layer3[20][31:24] = buffer_data_3[1191:1184];
        layer3[20][39:32] = buffer_data_3[1199:1192];
        layer3[20][47:40] = buffer_data_3[1207:1200];
        layer3[20][55:48] = buffer_data_3[1215:1208];
        layer4[20][7:0] = buffer_data_2[1167:1160];
        layer4[20][15:8] = buffer_data_2[1175:1168];
        layer4[20][23:16] = buffer_data_2[1183:1176];
        layer4[20][31:24] = buffer_data_2[1191:1184];
        layer4[20][39:32] = buffer_data_2[1199:1192];
        layer4[20][47:40] = buffer_data_2[1207:1200];
        layer4[20][55:48] = buffer_data_2[1215:1208];
        layer5[20][7:0] = buffer_data_1[1167:1160];
        layer5[20][15:8] = buffer_data_1[1175:1168];
        layer5[20][23:16] = buffer_data_1[1183:1176];
        layer5[20][31:24] = buffer_data_1[1191:1184];
        layer5[20][39:32] = buffer_data_1[1199:1192];
        layer5[20][47:40] = buffer_data_1[1207:1200];
        layer5[20][55:48] = buffer_data_1[1215:1208];
        layer6[20][7:0] = buffer_data_0[1167:1160];
        layer6[20][15:8] = buffer_data_0[1175:1168];
        layer6[20][23:16] = buffer_data_0[1183:1176];
        layer6[20][31:24] = buffer_data_0[1191:1184];
        layer6[20][39:32] = buffer_data_0[1199:1192];
        layer6[20][47:40] = buffer_data_0[1207:1200];
        layer6[20][55:48] = buffer_data_0[1215:1208];
        layer0[21][7:0] = buffer_data_6[1175:1168];
        layer0[21][15:8] = buffer_data_6[1183:1176];
        layer0[21][23:16] = buffer_data_6[1191:1184];
        layer0[21][31:24] = buffer_data_6[1199:1192];
        layer0[21][39:32] = buffer_data_6[1207:1200];
        layer0[21][47:40] = buffer_data_6[1215:1208];
        layer0[21][55:48] = buffer_data_6[1223:1216];
        layer1[21][7:0] = buffer_data_5[1175:1168];
        layer1[21][15:8] = buffer_data_5[1183:1176];
        layer1[21][23:16] = buffer_data_5[1191:1184];
        layer1[21][31:24] = buffer_data_5[1199:1192];
        layer1[21][39:32] = buffer_data_5[1207:1200];
        layer1[21][47:40] = buffer_data_5[1215:1208];
        layer1[21][55:48] = buffer_data_5[1223:1216];
        layer2[21][7:0] = buffer_data_4[1175:1168];
        layer2[21][15:8] = buffer_data_4[1183:1176];
        layer2[21][23:16] = buffer_data_4[1191:1184];
        layer2[21][31:24] = buffer_data_4[1199:1192];
        layer2[21][39:32] = buffer_data_4[1207:1200];
        layer2[21][47:40] = buffer_data_4[1215:1208];
        layer2[21][55:48] = buffer_data_4[1223:1216];
        layer3[21][7:0] = buffer_data_3[1175:1168];
        layer3[21][15:8] = buffer_data_3[1183:1176];
        layer3[21][23:16] = buffer_data_3[1191:1184];
        layer3[21][31:24] = buffer_data_3[1199:1192];
        layer3[21][39:32] = buffer_data_3[1207:1200];
        layer3[21][47:40] = buffer_data_3[1215:1208];
        layer3[21][55:48] = buffer_data_3[1223:1216];
        layer4[21][7:0] = buffer_data_2[1175:1168];
        layer4[21][15:8] = buffer_data_2[1183:1176];
        layer4[21][23:16] = buffer_data_2[1191:1184];
        layer4[21][31:24] = buffer_data_2[1199:1192];
        layer4[21][39:32] = buffer_data_2[1207:1200];
        layer4[21][47:40] = buffer_data_2[1215:1208];
        layer4[21][55:48] = buffer_data_2[1223:1216];
        layer5[21][7:0] = buffer_data_1[1175:1168];
        layer5[21][15:8] = buffer_data_1[1183:1176];
        layer5[21][23:16] = buffer_data_1[1191:1184];
        layer5[21][31:24] = buffer_data_1[1199:1192];
        layer5[21][39:32] = buffer_data_1[1207:1200];
        layer5[21][47:40] = buffer_data_1[1215:1208];
        layer5[21][55:48] = buffer_data_1[1223:1216];
        layer6[21][7:0] = buffer_data_0[1175:1168];
        layer6[21][15:8] = buffer_data_0[1183:1176];
        layer6[21][23:16] = buffer_data_0[1191:1184];
        layer6[21][31:24] = buffer_data_0[1199:1192];
        layer6[21][39:32] = buffer_data_0[1207:1200];
        layer6[21][47:40] = buffer_data_0[1215:1208];
        layer6[21][55:48] = buffer_data_0[1223:1216];
        layer0[22][7:0] = buffer_data_6[1183:1176];
        layer0[22][15:8] = buffer_data_6[1191:1184];
        layer0[22][23:16] = buffer_data_6[1199:1192];
        layer0[22][31:24] = buffer_data_6[1207:1200];
        layer0[22][39:32] = buffer_data_6[1215:1208];
        layer0[22][47:40] = buffer_data_6[1223:1216];
        layer0[22][55:48] = buffer_data_6[1231:1224];
        layer1[22][7:0] = buffer_data_5[1183:1176];
        layer1[22][15:8] = buffer_data_5[1191:1184];
        layer1[22][23:16] = buffer_data_5[1199:1192];
        layer1[22][31:24] = buffer_data_5[1207:1200];
        layer1[22][39:32] = buffer_data_5[1215:1208];
        layer1[22][47:40] = buffer_data_5[1223:1216];
        layer1[22][55:48] = buffer_data_5[1231:1224];
        layer2[22][7:0] = buffer_data_4[1183:1176];
        layer2[22][15:8] = buffer_data_4[1191:1184];
        layer2[22][23:16] = buffer_data_4[1199:1192];
        layer2[22][31:24] = buffer_data_4[1207:1200];
        layer2[22][39:32] = buffer_data_4[1215:1208];
        layer2[22][47:40] = buffer_data_4[1223:1216];
        layer2[22][55:48] = buffer_data_4[1231:1224];
        layer3[22][7:0] = buffer_data_3[1183:1176];
        layer3[22][15:8] = buffer_data_3[1191:1184];
        layer3[22][23:16] = buffer_data_3[1199:1192];
        layer3[22][31:24] = buffer_data_3[1207:1200];
        layer3[22][39:32] = buffer_data_3[1215:1208];
        layer3[22][47:40] = buffer_data_3[1223:1216];
        layer3[22][55:48] = buffer_data_3[1231:1224];
        layer4[22][7:0] = buffer_data_2[1183:1176];
        layer4[22][15:8] = buffer_data_2[1191:1184];
        layer4[22][23:16] = buffer_data_2[1199:1192];
        layer4[22][31:24] = buffer_data_2[1207:1200];
        layer4[22][39:32] = buffer_data_2[1215:1208];
        layer4[22][47:40] = buffer_data_2[1223:1216];
        layer4[22][55:48] = buffer_data_2[1231:1224];
        layer5[22][7:0] = buffer_data_1[1183:1176];
        layer5[22][15:8] = buffer_data_1[1191:1184];
        layer5[22][23:16] = buffer_data_1[1199:1192];
        layer5[22][31:24] = buffer_data_1[1207:1200];
        layer5[22][39:32] = buffer_data_1[1215:1208];
        layer5[22][47:40] = buffer_data_1[1223:1216];
        layer5[22][55:48] = buffer_data_1[1231:1224];
        layer6[22][7:0] = buffer_data_0[1183:1176];
        layer6[22][15:8] = buffer_data_0[1191:1184];
        layer6[22][23:16] = buffer_data_0[1199:1192];
        layer6[22][31:24] = buffer_data_0[1207:1200];
        layer6[22][39:32] = buffer_data_0[1215:1208];
        layer6[22][47:40] = buffer_data_0[1223:1216];
        layer6[22][55:48] = buffer_data_0[1231:1224];
        layer0[23][7:0] = buffer_data_6[1191:1184];
        layer0[23][15:8] = buffer_data_6[1199:1192];
        layer0[23][23:16] = buffer_data_6[1207:1200];
        layer0[23][31:24] = buffer_data_6[1215:1208];
        layer0[23][39:32] = buffer_data_6[1223:1216];
        layer0[23][47:40] = buffer_data_6[1231:1224];
        layer0[23][55:48] = buffer_data_6[1239:1232];
        layer1[23][7:0] = buffer_data_5[1191:1184];
        layer1[23][15:8] = buffer_data_5[1199:1192];
        layer1[23][23:16] = buffer_data_5[1207:1200];
        layer1[23][31:24] = buffer_data_5[1215:1208];
        layer1[23][39:32] = buffer_data_5[1223:1216];
        layer1[23][47:40] = buffer_data_5[1231:1224];
        layer1[23][55:48] = buffer_data_5[1239:1232];
        layer2[23][7:0] = buffer_data_4[1191:1184];
        layer2[23][15:8] = buffer_data_4[1199:1192];
        layer2[23][23:16] = buffer_data_4[1207:1200];
        layer2[23][31:24] = buffer_data_4[1215:1208];
        layer2[23][39:32] = buffer_data_4[1223:1216];
        layer2[23][47:40] = buffer_data_4[1231:1224];
        layer2[23][55:48] = buffer_data_4[1239:1232];
        layer3[23][7:0] = buffer_data_3[1191:1184];
        layer3[23][15:8] = buffer_data_3[1199:1192];
        layer3[23][23:16] = buffer_data_3[1207:1200];
        layer3[23][31:24] = buffer_data_3[1215:1208];
        layer3[23][39:32] = buffer_data_3[1223:1216];
        layer3[23][47:40] = buffer_data_3[1231:1224];
        layer3[23][55:48] = buffer_data_3[1239:1232];
        layer4[23][7:0] = buffer_data_2[1191:1184];
        layer4[23][15:8] = buffer_data_2[1199:1192];
        layer4[23][23:16] = buffer_data_2[1207:1200];
        layer4[23][31:24] = buffer_data_2[1215:1208];
        layer4[23][39:32] = buffer_data_2[1223:1216];
        layer4[23][47:40] = buffer_data_2[1231:1224];
        layer4[23][55:48] = buffer_data_2[1239:1232];
        layer5[23][7:0] = buffer_data_1[1191:1184];
        layer5[23][15:8] = buffer_data_1[1199:1192];
        layer5[23][23:16] = buffer_data_1[1207:1200];
        layer5[23][31:24] = buffer_data_1[1215:1208];
        layer5[23][39:32] = buffer_data_1[1223:1216];
        layer5[23][47:40] = buffer_data_1[1231:1224];
        layer5[23][55:48] = buffer_data_1[1239:1232];
        layer6[23][7:0] = buffer_data_0[1191:1184];
        layer6[23][15:8] = buffer_data_0[1199:1192];
        layer6[23][23:16] = buffer_data_0[1207:1200];
        layer6[23][31:24] = buffer_data_0[1215:1208];
        layer6[23][39:32] = buffer_data_0[1223:1216];
        layer6[23][47:40] = buffer_data_0[1231:1224];
        layer6[23][55:48] = buffer_data_0[1239:1232];
        layer0[24][7:0] = buffer_data_6[1199:1192];
        layer0[24][15:8] = buffer_data_6[1207:1200];
        layer0[24][23:16] = buffer_data_6[1215:1208];
        layer0[24][31:24] = buffer_data_6[1223:1216];
        layer0[24][39:32] = buffer_data_6[1231:1224];
        layer0[24][47:40] = buffer_data_6[1239:1232];
        layer0[24][55:48] = buffer_data_6[1247:1240];
        layer1[24][7:0] = buffer_data_5[1199:1192];
        layer1[24][15:8] = buffer_data_5[1207:1200];
        layer1[24][23:16] = buffer_data_5[1215:1208];
        layer1[24][31:24] = buffer_data_5[1223:1216];
        layer1[24][39:32] = buffer_data_5[1231:1224];
        layer1[24][47:40] = buffer_data_5[1239:1232];
        layer1[24][55:48] = buffer_data_5[1247:1240];
        layer2[24][7:0] = buffer_data_4[1199:1192];
        layer2[24][15:8] = buffer_data_4[1207:1200];
        layer2[24][23:16] = buffer_data_4[1215:1208];
        layer2[24][31:24] = buffer_data_4[1223:1216];
        layer2[24][39:32] = buffer_data_4[1231:1224];
        layer2[24][47:40] = buffer_data_4[1239:1232];
        layer2[24][55:48] = buffer_data_4[1247:1240];
        layer3[24][7:0] = buffer_data_3[1199:1192];
        layer3[24][15:8] = buffer_data_3[1207:1200];
        layer3[24][23:16] = buffer_data_3[1215:1208];
        layer3[24][31:24] = buffer_data_3[1223:1216];
        layer3[24][39:32] = buffer_data_3[1231:1224];
        layer3[24][47:40] = buffer_data_3[1239:1232];
        layer3[24][55:48] = buffer_data_3[1247:1240];
        layer4[24][7:0] = buffer_data_2[1199:1192];
        layer4[24][15:8] = buffer_data_2[1207:1200];
        layer4[24][23:16] = buffer_data_2[1215:1208];
        layer4[24][31:24] = buffer_data_2[1223:1216];
        layer4[24][39:32] = buffer_data_2[1231:1224];
        layer4[24][47:40] = buffer_data_2[1239:1232];
        layer4[24][55:48] = buffer_data_2[1247:1240];
        layer5[24][7:0] = buffer_data_1[1199:1192];
        layer5[24][15:8] = buffer_data_1[1207:1200];
        layer5[24][23:16] = buffer_data_1[1215:1208];
        layer5[24][31:24] = buffer_data_1[1223:1216];
        layer5[24][39:32] = buffer_data_1[1231:1224];
        layer5[24][47:40] = buffer_data_1[1239:1232];
        layer5[24][55:48] = buffer_data_1[1247:1240];
        layer6[24][7:0] = buffer_data_0[1199:1192];
        layer6[24][15:8] = buffer_data_0[1207:1200];
        layer6[24][23:16] = buffer_data_0[1215:1208];
        layer6[24][31:24] = buffer_data_0[1223:1216];
        layer6[24][39:32] = buffer_data_0[1231:1224];
        layer6[24][47:40] = buffer_data_0[1239:1232];
        layer6[24][55:48] = buffer_data_0[1247:1240];
        layer0[25][7:0] = buffer_data_6[1207:1200];
        layer0[25][15:8] = buffer_data_6[1215:1208];
        layer0[25][23:16] = buffer_data_6[1223:1216];
        layer0[25][31:24] = buffer_data_6[1231:1224];
        layer0[25][39:32] = buffer_data_6[1239:1232];
        layer0[25][47:40] = buffer_data_6[1247:1240];
        layer0[25][55:48] = buffer_data_6[1255:1248];
        layer1[25][7:0] = buffer_data_5[1207:1200];
        layer1[25][15:8] = buffer_data_5[1215:1208];
        layer1[25][23:16] = buffer_data_5[1223:1216];
        layer1[25][31:24] = buffer_data_5[1231:1224];
        layer1[25][39:32] = buffer_data_5[1239:1232];
        layer1[25][47:40] = buffer_data_5[1247:1240];
        layer1[25][55:48] = buffer_data_5[1255:1248];
        layer2[25][7:0] = buffer_data_4[1207:1200];
        layer2[25][15:8] = buffer_data_4[1215:1208];
        layer2[25][23:16] = buffer_data_4[1223:1216];
        layer2[25][31:24] = buffer_data_4[1231:1224];
        layer2[25][39:32] = buffer_data_4[1239:1232];
        layer2[25][47:40] = buffer_data_4[1247:1240];
        layer2[25][55:48] = buffer_data_4[1255:1248];
        layer3[25][7:0] = buffer_data_3[1207:1200];
        layer3[25][15:8] = buffer_data_3[1215:1208];
        layer3[25][23:16] = buffer_data_3[1223:1216];
        layer3[25][31:24] = buffer_data_3[1231:1224];
        layer3[25][39:32] = buffer_data_3[1239:1232];
        layer3[25][47:40] = buffer_data_3[1247:1240];
        layer3[25][55:48] = buffer_data_3[1255:1248];
        layer4[25][7:0] = buffer_data_2[1207:1200];
        layer4[25][15:8] = buffer_data_2[1215:1208];
        layer4[25][23:16] = buffer_data_2[1223:1216];
        layer4[25][31:24] = buffer_data_2[1231:1224];
        layer4[25][39:32] = buffer_data_2[1239:1232];
        layer4[25][47:40] = buffer_data_2[1247:1240];
        layer4[25][55:48] = buffer_data_2[1255:1248];
        layer5[25][7:0] = buffer_data_1[1207:1200];
        layer5[25][15:8] = buffer_data_1[1215:1208];
        layer5[25][23:16] = buffer_data_1[1223:1216];
        layer5[25][31:24] = buffer_data_1[1231:1224];
        layer5[25][39:32] = buffer_data_1[1239:1232];
        layer5[25][47:40] = buffer_data_1[1247:1240];
        layer5[25][55:48] = buffer_data_1[1255:1248];
        layer6[25][7:0] = buffer_data_0[1207:1200];
        layer6[25][15:8] = buffer_data_0[1215:1208];
        layer6[25][23:16] = buffer_data_0[1223:1216];
        layer6[25][31:24] = buffer_data_0[1231:1224];
        layer6[25][39:32] = buffer_data_0[1239:1232];
        layer6[25][47:40] = buffer_data_0[1247:1240];
        layer6[25][55:48] = buffer_data_0[1255:1248];
        layer0[26][7:0] = buffer_data_6[1215:1208];
        layer0[26][15:8] = buffer_data_6[1223:1216];
        layer0[26][23:16] = buffer_data_6[1231:1224];
        layer0[26][31:24] = buffer_data_6[1239:1232];
        layer0[26][39:32] = buffer_data_6[1247:1240];
        layer0[26][47:40] = buffer_data_6[1255:1248];
        layer0[26][55:48] = buffer_data_6[1263:1256];
        layer1[26][7:0] = buffer_data_5[1215:1208];
        layer1[26][15:8] = buffer_data_5[1223:1216];
        layer1[26][23:16] = buffer_data_5[1231:1224];
        layer1[26][31:24] = buffer_data_5[1239:1232];
        layer1[26][39:32] = buffer_data_5[1247:1240];
        layer1[26][47:40] = buffer_data_5[1255:1248];
        layer1[26][55:48] = buffer_data_5[1263:1256];
        layer2[26][7:0] = buffer_data_4[1215:1208];
        layer2[26][15:8] = buffer_data_4[1223:1216];
        layer2[26][23:16] = buffer_data_4[1231:1224];
        layer2[26][31:24] = buffer_data_4[1239:1232];
        layer2[26][39:32] = buffer_data_4[1247:1240];
        layer2[26][47:40] = buffer_data_4[1255:1248];
        layer2[26][55:48] = buffer_data_4[1263:1256];
        layer3[26][7:0] = buffer_data_3[1215:1208];
        layer3[26][15:8] = buffer_data_3[1223:1216];
        layer3[26][23:16] = buffer_data_3[1231:1224];
        layer3[26][31:24] = buffer_data_3[1239:1232];
        layer3[26][39:32] = buffer_data_3[1247:1240];
        layer3[26][47:40] = buffer_data_3[1255:1248];
        layer3[26][55:48] = buffer_data_3[1263:1256];
        layer4[26][7:0] = buffer_data_2[1215:1208];
        layer4[26][15:8] = buffer_data_2[1223:1216];
        layer4[26][23:16] = buffer_data_2[1231:1224];
        layer4[26][31:24] = buffer_data_2[1239:1232];
        layer4[26][39:32] = buffer_data_2[1247:1240];
        layer4[26][47:40] = buffer_data_2[1255:1248];
        layer4[26][55:48] = buffer_data_2[1263:1256];
        layer5[26][7:0] = buffer_data_1[1215:1208];
        layer5[26][15:8] = buffer_data_1[1223:1216];
        layer5[26][23:16] = buffer_data_1[1231:1224];
        layer5[26][31:24] = buffer_data_1[1239:1232];
        layer5[26][39:32] = buffer_data_1[1247:1240];
        layer5[26][47:40] = buffer_data_1[1255:1248];
        layer5[26][55:48] = buffer_data_1[1263:1256];
        layer6[26][7:0] = buffer_data_0[1215:1208];
        layer6[26][15:8] = buffer_data_0[1223:1216];
        layer6[26][23:16] = buffer_data_0[1231:1224];
        layer6[26][31:24] = buffer_data_0[1239:1232];
        layer6[26][39:32] = buffer_data_0[1247:1240];
        layer6[26][47:40] = buffer_data_0[1255:1248];
        layer6[26][55:48] = buffer_data_0[1263:1256];
        layer0[27][7:0] = buffer_data_6[1223:1216];
        layer0[27][15:8] = buffer_data_6[1231:1224];
        layer0[27][23:16] = buffer_data_6[1239:1232];
        layer0[27][31:24] = buffer_data_6[1247:1240];
        layer0[27][39:32] = buffer_data_6[1255:1248];
        layer0[27][47:40] = buffer_data_6[1263:1256];
        layer0[27][55:48] = buffer_data_6[1271:1264];
        layer1[27][7:0] = buffer_data_5[1223:1216];
        layer1[27][15:8] = buffer_data_5[1231:1224];
        layer1[27][23:16] = buffer_data_5[1239:1232];
        layer1[27][31:24] = buffer_data_5[1247:1240];
        layer1[27][39:32] = buffer_data_5[1255:1248];
        layer1[27][47:40] = buffer_data_5[1263:1256];
        layer1[27][55:48] = buffer_data_5[1271:1264];
        layer2[27][7:0] = buffer_data_4[1223:1216];
        layer2[27][15:8] = buffer_data_4[1231:1224];
        layer2[27][23:16] = buffer_data_4[1239:1232];
        layer2[27][31:24] = buffer_data_4[1247:1240];
        layer2[27][39:32] = buffer_data_4[1255:1248];
        layer2[27][47:40] = buffer_data_4[1263:1256];
        layer2[27][55:48] = buffer_data_4[1271:1264];
        layer3[27][7:0] = buffer_data_3[1223:1216];
        layer3[27][15:8] = buffer_data_3[1231:1224];
        layer3[27][23:16] = buffer_data_3[1239:1232];
        layer3[27][31:24] = buffer_data_3[1247:1240];
        layer3[27][39:32] = buffer_data_3[1255:1248];
        layer3[27][47:40] = buffer_data_3[1263:1256];
        layer3[27][55:48] = buffer_data_3[1271:1264];
        layer4[27][7:0] = buffer_data_2[1223:1216];
        layer4[27][15:8] = buffer_data_2[1231:1224];
        layer4[27][23:16] = buffer_data_2[1239:1232];
        layer4[27][31:24] = buffer_data_2[1247:1240];
        layer4[27][39:32] = buffer_data_2[1255:1248];
        layer4[27][47:40] = buffer_data_2[1263:1256];
        layer4[27][55:48] = buffer_data_2[1271:1264];
        layer5[27][7:0] = buffer_data_1[1223:1216];
        layer5[27][15:8] = buffer_data_1[1231:1224];
        layer5[27][23:16] = buffer_data_1[1239:1232];
        layer5[27][31:24] = buffer_data_1[1247:1240];
        layer5[27][39:32] = buffer_data_1[1255:1248];
        layer5[27][47:40] = buffer_data_1[1263:1256];
        layer5[27][55:48] = buffer_data_1[1271:1264];
        layer6[27][7:0] = buffer_data_0[1223:1216];
        layer6[27][15:8] = buffer_data_0[1231:1224];
        layer6[27][23:16] = buffer_data_0[1239:1232];
        layer6[27][31:24] = buffer_data_0[1247:1240];
        layer6[27][39:32] = buffer_data_0[1255:1248];
        layer6[27][47:40] = buffer_data_0[1263:1256];
        layer6[27][55:48] = buffer_data_0[1271:1264];
        layer0[28][7:0] = buffer_data_6[1231:1224];
        layer0[28][15:8] = buffer_data_6[1239:1232];
        layer0[28][23:16] = buffer_data_6[1247:1240];
        layer0[28][31:24] = buffer_data_6[1255:1248];
        layer0[28][39:32] = buffer_data_6[1263:1256];
        layer0[28][47:40] = buffer_data_6[1271:1264];
        layer0[28][55:48] = buffer_data_6[1279:1272];
        layer1[28][7:0] = buffer_data_5[1231:1224];
        layer1[28][15:8] = buffer_data_5[1239:1232];
        layer1[28][23:16] = buffer_data_5[1247:1240];
        layer1[28][31:24] = buffer_data_5[1255:1248];
        layer1[28][39:32] = buffer_data_5[1263:1256];
        layer1[28][47:40] = buffer_data_5[1271:1264];
        layer1[28][55:48] = buffer_data_5[1279:1272];
        layer2[28][7:0] = buffer_data_4[1231:1224];
        layer2[28][15:8] = buffer_data_4[1239:1232];
        layer2[28][23:16] = buffer_data_4[1247:1240];
        layer2[28][31:24] = buffer_data_4[1255:1248];
        layer2[28][39:32] = buffer_data_4[1263:1256];
        layer2[28][47:40] = buffer_data_4[1271:1264];
        layer2[28][55:48] = buffer_data_4[1279:1272];
        layer3[28][7:0] = buffer_data_3[1231:1224];
        layer3[28][15:8] = buffer_data_3[1239:1232];
        layer3[28][23:16] = buffer_data_3[1247:1240];
        layer3[28][31:24] = buffer_data_3[1255:1248];
        layer3[28][39:32] = buffer_data_3[1263:1256];
        layer3[28][47:40] = buffer_data_3[1271:1264];
        layer3[28][55:48] = buffer_data_3[1279:1272];
        layer4[28][7:0] = buffer_data_2[1231:1224];
        layer4[28][15:8] = buffer_data_2[1239:1232];
        layer4[28][23:16] = buffer_data_2[1247:1240];
        layer4[28][31:24] = buffer_data_2[1255:1248];
        layer4[28][39:32] = buffer_data_2[1263:1256];
        layer4[28][47:40] = buffer_data_2[1271:1264];
        layer4[28][55:48] = buffer_data_2[1279:1272];
        layer5[28][7:0] = buffer_data_1[1231:1224];
        layer5[28][15:8] = buffer_data_1[1239:1232];
        layer5[28][23:16] = buffer_data_1[1247:1240];
        layer5[28][31:24] = buffer_data_1[1255:1248];
        layer5[28][39:32] = buffer_data_1[1263:1256];
        layer5[28][47:40] = buffer_data_1[1271:1264];
        layer5[28][55:48] = buffer_data_1[1279:1272];
        layer6[28][7:0] = buffer_data_0[1231:1224];
        layer6[28][15:8] = buffer_data_0[1239:1232];
        layer6[28][23:16] = buffer_data_0[1247:1240];
        layer6[28][31:24] = buffer_data_0[1255:1248];
        layer6[28][39:32] = buffer_data_0[1263:1256];
        layer6[28][47:40] = buffer_data_0[1271:1264];
        layer6[28][55:48] = buffer_data_0[1279:1272];
        layer0[29][7:0] = buffer_data_6[1239:1232];
        layer0[29][15:8] = buffer_data_6[1247:1240];
        layer0[29][23:16] = buffer_data_6[1255:1248];
        layer0[29][31:24] = buffer_data_6[1263:1256];
        layer0[29][39:32] = buffer_data_6[1271:1264];
        layer0[29][47:40] = buffer_data_6[1279:1272];
        layer0[29][55:48] = buffer_data_6[1287:1280];
        layer1[29][7:0] = buffer_data_5[1239:1232];
        layer1[29][15:8] = buffer_data_5[1247:1240];
        layer1[29][23:16] = buffer_data_5[1255:1248];
        layer1[29][31:24] = buffer_data_5[1263:1256];
        layer1[29][39:32] = buffer_data_5[1271:1264];
        layer1[29][47:40] = buffer_data_5[1279:1272];
        layer1[29][55:48] = buffer_data_5[1287:1280];
        layer2[29][7:0] = buffer_data_4[1239:1232];
        layer2[29][15:8] = buffer_data_4[1247:1240];
        layer2[29][23:16] = buffer_data_4[1255:1248];
        layer2[29][31:24] = buffer_data_4[1263:1256];
        layer2[29][39:32] = buffer_data_4[1271:1264];
        layer2[29][47:40] = buffer_data_4[1279:1272];
        layer2[29][55:48] = buffer_data_4[1287:1280];
        layer3[29][7:0] = buffer_data_3[1239:1232];
        layer3[29][15:8] = buffer_data_3[1247:1240];
        layer3[29][23:16] = buffer_data_3[1255:1248];
        layer3[29][31:24] = buffer_data_3[1263:1256];
        layer3[29][39:32] = buffer_data_3[1271:1264];
        layer3[29][47:40] = buffer_data_3[1279:1272];
        layer3[29][55:48] = buffer_data_3[1287:1280];
        layer4[29][7:0] = buffer_data_2[1239:1232];
        layer4[29][15:8] = buffer_data_2[1247:1240];
        layer4[29][23:16] = buffer_data_2[1255:1248];
        layer4[29][31:24] = buffer_data_2[1263:1256];
        layer4[29][39:32] = buffer_data_2[1271:1264];
        layer4[29][47:40] = buffer_data_2[1279:1272];
        layer4[29][55:48] = buffer_data_2[1287:1280];
        layer5[29][7:0] = buffer_data_1[1239:1232];
        layer5[29][15:8] = buffer_data_1[1247:1240];
        layer5[29][23:16] = buffer_data_1[1255:1248];
        layer5[29][31:24] = buffer_data_1[1263:1256];
        layer5[29][39:32] = buffer_data_1[1271:1264];
        layer5[29][47:40] = buffer_data_1[1279:1272];
        layer5[29][55:48] = buffer_data_1[1287:1280];
        layer6[29][7:0] = buffer_data_0[1239:1232];
        layer6[29][15:8] = buffer_data_0[1247:1240];
        layer6[29][23:16] = buffer_data_0[1255:1248];
        layer6[29][31:24] = buffer_data_0[1263:1256];
        layer6[29][39:32] = buffer_data_0[1271:1264];
        layer6[29][47:40] = buffer_data_0[1279:1272];
        layer6[29][55:48] = buffer_data_0[1287:1280];
        layer0[30][7:0] = buffer_data_6[1247:1240];
        layer0[30][15:8] = buffer_data_6[1255:1248];
        layer0[30][23:16] = buffer_data_6[1263:1256];
        layer0[30][31:24] = buffer_data_6[1271:1264];
        layer0[30][39:32] = buffer_data_6[1279:1272];
        layer0[30][47:40] = buffer_data_6[1287:1280];
        layer0[30][55:48] = buffer_data_6[1295:1288];
        layer1[30][7:0] = buffer_data_5[1247:1240];
        layer1[30][15:8] = buffer_data_5[1255:1248];
        layer1[30][23:16] = buffer_data_5[1263:1256];
        layer1[30][31:24] = buffer_data_5[1271:1264];
        layer1[30][39:32] = buffer_data_5[1279:1272];
        layer1[30][47:40] = buffer_data_5[1287:1280];
        layer1[30][55:48] = buffer_data_5[1295:1288];
        layer2[30][7:0] = buffer_data_4[1247:1240];
        layer2[30][15:8] = buffer_data_4[1255:1248];
        layer2[30][23:16] = buffer_data_4[1263:1256];
        layer2[30][31:24] = buffer_data_4[1271:1264];
        layer2[30][39:32] = buffer_data_4[1279:1272];
        layer2[30][47:40] = buffer_data_4[1287:1280];
        layer2[30][55:48] = buffer_data_4[1295:1288];
        layer3[30][7:0] = buffer_data_3[1247:1240];
        layer3[30][15:8] = buffer_data_3[1255:1248];
        layer3[30][23:16] = buffer_data_3[1263:1256];
        layer3[30][31:24] = buffer_data_3[1271:1264];
        layer3[30][39:32] = buffer_data_3[1279:1272];
        layer3[30][47:40] = buffer_data_3[1287:1280];
        layer3[30][55:48] = buffer_data_3[1295:1288];
        layer4[30][7:0] = buffer_data_2[1247:1240];
        layer4[30][15:8] = buffer_data_2[1255:1248];
        layer4[30][23:16] = buffer_data_2[1263:1256];
        layer4[30][31:24] = buffer_data_2[1271:1264];
        layer4[30][39:32] = buffer_data_2[1279:1272];
        layer4[30][47:40] = buffer_data_2[1287:1280];
        layer4[30][55:48] = buffer_data_2[1295:1288];
        layer5[30][7:0] = buffer_data_1[1247:1240];
        layer5[30][15:8] = buffer_data_1[1255:1248];
        layer5[30][23:16] = buffer_data_1[1263:1256];
        layer5[30][31:24] = buffer_data_1[1271:1264];
        layer5[30][39:32] = buffer_data_1[1279:1272];
        layer5[30][47:40] = buffer_data_1[1287:1280];
        layer5[30][55:48] = buffer_data_1[1295:1288];
        layer6[30][7:0] = buffer_data_0[1247:1240];
        layer6[30][15:8] = buffer_data_0[1255:1248];
        layer6[30][23:16] = buffer_data_0[1263:1256];
        layer6[30][31:24] = buffer_data_0[1271:1264];
        layer6[30][39:32] = buffer_data_0[1279:1272];
        layer6[30][47:40] = buffer_data_0[1287:1280];
        layer6[30][55:48] = buffer_data_0[1295:1288];
        layer0[31][7:0] = buffer_data_6[1255:1248];
        layer0[31][15:8] = buffer_data_6[1263:1256];
        layer0[31][23:16] = buffer_data_6[1271:1264];
        layer0[31][31:24] = buffer_data_6[1279:1272];
        layer0[31][39:32] = buffer_data_6[1287:1280];
        layer0[31][47:40] = buffer_data_6[1295:1288];
        layer0[31][55:48] = buffer_data_6[1303:1296];
        layer1[31][7:0] = buffer_data_5[1255:1248];
        layer1[31][15:8] = buffer_data_5[1263:1256];
        layer1[31][23:16] = buffer_data_5[1271:1264];
        layer1[31][31:24] = buffer_data_5[1279:1272];
        layer1[31][39:32] = buffer_data_5[1287:1280];
        layer1[31][47:40] = buffer_data_5[1295:1288];
        layer1[31][55:48] = buffer_data_5[1303:1296];
        layer2[31][7:0] = buffer_data_4[1255:1248];
        layer2[31][15:8] = buffer_data_4[1263:1256];
        layer2[31][23:16] = buffer_data_4[1271:1264];
        layer2[31][31:24] = buffer_data_4[1279:1272];
        layer2[31][39:32] = buffer_data_4[1287:1280];
        layer2[31][47:40] = buffer_data_4[1295:1288];
        layer2[31][55:48] = buffer_data_4[1303:1296];
        layer3[31][7:0] = buffer_data_3[1255:1248];
        layer3[31][15:8] = buffer_data_3[1263:1256];
        layer3[31][23:16] = buffer_data_3[1271:1264];
        layer3[31][31:24] = buffer_data_3[1279:1272];
        layer3[31][39:32] = buffer_data_3[1287:1280];
        layer3[31][47:40] = buffer_data_3[1295:1288];
        layer3[31][55:48] = buffer_data_3[1303:1296];
        layer4[31][7:0] = buffer_data_2[1255:1248];
        layer4[31][15:8] = buffer_data_2[1263:1256];
        layer4[31][23:16] = buffer_data_2[1271:1264];
        layer4[31][31:24] = buffer_data_2[1279:1272];
        layer4[31][39:32] = buffer_data_2[1287:1280];
        layer4[31][47:40] = buffer_data_2[1295:1288];
        layer4[31][55:48] = buffer_data_2[1303:1296];
        layer5[31][7:0] = buffer_data_1[1255:1248];
        layer5[31][15:8] = buffer_data_1[1263:1256];
        layer5[31][23:16] = buffer_data_1[1271:1264];
        layer5[31][31:24] = buffer_data_1[1279:1272];
        layer5[31][39:32] = buffer_data_1[1287:1280];
        layer5[31][47:40] = buffer_data_1[1295:1288];
        layer5[31][55:48] = buffer_data_1[1303:1296];
        layer6[31][7:0] = buffer_data_0[1255:1248];
        layer6[31][15:8] = buffer_data_0[1263:1256];
        layer6[31][23:16] = buffer_data_0[1271:1264];
        layer6[31][31:24] = buffer_data_0[1279:1272];
        layer6[31][39:32] = buffer_data_0[1287:1280];
        layer6[31][47:40] = buffer_data_0[1295:1288];
        layer6[31][55:48] = buffer_data_0[1303:1296];
        layer0[32][7:0] = buffer_data_6[1263:1256];
        layer0[32][15:8] = buffer_data_6[1271:1264];
        layer0[32][23:16] = buffer_data_6[1279:1272];
        layer0[32][31:24] = buffer_data_6[1287:1280];
        layer0[32][39:32] = buffer_data_6[1295:1288];
        layer0[32][47:40] = buffer_data_6[1303:1296];
        layer0[32][55:48] = buffer_data_6[1311:1304];
        layer1[32][7:0] = buffer_data_5[1263:1256];
        layer1[32][15:8] = buffer_data_5[1271:1264];
        layer1[32][23:16] = buffer_data_5[1279:1272];
        layer1[32][31:24] = buffer_data_5[1287:1280];
        layer1[32][39:32] = buffer_data_5[1295:1288];
        layer1[32][47:40] = buffer_data_5[1303:1296];
        layer1[32][55:48] = buffer_data_5[1311:1304];
        layer2[32][7:0] = buffer_data_4[1263:1256];
        layer2[32][15:8] = buffer_data_4[1271:1264];
        layer2[32][23:16] = buffer_data_4[1279:1272];
        layer2[32][31:24] = buffer_data_4[1287:1280];
        layer2[32][39:32] = buffer_data_4[1295:1288];
        layer2[32][47:40] = buffer_data_4[1303:1296];
        layer2[32][55:48] = buffer_data_4[1311:1304];
        layer3[32][7:0] = buffer_data_3[1263:1256];
        layer3[32][15:8] = buffer_data_3[1271:1264];
        layer3[32][23:16] = buffer_data_3[1279:1272];
        layer3[32][31:24] = buffer_data_3[1287:1280];
        layer3[32][39:32] = buffer_data_3[1295:1288];
        layer3[32][47:40] = buffer_data_3[1303:1296];
        layer3[32][55:48] = buffer_data_3[1311:1304];
        layer4[32][7:0] = buffer_data_2[1263:1256];
        layer4[32][15:8] = buffer_data_2[1271:1264];
        layer4[32][23:16] = buffer_data_2[1279:1272];
        layer4[32][31:24] = buffer_data_2[1287:1280];
        layer4[32][39:32] = buffer_data_2[1295:1288];
        layer4[32][47:40] = buffer_data_2[1303:1296];
        layer4[32][55:48] = buffer_data_2[1311:1304];
        layer5[32][7:0] = buffer_data_1[1263:1256];
        layer5[32][15:8] = buffer_data_1[1271:1264];
        layer5[32][23:16] = buffer_data_1[1279:1272];
        layer5[32][31:24] = buffer_data_1[1287:1280];
        layer5[32][39:32] = buffer_data_1[1295:1288];
        layer5[32][47:40] = buffer_data_1[1303:1296];
        layer5[32][55:48] = buffer_data_1[1311:1304];
        layer6[32][7:0] = buffer_data_0[1263:1256];
        layer6[32][15:8] = buffer_data_0[1271:1264];
        layer6[32][23:16] = buffer_data_0[1279:1272];
        layer6[32][31:24] = buffer_data_0[1287:1280];
        layer6[32][39:32] = buffer_data_0[1295:1288];
        layer6[32][47:40] = buffer_data_0[1303:1296];
        layer6[32][55:48] = buffer_data_0[1311:1304];
        layer0[33][7:0] = buffer_data_6[1271:1264];
        layer0[33][15:8] = buffer_data_6[1279:1272];
        layer0[33][23:16] = buffer_data_6[1287:1280];
        layer0[33][31:24] = buffer_data_6[1295:1288];
        layer0[33][39:32] = buffer_data_6[1303:1296];
        layer0[33][47:40] = buffer_data_6[1311:1304];
        layer0[33][55:48] = buffer_data_6[1319:1312];
        layer1[33][7:0] = buffer_data_5[1271:1264];
        layer1[33][15:8] = buffer_data_5[1279:1272];
        layer1[33][23:16] = buffer_data_5[1287:1280];
        layer1[33][31:24] = buffer_data_5[1295:1288];
        layer1[33][39:32] = buffer_data_5[1303:1296];
        layer1[33][47:40] = buffer_data_5[1311:1304];
        layer1[33][55:48] = buffer_data_5[1319:1312];
        layer2[33][7:0] = buffer_data_4[1271:1264];
        layer2[33][15:8] = buffer_data_4[1279:1272];
        layer2[33][23:16] = buffer_data_4[1287:1280];
        layer2[33][31:24] = buffer_data_4[1295:1288];
        layer2[33][39:32] = buffer_data_4[1303:1296];
        layer2[33][47:40] = buffer_data_4[1311:1304];
        layer2[33][55:48] = buffer_data_4[1319:1312];
        layer3[33][7:0] = buffer_data_3[1271:1264];
        layer3[33][15:8] = buffer_data_3[1279:1272];
        layer3[33][23:16] = buffer_data_3[1287:1280];
        layer3[33][31:24] = buffer_data_3[1295:1288];
        layer3[33][39:32] = buffer_data_3[1303:1296];
        layer3[33][47:40] = buffer_data_3[1311:1304];
        layer3[33][55:48] = buffer_data_3[1319:1312];
        layer4[33][7:0] = buffer_data_2[1271:1264];
        layer4[33][15:8] = buffer_data_2[1279:1272];
        layer4[33][23:16] = buffer_data_2[1287:1280];
        layer4[33][31:24] = buffer_data_2[1295:1288];
        layer4[33][39:32] = buffer_data_2[1303:1296];
        layer4[33][47:40] = buffer_data_2[1311:1304];
        layer4[33][55:48] = buffer_data_2[1319:1312];
        layer5[33][7:0] = buffer_data_1[1271:1264];
        layer5[33][15:8] = buffer_data_1[1279:1272];
        layer5[33][23:16] = buffer_data_1[1287:1280];
        layer5[33][31:24] = buffer_data_1[1295:1288];
        layer5[33][39:32] = buffer_data_1[1303:1296];
        layer5[33][47:40] = buffer_data_1[1311:1304];
        layer5[33][55:48] = buffer_data_1[1319:1312];
        layer6[33][7:0] = buffer_data_0[1271:1264];
        layer6[33][15:8] = buffer_data_0[1279:1272];
        layer6[33][23:16] = buffer_data_0[1287:1280];
        layer6[33][31:24] = buffer_data_0[1295:1288];
        layer6[33][39:32] = buffer_data_0[1303:1296];
        layer6[33][47:40] = buffer_data_0[1311:1304];
        layer6[33][55:48] = buffer_data_0[1319:1312];
        layer0[34][7:0] = buffer_data_6[1279:1272];
        layer0[34][15:8] = buffer_data_6[1287:1280];
        layer0[34][23:16] = buffer_data_6[1295:1288];
        layer0[34][31:24] = buffer_data_6[1303:1296];
        layer0[34][39:32] = buffer_data_6[1311:1304];
        layer0[34][47:40] = buffer_data_6[1319:1312];
        layer0[34][55:48] = buffer_data_6[1327:1320];
        layer1[34][7:0] = buffer_data_5[1279:1272];
        layer1[34][15:8] = buffer_data_5[1287:1280];
        layer1[34][23:16] = buffer_data_5[1295:1288];
        layer1[34][31:24] = buffer_data_5[1303:1296];
        layer1[34][39:32] = buffer_data_5[1311:1304];
        layer1[34][47:40] = buffer_data_5[1319:1312];
        layer1[34][55:48] = buffer_data_5[1327:1320];
        layer2[34][7:0] = buffer_data_4[1279:1272];
        layer2[34][15:8] = buffer_data_4[1287:1280];
        layer2[34][23:16] = buffer_data_4[1295:1288];
        layer2[34][31:24] = buffer_data_4[1303:1296];
        layer2[34][39:32] = buffer_data_4[1311:1304];
        layer2[34][47:40] = buffer_data_4[1319:1312];
        layer2[34][55:48] = buffer_data_4[1327:1320];
        layer3[34][7:0] = buffer_data_3[1279:1272];
        layer3[34][15:8] = buffer_data_3[1287:1280];
        layer3[34][23:16] = buffer_data_3[1295:1288];
        layer3[34][31:24] = buffer_data_3[1303:1296];
        layer3[34][39:32] = buffer_data_3[1311:1304];
        layer3[34][47:40] = buffer_data_3[1319:1312];
        layer3[34][55:48] = buffer_data_3[1327:1320];
        layer4[34][7:0] = buffer_data_2[1279:1272];
        layer4[34][15:8] = buffer_data_2[1287:1280];
        layer4[34][23:16] = buffer_data_2[1295:1288];
        layer4[34][31:24] = buffer_data_2[1303:1296];
        layer4[34][39:32] = buffer_data_2[1311:1304];
        layer4[34][47:40] = buffer_data_2[1319:1312];
        layer4[34][55:48] = buffer_data_2[1327:1320];
        layer5[34][7:0] = buffer_data_1[1279:1272];
        layer5[34][15:8] = buffer_data_1[1287:1280];
        layer5[34][23:16] = buffer_data_1[1295:1288];
        layer5[34][31:24] = buffer_data_1[1303:1296];
        layer5[34][39:32] = buffer_data_1[1311:1304];
        layer5[34][47:40] = buffer_data_1[1319:1312];
        layer5[34][55:48] = buffer_data_1[1327:1320];
        layer6[34][7:0] = buffer_data_0[1279:1272];
        layer6[34][15:8] = buffer_data_0[1287:1280];
        layer6[34][23:16] = buffer_data_0[1295:1288];
        layer6[34][31:24] = buffer_data_0[1303:1296];
        layer6[34][39:32] = buffer_data_0[1311:1304];
        layer6[34][47:40] = buffer_data_0[1319:1312];
        layer6[34][55:48] = buffer_data_0[1327:1320];
        layer0[35][7:0] = buffer_data_6[1287:1280];
        layer0[35][15:8] = buffer_data_6[1295:1288];
        layer0[35][23:16] = buffer_data_6[1303:1296];
        layer0[35][31:24] = buffer_data_6[1311:1304];
        layer0[35][39:32] = buffer_data_6[1319:1312];
        layer0[35][47:40] = buffer_data_6[1327:1320];
        layer0[35][55:48] = buffer_data_6[1335:1328];
        layer1[35][7:0] = buffer_data_5[1287:1280];
        layer1[35][15:8] = buffer_data_5[1295:1288];
        layer1[35][23:16] = buffer_data_5[1303:1296];
        layer1[35][31:24] = buffer_data_5[1311:1304];
        layer1[35][39:32] = buffer_data_5[1319:1312];
        layer1[35][47:40] = buffer_data_5[1327:1320];
        layer1[35][55:48] = buffer_data_5[1335:1328];
        layer2[35][7:0] = buffer_data_4[1287:1280];
        layer2[35][15:8] = buffer_data_4[1295:1288];
        layer2[35][23:16] = buffer_data_4[1303:1296];
        layer2[35][31:24] = buffer_data_4[1311:1304];
        layer2[35][39:32] = buffer_data_4[1319:1312];
        layer2[35][47:40] = buffer_data_4[1327:1320];
        layer2[35][55:48] = buffer_data_4[1335:1328];
        layer3[35][7:0] = buffer_data_3[1287:1280];
        layer3[35][15:8] = buffer_data_3[1295:1288];
        layer3[35][23:16] = buffer_data_3[1303:1296];
        layer3[35][31:24] = buffer_data_3[1311:1304];
        layer3[35][39:32] = buffer_data_3[1319:1312];
        layer3[35][47:40] = buffer_data_3[1327:1320];
        layer3[35][55:48] = buffer_data_3[1335:1328];
        layer4[35][7:0] = buffer_data_2[1287:1280];
        layer4[35][15:8] = buffer_data_2[1295:1288];
        layer4[35][23:16] = buffer_data_2[1303:1296];
        layer4[35][31:24] = buffer_data_2[1311:1304];
        layer4[35][39:32] = buffer_data_2[1319:1312];
        layer4[35][47:40] = buffer_data_2[1327:1320];
        layer4[35][55:48] = buffer_data_2[1335:1328];
        layer5[35][7:0] = buffer_data_1[1287:1280];
        layer5[35][15:8] = buffer_data_1[1295:1288];
        layer5[35][23:16] = buffer_data_1[1303:1296];
        layer5[35][31:24] = buffer_data_1[1311:1304];
        layer5[35][39:32] = buffer_data_1[1319:1312];
        layer5[35][47:40] = buffer_data_1[1327:1320];
        layer5[35][55:48] = buffer_data_1[1335:1328];
        layer6[35][7:0] = buffer_data_0[1287:1280];
        layer6[35][15:8] = buffer_data_0[1295:1288];
        layer6[35][23:16] = buffer_data_0[1303:1296];
        layer6[35][31:24] = buffer_data_0[1311:1304];
        layer6[35][39:32] = buffer_data_0[1319:1312];
        layer6[35][47:40] = buffer_data_0[1327:1320];
        layer6[35][55:48] = buffer_data_0[1335:1328];
        layer0[36][7:0] = buffer_data_6[1295:1288];
        layer0[36][15:8] = buffer_data_6[1303:1296];
        layer0[36][23:16] = buffer_data_6[1311:1304];
        layer0[36][31:24] = buffer_data_6[1319:1312];
        layer0[36][39:32] = buffer_data_6[1327:1320];
        layer0[36][47:40] = buffer_data_6[1335:1328];
        layer0[36][55:48] = buffer_data_6[1343:1336];
        layer1[36][7:0] = buffer_data_5[1295:1288];
        layer1[36][15:8] = buffer_data_5[1303:1296];
        layer1[36][23:16] = buffer_data_5[1311:1304];
        layer1[36][31:24] = buffer_data_5[1319:1312];
        layer1[36][39:32] = buffer_data_5[1327:1320];
        layer1[36][47:40] = buffer_data_5[1335:1328];
        layer1[36][55:48] = buffer_data_5[1343:1336];
        layer2[36][7:0] = buffer_data_4[1295:1288];
        layer2[36][15:8] = buffer_data_4[1303:1296];
        layer2[36][23:16] = buffer_data_4[1311:1304];
        layer2[36][31:24] = buffer_data_4[1319:1312];
        layer2[36][39:32] = buffer_data_4[1327:1320];
        layer2[36][47:40] = buffer_data_4[1335:1328];
        layer2[36][55:48] = buffer_data_4[1343:1336];
        layer3[36][7:0] = buffer_data_3[1295:1288];
        layer3[36][15:8] = buffer_data_3[1303:1296];
        layer3[36][23:16] = buffer_data_3[1311:1304];
        layer3[36][31:24] = buffer_data_3[1319:1312];
        layer3[36][39:32] = buffer_data_3[1327:1320];
        layer3[36][47:40] = buffer_data_3[1335:1328];
        layer3[36][55:48] = buffer_data_3[1343:1336];
        layer4[36][7:0] = buffer_data_2[1295:1288];
        layer4[36][15:8] = buffer_data_2[1303:1296];
        layer4[36][23:16] = buffer_data_2[1311:1304];
        layer4[36][31:24] = buffer_data_2[1319:1312];
        layer4[36][39:32] = buffer_data_2[1327:1320];
        layer4[36][47:40] = buffer_data_2[1335:1328];
        layer4[36][55:48] = buffer_data_2[1343:1336];
        layer5[36][7:0] = buffer_data_1[1295:1288];
        layer5[36][15:8] = buffer_data_1[1303:1296];
        layer5[36][23:16] = buffer_data_1[1311:1304];
        layer5[36][31:24] = buffer_data_1[1319:1312];
        layer5[36][39:32] = buffer_data_1[1327:1320];
        layer5[36][47:40] = buffer_data_1[1335:1328];
        layer5[36][55:48] = buffer_data_1[1343:1336];
        layer6[36][7:0] = buffer_data_0[1295:1288];
        layer6[36][15:8] = buffer_data_0[1303:1296];
        layer6[36][23:16] = buffer_data_0[1311:1304];
        layer6[36][31:24] = buffer_data_0[1319:1312];
        layer6[36][39:32] = buffer_data_0[1327:1320];
        layer6[36][47:40] = buffer_data_0[1335:1328];
        layer6[36][55:48] = buffer_data_0[1343:1336];
        layer0[37][7:0] = buffer_data_6[1303:1296];
        layer0[37][15:8] = buffer_data_6[1311:1304];
        layer0[37][23:16] = buffer_data_6[1319:1312];
        layer0[37][31:24] = buffer_data_6[1327:1320];
        layer0[37][39:32] = buffer_data_6[1335:1328];
        layer0[37][47:40] = buffer_data_6[1343:1336];
        layer0[37][55:48] = buffer_data_6[1351:1344];
        layer1[37][7:0] = buffer_data_5[1303:1296];
        layer1[37][15:8] = buffer_data_5[1311:1304];
        layer1[37][23:16] = buffer_data_5[1319:1312];
        layer1[37][31:24] = buffer_data_5[1327:1320];
        layer1[37][39:32] = buffer_data_5[1335:1328];
        layer1[37][47:40] = buffer_data_5[1343:1336];
        layer1[37][55:48] = buffer_data_5[1351:1344];
        layer2[37][7:0] = buffer_data_4[1303:1296];
        layer2[37][15:8] = buffer_data_4[1311:1304];
        layer2[37][23:16] = buffer_data_4[1319:1312];
        layer2[37][31:24] = buffer_data_4[1327:1320];
        layer2[37][39:32] = buffer_data_4[1335:1328];
        layer2[37][47:40] = buffer_data_4[1343:1336];
        layer2[37][55:48] = buffer_data_4[1351:1344];
        layer3[37][7:0] = buffer_data_3[1303:1296];
        layer3[37][15:8] = buffer_data_3[1311:1304];
        layer3[37][23:16] = buffer_data_3[1319:1312];
        layer3[37][31:24] = buffer_data_3[1327:1320];
        layer3[37][39:32] = buffer_data_3[1335:1328];
        layer3[37][47:40] = buffer_data_3[1343:1336];
        layer3[37][55:48] = buffer_data_3[1351:1344];
        layer4[37][7:0] = buffer_data_2[1303:1296];
        layer4[37][15:8] = buffer_data_2[1311:1304];
        layer4[37][23:16] = buffer_data_2[1319:1312];
        layer4[37][31:24] = buffer_data_2[1327:1320];
        layer4[37][39:32] = buffer_data_2[1335:1328];
        layer4[37][47:40] = buffer_data_2[1343:1336];
        layer4[37][55:48] = buffer_data_2[1351:1344];
        layer5[37][7:0] = buffer_data_1[1303:1296];
        layer5[37][15:8] = buffer_data_1[1311:1304];
        layer5[37][23:16] = buffer_data_1[1319:1312];
        layer5[37][31:24] = buffer_data_1[1327:1320];
        layer5[37][39:32] = buffer_data_1[1335:1328];
        layer5[37][47:40] = buffer_data_1[1343:1336];
        layer5[37][55:48] = buffer_data_1[1351:1344];
        layer6[37][7:0] = buffer_data_0[1303:1296];
        layer6[37][15:8] = buffer_data_0[1311:1304];
        layer6[37][23:16] = buffer_data_0[1319:1312];
        layer6[37][31:24] = buffer_data_0[1327:1320];
        layer6[37][39:32] = buffer_data_0[1335:1328];
        layer6[37][47:40] = buffer_data_0[1343:1336];
        layer6[37][55:48] = buffer_data_0[1351:1344];
        layer0[38][7:0] = buffer_data_6[1311:1304];
        layer0[38][15:8] = buffer_data_6[1319:1312];
        layer0[38][23:16] = buffer_data_6[1327:1320];
        layer0[38][31:24] = buffer_data_6[1335:1328];
        layer0[38][39:32] = buffer_data_6[1343:1336];
        layer0[38][47:40] = buffer_data_6[1351:1344];
        layer0[38][55:48] = buffer_data_6[1359:1352];
        layer1[38][7:0] = buffer_data_5[1311:1304];
        layer1[38][15:8] = buffer_data_5[1319:1312];
        layer1[38][23:16] = buffer_data_5[1327:1320];
        layer1[38][31:24] = buffer_data_5[1335:1328];
        layer1[38][39:32] = buffer_data_5[1343:1336];
        layer1[38][47:40] = buffer_data_5[1351:1344];
        layer1[38][55:48] = buffer_data_5[1359:1352];
        layer2[38][7:0] = buffer_data_4[1311:1304];
        layer2[38][15:8] = buffer_data_4[1319:1312];
        layer2[38][23:16] = buffer_data_4[1327:1320];
        layer2[38][31:24] = buffer_data_4[1335:1328];
        layer2[38][39:32] = buffer_data_4[1343:1336];
        layer2[38][47:40] = buffer_data_4[1351:1344];
        layer2[38][55:48] = buffer_data_4[1359:1352];
        layer3[38][7:0] = buffer_data_3[1311:1304];
        layer3[38][15:8] = buffer_data_3[1319:1312];
        layer3[38][23:16] = buffer_data_3[1327:1320];
        layer3[38][31:24] = buffer_data_3[1335:1328];
        layer3[38][39:32] = buffer_data_3[1343:1336];
        layer3[38][47:40] = buffer_data_3[1351:1344];
        layer3[38][55:48] = buffer_data_3[1359:1352];
        layer4[38][7:0] = buffer_data_2[1311:1304];
        layer4[38][15:8] = buffer_data_2[1319:1312];
        layer4[38][23:16] = buffer_data_2[1327:1320];
        layer4[38][31:24] = buffer_data_2[1335:1328];
        layer4[38][39:32] = buffer_data_2[1343:1336];
        layer4[38][47:40] = buffer_data_2[1351:1344];
        layer4[38][55:48] = buffer_data_2[1359:1352];
        layer5[38][7:0] = buffer_data_1[1311:1304];
        layer5[38][15:8] = buffer_data_1[1319:1312];
        layer5[38][23:16] = buffer_data_1[1327:1320];
        layer5[38][31:24] = buffer_data_1[1335:1328];
        layer5[38][39:32] = buffer_data_1[1343:1336];
        layer5[38][47:40] = buffer_data_1[1351:1344];
        layer5[38][55:48] = buffer_data_1[1359:1352];
        layer6[38][7:0] = buffer_data_0[1311:1304];
        layer6[38][15:8] = buffer_data_0[1319:1312];
        layer6[38][23:16] = buffer_data_0[1327:1320];
        layer6[38][31:24] = buffer_data_0[1335:1328];
        layer6[38][39:32] = buffer_data_0[1343:1336];
        layer6[38][47:40] = buffer_data_0[1351:1344];
        layer6[38][55:48] = buffer_data_0[1359:1352];
        layer0[39][7:0] = buffer_data_6[1319:1312];
        layer0[39][15:8] = buffer_data_6[1327:1320];
        layer0[39][23:16] = buffer_data_6[1335:1328];
        layer0[39][31:24] = buffer_data_6[1343:1336];
        layer0[39][39:32] = buffer_data_6[1351:1344];
        layer0[39][47:40] = buffer_data_6[1359:1352];
        layer0[39][55:48] = buffer_data_6[1367:1360];
        layer1[39][7:0] = buffer_data_5[1319:1312];
        layer1[39][15:8] = buffer_data_5[1327:1320];
        layer1[39][23:16] = buffer_data_5[1335:1328];
        layer1[39][31:24] = buffer_data_5[1343:1336];
        layer1[39][39:32] = buffer_data_5[1351:1344];
        layer1[39][47:40] = buffer_data_5[1359:1352];
        layer1[39][55:48] = buffer_data_5[1367:1360];
        layer2[39][7:0] = buffer_data_4[1319:1312];
        layer2[39][15:8] = buffer_data_4[1327:1320];
        layer2[39][23:16] = buffer_data_4[1335:1328];
        layer2[39][31:24] = buffer_data_4[1343:1336];
        layer2[39][39:32] = buffer_data_4[1351:1344];
        layer2[39][47:40] = buffer_data_4[1359:1352];
        layer2[39][55:48] = buffer_data_4[1367:1360];
        layer3[39][7:0] = buffer_data_3[1319:1312];
        layer3[39][15:8] = buffer_data_3[1327:1320];
        layer3[39][23:16] = buffer_data_3[1335:1328];
        layer3[39][31:24] = buffer_data_3[1343:1336];
        layer3[39][39:32] = buffer_data_3[1351:1344];
        layer3[39][47:40] = buffer_data_3[1359:1352];
        layer3[39][55:48] = buffer_data_3[1367:1360];
        layer4[39][7:0] = buffer_data_2[1319:1312];
        layer4[39][15:8] = buffer_data_2[1327:1320];
        layer4[39][23:16] = buffer_data_2[1335:1328];
        layer4[39][31:24] = buffer_data_2[1343:1336];
        layer4[39][39:32] = buffer_data_2[1351:1344];
        layer4[39][47:40] = buffer_data_2[1359:1352];
        layer4[39][55:48] = buffer_data_2[1367:1360];
        layer5[39][7:0] = buffer_data_1[1319:1312];
        layer5[39][15:8] = buffer_data_1[1327:1320];
        layer5[39][23:16] = buffer_data_1[1335:1328];
        layer5[39][31:24] = buffer_data_1[1343:1336];
        layer5[39][39:32] = buffer_data_1[1351:1344];
        layer5[39][47:40] = buffer_data_1[1359:1352];
        layer5[39][55:48] = buffer_data_1[1367:1360];
        layer6[39][7:0] = buffer_data_0[1319:1312];
        layer6[39][15:8] = buffer_data_0[1327:1320];
        layer6[39][23:16] = buffer_data_0[1335:1328];
        layer6[39][31:24] = buffer_data_0[1343:1336];
        layer6[39][39:32] = buffer_data_0[1351:1344];
        layer6[39][47:40] = buffer_data_0[1359:1352];
        layer6[39][55:48] = buffer_data_0[1367:1360];
        layer0[40][7:0] = buffer_data_6[1327:1320];
        layer0[40][15:8] = buffer_data_6[1335:1328];
        layer0[40][23:16] = buffer_data_6[1343:1336];
        layer0[40][31:24] = buffer_data_6[1351:1344];
        layer0[40][39:32] = buffer_data_6[1359:1352];
        layer0[40][47:40] = buffer_data_6[1367:1360];
        layer0[40][55:48] = buffer_data_6[1375:1368];
        layer1[40][7:0] = buffer_data_5[1327:1320];
        layer1[40][15:8] = buffer_data_5[1335:1328];
        layer1[40][23:16] = buffer_data_5[1343:1336];
        layer1[40][31:24] = buffer_data_5[1351:1344];
        layer1[40][39:32] = buffer_data_5[1359:1352];
        layer1[40][47:40] = buffer_data_5[1367:1360];
        layer1[40][55:48] = buffer_data_5[1375:1368];
        layer2[40][7:0] = buffer_data_4[1327:1320];
        layer2[40][15:8] = buffer_data_4[1335:1328];
        layer2[40][23:16] = buffer_data_4[1343:1336];
        layer2[40][31:24] = buffer_data_4[1351:1344];
        layer2[40][39:32] = buffer_data_4[1359:1352];
        layer2[40][47:40] = buffer_data_4[1367:1360];
        layer2[40][55:48] = buffer_data_4[1375:1368];
        layer3[40][7:0] = buffer_data_3[1327:1320];
        layer3[40][15:8] = buffer_data_3[1335:1328];
        layer3[40][23:16] = buffer_data_3[1343:1336];
        layer3[40][31:24] = buffer_data_3[1351:1344];
        layer3[40][39:32] = buffer_data_3[1359:1352];
        layer3[40][47:40] = buffer_data_3[1367:1360];
        layer3[40][55:48] = buffer_data_3[1375:1368];
        layer4[40][7:0] = buffer_data_2[1327:1320];
        layer4[40][15:8] = buffer_data_2[1335:1328];
        layer4[40][23:16] = buffer_data_2[1343:1336];
        layer4[40][31:24] = buffer_data_2[1351:1344];
        layer4[40][39:32] = buffer_data_2[1359:1352];
        layer4[40][47:40] = buffer_data_2[1367:1360];
        layer4[40][55:48] = buffer_data_2[1375:1368];
        layer5[40][7:0] = buffer_data_1[1327:1320];
        layer5[40][15:8] = buffer_data_1[1335:1328];
        layer5[40][23:16] = buffer_data_1[1343:1336];
        layer5[40][31:24] = buffer_data_1[1351:1344];
        layer5[40][39:32] = buffer_data_1[1359:1352];
        layer5[40][47:40] = buffer_data_1[1367:1360];
        layer5[40][55:48] = buffer_data_1[1375:1368];
        layer6[40][7:0] = buffer_data_0[1327:1320];
        layer6[40][15:8] = buffer_data_0[1335:1328];
        layer6[40][23:16] = buffer_data_0[1343:1336];
        layer6[40][31:24] = buffer_data_0[1351:1344];
        layer6[40][39:32] = buffer_data_0[1359:1352];
        layer6[40][47:40] = buffer_data_0[1367:1360];
        layer6[40][55:48] = buffer_data_0[1375:1368];
        layer0[41][7:0] = buffer_data_6[1335:1328];
        layer0[41][15:8] = buffer_data_6[1343:1336];
        layer0[41][23:16] = buffer_data_6[1351:1344];
        layer0[41][31:24] = buffer_data_6[1359:1352];
        layer0[41][39:32] = buffer_data_6[1367:1360];
        layer0[41][47:40] = buffer_data_6[1375:1368];
        layer0[41][55:48] = buffer_data_6[1383:1376];
        layer1[41][7:0] = buffer_data_5[1335:1328];
        layer1[41][15:8] = buffer_data_5[1343:1336];
        layer1[41][23:16] = buffer_data_5[1351:1344];
        layer1[41][31:24] = buffer_data_5[1359:1352];
        layer1[41][39:32] = buffer_data_5[1367:1360];
        layer1[41][47:40] = buffer_data_5[1375:1368];
        layer1[41][55:48] = buffer_data_5[1383:1376];
        layer2[41][7:0] = buffer_data_4[1335:1328];
        layer2[41][15:8] = buffer_data_4[1343:1336];
        layer2[41][23:16] = buffer_data_4[1351:1344];
        layer2[41][31:24] = buffer_data_4[1359:1352];
        layer2[41][39:32] = buffer_data_4[1367:1360];
        layer2[41][47:40] = buffer_data_4[1375:1368];
        layer2[41][55:48] = buffer_data_4[1383:1376];
        layer3[41][7:0] = buffer_data_3[1335:1328];
        layer3[41][15:8] = buffer_data_3[1343:1336];
        layer3[41][23:16] = buffer_data_3[1351:1344];
        layer3[41][31:24] = buffer_data_3[1359:1352];
        layer3[41][39:32] = buffer_data_3[1367:1360];
        layer3[41][47:40] = buffer_data_3[1375:1368];
        layer3[41][55:48] = buffer_data_3[1383:1376];
        layer4[41][7:0] = buffer_data_2[1335:1328];
        layer4[41][15:8] = buffer_data_2[1343:1336];
        layer4[41][23:16] = buffer_data_2[1351:1344];
        layer4[41][31:24] = buffer_data_2[1359:1352];
        layer4[41][39:32] = buffer_data_2[1367:1360];
        layer4[41][47:40] = buffer_data_2[1375:1368];
        layer4[41][55:48] = buffer_data_2[1383:1376];
        layer5[41][7:0] = buffer_data_1[1335:1328];
        layer5[41][15:8] = buffer_data_1[1343:1336];
        layer5[41][23:16] = buffer_data_1[1351:1344];
        layer5[41][31:24] = buffer_data_1[1359:1352];
        layer5[41][39:32] = buffer_data_1[1367:1360];
        layer5[41][47:40] = buffer_data_1[1375:1368];
        layer5[41][55:48] = buffer_data_1[1383:1376];
        layer6[41][7:0] = buffer_data_0[1335:1328];
        layer6[41][15:8] = buffer_data_0[1343:1336];
        layer6[41][23:16] = buffer_data_0[1351:1344];
        layer6[41][31:24] = buffer_data_0[1359:1352];
        layer6[41][39:32] = buffer_data_0[1367:1360];
        layer6[41][47:40] = buffer_data_0[1375:1368];
        layer6[41][55:48] = buffer_data_0[1383:1376];
        layer0[42][7:0] = buffer_data_6[1343:1336];
        layer0[42][15:8] = buffer_data_6[1351:1344];
        layer0[42][23:16] = buffer_data_6[1359:1352];
        layer0[42][31:24] = buffer_data_6[1367:1360];
        layer0[42][39:32] = buffer_data_6[1375:1368];
        layer0[42][47:40] = buffer_data_6[1383:1376];
        layer0[42][55:48] = buffer_data_6[1391:1384];
        layer1[42][7:0] = buffer_data_5[1343:1336];
        layer1[42][15:8] = buffer_data_5[1351:1344];
        layer1[42][23:16] = buffer_data_5[1359:1352];
        layer1[42][31:24] = buffer_data_5[1367:1360];
        layer1[42][39:32] = buffer_data_5[1375:1368];
        layer1[42][47:40] = buffer_data_5[1383:1376];
        layer1[42][55:48] = buffer_data_5[1391:1384];
        layer2[42][7:0] = buffer_data_4[1343:1336];
        layer2[42][15:8] = buffer_data_4[1351:1344];
        layer2[42][23:16] = buffer_data_4[1359:1352];
        layer2[42][31:24] = buffer_data_4[1367:1360];
        layer2[42][39:32] = buffer_data_4[1375:1368];
        layer2[42][47:40] = buffer_data_4[1383:1376];
        layer2[42][55:48] = buffer_data_4[1391:1384];
        layer3[42][7:0] = buffer_data_3[1343:1336];
        layer3[42][15:8] = buffer_data_3[1351:1344];
        layer3[42][23:16] = buffer_data_3[1359:1352];
        layer3[42][31:24] = buffer_data_3[1367:1360];
        layer3[42][39:32] = buffer_data_3[1375:1368];
        layer3[42][47:40] = buffer_data_3[1383:1376];
        layer3[42][55:48] = buffer_data_3[1391:1384];
        layer4[42][7:0] = buffer_data_2[1343:1336];
        layer4[42][15:8] = buffer_data_2[1351:1344];
        layer4[42][23:16] = buffer_data_2[1359:1352];
        layer4[42][31:24] = buffer_data_2[1367:1360];
        layer4[42][39:32] = buffer_data_2[1375:1368];
        layer4[42][47:40] = buffer_data_2[1383:1376];
        layer4[42][55:48] = buffer_data_2[1391:1384];
        layer5[42][7:0] = buffer_data_1[1343:1336];
        layer5[42][15:8] = buffer_data_1[1351:1344];
        layer5[42][23:16] = buffer_data_1[1359:1352];
        layer5[42][31:24] = buffer_data_1[1367:1360];
        layer5[42][39:32] = buffer_data_1[1375:1368];
        layer5[42][47:40] = buffer_data_1[1383:1376];
        layer5[42][55:48] = buffer_data_1[1391:1384];
        layer6[42][7:0] = buffer_data_0[1343:1336];
        layer6[42][15:8] = buffer_data_0[1351:1344];
        layer6[42][23:16] = buffer_data_0[1359:1352];
        layer6[42][31:24] = buffer_data_0[1367:1360];
        layer6[42][39:32] = buffer_data_0[1375:1368];
        layer6[42][47:40] = buffer_data_0[1383:1376];
        layer6[42][55:48] = buffer_data_0[1391:1384];
        layer0[43][7:0] = buffer_data_6[1351:1344];
        layer0[43][15:8] = buffer_data_6[1359:1352];
        layer0[43][23:16] = buffer_data_6[1367:1360];
        layer0[43][31:24] = buffer_data_6[1375:1368];
        layer0[43][39:32] = buffer_data_6[1383:1376];
        layer0[43][47:40] = buffer_data_6[1391:1384];
        layer0[43][55:48] = buffer_data_6[1399:1392];
        layer1[43][7:0] = buffer_data_5[1351:1344];
        layer1[43][15:8] = buffer_data_5[1359:1352];
        layer1[43][23:16] = buffer_data_5[1367:1360];
        layer1[43][31:24] = buffer_data_5[1375:1368];
        layer1[43][39:32] = buffer_data_5[1383:1376];
        layer1[43][47:40] = buffer_data_5[1391:1384];
        layer1[43][55:48] = buffer_data_5[1399:1392];
        layer2[43][7:0] = buffer_data_4[1351:1344];
        layer2[43][15:8] = buffer_data_4[1359:1352];
        layer2[43][23:16] = buffer_data_4[1367:1360];
        layer2[43][31:24] = buffer_data_4[1375:1368];
        layer2[43][39:32] = buffer_data_4[1383:1376];
        layer2[43][47:40] = buffer_data_4[1391:1384];
        layer2[43][55:48] = buffer_data_4[1399:1392];
        layer3[43][7:0] = buffer_data_3[1351:1344];
        layer3[43][15:8] = buffer_data_3[1359:1352];
        layer3[43][23:16] = buffer_data_3[1367:1360];
        layer3[43][31:24] = buffer_data_3[1375:1368];
        layer3[43][39:32] = buffer_data_3[1383:1376];
        layer3[43][47:40] = buffer_data_3[1391:1384];
        layer3[43][55:48] = buffer_data_3[1399:1392];
        layer4[43][7:0] = buffer_data_2[1351:1344];
        layer4[43][15:8] = buffer_data_2[1359:1352];
        layer4[43][23:16] = buffer_data_2[1367:1360];
        layer4[43][31:24] = buffer_data_2[1375:1368];
        layer4[43][39:32] = buffer_data_2[1383:1376];
        layer4[43][47:40] = buffer_data_2[1391:1384];
        layer4[43][55:48] = buffer_data_2[1399:1392];
        layer5[43][7:0] = buffer_data_1[1351:1344];
        layer5[43][15:8] = buffer_data_1[1359:1352];
        layer5[43][23:16] = buffer_data_1[1367:1360];
        layer5[43][31:24] = buffer_data_1[1375:1368];
        layer5[43][39:32] = buffer_data_1[1383:1376];
        layer5[43][47:40] = buffer_data_1[1391:1384];
        layer5[43][55:48] = buffer_data_1[1399:1392];
        layer6[43][7:0] = buffer_data_0[1351:1344];
        layer6[43][15:8] = buffer_data_0[1359:1352];
        layer6[43][23:16] = buffer_data_0[1367:1360];
        layer6[43][31:24] = buffer_data_0[1375:1368];
        layer6[43][39:32] = buffer_data_0[1383:1376];
        layer6[43][47:40] = buffer_data_0[1391:1384];
        layer6[43][55:48] = buffer_data_0[1399:1392];
        layer0[44][7:0] = buffer_data_6[1359:1352];
        layer0[44][15:8] = buffer_data_6[1367:1360];
        layer0[44][23:16] = buffer_data_6[1375:1368];
        layer0[44][31:24] = buffer_data_6[1383:1376];
        layer0[44][39:32] = buffer_data_6[1391:1384];
        layer0[44][47:40] = buffer_data_6[1399:1392];
        layer0[44][55:48] = buffer_data_6[1407:1400];
        layer1[44][7:0] = buffer_data_5[1359:1352];
        layer1[44][15:8] = buffer_data_5[1367:1360];
        layer1[44][23:16] = buffer_data_5[1375:1368];
        layer1[44][31:24] = buffer_data_5[1383:1376];
        layer1[44][39:32] = buffer_data_5[1391:1384];
        layer1[44][47:40] = buffer_data_5[1399:1392];
        layer1[44][55:48] = buffer_data_5[1407:1400];
        layer2[44][7:0] = buffer_data_4[1359:1352];
        layer2[44][15:8] = buffer_data_4[1367:1360];
        layer2[44][23:16] = buffer_data_4[1375:1368];
        layer2[44][31:24] = buffer_data_4[1383:1376];
        layer2[44][39:32] = buffer_data_4[1391:1384];
        layer2[44][47:40] = buffer_data_4[1399:1392];
        layer2[44][55:48] = buffer_data_4[1407:1400];
        layer3[44][7:0] = buffer_data_3[1359:1352];
        layer3[44][15:8] = buffer_data_3[1367:1360];
        layer3[44][23:16] = buffer_data_3[1375:1368];
        layer3[44][31:24] = buffer_data_3[1383:1376];
        layer3[44][39:32] = buffer_data_3[1391:1384];
        layer3[44][47:40] = buffer_data_3[1399:1392];
        layer3[44][55:48] = buffer_data_3[1407:1400];
        layer4[44][7:0] = buffer_data_2[1359:1352];
        layer4[44][15:8] = buffer_data_2[1367:1360];
        layer4[44][23:16] = buffer_data_2[1375:1368];
        layer4[44][31:24] = buffer_data_2[1383:1376];
        layer4[44][39:32] = buffer_data_2[1391:1384];
        layer4[44][47:40] = buffer_data_2[1399:1392];
        layer4[44][55:48] = buffer_data_2[1407:1400];
        layer5[44][7:0] = buffer_data_1[1359:1352];
        layer5[44][15:8] = buffer_data_1[1367:1360];
        layer5[44][23:16] = buffer_data_1[1375:1368];
        layer5[44][31:24] = buffer_data_1[1383:1376];
        layer5[44][39:32] = buffer_data_1[1391:1384];
        layer5[44][47:40] = buffer_data_1[1399:1392];
        layer5[44][55:48] = buffer_data_1[1407:1400];
        layer6[44][7:0] = buffer_data_0[1359:1352];
        layer6[44][15:8] = buffer_data_0[1367:1360];
        layer6[44][23:16] = buffer_data_0[1375:1368];
        layer6[44][31:24] = buffer_data_0[1383:1376];
        layer6[44][39:32] = buffer_data_0[1391:1384];
        layer6[44][47:40] = buffer_data_0[1399:1392];
        layer6[44][55:48] = buffer_data_0[1407:1400];
        layer0[45][7:0] = buffer_data_6[1367:1360];
        layer0[45][15:8] = buffer_data_6[1375:1368];
        layer0[45][23:16] = buffer_data_6[1383:1376];
        layer0[45][31:24] = buffer_data_6[1391:1384];
        layer0[45][39:32] = buffer_data_6[1399:1392];
        layer0[45][47:40] = buffer_data_6[1407:1400];
        layer0[45][55:48] = buffer_data_6[1415:1408];
        layer1[45][7:0] = buffer_data_5[1367:1360];
        layer1[45][15:8] = buffer_data_5[1375:1368];
        layer1[45][23:16] = buffer_data_5[1383:1376];
        layer1[45][31:24] = buffer_data_5[1391:1384];
        layer1[45][39:32] = buffer_data_5[1399:1392];
        layer1[45][47:40] = buffer_data_5[1407:1400];
        layer1[45][55:48] = buffer_data_5[1415:1408];
        layer2[45][7:0] = buffer_data_4[1367:1360];
        layer2[45][15:8] = buffer_data_4[1375:1368];
        layer2[45][23:16] = buffer_data_4[1383:1376];
        layer2[45][31:24] = buffer_data_4[1391:1384];
        layer2[45][39:32] = buffer_data_4[1399:1392];
        layer2[45][47:40] = buffer_data_4[1407:1400];
        layer2[45][55:48] = buffer_data_4[1415:1408];
        layer3[45][7:0] = buffer_data_3[1367:1360];
        layer3[45][15:8] = buffer_data_3[1375:1368];
        layer3[45][23:16] = buffer_data_3[1383:1376];
        layer3[45][31:24] = buffer_data_3[1391:1384];
        layer3[45][39:32] = buffer_data_3[1399:1392];
        layer3[45][47:40] = buffer_data_3[1407:1400];
        layer3[45][55:48] = buffer_data_3[1415:1408];
        layer4[45][7:0] = buffer_data_2[1367:1360];
        layer4[45][15:8] = buffer_data_2[1375:1368];
        layer4[45][23:16] = buffer_data_2[1383:1376];
        layer4[45][31:24] = buffer_data_2[1391:1384];
        layer4[45][39:32] = buffer_data_2[1399:1392];
        layer4[45][47:40] = buffer_data_2[1407:1400];
        layer4[45][55:48] = buffer_data_2[1415:1408];
        layer5[45][7:0] = buffer_data_1[1367:1360];
        layer5[45][15:8] = buffer_data_1[1375:1368];
        layer5[45][23:16] = buffer_data_1[1383:1376];
        layer5[45][31:24] = buffer_data_1[1391:1384];
        layer5[45][39:32] = buffer_data_1[1399:1392];
        layer5[45][47:40] = buffer_data_1[1407:1400];
        layer5[45][55:48] = buffer_data_1[1415:1408];
        layer6[45][7:0] = buffer_data_0[1367:1360];
        layer6[45][15:8] = buffer_data_0[1375:1368];
        layer6[45][23:16] = buffer_data_0[1383:1376];
        layer6[45][31:24] = buffer_data_0[1391:1384];
        layer6[45][39:32] = buffer_data_0[1399:1392];
        layer6[45][47:40] = buffer_data_0[1407:1400];
        layer6[45][55:48] = buffer_data_0[1415:1408];
        layer0[46][7:0] = buffer_data_6[1375:1368];
        layer0[46][15:8] = buffer_data_6[1383:1376];
        layer0[46][23:16] = buffer_data_6[1391:1384];
        layer0[46][31:24] = buffer_data_6[1399:1392];
        layer0[46][39:32] = buffer_data_6[1407:1400];
        layer0[46][47:40] = buffer_data_6[1415:1408];
        layer0[46][55:48] = buffer_data_6[1423:1416];
        layer1[46][7:0] = buffer_data_5[1375:1368];
        layer1[46][15:8] = buffer_data_5[1383:1376];
        layer1[46][23:16] = buffer_data_5[1391:1384];
        layer1[46][31:24] = buffer_data_5[1399:1392];
        layer1[46][39:32] = buffer_data_5[1407:1400];
        layer1[46][47:40] = buffer_data_5[1415:1408];
        layer1[46][55:48] = buffer_data_5[1423:1416];
        layer2[46][7:0] = buffer_data_4[1375:1368];
        layer2[46][15:8] = buffer_data_4[1383:1376];
        layer2[46][23:16] = buffer_data_4[1391:1384];
        layer2[46][31:24] = buffer_data_4[1399:1392];
        layer2[46][39:32] = buffer_data_4[1407:1400];
        layer2[46][47:40] = buffer_data_4[1415:1408];
        layer2[46][55:48] = buffer_data_4[1423:1416];
        layer3[46][7:0] = buffer_data_3[1375:1368];
        layer3[46][15:8] = buffer_data_3[1383:1376];
        layer3[46][23:16] = buffer_data_3[1391:1384];
        layer3[46][31:24] = buffer_data_3[1399:1392];
        layer3[46][39:32] = buffer_data_3[1407:1400];
        layer3[46][47:40] = buffer_data_3[1415:1408];
        layer3[46][55:48] = buffer_data_3[1423:1416];
        layer4[46][7:0] = buffer_data_2[1375:1368];
        layer4[46][15:8] = buffer_data_2[1383:1376];
        layer4[46][23:16] = buffer_data_2[1391:1384];
        layer4[46][31:24] = buffer_data_2[1399:1392];
        layer4[46][39:32] = buffer_data_2[1407:1400];
        layer4[46][47:40] = buffer_data_2[1415:1408];
        layer4[46][55:48] = buffer_data_2[1423:1416];
        layer5[46][7:0] = buffer_data_1[1375:1368];
        layer5[46][15:8] = buffer_data_1[1383:1376];
        layer5[46][23:16] = buffer_data_1[1391:1384];
        layer5[46][31:24] = buffer_data_1[1399:1392];
        layer5[46][39:32] = buffer_data_1[1407:1400];
        layer5[46][47:40] = buffer_data_1[1415:1408];
        layer5[46][55:48] = buffer_data_1[1423:1416];
        layer6[46][7:0] = buffer_data_0[1375:1368];
        layer6[46][15:8] = buffer_data_0[1383:1376];
        layer6[46][23:16] = buffer_data_0[1391:1384];
        layer6[46][31:24] = buffer_data_0[1399:1392];
        layer6[46][39:32] = buffer_data_0[1407:1400];
        layer6[46][47:40] = buffer_data_0[1415:1408];
        layer6[46][55:48] = buffer_data_0[1423:1416];
        layer0[47][7:0] = buffer_data_6[1383:1376];
        layer0[47][15:8] = buffer_data_6[1391:1384];
        layer0[47][23:16] = buffer_data_6[1399:1392];
        layer0[47][31:24] = buffer_data_6[1407:1400];
        layer0[47][39:32] = buffer_data_6[1415:1408];
        layer0[47][47:40] = buffer_data_6[1423:1416];
        layer0[47][55:48] = buffer_data_6[1431:1424];
        layer1[47][7:0] = buffer_data_5[1383:1376];
        layer1[47][15:8] = buffer_data_5[1391:1384];
        layer1[47][23:16] = buffer_data_5[1399:1392];
        layer1[47][31:24] = buffer_data_5[1407:1400];
        layer1[47][39:32] = buffer_data_5[1415:1408];
        layer1[47][47:40] = buffer_data_5[1423:1416];
        layer1[47][55:48] = buffer_data_5[1431:1424];
        layer2[47][7:0] = buffer_data_4[1383:1376];
        layer2[47][15:8] = buffer_data_4[1391:1384];
        layer2[47][23:16] = buffer_data_4[1399:1392];
        layer2[47][31:24] = buffer_data_4[1407:1400];
        layer2[47][39:32] = buffer_data_4[1415:1408];
        layer2[47][47:40] = buffer_data_4[1423:1416];
        layer2[47][55:48] = buffer_data_4[1431:1424];
        layer3[47][7:0] = buffer_data_3[1383:1376];
        layer3[47][15:8] = buffer_data_3[1391:1384];
        layer3[47][23:16] = buffer_data_3[1399:1392];
        layer3[47][31:24] = buffer_data_3[1407:1400];
        layer3[47][39:32] = buffer_data_3[1415:1408];
        layer3[47][47:40] = buffer_data_3[1423:1416];
        layer3[47][55:48] = buffer_data_3[1431:1424];
        layer4[47][7:0] = buffer_data_2[1383:1376];
        layer4[47][15:8] = buffer_data_2[1391:1384];
        layer4[47][23:16] = buffer_data_2[1399:1392];
        layer4[47][31:24] = buffer_data_2[1407:1400];
        layer4[47][39:32] = buffer_data_2[1415:1408];
        layer4[47][47:40] = buffer_data_2[1423:1416];
        layer4[47][55:48] = buffer_data_2[1431:1424];
        layer5[47][7:0] = buffer_data_1[1383:1376];
        layer5[47][15:8] = buffer_data_1[1391:1384];
        layer5[47][23:16] = buffer_data_1[1399:1392];
        layer5[47][31:24] = buffer_data_1[1407:1400];
        layer5[47][39:32] = buffer_data_1[1415:1408];
        layer5[47][47:40] = buffer_data_1[1423:1416];
        layer5[47][55:48] = buffer_data_1[1431:1424];
        layer6[47][7:0] = buffer_data_0[1383:1376];
        layer6[47][15:8] = buffer_data_0[1391:1384];
        layer6[47][23:16] = buffer_data_0[1399:1392];
        layer6[47][31:24] = buffer_data_0[1407:1400];
        layer6[47][39:32] = buffer_data_0[1415:1408];
        layer6[47][47:40] = buffer_data_0[1423:1416];
        layer6[47][55:48] = buffer_data_0[1431:1424];
        layer0[48][7:0] = buffer_data_6[1391:1384];
        layer0[48][15:8] = buffer_data_6[1399:1392];
        layer0[48][23:16] = buffer_data_6[1407:1400];
        layer0[48][31:24] = buffer_data_6[1415:1408];
        layer0[48][39:32] = buffer_data_6[1423:1416];
        layer0[48][47:40] = buffer_data_6[1431:1424];
        layer0[48][55:48] = buffer_data_6[1439:1432];
        layer1[48][7:0] = buffer_data_5[1391:1384];
        layer1[48][15:8] = buffer_data_5[1399:1392];
        layer1[48][23:16] = buffer_data_5[1407:1400];
        layer1[48][31:24] = buffer_data_5[1415:1408];
        layer1[48][39:32] = buffer_data_5[1423:1416];
        layer1[48][47:40] = buffer_data_5[1431:1424];
        layer1[48][55:48] = buffer_data_5[1439:1432];
        layer2[48][7:0] = buffer_data_4[1391:1384];
        layer2[48][15:8] = buffer_data_4[1399:1392];
        layer2[48][23:16] = buffer_data_4[1407:1400];
        layer2[48][31:24] = buffer_data_4[1415:1408];
        layer2[48][39:32] = buffer_data_4[1423:1416];
        layer2[48][47:40] = buffer_data_4[1431:1424];
        layer2[48][55:48] = buffer_data_4[1439:1432];
        layer3[48][7:0] = buffer_data_3[1391:1384];
        layer3[48][15:8] = buffer_data_3[1399:1392];
        layer3[48][23:16] = buffer_data_3[1407:1400];
        layer3[48][31:24] = buffer_data_3[1415:1408];
        layer3[48][39:32] = buffer_data_3[1423:1416];
        layer3[48][47:40] = buffer_data_3[1431:1424];
        layer3[48][55:48] = buffer_data_3[1439:1432];
        layer4[48][7:0] = buffer_data_2[1391:1384];
        layer4[48][15:8] = buffer_data_2[1399:1392];
        layer4[48][23:16] = buffer_data_2[1407:1400];
        layer4[48][31:24] = buffer_data_2[1415:1408];
        layer4[48][39:32] = buffer_data_2[1423:1416];
        layer4[48][47:40] = buffer_data_2[1431:1424];
        layer4[48][55:48] = buffer_data_2[1439:1432];
        layer5[48][7:0] = buffer_data_1[1391:1384];
        layer5[48][15:8] = buffer_data_1[1399:1392];
        layer5[48][23:16] = buffer_data_1[1407:1400];
        layer5[48][31:24] = buffer_data_1[1415:1408];
        layer5[48][39:32] = buffer_data_1[1423:1416];
        layer5[48][47:40] = buffer_data_1[1431:1424];
        layer5[48][55:48] = buffer_data_1[1439:1432];
        layer6[48][7:0] = buffer_data_0[1391:1384];
        layer6[48][15:8] = buffer_data_0[1399:1392];
        layer6[48][23:16] = buffer_data_0[1407:1400];
        layer6[48][31:24] = buffer_data_0[1415:1408];
        layer6[48][39:32] = buffer_data_0[1423:1416];
        layer6[48][47:40] = buffer_data_0[1431:1424];
        layer6[48][55:48] = buffer_data_0[1439:1432];
        layer0[49][7:0] = buffer_data_6[1399:1392];
        layer0[49][15:8] = buffer_data_6[1407:1400];
        layer0[49][23:16] = buffer_data_6[1415:1408];
        layer0[49][31:24] = buffer_data_6[1423:1416];
        layer0[49][39:32] = buffer_data_6[1431:1424];
        layer0[49][47:40] = buffer_data_6[1439:1432];
        layer0[49][55:48] = buffer_data_6[1447:1440];
        layer1[49][7:0] = buffer_data_5[1399:1392];
        layer1[49][15:8] = buffer_data_5[1407:1400];
        layer1[49][23:16] = buffer_data_5[1415:1408];
        layer1[49][31:24] = buffer_data_5[1423:1416];
        layer1[49][39:32] = buffer_data_5[1431:1424];
        layer1[49][47:40] = buffer_data_5[1439:1432];
        layer1[49][55:48] = buffer_data_5[1447:1440];
        layer2[49][7:0] = buffer_data_4[1399:1392];
        layer2[49][15:8] = buffer_data_4[1407:1400];
        layer2[49][23:16] = buffer_data_4[1415:1408];
        layer2[49][31:24] = buffer_data_4[1423:1416];
        layer2[49][39:32] = buffer_data_4[1431:1424];
        layer2[49][47:40] = buffer_data_4[1439:1432];
        layer2[49][55:48] = buffer_data_4[1447:1440];
        layer3[49][7:0] = buffer_data_3[1399:1392];
        layer3[49][15:8] = buffer_data_3[1407:1400];
        layer3[49][23:16] = buffer_data_3[1415:1408];
        layer3[49][31:24] = buffer_data_3[1423:1416];
        layer3[49][39:32] = buffer_data_3[1431:1424];
        layer3[49][47:40] = buffer_data_3[1439:1432];
        layer3[49][55:48] = buffer_data_3[1447:1440];
        layer4[49][7:0] = buffer_data_2[1399:1392];
        layer4[49][15:8] = buffer_data_2[1407:1400];
        layer4[49][23:16] = buffer_data_2[1415:1408];
        layer4[49][31:24] = buffer_data_2[1423:1416];
        layer4[49][39:32] = buffer_data_2[1431:1424];
        layer4[49][47:40] = buffer_data_2[1439:1432];
        layer4[49][55:48] = buffer_data_2[1447:1440];
        layer5[49][7:0] = buffer_data_1[1399:1392];
        layer5[49][15:8] = buffer_data_1[1407:1400];
        layer5[49][23:16] = buffer_data_1[1415:1408];
        layer5[49][31:24] = buffer_data_1[1423:1416];
        layer5[49][39:32] = buffer_data_1[1431:1424];
        layer5[49][47:40] = buffer_data_1[1439:1432];
        layer5[49][55:48] = buffer_data_1[1447:1440];
        layer6[49][7:0] = buffer_data_0[1399:1392];
        layer6[49][15:8] = buffer_data_0[1407:1400];
        layer6[49][23:16] = buffer_data_0[1415:1408];
        layer6[49][31:24] = buffer_data_0[1423:1416];
        layer6[49][39:32] = buffer_data_0[1431:1424];
        layer6[49][47:40] = buffer_data_0[1439:1432];
        layer6[49][55:48] = buffer_data_0[1447:1440];
        layer0[50][7:0] = buffer_data_6[1407:1400];
        layer0[50][15:8] = buffer_data_6[1415:1408];
        layer0[50][23:16] = buffer_data_6[1423:1416];
        layer0[50][31:24] = buffer_data_6[1431:1424];
        layer0[50][39:32] = buffer_data_6[1439:1432];
        layer0[50][47:40] = buffer_data_6[1447:1440];
        layer0[50][55:48] = buffer_data_6[1455:1448];
        layer1[50][7:0] = buffer_data_5[1407:1400];
        layer1[50][15:8] = buffer_data_5[1415:1408];
        layer1[50][23:16] = buffer_data_5[1423:1416];
        layer1[50][31:24] = buffer_data_5[1431:1424];
        layer1[50][39:32] = buffer_data_5[1439:1432];
        layer1[50][47:40] = buffer_data_5[1447:1440];
        layer1[50][55:48] = buffer_data_5[1455:1448];
        layer2[50][7:0] = buffer_data_4[1407:1400];
        layer2[50][15:8] = buffer_data_4[1415:1408];
        layer2[50][23:16] = buffer_data_4[1423:1416];
        layer2[50][31:24] = buffer_data_4[1431:1424];
        layer2[50][39:32] = buffer_data_4[1439:1432];
        layer2[50][47:40] = buffer_data_4[1447:1440];
        layer2[50][55:48] = buffer_data_4[1455:1448];
        layer3[50][7:0] = buffer_data_3[1407:1400];
        layer3[50][15:8] = buffer_data_3[1415:1408];
        layer3[50][23:16] = buffer_data_3[1423:1416];
        layer3[50][31:24] = buffer_data_3[1431:1424];
        layer3[50][39:32] = buffer_data_3[1439:1432];
        layer3[50][47:40] = buffer_data_3[1447:1440];
        layer3[50][55:48] = buffer_data_3[1455:1448];
        layer4[50][7:0] = buffer_data_2[1407:1400];
        layer4[50][15:8] = buffer_data_2[1415:1408];
        layer4[50][23:16] = buffer_data_2[1423:1416];
        layer4[50][31:24] = buffer_data_2[1431:1424];
        layer4[50][39:32] = buffer_data_2[1439:1432];
        layer4[50][47:40] = buffer_data_2[1447:1440];
        layer4[50][55:48] = buffer_data_2[1455:1448];
        layer5[50][7:0] = buffer_data_1[1407:1400];
        layer5[50][15:8] = buffer_data_1[1415:1408];
        layer5[50][23:16] = buffer_data_1[1423:1416];
        layer5[50][31:24] = buffer_data_1[1431:1424];
        layer5[50][39:32] = buffer_data_1[1439:1432];
        layer5[50][47:40] = buffer_data_1[1447:1440];
        layer5[50][55:48] = buffer_data_1[1455:1448];
        layer6[50][7:0] = buffer_data_0[1407:1400];
        layer6[50][15:8] = buffer_data_0[1415:1408];
        layer6[50][23:16] = buffer_data_0[1423:1416];
        layer6[50][31:24] = buffer_data_0[1431:1424];
        layer6[50][39:32] = buffer_data_0[1439:1432];
        layer6[50][47:40] = buffer_data_0[1447:1440];
        layer6[50][55:48] = buffer_data_0[1455:1448];
        layer0[51][7:0] = buffer_data_6[1415:1408];
        layer0[51][15:8] = buffer_data_6[1423:1416];
        layer0[51][23:16] = buffer_data_6[1431:1424];
        layer0[51][31:24] = buffer_data_6[1439:1432];
        layer0[51][39:32] = buffer_data_6[1447:1440];
        layer0[51][47:40] = buffer_data_6[1455:1448];
        layer0[51][55:48] = buffer_data_6[1463:1456];
        layer1[51][7:0] = buffer_data_5[1415:1408];
        layer1[51][15:8] = buffer_data_5[1423:1416];
        layer1[51][23:16] = buffer_data_5[1431:1424];
        layer1[51][31:24] = buffer_data_5[1439:1432];
        layer1[51][39:32] = buffer_data_5[1447:1440];
        layer1[51][47:40] = buffer_data_5[1455:1448];
        layer1[51][55:48] = buffer_data_5[1463:1456];
        layer2[51][7:0] = buffer_data_4[1415:1408];
        layer2[51][15:8] = buffer_data_4[1423:1416];
        layer2[51][23:16] = buffer_data_4[1431:1424];
        layer2[51][31:24] = buffer_data_4[1439:1432];
        layer2[51][39:32] = buffer_data_4[1447:1440];
        layer2[51][47:40] = buffer_data_4[1455:1448];
        layer2[51][55:48] = buffer_data_4[1463:1456];
        layer3[51][7:0] = buffer_data_3[1415:1408];
        layer3[51][15:8] = buffer_data_3[1423:1416];
        layer3[51][23:16] = buffer_data_3[1431:1424];
        layer3[51][31:24] = buffer_data_3[1439:1432];
        layer3[51][39:32] = buffer_data_3[1447:1440];
        layer3[51][47:40] = buffer_data_3[1455:1448];
        layer3[51][55:48] = buffer_data_3[1463:1456];
        layer4[51][7:0] = buffer_data_2[1415:1408];
        layer4[51][15:8] = buffer_data_2[1423:1416];
        layer4[51][23:16] = buffer_data_2[1431:1424];
        layer4[51][31:24] = buffer_data_2[1439:1432];
        layer4[51][39:32] = buffer_data_2[1447:1440];
        layer4[51][47:40] = buffer_data_2[1455:1448];
        layer4[51][55:48] = buffer_data_2[1463:1456];
        layer5[51][7:0] = buffer_data_1[1415:1408];
        layer5[51][15:8] = buffer_data_1[1423:1416];
        layer5[51][23:16] = buffer_data_1[1431:1424];
        layer5[51][31:24] = buffer_data_1[1439:1432];
        layer5[51][39:32] = buffer_data_1[1447:1440];
        layer5[51][47:40] = buffer_data_1[1455:1448];
        layer5[51][55:48] = buffer_data_1[1463:1456];
        layer6[51][7:0] = buffer_data_0[1415:1408];
        layer6[51][15:8] = buffer_data_0[1423:1416];
        layer6[51][23:16] = buffer_data_0[1431:1424];
        layer6[51][31:24] = buffer_data_0[1439:1432];
        layer6[51][39:32] = buffer_data_0[1447:1440];
        layer6[51][47:40] = buffer_data_0[1455:1448];
        layer6[51][55:48] = buffer_data_0[1463:1456];
        layer0[52][7:0] = buffer_data_6[1423:1416];
        layer0[52][15:8] = buffer_data_6[1431:1424];
        layer0[52][23:16] = buffer_data_6[1439:1432];
        layer0[52][31:24] = buffer_data_6[1447:1440];
        layer0[52][39:32] = buffer_data_6[1455:1448];
        layer0[52][47:40] = buffer_data_6[1463:1456];
        layer0[52][55:48] = buffer_data_6[1471:1464];
        layer1[52][7:0] = buffer_data_5[1423:1416];
        layer1[52][15:8] = buffer_data_5[1431:1424];
        layer1[52][23:16] = buffer_data_5[1439:1432];
        layer1[52][31:24] = buffer_data_5[1447:1440];
        layer1[52][39:32] = buffer_data_5[1455:1448];
        layer1[52][47:40] = buffer_data_5[1463:1456];
        layer1[52][55:48] = buffer_data_5[1471:1464];
        layer2[52][7:0] = buffer_data_4[1423:1416];
        layer2[52][15:8] = buffer_data_4[1431:1424];
        layer2[52][23:16] = buffer_data_4[1439:1432];
        layer2[52][31:24] = buffer_data_4[1447:1440];
        layer2[52][39:32] = buffer_data_4[1455:1448];
        layer2[52][47:40] = buffer_data_4[1463:1456];
        layer2[52][55:48] = buffer_data_4[1471:1464];
        layer3[52][7:0] = buffer_data_3[1423:1416];
        layer3[52][15:8] = buffer_data_3[1431:1424];
        layer3[52][23:16] = buffer_data_3[1439:1432];
        layer3[52][31:24] = buffer_data_3[1447:1440];
        layer3[52][39:32] = buffer_data_3[1455:1448];
        layer3[52][47:40] = buffer_data_3[1463:1456];
        layer3[52][55:48] = buffer_data_3[1471:1464];
        layer4[52][7:0] = buffer_data_2[1423:1416];
        layer4[52][15:8] = buffer_data_2[1431:1424];
        layer4[52][23:16] = buffer_data_2[1439:1432];
        layer4[52][31:24] = buffer_data_2[1447:1440];
        layer4[52][39:32] = buffer_data_2[1455:1448];
        layer4[52][47:40] = buffer_data_2[1463:1456];
        layer4[52][55:48] = buffer_data_2[1471:1464];
        layer5[52][7:0] = buffer_data_1[1423:1416];
        layer5[52][15:8] = buffer_data_1[1431:1424];
        layer5[52][23:16] = buffer_data_1[1439:1432];
        layer5[52][31:24] = buffer_data_1[1447:1440];
        layer5[52][39:32] = buffer_data_1[1455:1448];
        layer5[52][47:40] = buffer_data_1[1463:1456];
        layer5[52][55:48] = buffer_data_1[1471:1464];
        layer6[52][7:0] = buffer_data_0[1423:1416];
        layer6[52][15:8] = buffer_data_0[1431:1424];
        layer6[52][23:16] = buffer_data_0[1439:1432];
        layer6[52][31:24] = buffer_data_0[1447:1440];
        layer6[52][39:32] = buffer_data_0[1455:1448];
        layer6[52][47:40] = buffer_data_0[1463:1456];
        layer6[52][55:48] = buffer_data_0[1471:1464];
        layer0[53][7:0] = buffer_data_6[1431:1424];
        layer0[53][15:8] = buffer_data_6[1439:1432];
        layer0[53][23:16] = buffer_data_6[1447:1440];
        layer0[53][31:24] = buffer_data_6[1455:1448];
        layer0[53][39:32] = buffer_data_6[1463:1456];
        layer0[53][47:40] = buffer_data_6[1471:1464];
        layer0[53][55:48] = buffer_data_6[1479:1472];
        layer1[53][7:0] = buffer_data_5[1431:1424];
        layer1[53][15:8] = buffer_data_5[1439:1432];
        layer1[53][23:16] = buffer_data_5[1447:1440];
        layer1[53][31:24] = buffer_data_5[1455:1448];
        layer1[53][39:32] = buffer_data_5[1463:1456];
        layer1[53][47:40] = buffer_data_5[1471:1464];
        layer1[53][55:48] = buffer_data_5[1479:1472];
        layer2[53][7:0] = buffer_data_4[1431:1424];
        layer2[53][15:8] = buffer_data_4[1439:1432];
        layer2[53][23:16] = buffer_data_4[1447:1440];
        layer2[53][31:24] = buffer_data_4[1455:1448];
        layer2[53][39:32] = buffer_data_4[1463:1456];
        layer2[53][47:40] = buffer_data_4[1471:1464];
        layer2[53][55:48] = buffer_data_4[1479:1472];
        layer3[53][7:0] = buffer_data_3[1431:1424];
        layer3[53][15:8] = buffer_data_3[1439:1432];
        layer3[53][23:16] = buffer_data_3[1447:1440];
        layer3[53][31:24] = buffer_data_3[1455:1448];
        layer3[53][39:32] = buffer_data_3[1463:1456];
        layer3[53][47:40] = buffer_data_3[1471:1464];
        layer3[53][55:48] = buffer_data_3[1479:1472];
        layer4[53][7:0] = buffer_data_2[1431:1424];
        layer4[53][15:8] = buffer_data_2[1439:1432];
        layer4[53][23:16] = buffer_data_2[1447:1440];
        layer4[53][31:24] = buffer_data_2[1455:1448];
        layer4[53][39:32] = buffer_data_2[1463:1456];
        layer4[53][47:40] = buffer_data_2[1471:1464];
        layer4[53][55:48] = buffer_data_2[1479:1472];
        layer5[53][7:0] = buffer_data_1[1431:1424];
        layer5[53][15:8] = buffer_data_1[1439:1432];
        layer5[53][23:16] = buffer_data_1[1447:1440];
        layer5[53][31:24] = buffer_data_1[1455:1448];
        layer5[53][39:32] = buffer_data_1[1463:1456];
        layer5[53][47:40] = buffer_data_1[1471:1464];
        layer5[53][55:48] = buffer_data_1[1479:1472];
        layer6[53][7:0] = buffer_data_0[1431:1424];
        layer6[53][15:8] = buffer_data_0[1439:1432];
        layer6[53][23:16] = buffer_data_0[1447:1440];
        layer6[53][31:24] = buffer_data_0[1455:1448];
        layer6[53][39:32] = buffer_data_0[1463:1456];
        layer6[53][47:40] = buffer_data_0[1471:1464];
        layer6[53][55:48] = buffer_data_0[1479:1472];
        layer0[54][7:0] = buffer_data_6[1439:1432];
        layer0[54][15:8] = buffer_data_6[1447:1440];
        layer0[54][23:16] = buffer_data_6[1455:1448];
        layer0[54][31:24] = buffer_data_6[1463:1456];
        layer0[54][39:32] = buffer_data_6[1471:1464];
        layer0[54][47:40] = buffer_data_6[1479:1472];
        layer0[54][55:48] = buffer_data_6[1487:1480];
        layer1[54][7:0] = buffer_data_5[1439:1432];
        layer1[54][15:8] = buffer_data_5[1447:1440];
        layer1[54][23:16] = buffer_data_5[1455:1448];
        layer1[54][31:24] = buffer_data_5[1463:1456];
        layer1[54][39:32] = buffer_data_5[1471:1464];
        layer1[54][47:40] = buffer_data_5[1479:1472];
        layer1[54][55:48] = buffer_data_5[1487:1480];
        layer2[54][7:0] = buffer_data_4[1439:1432];
        layer2[54][15:8] = buffer_data_4[1447:1440];
        layer2[54][23:16] = buffer_data_4[1455:1448];
        layer2[54][31:24] = buffer_data_4[1463:1456];
        layer2[54][39:32] = buffer_data_4[1471:1464];
        layer2[54][47:40] = buffer_data_4[1479:1472];
        layer2[54][55:48] = buffer_data_4[1487:1480];
        layer3[54][7:0] = buffer_data_3[1439:1432];
        layer3[54][15:8] = buffer_data_3[1447:1440];
        layer3[54][23:16] = buffer_data_3[1455:1448];
        layer3[54][31:24] = buffer_data_3[1463:1456];
        layer3[54][39:32] = buffer_data_3[1471:1464];
        layer3[54][47:40] = buffer_data_3[1479:1472];
        layer3[54][55:48] = buffer_data_3[1487:1480];
        layer4[54][7:0] = buffer_data_2[1439:1432];
        layer4[54][15:8] = buffer_data_2[1447:1440];
        layer4[54][23:16] = buffer_data_2[1455:1448];
        layer4[54][31:24] = buffer_data_2[1463:1456];
        layer4[54][39:32] = buffer_data_2[1471:1464];
        layer4[54][47:40] = buffer_data_2[1479:1472];
        layer4[54][55:48] = buffer_data_2[1487:1480];
        layer5[54][7:0] = buffer_data_1[1439:1432];
        layer5[54][15:8] = buffer_data_1[1447:1440];
        layer5[54][23:16] = buffer_data_1[1455:1448];
        layer5[54][31:24] = buffer_data_1[1463:1456];
        layer5[54][39:32] = buffer_data_1[1471:1464];
        layer5[54][47:40] = buffer_data_1[1479:1472];
        layer5[54][55:48] = buffer_data_1[1487:1480];
        layer6[54][7:0] = buffer_data_0[1439:1432];
        layer6[54][15:8] = buffer_data_0[1447:1440];
        layer6[54][23:16] = buffer_data_0[1455:1448];
        layer6[54][31:24] = buffer_data_0[1463:1456];
        layer6[54][39:32] = buffer_data_0[1471:1464];
        layer6[54][47:40] = buffer_data_0[1479:1472];
        layer6[54][55:48] = buffer_data_0[1487:1480];
        layer0[55][7:0] = buffer_data_6[1447:1440];
        layer0[55][15:8] = buffer_data_6[1455:1448];
        layer0[55][23:16] = buffer_data_6[1463:1456];
        layer0[55][31:24] = buffer_data_6[1471:1464];
        layer0[55][39:32] = buffer_data_6[1479:1472];
        layer0[55][47:40] = buffer_data_6[1487:1480];
        layer0[55][55:48] = buffer_data_6[1495:1488];
        layer1[55][7:0] = buffer_data_5[1447:1440];
        layer1[55][15:8] = buffer_data_5[1455:1448];
        layer1[55][23:16] = buffer_data_5[1463:1456];
        layer1[55][31:24] = buffer_data_5[1471:1464];
        layer1[55][39:32] = buffer_data_5[1479:1472];
        layer1[55][47:40] = buffer_data_5[1487:1480];
        layer1[55][55:48] = buffer_data_5[1495:1488];
        layer2[55][7:0] = buffer_data_4[1447:1440];
        layer2[55][15:8] = buffer_data_4[1455:1448];
        layer2[55][23:16] = buffer_data_4[1463:1456];
        layer2[55][31:24] = buffer_data_4[1471:1464];
        layer2[55][39:32] = buffer_data_4[1479:1472];
        layer2[55][47:40] = buffer_data_4[1487:1480];
        layer2[55][55:48] = buffer_data_4[1495:1488];
        layer3[55][7:0] = buffer_data_3[1447:1440];
        layer3[55][15:8] = buffer_data_3[1455:1448];
        layer3[55][23:16] = buffer_data_3[1463:1456];
        layer3[55][31:24] = buffer_data_3[1471:1464];
        layer3[55][39:32] = buffer_data_3[1479:1472];
        layer3[55][47:40] = buffer_data_3[1487:1480];
        layer3[55][55:48] = buffer_data_3[1495:1488];
        layer4[55][7:0] = buffer_data_2[1447:1440];
        layer4[55][15:8] = buffer_data_2[1455:1448];
        layer4[55][23:16] = buffer_data_2[1463:1456];
        layer4[55][31:24] = buffer_data_2[1471:1464];
        layer4[55][39:32] = buffer_data_2[1479:1472];
        layer4[55][47:40] = buffer_data_2[1487:1480];
        layer4[55][55:48] = buffer_data_2[1495:1488];
        layer5[55][7:0] = buffer_data_1[1447:1440];
        layer5[55][15:8] = buffer_data_1[1455:1448];
        layer5[55][23:16] = buffer_data_1[1463:1456];
        layer5[55][31:24] = buffer_data_1[1471:1464];
        layer5[55][39:32] = buffer_data_1[1479:1472];
        layer5[55][47:40] = buffer_data_1[1487:1480];
        layer5[55][55:48] = buffer_data_1[1495:1488];
        layer6[55][7:0] = buffer_data_0[1447:1440];
        layer6[55][15:8] = buffer_data_0[1455:1448];
        layer6[55][23:16] = buffer_data_0[1463:1456];
        layer6[55][31:24] = buffer_data_0[1471:1464];
        layer6[55][39:32] = buffer_data_0[1479:1472];
        layer6[55][47:40] = buffer_data_0[1487:1480];
        layer6[55][55:48] = buffer_data_0[1495:1488];
        layer0[56][7:0] = buffer_data_6[1455:1448];
        layer0[56][15:8] = buffer_data_6[1463:1456];
        layer0[56][23:16] = buffer_data_6[1471:1464];
        layer0[56][31:24] = buffer_data_6[1479:1472];
        layer0[56][39:32] = buffer_data_6[1487:1480];
        layer0[56][47:40] = buffer_data_6[1495:1488];
        layer0[56][55:48] = buffer_data_6[1503:1496];
        layer1[56][7:0] = buffer_data_5[1455:1448];
        layer1[56][15:8] = buffer_data_5[1463:1456];
        layer1[56][23:16] = buffer_data_5[1471:1464];
        layer1[56][31:24] = buffer_data_5[1479:1472];
        layer1[56][39:32] = buffer_data_5[1487:1480];
        layer1[56][47:40] = buffer_data_5[1495:1488];
        layer1[56][55:48] = buffer_data_5[1503:1496];
        layer2[56][7:0] = buffer_data_4[1455:1448];
        layer2[56][15:8] = buffer_data_4[1463:1456];
        layer2[56][23:16] = buffer_data_4[1471:1464];
        layer2[56][31:24] = buffer_data_4[1479:1472];
        layer2[56][39:32] = buffer_data_4[1487:1480];
        layer2[56][47:40] = buffer_data_4[1495:1488];
        layer2[56][55:48] = buffer_data_4[1503:1496];
        layer3[56][7:0] = buffer_data_3[1455:1448];
        layer3[56][15:8] = buffer_data_3[1463:1456];
        layer3[56][23:16] = buffer_data_3[1471:1464];
        layer3[56][31:24] = buffer_data_3[1479:1472];
        layer3[56][39:32] = buffer_data_3[1487:1480];
        layer3[56][47:40] = buffer_data_3[1495:1488];
        layer3[56][55:48] = buffer_data_3[1503:1496];
        layer4[56][7:0] = buffer_data_2[1455:1448];
        layer4[56][15:8] = buffer_data_2[1463:1456];
        layer4[56][23:16] = buffer_data_2[1471:1464];
        layer4[56][31:24] = buffer_data_2[1479:1472];
        layer4[56][39:32] = buffer_data_2[1487:1480];
        layer4[56][47:40] = buffer_data_2[1495:1488];
        layer4[56][55:48] = buffer_data_2[1503:1496];
        layer5[56][7:0] = buffer_data_1[1455:1448];
        layer5[56][15:8] = buffer_data_1[1463:1456];
        layer5[56][23:16] = buffer_data_1[1471:1464];
        layer5[56][31:24] = buffer_data_1[1479:1472];
        layer5[56][39:32] = buffer_data_1[1487:1480];
        layer5[56][47:40] = buffer_data_1[1495:1488];
        layer5[56][55:48] = buffer_data_1[1503:1496];
        layer6[56][7:0] = buffer_data_0[1455:1448];
        layer6[56][15:8] = buffer_data_0[1463:1456];
        layer6[56][23:16] = buffer_data_0[1471:1464];
        layer6[56][31:24] = buffer_data_0[1479:1472];
        layer6[56][39:32] = buffer_data_0[1487:1480];
        layer6[56][47:40] = buffer_data_0[1495:1488];
        layer6[56][55:48] = buffer_data_0[1503:1496];
        layer0[57][7:0] = buffer_data_6[1463:1456];
        layer0[57][15:8] = buffer_data_6[1471:1464];
        layer0[57][23:16] = buffer_data_6[1479:1472];
        layer0[57][31:24] = buffer_data_6[1487:1480];
        layer0[57][39:32] = buffer_data_6[1495:1488];
        layer0[57][47:40] = buffer_data_6[1503:1496];
        layer0[57][55:48] = buffer_data_6[1511:1504];
        layer1[57][7:0] = buffer_data_5[1463:1456];
        layer1[57][15:8] = buffer_data_5[1471:1464];
        layer1[57][23:16] = buffer_data_5[1479:1472];
        layer1[57][31:24] = buffer_data_5[1487:1480];
        layer1[57][39:32] = buffer_data_5[1495:1488];
        layer1[57][47:40] = buffer_data_5[1503:1496];
        layer1[57][55:48] = buffer_data_5[1511:1504];
        layer2[57][7:0] = buffer_data_4[1463:1456];
        layer2[57][15:8] = buffer_data_4[1471:1464];
        layer2[57][23:16] = buffer_data_4[1479:1472];
        layer2[57][31:24] = buffer_data_4[1487:1480];
        layer2[57][39:32] = buffer_data_4[1495:1488];
        layer2[57][47:40] = buffer_data_4[1503:1496];
        layer2[57][55:48] = buffer_data_4[1511:1504];
        layer3[57][7:0] = buffer_data_3[1463:1456];
        layer3[57][15:8] = buffer_data_3[1471:1464];
        layer3[57][23:16] = buffer_data_3[1479:1472];
        layer3[57][31:24] = buffer_data_3[1487:1480];
        layer3[57][39:32] = buffer_data_3[1495:1488];
        layer3[57][47:40] = buffer_data_3[1503:1496];
        layer3[57][55:48] = buffer_data_3[1511:1504];
        layer4[57][7:0] = buffer_data_2[1463:1456];
        layer4[57][15:8] = buffer_data_2[1471:1464];
        layer4[57][23:16] = buffer_data_2[1479:1472];
        layer4[57][31:24] = buffer_data_2[1487:1480];
        layer4[57][39:32] = buffer_data_2[1495:1488];
        layer4[57][47:40] = buffer_data_2[1503:1496];
        layer4[57][55:48] = buffer_data_2[1511:1504];
        layer5[57][7:0] = buffer_data_1[1463:1456];
        layer5[57][15:8] = buffer_data_1[1471:1464];
        layer5[57][23:16] = buffer_data_1[1479:1472];
        layer5[57][31:24] = buffer_data_1[1487:1480];
        layer5[57][39:32] = buffer_data_1[1495:1488];
        layer5[57][47:40] = buffer_data_1[1503:1496];
        layer5[57][55:48] = buffer_data_1[1511:1504];
        layer6[57][7:0] = buffer_data_0[1463:1456];
        layer6[57][15:8] = buffer_data_0[1471:1464];
        layer6[57][23:16] = buffer_data_0[1479:1472];
        layer6[57][31:24] = buffer_data_0[1487:1480];
        layer6[57][39:32] = buffer_data_0[1495:1488];
        layer6[57][47:40] = buffer_data_0[1503:1496];
        layer6[57][55:48] = buffer_data_0[1511:1504];
        layer0[58][7:0] = buffer_data_6[1471:1464];
        layer0[58][15:8] = buffer_data_6[1479:1472];
        layer0[58][23:16] = buffer_data_6[1487:1480];
        layer0[58][31:24] = buffer_data_6[1495:1488];
        layer0[58][39:32] = buffer_data_6[1503:1496];
        layer0[58][47:40] = buffer_data_6[1511:1504];
        layer0[58][55:48] = buffer_data_6[1519:1512];
        layer1[58][7:0] = buffer_data_5[1471:1464];
        layer1[58][15:8] = buffer_data_5[1479:1472];
        layer1[58][23:16] = buffer_data_5[1487:1480];
        layer1[58][31:24] = buffer_data_5[1495:1488];
        layer1[58][39:32] = buffer_data_5[1503:1496];
        layer1[58][47:40] = buffer_data_5[1511:1504];
        layer1[58][55:48] = buffer_data_5[1519:1512];
        layer2[58][7:0] = buffer_data_4[1471:1464];
        layer2[58][15:8] = buffer_data_4[1479:1472];
        layer2[58][23:16] = buffer_data_4[1487:1480];
        layer2[58][31:24] = buffer_data_4[1495:1488];
        layer2[58][39:32] = buffer_data_4[1503:1496];
        layer2[58][47:40] = buffer_data_4[1511:1504];
        layer2[58][55:48] = buffer_data_4[1519:1512];
        layer3[58][7:0] = buffer_data_3[1471:1464];
        layer3[58][15:8] = buffer_data_3[1479:1472];
        layer3[58][23:16] = buffer_data_3[1487:1480];
        layer3[58][31:24] = buffer_data_3[1495:1488];
        layer3[58][39:32] = buffer_data_3[1503:1496];
        layer3[58][47:40] = buffer_data_3[1511:1504];
        layer3[58][55:48] = buffer_data_3[1519:1512];
        layer4[58][7:0] = buffer_data_2[1471:1464];
        layer4[58][15:8] = buffer_data_2[1479:1472];
        layer4[58][23:16] = buffer_data_2[1487:1480];
        layer4[58][31:24] = buffer_data_2[1495:1488];
        layer4[58][39:32] = buffer_data_2[1503:1496];
        layer4[58][47:40] = buffer_data_2[1511:1504];
        layer4[58][55:48] = buffer_data_2[1519:1512];
        layer5[58][7:0] = buffer_data_1[1471:1464];
        layer5[58][15:8] = buffer_data_1[1479:1472];
        layer5[58][23:16] = buffer_data_1[1487:1480];
        layer5[58][31:24] = buffer_data_1[1495:1488];
        layer5[58][39:32] = buffer_data_1[1503:1496];
        layer5[58][47:40] = buffer_data_1[1511:1504];
        layer5[58][55:48] = buffer_data_1[1519:1512];
        layer6[58][7:0] = buffer_data_0[1471:1464];
        layer6[58][15:8] = buffer_data_0[1479:1472];
        layer6[58][23:16] = buffer_data_0[1487:1480];
        layer6[58][31:24] = buffer_data_0[1495:1488];
        layer6[58][39:32] = buffer_data_0[1503:1496];
        layer6[58][47:40] = buffer_data_0[1511:1504];
        layer6[58][55:48] = buffer_data_0[1519:1512];
        layer0[59][7:0] = buffer_data_6[1479:1472];
        layer0[59][15:8] = buffer_data_6[1487:1480];
        layer0[59][23:16] = buffer_data_6[1495:1488];
        layer0[59][31:24] = buffer_data_6[1503:1496];
        layer0[59][39:32] = buffer_data_6[1511:1504];
        layer0[59][47:40] = buffer_data_6[1519:1512];
        layer0[59][55:48] = buffer_data_6[1527:1520];
        layer1[59][7:0] = buffer_data_5[1479:1472];
        layer1[59][15:8] = buffer_data_5[1487:1480];
        layer1[59][23:16] = buffer_data_5[1495:1488];
        layer1[59][31:24] = buffer_data_5[1503:1496];
        layer1[59][39:32] = buffer_data_5[1511:1504];
        layer1[59][47:40] = buffer_data_5[1519:1512];
        layer1[59][55:48] = buffer_data_5[1527:1520];
        layer2[59][7:0] = buffer_data_4[1479:1472];
        layer2[59][15:8] = buffer_data_4[1487:1480];
        layer2[59][23:16] = buffer_data_4[1495:1488];
        layer2[59][31:24] = buffer_data_4[1503:1496];
        layer2[59][39:32] = buffer_data_4[1511:1504];
        layer2[59][47:40] = buffer_data_4[1519:1512];
        layer2[59][55:48] = buffer_data_4[1527:1520];
        layer3[59][7:0] = buffer_data_3[1479:1472];
        layer3[59][15:8] = buffer_data_3[1487:1480];
        layer3[59][23:16] = buffer_data_3[1495:1488];
        layer3[59][31:24] = buffer_data_3[1503:1496];
        layer3[59][39:32] = buffer_data_3[1511:1504];
        layer3[59][47:40] = buffer_data_3[1519:1512];
        layer3[59][55:48] = buffer_data_3[1527:1520];
        layer4[59][7:0] = buffer_data_2[1479:1472];
        layer4[59][15:8] = buffer_data_2[1487:1480];
        layer4[59][23:16] = buffer_data_2[1495:1488];
        layer4[59][31:24] = buffer_data_2[1503:1496];
        layer4[59][39:32] = buffer_data_2[1511:1504];
        layer4[59][47:40] = buffer_data_2[1519:1512];
        layer4[59][55:48] = buffer_data_2[1527:1520];
        layer5[59][7:0] = buffer_data_1[1479:1472];
        layer5[59][15:8] = buffer_data_1[1487:1480];
        layer5[59][23:16] = buffer_data_1[1495:1488];
        layer5[59][31:24] = buffer_data_1[1503:1496];
        layer5[59][39:32] = buffer_data_1[1511:1504];
        layer5[59][47:40] = buffer_data_1[1519:1512];
        layer5[59][55:48] = buffer_data_1[1527:1520];
        layer6[59][7:0] = buffer_data_0[1479:1472];
        layer6[59][15:8] = buffer_data_0[1487:1480];
        layer6[59][23:16] = buffer_data_0[1495:1488];
        layer6[59][31:24] = buffer_data_0[1503:1496];
        layer6[59][39:32] = buffer_data_0[1511:1504];
        layer6[59][47:40] = buffer_data_0[1519:1512];
        layer6[59][55:48] = buffer_data_0[1527:1520];
        layer0[60][7:0] = buffer_data_6[1487:1480];
        layer0[60][15:8] = buffer_data_6[1495:1488];
        layer0[60][23:16] = buffer_data_6[1503:1496];
        layer0[60][31:24] = buffer_data_6[1511:1504];
        layer0[60][39:32] = buffer_data_6[1519:1512];
        layer0[60][47:40] = buffer_data_6[1527:1520];
        layer0[60][55:48] = buffer_data_6[1535:1528];
        layer1[60][7:0] = buffer_data_5[1487:1480];
        layer1[60][15:8] = buffer_data_5[1495:1488];
        layer1[60][23:16] = buffer_data_5[1503:1496];
        layer1[60][31:24] = buffer_data_5[1511:1504];
        layer1[60][39:32] = buffer_data_5[1519:1512];
        layer1[60][47:40] = buffer_data_5[1527:1520];
        layer1[60][55:48] = buffer_data_5[1535:1528];
        layer2[60][7:0] = buffer_data_4[1487:1480];
        layer2[60][15:8] = buffer_data_4[1495:1488];
        layer2[60][23:16] = buffer_data_4[1503:1496];
        layer2[60][31:24] = buffer_data_4[1511:1504];
        layer2[60][39:32] = buffer_data_4[1519:1512];
        layer2[60][47:40] = buffer_data_4[1527:1520];
        layer2[60][55:48] = buffer_data_4[1535:1528];
        layer3[60][7:0] = buffer_data_3[1487:1480];
        layer3[60][15:8] = buffer_data_3[1495:1488];
        layer3[60][23:16] = buffer_data_3[1503:1496];
        layer3[60][31:24] = buffer_data_3[1511:1504];
        layer3[60][39:32] = buffer_data_3[1519:1512];
        layer3[60][47:40] = buffer_data_3[1527:1520];
        layer3[60][55:48] = buffer_data_3[1535:1528];
        layer4[60][7:0] = buffer_data_2[1487:1480];
        layer4[60][15:8] = buffer_data_2[1495:1488];
        layer4[60][23:16] = buffer_data_2[1503:1496];
        layer4[60][31:24] = buffer_data_2[1511:1504];
        layer4[60][39:32] = buffer_data_2[1519:1512];
        layer4[60][47:40] = buffer_data_2[1527:1520];
        layer4[60][55:48] = buffer_data_2[1535:1528];
        layer5[60][7:0] = buffer_data_1[1487:1480];
        layer5[60][15:8] = buffer_data_1[1495:1488];
        layer5[60][23:16] = buffer_data_1[1503:1496];
        layer5[60][31:24] = buffer_data_1[1511:1504];
        layer5[60][39:32] = buffer_data_1[1519:1512];
        layer5[60][47:40] = buffer_data_1[1527:1520];
        layer5[60][55:48] = buffer_data_1[1535:1528];
        layer6[60][7:0] = buffer_data_0[1487:1480];
        layer6[60][15:8] = buffer_data_0[1495:1488];
        layer6[60][23:16] = buffer_data_0[1503:1496];
        layer6[60][31:24] = buffer_data_0[1511:1504];
        layer6[60][39:32] = buffer_data_0[1519:1512];
        layer6[60][47:40] = buffer_data_0[1527:1520];
        layer6[60][55:48] = buffer_data_0[1535:1528];
        layer0[61][7:0] = buffer_data_6[1495:1488];
        layer0[61][15:8] = buffer_data_6[1503:1496];
        layer0[61][23:16] = buffer_data_6[1511:1504];
        layer0[61][31:24] = buffer_data_6[1519:1512];
        layer0[61][39:32] = buffer_data_6[1527:1520];
        layer0[61][47:40] = buffer_data_6[1535:1528];
        layer0[61][55:48] = buffer_data_6[1543:1536];
        layer1[61][7:0] = buffer_data_5[1495:1488];
        layer1[61][15:8] = buffer_data_5[1503:1496];
        layer1[61][23:16] = buffer_data_5[1511:1504];
        layer1[61][31:24] = buffer_data_5[1519:1512];
        layer1[61][39:32] = buffer_data_5[1527:1520];
        layer1[61][47:40] = buffer_data_5[1535:1528];
        layer1[61][55:48] = buffer_data_5[1543:1536];
        layer2[61][7:0] = buffer_data_4[1495:1488];
        layer2[61][15:8] = buffer_data_4[1503:1496];
        layer2[61][23:16] = buffer_data_4[1511:1504];
        layer2[61][31:24] = buffer_data_4[1519:1512];
        layer2[61][39:32] = buffer_data_4[1527:1520];
        layer2[61][47:40] = buffer_data_4[1535:1528];
        layer2[61][55:48] = buffer_data_4[1543:1536];
        layer3[61][7:0] = buffer_data_3[1495:1488];
        layer3[61][15:8] = buffer_data_3[1503:1496];
        layer3[61][23:16] = buffer_data_3[1511:1504];
        layer3[61][31:24] = buffer_data_3[1519:1512];
        layer3[61][39:32] = buffer_data_3[1527:1520];
        layer3[61][47:40] = buffer_data_3[1535:1528];
        layer3[61][55:48] = buffer_data_3[1543:1536];
        layer4[61][7:0] = buffer_data_2[1495:1488];
        layer4[61][15:8] = buffer_data_2[1503:1496];
        layer4[61][23:16] = buffer_data_2[1511:1504];
        layer4[61][31:24] = buffer_data_2[1519:1512];
        layer4[61][39:32] = buffer_data_2[1527:1520];
        layer4[61][47:40] = buffer_data_2[1535:1528];
        layer4[61][55:48] = buffer_data_2[1543:1536];
        layer5[61][7:0] = buffer_data_1[1495:1488];
        layer5[61][15:8] = buffer_data_1[1503:1496];
        layer5[61][23:16] = buffer_data_1[1511:1504];
        layer5[61][31:24] = buffer_data_1[1519:1512];
        layer5[61][39:32] = buffer_data_1[1527:1520];
        layer5[61][47:40] = buffer_data_1[1535:1528];
        layer5[61][55:48] = buffer_data_1[1543:1536];
        layer6[61][7:0] = buffer_data_0[1495:1488];
        layer6[61][15:8] = buffer_data_0[1503:1496];
        layer6[61][23:16] = buffer_data_0[1511:1504];
        layer6[61][31:24] = buffer_data_0[1519:1512];
        layer6[61][39:32] = buffer_data_0[1527:1520];
        layer6[61][47:40] = buffer_data_0[1535:1528];
        layer6[61][55:48] = buffer_data_0[1543:1536];
        layer0[62][7:0] = buffer_data_6[1503:1496];
        layer0[62][15:8] = buffer_data_6[1511:1504];
        layer0[62][23:16] = buffer_data_6[1519:1512];
        layer0[62][31:24] = buffer_data_6[1527:1520];
        layer0[62][39:32] = buffer_data_6[1535:1528];
        layer0[62][47:40] = buffer_data_6[1543:1536];
        layer0[62][55:48] = buffer_data_6[1551:1544];
        layer1[62][7:0] = buffer_data_5[1503:1496];
        layer1[62][15:8] = buffer_data_5[1511:1504];
        layer1[62][23:16] = buffer_data_5[1519:1512];
        layer1[62][31:24] = buffer_data_5[1527:1520];
        layer1[62][39:32] = buffer_data_5[1535:1528];
        layer1[62][47:40] = buffer_data_5[1543:1536];
        layer1[62][55:48] = buffer_data_5[1551:1544];
        layer2[62][7:0] = buffer_data_4[1503:1496];
        layer2[62][15:8] = buffer_data_4[1511:1504];
        layer2[62][23:16] = buffer_data_4[1519:1512];
        layer2[62][31:24] = buffer_data_4[1527:1520];
        layer2[62][39:32] = buffer_data_4[1535:1528];
        layer2[62][47:40] = buffer_data_4[1543:1536];
        layer2[62][55:48] = buffer_data_4[1551:1544];
        layer3[62][7:0] = buffer_data_3[1503:1496];
        layer3[62][15:8] = buffer_data_3[1511:1504];
        layer3[62][23:16] = buffer_data_3[1519:1512];
        layer3[62][31:24] = buffer_data_3[1527:1520];
        layer3[62][39:32] = buffer_data_3[1535:1528];
        layer3[62][47:40] = buffer_data_3[1543:1536];
        layer3[62][55:48] = buffer_data_3[1551:1544];
        layer4[62][7:0] = buffer_data_2[1503:1496];
        layer4[62][15:8] = buffer_data_2[1511:1504];
        layer4[62][23:16] = buffer_data_2[1519:1512];
        layer4[62][31:24] = buffer_data_2[1527:1520];
        layer4[62][39:32] = buffer_data_2[1535:1528];
        layer4[62][47:40] = buffer_data_2[1543:1536];
        layer4[62][55:48] = buffer_data_2[1551:1544];
        layer5[62][7:0] = buffer_data_1[1503:1496];
        layer5[62][15:8] = buffer_data_1[1511:1504];
        layer5[62][23:16] = buffer_data_1[1519:1512];
        layer5[62][31:24] = buffer_data_1[1527:1520];
        layer5[62][39:32] = buffer_data_1[1535:1528];
        layer5[62][47:40] = buffer_data_1[1543:1536];
        layer5[62][55:48] = buffer_data_1[1551:1544];
        layer6[62][7:0] = buffer_data_0[1503:1496];
        layer6[62][15:8] = buffer_data_0[1511:1504];
        layer6[62][23:16] = buffer_data_0[1519:1512];
        layer6[62][31:24] = buffer_data_0[1527:1520];
        layer6[62][39:32] = buffer_data_0[1535:1528];
        layer6[62][47:40] = buffer_data_0[1543:1536];
        layer6[62][55:48] = buffer_data_0[1551:1544];
        layer0[63][7:0] = buffer_data_6[1511:1504];
        layer0[63][15:8] = buffer_data_6[1519:1512];
        layer0[63][23:16] = buffer_data_6[1527:1520];
        layer0[63][31:24] = buffer_data_6[1535:1528];
        layer0[63][39:32] = buffer_data_6[1543:1536];
        layer0[63][47:40] = buffer_data_6[1551:1544];
        layer0[63][55:48] = buffer_data_6[1559:1552];
        layer1[63][7:0] = buffer_data_5[1511:1504];
        layer1[63][15:8] = buffer_data_5[1519:1512];
        layer1[63][23:16] = buffer_data_5[1527:1520];
        layer1[63][31:24] = buffer_data_5[1535:1528];
        layer1[63][39:32] = buffer_data_5[1543:1536];
        layer1[63][47:40] = buffer_data_5[1551:1544];
        layer1[63][55:48] = buffer_data_5[1559:1552];
        layer2[63][7:0] = buffer_data_4[1511:1504];
        layer2[63][15:8] = buffer_data_4[1519:1512];
        layer2[63][23:16] = buffer_data_4[1527:1520];
        layer2[63][31:24] = buffer_data_4[1535:1528];
        layer2[63][39:32] = buffer_data_4[1543:1536];
        layer2[63][47:40] = buffer_data_4[1551:1544];
        layer2[63][55:48] = buffer_data_4[1559:1552];
        layer3[63][7:0] = buffer_data_3[1511:1504];
        layer3[63][15:8] = buffer_data_3[1519:1512];
        layer3[63][23:16] = buffer_data_3[1527:1520];
        layer3[63][31:24] = buffer_data_3[1535:1528];
        layer3[63][39:32] = buffer_data_3[1543:1536];
        layer3[63][47:40] = buffer_data_3[1551:1544];
        layer3[63][55:48] = buffer_data_3[1559:1552];
        layer4[63][7:0] = buffer_data_2[1511:1504];
        layer4[63][15:8] = buffer_data_2[1519:1512];
        layer4[63][23:16] = buffer_data_2[1527:1520];
        layer4[63][31:24] = buffer_data_2[1535:1528];
        layer4[63][39:32] = buffer_data_2[1543:1536];
        layer4[63][47:40] = buffer_data_2[1551:1544];
        layer4[63][55:48] = buffer_data_2[1559:1552];
        layer5[63][7:0] = buffer_data_1[1511:1504];
        layer5[63][15:8] = buffer_data_1[1519:1512];
        layer5[63][23:16] = buffer_data_1[1527:1520];
        layer5[63][31:24] = buffer_data_1[1535:1528];
        layer5[63][39:32] = buffer_data_1[1543:1536];
        layer5[63][47:40] = buffer_data_1[1551:1544];
        layer5[63][55:48] = buffer_data_1[1559:1552];
        layer6[63][7:0] = buffer_data_0[1511:1504];
        layer6[63][15:8] = buffer_data_0[1519:1512];
        layer6[63][23:16] = buffer_data_0[1527:1520];
        layer6[63][31:24] = buffer_data_0[1535:1528];
        layer6[63][39:32] = buffer_data_0[1543:1536];
        layer6[63][47:40] = buffer_data_0[1551:1544];
        layer6[63][55:48] = buffer_data_0[1559:1552];
    end
    ST_GAUSSIAN_3: begin
        layer0[0][7:0] = buffer_data_6[1519:1512];
        layer0[0][15:8] = buffer_data_6[1527:1520];
        layer0[0][23:16] = buffer_data_6[1535:1528];
        layer0[0][31:24] = buffer_data_6[1543:1536];
        layer0[0][39:32] = buffer_data_6[1551:1544];
        layer0[0][47:40] = buffer_data_6[1559:1552];
        layer0[0][55:48] = buffer_data_6[1567:1560];
        layer1[0][7:0] = buffer_data_5[1519:1512];
        layer1[0][15:8] = buffer_data_5[1527:1520];
        layer1[0][23:16] = buffer_data_5[1535:1528];
        layer1[0][31:24] = buffer_data_5[1543:1536];
        layer1[0][39:32] = buffer_data_5[1551:1544];
        layer1[0][47:40] = buffer_data_5[1559:1552];
        layer1[0][55:48] = buffer_data_5[1567:1560];
        layer2[0][7:0] = buffer_data_4[1519:1512];
        layer2[0][15:8] = buffer_data_4[1527:1520];
        layer2[0][23:16] = buffer_data_4[1535:1528];
        layer2[0][31:24] = buffer_data_4[1543:1536];
        layer2[0][39:32] = buffer_data_4[1551:1544];
        layer2[0][47:40] = buffer_data_4[1559:1552];
        layer2[0][55:48] = buffer_data_4[1567:1560];
        layer3[0][7:0] = buffer_data_3[1519:1512];
        layer3[0][15:8] = buffer_data_3[1527:1520];
        layer3[0][23:16] = buffer_data_3[1535:1528];
        layer3[0][31:24] = buffer_data_3[1543:1536];
        layer3[0][39:32] = buffer_data_3[1551:1544];
        layer3[0][47:40] = buffer_data_3[1559:1552];
        layer3[0][55:48] = buffer_data_3[1567:1560];
        layer4[0][7:0] = buffer_data_2[1519:1512];
        layer4[0][15:8] = buffer_data_2[1527:1520];
        layer4[0][23:16] = buffer_data_2[1535:1528];
        layer4[0][31:24] = buffer_data_2[1543:1536];
        layer4[0][39:32] = buffer_data_2[1551:1544];
        layer4[0][47:40] = buffer_data_2[1559:1552];
        layer4[0][55:48] = buffer_data_2[1567:1560];
        layer5[0][7:0] = buffer_data_1[1519:1512];
        layer5[0][15:8] = buffer_data_1[1527:1520];
        layer5[0][23:16] = buffer_data_1[1535:1528];
        layer5[0][31:24] = buffer_data_1[1543:1536];
        layer5[0][39:32] = buffer_data_1[1551:1544];
        layer5[0][47:40] = buffer_data_1[1559:1552];
        layer5[0][55:48] = buffer_data_1[1567:1560];
        layer6[0][7:0] = buffer_data_0[1519:1512];
        layer6[0][15:8] = buffer_data_0[1527:1520];
        layer6[0][23:16] = buffer_data_0[1535:1528];
        layer6[0][31:24] = buffer_data_0[1543:1536];
        layer6[0][39:32] = buffer_data_0[1551:1544];
        layer6[0][47:40] = buffer_data_0[1559:1552];
        layer6[0][55:48] = buffer_data_0[1567:1560];
        layer0[1][7:0] = buffer_data_6[1527:1520];
        layer0[1][15:8] = buffer_data_6[1535:1528];
        layer0[1][23:16] = buffer_data_6[1543:1536];
        layer0[1][31:24] = buffer_data_6[1551:1544];
        layer0[1][39:32] = buffer_data_6[1559:1552];
        layer0[1][47:40] = buffer_data_6[1567:1560];
        layer0[1][55:48] = buffer_data_6[1575:1568];
        layer1[1][7:0] = buffer_data_5[1527:1520];
        layer1[1][15:8] = buffer_data_5[1535:1528];
        layer1[1][23:16] = buffer_data_5[1543:1536];
        layer1[1][31:24] = buffer_data_5[1551:1544];
        layer1[1][39:32] = buffer_data_5[1559:1552];
        layer1[1][47:40] = buffer_data_5[1567:1560];
        layer1[1][55:48] = buffer_data_5[1575:1568];
        layer2[1][7:0] = buffer_data_4[1527:1520];
        layer2[1][15:8] = buffer_data_4[1535:1528];
        layer2[1][23:16] = buffer_data_4[1543:1536];
        layer2[1][31:24] = buffer_data_4[1551:1544];
        layer2[1][39:32] = buffer_data_4[1559:1552];
        layer2[1][47:40] = buffer_data_4[1567:1560];
        layer2[1][55:48] = buffer_data_4[1575:1568];
        layer3[1][7:0] = buffer_data_3[1527:1520];
        layer3[1][15:8] = buffer_data_3[1535:1528];
        layer3[1][23:16] = buffer_data_3[1543:1536];
        layer3[1][31:24] = buffer_data_3[1551:1544];
        layer3[1][39:32] = buffer_data_3[1559:1552];
        layer3[1][47:40] = buffer_data_3[1567:1560];
        layer3[1][55:48] = buffer_data_3[1575:1568];
        layer4[1][7:0] = buffer_data_2[1527:1520];
        layer4[1][15:8] = buffer_data_2[1535:1528];
        layer4[1][23:16] = buffer_data_2[1543:1536];
        layer4[1][31:24] = buffer_data_2[1551:1544];
        layer4[1][39:32] = buffer_data_2[1559:1552];
        layer4[1][47:40] = buffer_data_2[1567:1560];
        layer4[1][55:48] = buffer_data_2[1575:1568];
        layer5[1][7:0] = buffer_data_1[1527:1520];
        layer5[1][15:8] = buffer_data_1[1535:1528];
        layer5[1][23:16] = buffer_data_1[1543:1536];
        layer5[1][31:24] = buffer_data_1[1551:1544];
        layer5[1][39:32] = buffer_data_1[1559:1552];
        layer5[1][47:40] = buffer_data_1[1567:1560];
        layer5[1][55:48] = buffer_data_1[1575:1568];
        layer6[1][7:0] = buffer_data_0[1527:1520];
        layer6[1][15:8] = buffer_data_0[1535:1528];
        layer6[1][23:16] = buffer_data_0[1543:1536];
        layer6[1][31:24] = buffer_data_0[1551:1544];
        layer6[1][39:32] = buffer_data_0[1559:1552];
        layer6[1][47:40] = buffer_data_0[1567:1560];
        layer6[1][55:48] = buffer_data_0[1575:1568];
        layer0[2][7:0] = buffer_data_6[1535:1528];
        layer0[2][15:8] = buffer_data_6[1543:1536];
        layer0[2][23:16] = buffer_data_6[1551:1544];
        layer0[2][31:24] = buffer_data_6[1559:1552];
        layer0[2][39:32] = buffer_data_6[1567:1560];
        layer0[2][47:40] = buffer_data_6[1575:1568];
        layer0[2][55:48] = buffer_data_6[1583:1576];
        layer1[2][7:0] = buffer_data_5[1535:1528];
        layer1[2][15:8] = buffer_data_5[1543:1536];
        layer1[2][23:16] = buffer_data_5[1551:1544];
        layer1[2][31:24] = buffer_data_5[1559:1552];
        layer1[2][39:32] = buffer_data_5[1567:1560];
        layer1[2][47:40] = buffer_data_5[1575:1568];
        layer1[2][55:48] = buffer_data_5[1583:1576];
        layer2[2][7:0] = buffer_data_4[1535:1528];
        layer2[2][15:8] = buffer_data_4[1543:1536];
        layer2[2][23:16] = buffer_data_4[1551:1544];
        layer2[2][31:24] = buffer_data_4[1559:1552];
        layer2[2][39:32] = buffer_data_4[1567:1560];
        layer2[2][47:40] = buffer_data_4[1575:1568];
        layer2[2][55:48] = buffer_data_4[1583:1576];
        layer3[2][7:0] = buffer_data_3[1535:1528];
        layer3[2][15:8] = buffer_data_3[1543:1536];
        layer3[2][23:16] = buffer_data_3[1551:1544];
        layer3[2][31:24] = buffer_data_3[1559:1552];
        layer3[2][39:32] = buffer_data_3[1567:1560];
        layer3[2][47:40] = buffer_data_3[1575:1568];
        layer3[2][55:48] = buffer_data_3[1583:1576];
        layer4[2][7:0] = buffer_data_2[1535:1528];
        layer4[2][15:8] = buffer_data_2[1543:1536];
        layer4[2][23:16] = buffer_data_2[1551:1544];
        layer4[2][31:24] = buffer_data_2[1559:1552];
        layer4[2][39:32] = buffer_data_2[1567:1560];
        layer4[2][47:40] = buffer_data_2[1575:1568];
        layer4[2][55:48] = buffer_data_2[1583:1576];
        layer5[2][7:0] = buffer_data_1[1535:1528];
        layer5[2][15:8] = buffer_data_1[1543:1536];
        layer5[2][23:16] = buffer_data_1[1551:1544];
        layer5[2][31:24] = buffer_data_1[1559:1552];
        layer5[2][39:32] = buffer_data_1[1567:1560];
        layer5[2][47:40] = buffer_data_1[1575:1568];
        layer5[2][55:48] = buffer_data_1[1583:1576];
        layer6[2][7:0] = buffer_data_0[1535:1528];
        layer6[2][15:8] = buffer_data_0[1543:1536];
        layer6[2][23:16] = buffer_data_0[1551:1544];
        layer6[2][31:24] = buffer_data_0[1559:1552];
        layer6[2][39:32] = buffer_data_0[1567:1560];
        layer6[2][47:40] = buffer_data_0[1575:1568];
        layer6[2][55:48] = buffer_data_0[1583:1576];
        layer0[3][7:0] = buffer_data_6[1543:1536];
        layer0[3][15:8] = buffer_data_6[1551:1544];
        layer0[3][23:16] = buffer_data_6[1559:1552];
        layer0[3][31:24] = buffer_data_6[1567:1560];
        layer0[3][39:32] = buffer_data_6[1575:1568];
        layer0[3][47:40] = buffer_data_6[1583:1576];
        layer0[3][55:48] = buffer_data_6[1591:1584];
        layer1[3][7:0] = buffer_data_5[1543:1536];
        layer1[3][15:8] = buffer_data_5[1551:1544];
        layer1[3][23:16] = buffer_data_5[1559:1552];
        layer1[3][31:24] = buffer_data_5[1567:1560];
        layer1[3][39:32] = buffer_data_5[1575:1568];
        layer1[3][47:40] = buffer_data_5[1583:1576];
        layer1[3][55:48] = buffer_data_5[1591:1584];
        layer2[3][7:0] = buffer_data_4[1543:1536];
        layer2[3][15:8] = buffer_data_4[1551:1544];
        layer2[3][23:16] = buffer_data_4[1559:1552];
        layer2[3][31:24] = buffer_data_4[1567:1560];
        layer2[3][39:32] = buffer_data_4[1575:1568];
        layer2[3][47:40] = buffer_data_4[1583:1576];
        layer2[3][55:48] = buffer_data_4[1591:1584];
        layer3[3][7:0] = buffer_data_3[1543:1536];
        layer3[3][15:8] = buffer_data_3[1551:1544];
        layer3[3][23:16] = buffer_data_3[1559:1552];
        layer3[3][31:24] = buffer_data_3[1567:1560];
        layer3[3][39:32] = buffer_data_3[1575:1568];
        layer3[3][47:40] = buffer_data_3[1583:1576];
        layer3[3][55:48] = buffer_data_3[1591:1584];
        layer4[3][7:0] = buffer_data_2[1543:1536];
        layer4[3][15:8] = buffer_data_2[1551:1544];
        layer4[3][23:16] = buffer_data_2[1559:1552];
        layer4[3][31:24] = buffer_data_2[1567:1560];
        layer4[3][39:32] = buffer_data_2[1575:1568];
        layer4[3][47:40] = buffer_data_2[1583:1576];
        layer4[3][55:48] = buffer_data_2[1591:1584];
        layer5[3][7:0] = buffer_data_1[1543:1536];
        layer5[3][15:8] = buffer_data_1[1551:1544];
        layer5[3][23:16] = buffer_data_1[1559:1552];
        layer5[3][31:24] = buffer_data_1[1567:1560];
        layer5[3][39:32] = buffer_data_1[1575:1568];
        layer5[3][47:40] = buffer_data_1[1583:1576];
        layer5[3][55:48] = buffer_data_1[1591:1584];
        layer6[3][7:0] = buffer_data_0[1543:1536];
        layer6[3][15:8] = buffer_data_0[1551:1544];
        layer6[3][23:16] = buffer_data_0[1559:1552];
        layer6[3][31:24] = buffer_data_0[1567:1560];
        layer6[3][39:32] = buffer_data_0[1575:1568];
        layer6[3][47:40] = buffer_data_0[1583:1576];
        layer6[3][55:48] = buffer_data_0[1591:1584];
        layer0[4][7:0] = buffer_data_6[1551:1544];
        layer0[4][15:8] = buffer_data_6[1559:1552];
        layer0[4][23:16] = buffer_data_6[1567:1560];
        layer0[4][31:24] = buffer_data_6[1575:1568];
        layer0[4][39:32] = buffer_data_6[1583:1576];
        layer0[4][47:40] = buffer_data_6[1591:1584];
        layer0[4][55:48] = buffer_data_6[1599:1592];
        layer1[4][7:0] = buffer_data_5[1551:1544];
        layer1[4][15:8] = buffer_data_5[1559:1552];
        layer1[4][23:16] = buffer_data_5[1567:1560];
        layer1[4][31:24] = buffer_data_5[1575:1568];
        layer1[4][39:32] = buffer_data_5[1583:1576];
        layer1[4][47:40] = buffer_data_5[1591:1584];
        layer1[4][55:48] = buffer_data_5[1599:1592];
        layer2[4][7:0] = buffer_data_4[1551:1544];
        layer2[4][15:8] = buffer_data_4[1559:1552];
        layer2[4][23:16] = buffer_data_4[1567:1560];
        layer2[4][31:24] = buffer_data_4[1575:1568];
        layer2[4][39:32] = buffer_data_4[1583:1576];
        layer2[4][47:40] = buffer_data_4[1591:1584];
        layer2[4][55:48] = buffer_data_4[1599:1592];
        layer3[4][7:0] = buffer_data_3[1551:1544];
        layer3[4][15:8] = buffer_data_3[1559:1552];
        layer3[4][23:16] = buffer_data_3[1567:1560];
        layer3[4][31:24] = buffer_data_3[1575:1568];
        layer3[4][39:32] = buffer_data_3[1583:1576];
        layer3[4][47:40] = buffer_data_3[1591:1584];
        layer3[4][55:48] = buffer_data_3[1599:1592];
        layer4[4][7:0] = buffer_data_2[1551:1544];
        layer4[4][15:8] = buffer_data_2[1559:1552];
        layer4[4][23:16] = buffer_data_2[1567:1560];
        layer4[4][31:24] = buffer_data_2[1575:1568];
        layer4[4][39:32] = buffer_data_2[1583:1576];
        layer4[4][47:40] = buffer_data_2[1591:1584];
        layer4[4][55:48] = buffer_data_2[1599:1592];
        layer5[4][7:0] = buffer_data_1[1551:1544];
        layer5[4][15:8] = buffer_data_1[1559:1552];
        layer5[4][23:16] = buffer_data_1[1567:1560];
        layer5[4][31:24] = buffer_data_1[1575:1568];
        layer5[4][39:32] = buffer_data_1[1583:1576];
        layer5[4][47:40] = buffer_data_1[1591:1584];
        layer5[4][55:48] = buffer_data_1[1599:1592];
        layer6[4][7:0] = buffer_data_0[1551:1544];
        layer6[4][15:8] = buffer_data_0[1559:1552];
        layer6[4][23:16] = buffer_data_0[1567:1560];
        layer6[4][31:24] = buffer_data_0[1575:1568];
        layer6[4][39:32] = buffer_data_0[1583:1576];
        layer6[4][47:40] = buffer_data_0[1591:1584];
        layer6[4][55:48] = buffer_data_0[1599:1592];
        layer0[5][7:0] = buffer_data_6[1559:1552];
        layer0[5][15:8] = buffer_data_6[1567:1560];
        layer0[5][23:16] = buffer_data_6[1575:1568];
        layer0[5][31:24] = buffer_data_6[1583:1576];
        layer0[5][39:32] = buffer_data_6[1591:1584];
        layer0[5][47:40] = buffer_data_6[1599:1592];
        layer0[5][55:48] = buffer_data_6[1607:1600];
        layer1[5][7:0] = buffer_data_5[1559:1552];
        layer1[5][15:8] = buffer_data_5[1567:1560];
        layer1[5][23:16] = buffer_data_5[1575:1568];
        layer1[5][31:24] = buffer_data_5[1583:1576];
        layer1[5][39:32] = buffer_data_5[1591:1584];
        layer1[5][47:40] = buffer_data_5[1599:1592];
        layer1[5][55:48] = buffer_data_5[1607:1600];
        layer2[5][7:0] = buffer_data_4[1559:1552];
        layer2[5][15:8] = buffer_data_4[1567:1560];
        layer2[5][23:16] = buffer_data_4[1575:1568];
        layer2[5][31:24] = buffer_data_4[1583:1576];
        layer2[5][39:32] = buffer_data_4[1591:1584];
        layer2[5][47:40] = buffer_data_4[1599:1592];
        layer2[5][55:48] = buffer_data_4[1607:1600];
        layer3[5][7:0] = buffer_data_3[1559:1552];
        layer3[5][15:8] = buffer_data_3[1567:1560];
        layer3[5][23:16] = buffer_data_3[1575:1568];
        layer3[5][31:24] = buffer_data_3[1583:1576];
        layer3[5][39:32] = buffer_data_3[1591:1584];
        layer3[5][47:40] = buffer_data_3[1599:1592];
        layer3[5][55:48] = buffer_data_3[1607:1600];
        layer4[5][7:0] = buffer_data_2[1559:1552];
        layer4[5][15:8] = buffer_data_2[1567:1560];
        layer4[5][23:16] = buffer_data_2[1575:1568];
        layer4[5][31:24] = buffer_data_2[1583:1576];
        layer4[5][39:32] = buffer_data_2[1591:1584];
        layer4[5][47:40] = buffer_data_2[1599:1592];
        layer4[5][55:48] = buffer_data_2[1607:1600];
        layer5[5][7:0] = buffer_data_1[1559:1552];
        layer5[5][15:8] = buffer_data_1[1567:1560];
        layer5[5][23:16] = buffer_data_1[1575:1568];
        layer5[5][31:24] = buffer_data_1[1583:1576];
        layer5[5][39:32] = buffer_data_1[1591:1584];
        layer5[5][47:40] = buffer_data_1[1599:1592];
        layer5[5][55:48] = buffer_data_1[1607:1600];
        layer6[5][7:0] = buffer_data_0[1559:1552];
        layer6[5][15:8] = buffer_data_0[1567:1560];
        layer6[5][23:16] = buffer_data_0[1575:1568];
        layer6[5][31:24] = buffer_data_0[1583:1576];
        layer6[5][39:32] = buffer_data_0[1591:1584];
        layer6[5][47:40] = buffer_data_0[1599:1592];
        layer6[5][55:48] = buffer_data_0[1607:1600];
        layer0[6][7:0] = buffer_data_6[1567:1560];
        layer0[6][15:8] = buffer_data_6[1575:1568];
        layer0[6][23:16] = buffer_data_6[1583:1576];
        layer0[6][31:24] = buffer_data_6[1591:1584];
        layer0[6][39:32] = buffer_data_6[1599:1592];
        layer0[6][47:40] = buffer_data_6[1607:1600];
        layer0[6][55:48] = buffer_data_6[1615:1608];
        layer1[6][7:0] = buffer_data_5[1567:1560];
        layer1[6][15:8] = buffer_data_5[1575:1568];
        layer1[6][23:16] = buffer_data_5[1583:1576];
        layer1[6][31:24] = buffer_data_5[1591:1584];
        layer1[6][39:32] = buffer_data_5[1599:1592];
        layer1[6][47:40] = buffer_data_5[1607:1600];
        layer1[6][55:48] = buffer_data_5[1615:1608];
        layer2[6][7:0] = buffer_data_4[1567:1560];
        layer2[6][15:8] = buffer_data_4[1575:1568];
        layer2[6][23:16] = buffer_data_4[1583:1576];
        layer2[6][31:24] = buffer_data_4[1591:1584];
        layer2[6][39:32] = buffer_data_4[1599:1592];
        layer2[6][47:40] = buffer_data_4[1607:1600];
        layer2[6][55:48] = buffer_data_4[1615:1608];
        layer3[6][7:0] = buffer_data_3[1567:1560];
        layer3[6][15:8] = buffer_data_3[1575:1568];
        layer3[6][23:16] = buffer_data_3[1583:1576];
        layer3[6][31:24] = buffer_data_3[1591:1584];
        layer3[6][39:32] = buffer_data_3[1599:1592];
        layer3[6][47:40] = buffer_data_3[1607:1600];
        layer3[6][55:48] = buffer_data_3[1615:1608];
        layer4[6][7:0] = buffer_data_2[1567:1560];
        layer4[6][15:8] = buffer_data_2[1575:1568];
        layer4[6][23:16] = buffer_data_2[1583:1576];
        layer4[6][31:24] = buffer_data_2[1591:1584];
        layer4[6][39:32] = buffer_data_2[1599:1592];
        layer4[6][47:40] = buffer_data_2[1607:1600];
        layer4[6][55:48] = buffer_data_2[1615:1608];
        layer5[6][7:0] = buffer_data_1[1567:1560];
        layer5[6][15:8] = buffer_data_1[1575:1568];
        layer5[6][23:16] = buffer_data_1[1583:1576];
        layer5[6][31:24] = buffer_data_1[1591:1584];
        layer5[6][39:32] = buffer_data_1[1599:1592];
        layer5[6][47:40] = buffer_data_1[1607:1600];
        layer5[6][55:48] = buffer_data_1[1615:1608];
        layer6[6][7:0] = buffer_data_0[1567:1560];
        layer6[6][15:8] = buffer_data_0[1575:1568];
        layer6[6][23:16] = buffer_data_0[1583:1576];
        layer6[6][31:24] = buffer_data_0[1591:1584];
        layer6[6][39:32] = buffer_data_0[1599:1592];
        layer6[6][47:40] = buffer_data_0[1607:1600];
        layer6[6][55:48] = buffer_data_0[1615:1608];
        layer0[7][7:0] = buffer_data_6[1575:1568];
        layer0[7][15:8] = buffer_data_6[1583:1576];
        layer0[7][23:16] = buffer_data_6[1591:1584];
        layer0[7][31:24] = buffer_data_6[1599:1592];
        layer0[7][39:32] = buffer_data_6[1607:1600];
        layer0[7][47:40] = buffer_data_6[1615:1608];
        layer0[7][55:48] = buffer_data_6[1623:1616];
        layer1[7][7:0] = buffer_data_5[1575:1568];
        layer1[7][15:8] = buffer_data_5[1583:1576];
        layer1[7][23:16] = buffer_data_5[1591:1584];
        layer1[7][31:24] = buffer_data_5[1599:1592];
        layer1[7][39:32] = buffer_data_5[1607:1600];
        layer1[7][47:40] = buffer_data_5[1615:1608];
        layer1[7][55:48] = buffer_data_5[1623:1616];
        layer2[7][7:0] = buffer_data_4[1575:1568];
        layer2[7][15:8] = buffer_data_4[1583:1576];
        layer2[7][23:16] = buffer_data_4[1591:1584];
        layer2[7][31:24] = buffer_data_4[1599:1592];
        layer2[7][39:32] = buffer_data_4[1607:1600];
        layer2[7][47:40] = buffer_data_4[1615:1608];
        layer2[7][55:48] = buffer_data_4[1623:1616];
        layer3[7][7:0] = buffer_data_3[1575:1568];
        layer3[7][15:8] = buffer_data_3[1583:1576];
        layer3[7][23:16] = buffer_data_3[1591:1584];
        layer3[7][31:24] = buffer_data_3[1599:1592];
        layer3[7][39:32] = buffer_data_3[1607:1600];
        layer3[7][47:40] = buffer_data_3[1615:1608];
        layer3[7][55:48] = buffer_data_3[1623:1616];
        layer4[7][7:0] = buffer_data_2[1575:1568];
        layer4[7][15:8] = buffer_data_2[1583:1576];
        layer4[7][23:16] = buffer_data_2[1591:1584];
        layer4[7][31:24] = buffer_data_2[1599:1592];
        layer4[7][39:32] = buffer_data_2[1607:1600];
        layer4[7][47:40] = buffer_data_2[1615:1608];
        layer4[7][55:48] = buffer_data_2[1623:1616];
        layer5[7][7:0] = buffer_data_1[1575:1568];
        layer5[7][15:8] = buffer_data_1[1583:1576];
        layer5[7][23:16] = buffer_data_1[1591:1584];
        layer5[7][31:24] = buffer_data_1[1599:1592];
        layer5[7][39:32] = buffer_data_1[1607:1600];
        layer5[7][47:40] = buffer_data_1[1615:1608];
        layer5[7][55:48] = buffer_data_1[1623:1616];
        layer6[7][7:0] = buffer_data_0[1575:1568];
        layer6[7][15:8] = buffer_data_0[1583:1576];
        layer6[7][23:16] = buffer_data_0[1591:1584];
        layer6[7][31:24] = buffer_data_0[1599:1592];
        layer6[7][39:32] = buffer_data_0[1607:1600];
        layer6[7][47:40] = buffer_data_0[1615:1608];
        layer6[7][55:48] = buffer_data_0[1623:1616];
        layer0[8][7:0] = buffer_data_6[1583:1576];
        layer0[8][15:8] = buffer_data_6[1591:1584];
        layer0[8][23:16] = buffer_data_6[1599:1592];
        layer0[8][31:24] = buffer_data_6[1607:1600];
        layer0[8][39:32] = buffer_data_6[1615:1608];
        layer0[8][47:40] = buffer_data_6[1623:1616];
        layer0[8][55:48] = buffer_data_6[1631:1624];
        layer1[8][7:0] = buffer_data_5[1583:1576];
        layer1[8][15:8] = buffer_data_5[1591:1584];
        layer1[8][23:16] = buffer_data_5[1599:1592];
        layer1[8][31:24] = buffer_data_5[1607:1600];
        layer1[8][39:32] = buffer_data_5[1615:1608];
        layer1[8][47:40] = buffer_data_5[1623:1616];
        layer1[8][55:48] = buffer_data_5[1631:1624];
        layer2[8][7:0] = buffer_data_4[1583:1576];
        layer2[8][15:8] = buffer_data_4[1591:1584];
        layer2[8][23:16] = buffer_data_4[1599:1592];
        layer2[8][31:24] = buffer_data_4[1607:1600];
        layer2[8][39:32] = buffer_data_4[1615:1608];
        layer2[8][47:40] = buffer_data_4[1623:1616];
        layer2[8][55:48] = buffer_data_4[1631:1624];
        layer3[8][7:0] = buffer_data_3[1583:1576];
        layer3[8][15:8] = buffer_data_3[1591:1584];
        layer3[8][23:16] = buffer_data_3[1599:1592];
        layer3[8][31:24] = buffer_data_3[1607:1600];
        layer3[8][39:32] = buffer_data_3[1615:1608];
        layer3[8][47:40] = buffer_data_3[1623:1616];
        layer3[8][55:48] = buffer_data_3[1631:1624];
        layer4[8][7:0] = buffer_data_2[1583:1576];
        layer4[8][15:8] = buffer_data_2[1591:1584];
        layer4[8][23:16] = buffer_data_2[1599:1592];
        layer4[8][31:24] = buffer_data_2[1607:1600];
        layer4[8][39:32] = buffer_data_2[1615:1608];
        layer4[8][47:40] = buffer_data_2[1623:1616];
        layer4[8][55:48] = buffer_data_2[1631:1624];
        layer5[8][7:0] = buffer_data_1[1583:1576];
        layer5[8][15:8] = buffer_data_1[1591:1584];
        layer5[8][23:16] = buffer_data_1[1599:1592];
        layer5[8][31:24] = buffer_data_1[1607:1600];
        layer5[8][39:32] = buffer_data_1[1615:1608];
        layer5[8][47:40] = buffer_data_1[1623:1616];
        layer5[8][55:48] = buffer_data_1[1631:1624];
        layer6[8][7:0] = buffer_data_0[1583:1576];
        layer6[8][15:8] = buffer_data_0[1591:1584];
        layer6[8][23:16] = buffer_data_0[1599:1592];
        layer6[8][31:24] = buffer_data_0[1607:1600];
        layer6[8][39:32] = buffer_data_0[1615:1608];
        layer6[8][47:40] = buffer_data_0[1623:1616];
        layer6[8][55:48] = buffer_data_0[1631:1624];
        layer0[9][7:0] = buffer_data_6[1591:1584];
        layer0[9][15:8] = buffer_data_6[1599:1592];
        layer0[9][23:16] = buffer_data_6[1607:1600];
        layer0[9][31:24] = buffer_data_6[1615:1608];
        layer0[9][39:32] = buffer_data_6[1623:1616];
        layer0[9][47:40] = buffer_data_6[1631:1624];
        layer0[9][55:48] = buffer_data_6[1639:1632];
        layer1[9][7:0] = buffer_data_5[1591:1584];
        layer1[9][15:8] = buffer_data_5[1599:1592];
        layer1[9][23:16] = buffer_data_5[1607:1600];
        layer1[9][31:24] = buffer_data_5[1615:1608];
        layer1[9][39:32] = buffer_data_5[1623:1616];
        layer1[9][47:40] = buffer_data_5[1631:1624];
        layer1[9][55:48] = buffer_data_5[1639:1632];
        layer2[9][7:0] = buffer_data_4[1591:1584];
        layer2[9][15:8] = buffer_data_4[1599:1592];
        layer2[9][23:16] = buffer_data_4[1607:1600];
        layer2[9][31:24] = buffer_data_4[1615:1608];
        layer2[9][39:32] = buffer_data_4[1623:1616];
        layer2[9][47:40] = buffer_data_4[1631:1624];
        layer2[9][55:48] = buffer_data_4[1639:1632];
        layer3[9][7:0] = buffer_data_3[1591:1584];
        layer3[9][15:8] = buffer_data_3[1599:1592];
        layer3[9][23:16] = buffer_data_3[1607:1600];
        layer3[9][31:24] = buffer_data_3[1615:1608];
        layer3[9][39:32] = buffer_data_3[1623:1616];
        layer3[9][47:40] = buffer_data_3[1631:1624];
        layer3[9][55:48] = buffer_data_3[1639:1632];
        layer4[9][7:0] = buffer_data_2[1591:1584];
        layer4[9][15:8] = buffer_data_2[1599:1592];
        layer4[9][23:16] = buffer_data_2[1607:1600];
        layer4[9][31:24] = buffer_data_2[1615:1608];
        layer4[9][39:32] = buffer_data_2[1623:1616];
        layer4[9][47:40] = buffer_data_2[1631:1624];
        layer4[9][55:48] = buffer_data_2[1639:1632];
        layer5[9][7:0] = buffer_data_1[1591:1584];
        layer5[9][15:8] = buffer_data_1[1599:1592];
        layer5[9][23:16] = buffer_data_1[1607:1600];
        layer5[9][31:24] = buffer_data_1[1615:1608];
        layer5[9][39:32] = buffer_data_1[1623:1616];
        layer5[9][47:40] = buffer_data_1[1631:1624];
        layer5[9][55:48] = buffer_data_1[1639:1632];
        layer6[9][7:0] = buffer_data_0[1591:1584];
        layer6[9][15:8] = buffer_data_0[1599:1592];
        layer6[9][23:16] = buffer_data_0[1607:1600];
        layer6[9][31:24] = buffer_data_0[1615:1608];
        layer6[9][39:32] = buffer_data_0[1623:1616];
        layer6[9][47:40] = buffer_data_0[1631:1624];
        layer6[9][55:48] = buffer_data_0[1639:1632];
        layer0[10][7:0] = buffer_data_6[1599:1592];
        layer0[10][15:8] = buffer_data_6[1607:1600];
        layer0[10][23:16] = buffer_data_6[1615:1608];
        layer0[10][31:24] = buffer_data_6[1623:1616];
        layer0[10][39:32] = buffer_data_6[1631:1624];
        layer0[10][47:40] = buffer_data_6[1639:1632];
        layer0[10][55:48] = buffer_data_6[1647:1640];
        layer1[10][7:0] = buffer_data_5[1599:1592];
        layer1[10][15:8] = buffer_data_5[1607:1600];
        layer1[10][23:16] = buffer_data_5[1615:1608];
        layer1[10][31:24] = buffer_data_5[1623:1616];
        layer1[10][39:32] = buffer_data_5[1631:1624];
        layer1[10][47:40] = buffer_data_5[1639:1632];
        layer1[10][55:48] = buffer_data_5[1647:1640];
        layer2[10][7:0] = buffer_data_4[1599:1592];
        layer2[10][15:8] = buffer_data_4[1607:1600];
        layer2[10][23:16] = buffer_data_4[1615:1608];
        layer2[10][31:24] = buffer_data_4[1623:1616];
        layer2[10][39:32] = buffer_data_4[1631:1624];
        layer2[10][47:40] = buffer_data_4[1639:1632];
        layer2[10][55:48] = buffer_data_4[1647:1640];
        layer3[10][7:0] = buffer_data_3[1599:1592];
        layer3[10][15:8] = buffer_data_3[1607:1600];
        layer3[10][23:16] = buffer_data_3[1615:1608];
        layer3[10][31:24] = buffer_data_3[1623:1616];
        layer3[10][39:32] = buffer_data_3[1631:1624];
        layer3[10][47:40] = buffer_data_3[1639:1632];
        layer3[10][55:48] = buffer_data_3[1647:1640];
        layer4[10][7:0] = buffer_data_2[1599:1592];
        layer4[10][15:8] = buffer_data_2[1607:1600];
        layer4[10][23:16] = buffer_data_2[1615:1608];
        layer4[10][31:24] = buffer_data_2[1623:1616];
        layer4[10][39:32] = buffer_data_2[1631:1624];
        layer4[10][47:40] = buffer_data_2[1639:1632];
        layer4[10][55:48] = buffer_data_2[1647:1640];
        layer5[10][7:0] = buffer_data_1[1599:1592];
        layer5[10][15:8] = buffer_data_1[1607:1600];
        layer5[10][23:16] = buffer_data_1[1615:1608];
        layer5[10][31:24] = buffer_data_1[1623:1616];
        layer5[10][39:32] = buffer_data_1[1631:1624];
        layer5[10][47:40] = buffer_data_1[1639:1632];
        layer5[10][55:48] = buffer_data_1[1647:1640];
        layer6[10][7:0] = buffer_data_0[1599:1592];
        layer6[10][15:8] = buffer_data_0[1607:1600];
        layer6[10][23:16] = buffer_data_0[1615:1608];
        layer6[10][31:24] = buffer_data_0[1623:1616];
        layer6[10][39:32] = buffer_data_0[1631:1624];
        layer6[10][47:40] = buffer_data_0[1639:1632];
        layer6[10][55:48] = buffer_data_0[1647:1640];
        layer0[11][7:0] = buffer_data_6[1607:1600];
        layer0[11][15:8] = buffer_data_6[1615:1608];
        layer0[11][23:16] = buffer_data_6[1623:1616];
        layer0[11][31:24] = buffer_data_6[1631:1624];
        layer0[11][39:32] = buffer_data_6[1639:1632];
        layer0[11][47:40] = buffer_data_6[1647:1640];
        layer0[11][55:48] = buffer_data_6[1655:1648];
        layer1[11][7:0] = buffer_data_5[1607:1600];
        layer1[11][15:8] = buffer_data_5[1615:1608];
        layer1[11][23:16] = buffer_data_5[1623:1616];
        layer1[11][31:24] = buffer_data_5[1631:1624];
        layer1[11][39:32] = buffer_data_5[1639:1632];
        layer1[11][47:40] = buffer_data_5[1647:1640];
        layer1[11][55:48] = buffer_data_5[1655:1648];
        layer2[11][7:0] = buffer_data_4[1607:1600];
        layer2[11][15:8] = buffer_data_4[1615:1608];
        layer2[11][23:16] = buffer_data_4[1623:1616];
        layer2[11][31:24] = buffer_data_4[1631:1624];
        layer2[11][39:32] = buffer_data_4[1639:1632];
        layer2[11][47:40] = buffer_data_4[1647:1640];
        layer2[11][55:48] = buffer_data_4[1655:1648];
        layer3[11][7:0] = buffer_data_3[1607:1600];
        layer3[11][15:8] = buffer_data_3[1615:1608];
        layer3[11][23:16] = buffer_data_3[1623:1616];
        layer3[11][31:24] = buffer_data_3[1631:1624];
        layer3[11][39:32] = buffer_data_3[1639:1632];
        layer3[11][47:40] = buffer_data_3[1647:1640];
        layer3[11][55:48] = buffer_data_3[1655:1648];
        layer4[11][7:0] = buffer_data_2[1607:1600];
        layer4[11][15:8] = buffer_data_2[1615:1608];
        layer4[11][23:16] = buffer_data_2[1623:1616];
        layer4[11][31:24] = buffer_data_2[1631:1624];
        layer4[11][39:32] = buffer_data_2[1639:1632];
        layer4[11][47:40] = buffer_data_2[1647:1640];
        layer4[11][55:48] = buffer_data_2[1655:1648];
        layer5[11][7:0] = buffer_data_1[1607:1600];
        layer5[11][15:8] = buffer_data_1[1615:1608];
        layer5[11][23:16] = buffer_data_1[1623:1616];
        layer5[11][31:24] = buffer_data_1[1631:1624];
        layer5[11][39:32] = buffer_data_1[1639:1632];
        layer5[11][47:40] = buffer_data_1[1647:1640];
        layer5[11][55:48] = buffer_data_1[1655:1648];
        layer6[11][7:0] = buffer_data_0[1607:1600];
        layer6[11][15:8] = buffer_data_0[1615:1608];
        layer6[11][23:16] = buffer_data_0[1623:1616];
        layer6[11][31:24] = buffer_data_0[1631:1624];
        layer6[11][39:32] = buffer_data_0[1639:1632];
        layer6[11][47:40] = buffer_data_0[1647:1640];
        layer6[11][55:48] = buffer_data_0[1655:1648];
        layer0[12][7:0] = buffer_data_6[1615:1608];
        layer0[12][15:8] = buffer_data_6[1623:1616];
        layer0[12][23:16] = buffer_data_6[1631:1624];
        layer0[12][31:24] = buffer_data_6[1639:1632];
        layer0[12][39:32] = buffer_data_6[1647:1640];
        layer0[12][47:40] = buffer_data_6[1655:1648];
        layer0[12][55:48] = buffer_data_6[1663:1656];
        layer1[12][7:0] = buffer_data_5[1615:1608];
        layer1[12][15:8] = buffer_data_5[1623:1616];
        layer1[12][23:16] = buffer_data_5[1631:1624];
        layer1[12][31:24] = buffer_data_5[1639:1632];
        layer1[12][39:32] = buffer_data_5[1647:1640];
        layer1[12][47:40] = buffer_data_5[1655:1648];
        layer1[12][55:48] = buffer_data_5[1663:1656];
        layer2[12][7:0] = buffer_data_4[1615:1608];
        layer2[12][15:8] = buffer_data_4[1623:1616];
        layer2[12][23:16] = buffer_data_4[1631:1624];
        layer2[12][31:24] = buffer_data_4[1639:1632];
        layer2[12][39:32] = buffer_data_4[1647:1640];
        layer2[12][47:40] = buffer_data_4[1655:1648];
        layer2[12][55:48] = buffer_data_4[1663:1656];
        layer3[12][7:0] = buffer_data_3[1615:1608];
        layer3[12][15:8] = buffer_data_3[1623:1616];
        layer3[12][23:16] = buffer_data_3[1631:1624];
        layer3[12][31:24] = buffer_data_3[1639:1632];
        layer3[12][39:32] = buffer_data_3[1647:1640];
        layer3[12][47:40] = buffer_data_3[1655:1648];
        layer3[12][55:48] = buffer_data_3[1663:1656];
        layer4[12][7:0] = buffer_data_2[1615:1608];
        layer4[12][15:8] = buffer_data_2[1623:1616];
        layer4[12][23:16] = buffer_data_2[1631:1624];
        layer4[12][31:24] = buffer_data_2[1639:1632];
        layer4[12][39:32] = buffer_data_2[1647:1640];
        layer4[12][47:40] = buffer_data_2[1655:1648];
        layer4[12][55:48] = buffer_data_2[1663:1656];
        layer5[12][7:0] = buffer_data_1[1615:1608];
        layer5[12][15:8] = buffer_data_1[1623:1616];
        layer5[12][23:16] = buffer_data_1[1631:1624];
        layer5[12][31:24] = buffer_data_1[1639:1632];
        layer5[12][39:32] = buffer_data_1[1647:1640];
        layer5[12][47:40] = buffer_data_1[1655:1648];
        layer5[12][55:48] = buffer_data_1[1663:1656];
        layer6[12][7:0] = buffer_data_0[1615:1608];
        layer6[12][15:8] = buffer_data_0[1623:1616];
        layer6[12][23:16] = buffer_data_0[1631:1624];
        layer6[12][31:24] = buffer_data_0[1639:1632];
        layer6[12][39:32] = buffer_data_0[1647:1640];
        layer6[12][47:40] = buffer_data_0[1655:1648];
        layer6[12][55:48] = buffer_data_0[1663:1656];
        layer0[13][7:0] = buffer_data_6[1623:1616];
        layer0[13][15:8] = buffer_data_6[1631:1624];
        layer0[13][23:16] = buffer_data_6[1639:1632];
        layer0[13][31:24] = buffer_data_6[1647:1640];
        layer0[13][39:32] = buffer_data_6[1655:1648];
        layer0[13][47:40] = buffer_data_6[1663:1656];
        layer0[13][55:48] = buffer_data_6[1671:1664];
        layer1[13][7:0] = buffer_data_5[1623:1616];
        layer1[13][15:8] = buffer_data_5[1631:1624];
        layer1[13][23:16] = buffer_data_5[1639:1632];
        layer1[13][31:24] = buffer_data_5[1647:1640];
        layer1[13][39:32] = buffer_data_5[1655:1648];
        layer1[13][47:40] = buffer_data_5[1663:1656];
        layer1[13][55:48] = buffer_data_5[1671:1664];
        layer2[13][7:0] = buffer_data_4[1623:1616];
        layer2[13][15:8] = buffer_data_4[1631:1624];
        layer2[13][23:16] = buffer_data_4[1639:1632];
        layer2[13][31:24] = buffer_data_4[1647:1640];
        layer2[13][39:32] = buffer_data_4[1655:1648];
        layer2[13][47:40] = buffer_data_4[1663:1656];
        layer2[13][55:48] = buffer_data_4[1671:1664];
        layer3[13][7:0] = buffer_data_3[1623:1616];
        layer3[13][15:8] = buffer_data_3[1631:1624];
        layer3[13][23:16] = buffer_data_3[1639:1632];
        layer3[13][31:24] = buffer_data_3[1647:1640];
        layer3[13][39:32] = buffer_data_3[1655:1648];
        layer3[13][47:40] = buffer_data_3[1663:1656];
        layer3[13][55:48] = buffer_data_3[1671:1664];
        layer4[13][7:0] = buffer_data_2[1623:1616];
        layer4[13][15:8] = buffer_data_2[1631:1624];
        layer4[13][23:16] = buffer_data_2[1639:1632];
        layer4[13][31:24] = buffer_data_2[1647:1640];
        layer4[13][39:32] = buffer_data_2[1655:1648];
        layer4[13][47:40] = buffer_data_2[1663:1656];
        layer4[13][55:48] = buffer_data_2[1671:1664];
        layer5[13][7:0] = buffer_data_1[1623:1616];
        layer5[13][15:8] = buffer_data_1[1631:1624];
        layer5[13][23:16] = buffer_data_1[1639:1632];
        layer5[13][31:24] = buffer_data_1[1647:1640];
        layer5[13][39:32] = buffer_data_1[1655:1648];
        layer5[13][47:40] = buffer_data_1[1663:1656];
        layer5[13][55:48] = buffer_data_1[1671:1664];
        layer6[13][7:0] = buffer_data_0[1623:1616];
        layer6[13][15:8] = buffer_data_0[1631:1624];
        layer6[13][23:16] = buffer_data_0[1639:1632];
        layer6[13][31:24] = buffer_data_0[1647:1640];
        layer6[13][39:32] = buffer_data_0[1655:1648];
        layer6[13][47:40] = buffer_data_0[1663:1656];
        layer6[13][55:48] = buffer_data_0[1671:1664];
        layer0[14][7:0] = buffer_data_6[1631:1624];
        layer0[14][15:8] = buffer_data_6[1639:1632];
        layer0[14][23:16] = buffer_data_6[1647:1640];
        layer0[14][31:24] = buffer_data_6[1655:1648];
        layer0[14][39:32] = buffer_data_6[1663:1656];
        layer0[14][47:40] = buffer_data_6[1671:1664];
        layer0[14][55:48] = buffer_data_6[1679:1672];
        layer1[14][7:0] = buffer_data_5[1631:1624];
        layer1[14][15:8] = buffer_data_5[1639:1632];
        layer1[14][23:16] = buffer_data_5[1647:1640];
        layer1[14][31:24] = buffer_data_5[1655:1648];
        layer1[14][39:32] = buffer_data_5[1663:1656];
        layer1[14][47:40] = buffer_data_5[1671:1664];
        layer1[14][55:48] = buffer_data_5[1679:1672];
        layer2[14][7:0] = buffer_data_4[1631:1624];
        layer2[14][15:8] = buffer_data_4[1639:1632];
        layer2[14][23:16] = buffer_data_4[1647:1640];
        layer2[14][31:24] = buffer_data_4[1655:1648];
        layer2[14][39:32] = buffer_data_4[1663:1656];
        layer2[14][47:40] = buffer_data_4[1671:1664];
        layer2[14][55:48] = buffer_data_4[1679:1672];
        layer3[14][7:0] = buffer_data_3[1631:1624];
        layer3[14][15:8] = buffer_data_3[1639:1632];
        layer3[14][23:16] = buffer_data_3[1647:1640];
        layer3[14][31:24] = buffer_data_3[1655:1648];
        layer3[14][39:32] = buffer_data_3[1663:1656];
        layer3[14][47:40] = buffer_data_3[1671:1664];
        layer3[14][55:48] = buffer_data_3[1679:1672];
        layer4[14][7:0] = buffer_data_2[1631:1624];
        layer4[14][15:8] = buffer_data_2[1639:1632];
        layer4[14][23:16] = buffer_data_2[1647:1640];
        layer4[14][31:24] = buffer_data_2[1655:1648];
        layer4[14][39:32] = buffer_data_2[1663:1656];
        layer4[14][47:40] = buffer_data_2[1671:1664];
        layer4[14][55:48] = buffer_data_2[1679:1672];
        layer5[14][7:0] = buffer_data_1[1631:1624];
        layer5[14][15:8] = buffer_data_1[1639:1632];
        layer5[14][23:16] = buffer_data_1[1647:1640];
        layer5[14][31:24] = buffer_data_1[1655:1648];
        layer5[14][39:32] = buffer_data_1[1663:1656];
        layer5[14][47:40] = buffer_data_1[1671:1664];
        layer5[14][55:48] = buffer_data_1[1679:1672];
        layer6[14][7:0] = buffer_data_0[1631:1624];
        layer6[14][15:8] = buffer_data_0[1639:1632];
        layer6[14][23:16] = buffer_data_0[1647:1640];
        layer6[14][31:24] = buffer_data_0[1655:1648];
        layer6[14][39:32] = buffer_data_0[1663:1656];
        layer6[14][47:40] = buffer_data_0[1671:1664];
        layer6[14][55:48] = buffer_data_0[1679:1672];
        layer0[15][7:0] = buffer_data_6[1639:1632];
        layer0[15][15:8] = buffer_data_6[1647:1640];
        layer0[15][23:16] = buffer_data_6[1655:1648];
        layer0[15][31:24] = buffer_data_6[1663:1656];
        layer0[15][39:32] = buffer_data_6[1671:1664];
        layer0[15][47:40] = buffer_data_6[1679:1672];
        layer0[15][55:48] = buffer_data_6[1687:1680];
        layer1[15][7:0] = buffer_data_5[1639:1632];
        layer1[15][15:8] = buffer_data_5[1647:1640];
        layer1[15][23:16] = buffer_data_5[1655:1648];
        layer1[15][31:24] = buffer_data_5[1663:1656];
        layer1[15][39:32] = buffer_data_5[1671:1664];
        layer1[15][47:40] = buffer_data_5[1679:1672];
        layer1[15][55:48] = buffer_data_5[1687:1680];
        layer2[15][7:0] = buffer_data_4[1639:1632];
        layer2[15][15:8] = buffer_data_4[1647:1640];
        layer2[15][23:16] = buffer_data_4[1655:1648];
        layer2[15][31:24] = buffer_data_4[1663:1656];
        layer2[15][39:32] = buffer_data_4[1671:1664];
        layer2[15][47:40] = buffer_data_4[1679:1672];
        layer2[15][55:48] = buffer_data_4[1687:1680];
        layer3[15][7:0] = buffer_data_3[1639:1632];
        layer3[15][15:8] = buffer_data_3[1647:1640];
        layer3[15][23:16] = buffer_data_3[1655:1648];
        layer3[15][31:24] = buffer_data_3[1663:1656];
        layer3[15][39:32] = buffer_data_3[1671:1664];
        layer3[15][47:40] = buffer_data_3[1679:1672];
        layer3[15][55:48] = buffer_data_3[1687:1680];
        layer4[15][7:0] = buffer_data_2[1639:1632];
        layer4[15][15:8] = buffer_data_2[1647:1640];
        layer4[15][23:16] = buffer_data_2[1655:1648];
        layer4[15][31:24] = buffer_data_2[1663:1656];
        layer4[15][39:32] = buffer_data_2[1671:1664];
        layer4[15][47:40] = buffer_data_2[1679:1672];
        layer4[15][55:48] = buffer_data_2[1687:1680];
        layer5[15][7:0] = buffer_data_1[1639:1632];
        layer5[15][15:8] = buffer_data_1[1647:1640];
        layer5[15][23:16] = buffer_data_1[1655:1648];
        layer5[15][31:24] = buffer_data_1[1663:1656];
        layer5[15][39:32] = buffer_data_1[1671:1664];
        layer5[15][47:40] = buffer_data_1[1679:1672];
        layer5[15][55:48] = buffer_data_1[1687:1680];
        layer6[15][7:0] = buffer_data_0[1639:1632];
        layer6[15][15:8] = buffer_data_0[1647:1640];
        layer6[15][23:16] = buffer_data_0[1655:1648];
        layer6[15][31:24] = buffer_data_0[1663:1656];
        layer6[15][39:32] = buffer_data_0[1671:1664];
        layer6[15][47:40] = buffer_data_0[1679:1672];
        layer6[15][55:48] = buffer_data_0[1687:1680];
        layer0[16][7:0] = buffer_data_6[1647:1640];
        layer0[16][15:8] = buffer_data_6[1655:1648];
        layer0[16][23:16] = buffer_data_6[1663:1656];
        layer0[16][31:24] = buffer_data_6[1671:1664];
        layer0[16][39:32] = buffer_data_6[1679:1672];
        layer0[16][47:40] = buffer_data_6[1687:1680];
        layer0[16][55:48] = buffer_data_6[1695:1688];
        layer1[16][7:0] = buffer_data_5[1647:1640];
        layer1[16][15:8] = buffer_data_5[1655:1648];
        layer1[16][23:16] = buffer_data_5[1663:1656];
        layer1[16][31:24] = buffer_data_5[1671:1664];
        layer1[16][39:32] = buffer_data_5[1679:1672];
        layer1[16][47:40] = buffer_data_5[1687:1680];
        layer1[16][55:48] = buffer_data_5[1695:1688];
        layer2[16][7:0] = buffer_data_4[1647:1640];
        layer2[16][15:8] = buffer_data_4[1655:1648];
        layer2[16][23:16] = buffer_data_4[1663:1656];
        layer2[16][31:24] = buffer_data_4[1671:1664];
        layer2[16][39:32] = buffer_data_4[1679:1672];
        layer2[16][47:40] = buffer_data_4[1687:1680];
        layer2[16][55:48] = buffer_data_4[1695:1688];
        layer3[16][7:0] = buffer_data_3[1647:1640];
        layer3[16][15:8] = buffer_data_3[1655:1648];
        layer3[16][23:16] = buffer_data_3[1663:1656];
        layer3[16][31:24] = buffer_data_3[1671:1664];
        layer3[16][39:32] = buffer_data_3[1679:1672];
        layer3[16][47:40] = buffer_data_3[1687:1680];
        layer3[16][55:48] = buffer_data_3[1695:1688];
        layer4[16][7:0] = buffer_data_2[1647:1640];
        layer4[16][15:8] = buffer_data_2[1655:1648];
        layer4[16][23:16] = buffer_data_2[1663:1656];
        layer4[16][31:24] = buffer_data_2[1671:1664];
        layer4[16][39:32] = buffer_data_2[1679:1672];
        layer4[16][47:40] = buffer_data_2[1687:1680];
        layer4[16][55:48] = buffer_data_2[1695:1688];
        layer5[16][7:0] = buffer_data_1[1647:1640];
        layer5[16][15:8] = buffer_data_1[1655:1648];
        layer5[16][23:16] = buffer_data_1[1663:1656];
        layer5[16][31:24] = buffer_data_1[1671:1664];
        layer5[16][39:32] = buffer_data_1[1679:1672];
        layer5[16][47:40] = buffer_data_1[1687:1680];
        layer5[16][55:48] = buffer_data_1[1695:1688];
        layer6[16][7:0] = buffer_data_0[1647:1640];
        layer6[16][15:8] = buffer_data_0[1655:1648];
        layer6[16][23:16] = buffer_data_0[1663:1656];
        layer6[16][31:24] = buffer_data_0[1671:1664];
        layer6[16][39:32] = buffer_data_0[1679:1672];
        layer6[16][47:40] = buffer_data_0[1687:1680];
        layer6[16][55:48] = buffer_data_0[1695:1688];
        layer0[17][7:0] = buffer_data_6[1655:1648];
        layer0[17][15:8] = buffer_data_6[1663:1656];
        layer0[17][23:16] = buffer_data_6[1671:1664];
        layer0[17][31:24] = buffer_data_6[1679:1672];
        layer0[17][39:32] = buffer_data_6[1687:1680];
        layer0[17][47:40] = buffer_data_6[1695:1688];
        layer0[17][55:48] = buffer_data_6[1703:1696];
        layer1[17][7:0] = buffer_data_5[1655:1648];
        layer1[17][15:8] = buffer_data_5[1663:1656];
        layer1[17][23:16] = buffer_data_5[1671:1664];
        layer1[17][31:24] = buffer_data_5[1679:1672];
        layer1[17][39:32] = buffer_data_5[1687:1680];
        layer1[17][47:40] = buffer_data_5[1695:1688];
        layer1[17][55:48] = buffer_data_5[1703:1696];
        layer2[17][7:0] = buffer_data_4[1655:1648];
        layer2[17][15:8] = buffer_data_4[1663:1656];
        layer2[17][23:16] = buffer_data_4[1671:1664];
        layer2[17][31:24] = buffer_data_4[1679:1672];
        layer2[17][39:32] = buffer_data_4[1687:1680];
        layer2[17][47:40] = buffer_data_4[1695:1688];
        layer2[17][55:48] = buffer_data_4[1703:1696];
        layer3[17][7:0] = buffer_data_3[1655:1648];
        layer3[17][15:8] = buffer_data_3[1663:1656];
        layer3[17][23:16] = buffer_data_3[1671:1664];
        layer3[17][31:24] = buffer_data_3[1679:1672];
        layer3[17][39:32] = buffer_data_3[1687:1680];
        layer3[17][47:40] = buffer_data_3[1695:1688];
        layer3[17][55:48] = buffer_data_3[1703:1696];
        layer4[17][7:0] = buffer_data_2[1655:1648];
        layer4[17][15:8] = buffer_data_2[1663:1656];
        layer4[17][23:16] = buffer_data_2[1671:1664];
        layer4[17][31:24] = buffer_data_2[1679:1672];
        layer4[17][39:32] = buffer_data_2[1687:1680];
        layer4[17][47:40] = buffer_data_2[1695:1688];
        layer4[17][55:48] = buffer_data_2[1703:1696];
        layer5[17][7:0] = buffer_data_1[1655:1648];
        layer5[17][15:8] = buffer_data_1[1663:1656];
        layer5[17][23:16] = buffer_data_1[1671:1664];
        layer5[17][31:24] = buffer_data_1[1679:1672];
        layer5[17][39:32] = buffer_data_1[1687:1680];
        layer5[17][47:40] = buffer_data_1[1695:1688];
        layer5[17][55:48] = buffer_data_1[1703:1696];
        layer6[17][7:0] = buffer_data_0[1655:1648];
        layer6[17][15:8] = buffer_data_0[1663:1656];
        layer6[17][23:16] = buffer_data_0[1671:1664];
        layer6[17][31:24] = buffer_data_0[1679:1672];
        layer6[17][39:32] = buffer_data_0[1687:1680];
        layer6[17][47:40] = buffer_data_0[1695:1688];
        layer6[17][55:48] = buffer_data_0[1703:1696];
        layer0[18][7:0] = buffer_data_6[1663:1656];
        layer0[18][15:8] = buffer_data_6[1671:1664];
        layer0[18][23:16] = buffer_data_6[1679:1672];
        layer0[18][31:24] = buffer_data_6[1687:1680];
        layer0[18][39:32] = buffer_data_6[1695:1688];
        layer0[18][47:40] = buffer_data_6[1703:1696];
        layer0[18][55:48] = buffer_data_6[1711:1704];
        layer1[18][7:0] = buffer_data_5[1663:1656];
        layer1[18][15:8] = buffer_data_5[1671:1664];
        layer1[18][23:16] = buffer_data_5[1679:1672];
        layer1[18][31:24] = buffer_data_5[1687:1680];
        layer1[18][39:32] = buffer_data_5[1695:1688];
        layer1[18][47:40] = buffer_data_5[1703:1696];
        layer1[18][55:48] = buffer_data_5[1711:1704];
        layer2[18][7:0] = buffer_data_4[1663:1656];
        layer2[18][15:8] = buffer_data_4[1671:1664];
        layer2[18][23:16] = buffer_data_4[1679:1672];
        layer2[18][31:24] = buffer_data_4[1687:1680];
        layer2[18][39:32] = buffer_data_4[1695:1688];
        layer2[18][47:40] = buffer_data_4[1703:1696];
        layer2[18][55:48] = buffer_data_4[1711:1704];
        layer3[18][7:0] = buffer_data_3[1663:1656];
        layer3[18][15:8] = buffer_data_3[1671:1664];
        layer3[18][23:16] = buffer_data_3[1679:1672];
        layer3[18][31:24] = buffer_data_3[1687:1680];
        layer3[18][39:32] = buffer_data_3[1695:1688];
        layer3[18][47:40] = buffer_data_3[1703:1696];
        layer3[18][55:48] = buffer_data_3[1711:1704];
        layer4[18][7:0] = buffer_data_2[1663:1656];
        layer4[18][15:8] = buffer_data_2[1671:1664];
        layer4[18][23:16] = buffer_data_2[1679:1672];
        layer4[18][31:24] = buffer_data_2[1687:1680];
        layer4[18][39:32] = buffer_data_2[1695:1688];
        layer4[18][47:40] = buffer_data_2[1703:1696];
        layer4[18][55:48] = buffer_data_2[1711:1704];
        layer5[18][7:0] = buffer_data_1[1663:1656];
        layer5[18][15:8] = buffer_data_1[1671:1664];
        layer5[18][23:16] = buffer_data_1[1679:1672];
        layer5[18][31:24] = buffer_data_1[1687:1680];
        layer5[18][39:32] = buffer_data_1[1695:1688];
        layer5[18][47:40] = buffer_data_1[1703:1696];
        layer5[18][55:48] = buffer_data_1[1711:1704];
        layer6[18][7:0] = buffer_data_0[1663:1656];
        layer6[18][15:8] = buffer_data_0[1671:1664];
        layer6[18][23:16] = buffer_data_0[1679:1672];
        layer6[18][31:24] = buffer_data_0[1687:1680];
        layer6[18][39:32] = buffer_data_0[1695:1688];
        layer6[18][47:40] = buffer_data_0[1703:1696];
        layer6[18][55:48] = buffer_data_0[1711:1704];
        layer0[19][7:0] = buffer_data_6[1671:1664];
        layer0[19][15:8] = buffer_data_6[1679:1672];
        layer0[19][23:16] = buffer_data_6[1687:1680];
        layer0[19][31:24] = buffer_data_6[1695:1688];
        layer0[19][39:32] = buffer_data_6[1703:1696];
        layer0[19][47:40] = buffer_data_6[1711:1704];
        layer0[19][55:48] = buffer_data_6[1719:1712];
        layer1[19][7:0] = buffer_data_5[1671:1664];
        layer1[19][15:8] = buffer_data_5[1679:1672];
        layer1[19][23:16] = buffer_data_5[1687:1680];
        layer1[19][31:24] = buffer_data_5[1695:1688];
        layer1[19][39:32] = buffer_data_5[1703:1696];
        layer1[19][47:40] = buffer_data_5[1711:1704];
        layer1[19][55:48] = buffer_data_5[1719:1712];
        layer2[19][7:0] = buffer_data_4[1671:1664];
        layer2[19][15:8] = buffer_data_4[1679:1672];
        layer2[19][23:16] = buffer_data_4[1687:1680];
        layer2[19][31:24] = buffer_data_4[1695:1688];
        layer2[19][39:32] = buffer_data_4[1703:1696];
        layer2[19][47:40] = buffer_data_4[1711:1704];
        layer2[19][55:48] = buffer_data_4[1719:1712];
        layer3[19][7:0] = buffer_data_3[1671:1664];
        layer3[19][15:8] = buffer_data_3[1679:1672];
        layer3[19][23:16] = buffer_data_3[1687:1680];
        layer3[19][31:24] = buffer_data_3[1695:1688];
        layer3[19][39:32] = buffer_data_3[1703:1696];
        layer3[19][47:40] = buffer_data_3[1711:1704];
        layer3[19][55:48] = buffer_data_3[1719:1712];
        layer4[19][7:0] = buffer_data_2[1671:1664];
        layer4[19][15:8] = buffer_data_2[1679:1672];
        layer4[19][23:16] = buffer_data_2[1687:1680];
        layer4[19][31:24] = buffer_data_2[1695:1688];
        layer4[19][39:32] = buffer_data_2[1703:1696];
        layer4[19][47:40] = buffer_data_2[1711:1704];
        layer4[19][55:48] = buffer_data_2[1719:1712];
        layer5[19][7:0] = buffer_data_1[1671:1664];
        layer5[19][15:8] = buffer_data_1[1679:1672];
        layer5[19][23:16] = buffer_data_1[1687:1680];
        layer5[19][31:24] = buffer_data_1[1695:1688];
        layer5[19][39:32] = buffer_data_1[1703:1696];
        layer5[19][47:40] = buffer_data_1[1711:1704];
        layer5[19][55:48] = buffer_data_1[1719:1712];
        layer6[19][7:0] = buffer_data_0[1671:1664];
        layer6[19][15:8] = buffer_data_0[1679:1672];
        layer6[19][23:16] = buffer_data_0[1687:1680];
        layer6[19][31:24] = buffer_data_0[1695:1688];
        layer6[19][39:32] = buffer_data_0[1703:1696];
        layer6[19][47:40] = buffer_data_0[1711:1704];
        layer6[19][55:48] = buffer_data_0[1719:1712];
        layer0[20][7:0] = buffer_data_6[1679:1672];
        layer0[20][15:8] = buffer_data_6[1687:1680];
        layer0[20][23:16] = buffer_data_6[1695:1688];
        layer0[20][31:24] = buffer_data_6[1703:1696];
        layer0[20][39:32] = buffer_data_6[1711:1704];
        layer0[20][47:40] = buffer_data_6[1719:1712];
        layer0[20][55:48] = buffer_data_6[1727:1720];
        layer1[20][7:0] = buffer_data_5[1679:1672];
        layer1[20][15:8] = buffer_data_5[1687:1680];
        layer1[20][23:16] = buffer_data_5[1695:1688];
        layer1[20][31:24] = buffer_data_5[1703:1696];
        layer1[20][39:32] = buffer_data_5[1711:1704];
        layer1[20][47:40] = buffer_data_5[1719:1712];
        layer1[20][55:48] = buffer_data_5[1727:1720];
        layer2[20][7:0] = buffer_data_4[1679:1672];
        layer2[20][15:8] = buffer_data_4[1687:1680];
        layer2[20][23:16] = buffer_data_4[1695:1688];
        layer2[20][31:24] = buffer_data_4[1703:1696];
        layer2[20][39:32] = buffer_data_4[1711:1704];
        layer2[20][47:40] = buffer_data_4[1719:1712];
        layer2[20][55:48] = buffer_data_4[1727:1720];
        layer3[20][7:0] = buffer_data_3[1679:1672];
        layer3[20][15:8] = buffer_data_3[1687:1680];
        layer3[20][23:16] = buffer_data_3[1695:1688];
        layer3[20][31:24] = buffer_data_3[1703:1696];
        layer3[20][39:32] = buffer_data_3[1711:1704];
        layer3[20][47:40] = buffer_data_3[1719:1712];
        layer3[20][55:48] = buffer_data_3[1727:1720];
        layer4[20][7:0] = buffer_data_2[1679:1672];
        layer4[20][15:8] = buffer_data_2[1687:1680];
        layer4[20][23:16] = buffer_data_2[1695:1688];
        layer4[20][31:24] = buffer_data_2[1703:1696];
        layer4[20][39:32] = buffer_data_2[1711:1704];
        layer4[20][47:40] = buffer_data_2[1719:1712];
        layer4[20][55:48] = buffer_data_2[1727:1720];
        layer5[20][7:0] = buffer_data_1[1679:1672];
        layer5[20][15:8] = buffer_data_1[1687:1680];
        layer5[20][23:16] = buffer_data_1[1695:1688];
        layer5[20][31:24] = buffer_data_1[1703:1696];
        layer5[20][39:32] = buffer_data_1[1711:1704];
        layer5[20][47:40] = buffer_data_1[1719:1712];
        layer5[20][55:48] = buffer_data_1[1727:1720];
        layer6[20][7:0] = buffer_data_0[1679:1672];
        layer6[20][15:8] = buffer_data_0[1687:1680];
        layer6[20][23:16] = buffer_data_0[1695:1688];
        layer6[20][31:24] = buffer_data_0[1703:1696];
        layer6[20][39:32] = buffer_data_0[1711:1704];
        layer6[20][47:40] = buffer_data_0[1719:1712];
        layer6[20][55:48] = buffer_data_0[1727:1720];
        layer0[21][7:0] = buffer_data_6[1687:1680];
        layer0[21][15:8] = buffer_data_6[1695:1688];
        layer0[21][23:16] = buffer_data_6[1703:1696];
        layer0[21][31:24] = buffer_data_6[1711:1704];
        layer0[21][39:32] = buffer_data_6[1719:1712];
        layer0[21][47:40] = buffer_data_6[1727:1720];
        layer0[21][55:48] = buffer_data_6[1735:1728];
        layer1[21][7:0] = buffer_data_5[1687:1680];
        layer1[21][15:8] = buffer_data_5[1695:1688];
        layer1[21][23:16] = buffer_data_5[1703:1696];
        layer1[21][31:24] = buffer_data_5[1711:1704];
        layer1[21][39:32] = buffer_data_5[1719:1712];
        layer1[21][47:40] = buffer_data_5[1727:1720];
        layer1[21][55:48] = buffer_data_5[1735:1728];
        layer2[21][7:0] = buffer_data_4[1687:1680];
        layer2[21][15:8] = buffer_data_4[1695:1688];
        layer2[21][23:16] = buffer_data_4[1703:1696];
        layer2[21][31:24] = buffer_data_4[1711:1704];
        layer2[21][39:32] = buffer_data_4[1719:1712];
        layer2[21][47:40] = buffer_data_4[1727:1720];
        layer2[21][55:48] = buffer_data_4[1735:1728];
        layer3[21][7:0] = buffer_data_3[1687:1680];
        layer3[21][15:8] = buffer_data_3[1695:1688];
        layer3[21][23:16] = buffer_data_3[1703:1696];
        layer3[21][31:24] = buffer_data_3[1711:1704];
        layer3[21][39:32] = buffer_data_3[1719:1712];
        layer3[21][47:40] = buffer_data_3[1727:1720];
        layer3[21][55:48] = buffer_data_3[1735:1728];
        layer4[21][7:0] = buffer_data_2[1687:1680];
        layer4[21][15:8] = buffer_data_2[1695:1688];
        layer4[21][23:16] = buffer_data_2[1703:1696];
        layer4[21][31:24] = buffer_data_2[1711:1704];
        layer4[21][39:32] = buffer_data_2[1719:1712];
        layer4[21][47:40] = buffer_data_2[1727:1720];
        layer4[21][55:48] = buffer_data_2[1735:1728];
        layer5[21][7:0] = buffer_data_1[1687:1680];
        layer5[21][15:8] = buffer_data_1[1695:1688];
        layer5[21][23:16] = buffer_data_1[1703:1696];
        layer5[21][31:24] = buffer_data_1[1711:1704];
        layer5[21][39:32] = buffer_data_1[1719:1712];
        layer5[21][47:40] = buffer_data_1[1727:1720];
        layer5[21][55:48] = buffer_data_1[1735:1728];
        layer6[21][7:0] = buffer_data_0[1687:1680];
        layer6[21][15:8] = buffer_data_0[1695:1688];
        layer6[21][23:16] = buffer_data_0[1703:1696];
        layer6[21][31:24] = buffer_data_0[1711:1704];
        layer6[21][39:32] = buffer_data_0[1719:1712];
        layer6[21][47:40] = buffer_data_0[1727:1720];
        layer6[21][55:48] = buffer_data_0[1735:1728];
        layer0[22][7:0] = buffer_data_6[1695:1688];
        layer0[22][15:8] = buffer_data_6[1703:1696];
        layer0[22][23:16] = buffer_data_6[1711:1704];
        layer0[22][31:24] = buffer_data_6[1719:1712];
        layer0[22][39:32] = buffer_data_6[1727:1720];
        layer0[22][47:40] = buffer_data_6[1735:1728];
        layer0[22][55:48] = buffer_data_6[1743:1736];
        layer1[22][7:0] = buffer_data_5[1695:1688];
        layer1[22][15:8] = buffer_data_5[1703:1696];
        layer1[22][23:16] = buffer_data_5[1711:1704];
        layer1[22][31:24] = buffer_data_5[1719:1712];
        layer1[22][39:32] = buffer_data_5[1727:1720];
        layer1[22][47:40] = buffer_data_5[1735:1728];
        layer1[22][55:48] = buffer_data_5[1743:1736];
        layer2[22][7:0] = buffer_data_4[1695:1688];
        layer2[22][15:8] = buffer_data_4[1703:1696];
        layer2[22][23:16] = buffer_data_4[1711:1704];
        layer2[22][31:24] = buffer_data_4[1719:1712];
        layer2[22][39:32] = buffer_data_4[1727:1720];
        layer2[22][47:40] = buffer_data_4[1735:1728];
        layer2[22][55:48] = buffer_data_4[1743:1736];
        layer3[22][7:0] = buffer_data_3[1695:1688];
        layer3[22][15:8] = buffer_data_3[1703:1696];
        layer3[22][23:16] = buffer_data_3[1711:1704];
        layer3[22][31:24] = buffer_data_3[1719:1712];
        layer3[22][39:32] = buffer_data_3[1727:1720];
        layer3[22][47:40] = buffer_data_3[1735:1728];
        layer3[22][55:48] = buffer_data_3[1743:1736];
        layer4[22][7:0] = buffer_data_2[1695:1688];
        layer4[22][15:8] = buffer_data_2[1703:1696];
        layer4[22][23:16] = buffer_data_2[1711:1704];
        layer4[22][31:24] = buffer_data_2[1719:1712];
        layer4[22][39:32] = buffer_data_2[1727:1720];
        layer4[22][47:40] = buffer_data_2[1735:1728];
        layer4[22][55:48] = buffer_data_2[1743:1736];
        layer5[22][7:0] = buffer_data_1[1695:1688];
        layer5[22][15:8] = buffer_data_1[1703:1696];
        layer5[22][23:16] = buffer_data_1[1711:1704];
        layer5[22][31:24] = buffer_data_1[1719:1712];
        layer5[22][39:32] = buffer_data_1[1727:1720];
        layer5[22][47:40] = buffer_data_1[1735:1728];
        layer5[22][55:48] = buffer_data_1[1743:1736];
        layer6[22][7:0] = buffer_data_0[1695:1688];
        layer6[22][15:8] = buffer_data_0[1703:1696];
        layer6[22][23:16] = buffer_data_0[1711:1704];
        layer6[22][31:24] = buffer_data_0[1719:1712];
        layer6[22][39:32] = buffer_data_0[1727:1720];
        layer6[22][47:40] = buffer_data_0[1735:1728];
        layer6[22][55:48] = buffer_data_0[1743:1736];
        layer0[23][7:0] = buffer_data_6[1703:1696];
        layer0[23][15:8] = buffer_data_6[1711:1704];
        layer0[23][23:16] = buffer_data_6[1719:1712];
        layer0[23][31:24] = buffer_data_6[1727:1720];
        layer0[23][39:32] = buffer_data_6[1735:1728];
        layer0[23][47:40] = buffer_data_6[1743:1736];
        layer0[23][55:48] = buffer_data_6[1751:1744];
        layer1[23][7:0] = buffer_data_5[1703:1696];
        layer1[23][15:8] = buffer_data_5[1711:1704];
        layer1[23][23:16] = buffer_data_5[1719:1712];
        layer1[23][31:24] = buffer_data_5[1727:1720];
        layer1[23][39:32] = buffer_data_5[1735:1728];
        layer1[23][47:40] = buffer_data_5[1743:1736];
        layer1[23][55:48] = buffer_data_5[1751:1744];
        layer2[23][7:0] = buffer_data_4[1703:1696];
        layer2[23][15:8] = buffer_data_4[1711:1704];
        layer2[23][23:16] = buffer_data_4[1719:1712];
        layer2[23][31:24] = buffer_data_4[1727:1720];
        layer2[23][39:32] = buffer_data_4[1735:1728];
        layer2[23][47:40] = buffer_data_4[1743:1736];
        layer2[23][55:48] = buffer_data_4[1751:1744];
        layer3[23][7:0] = buffer_data_3[1703:1696];
        layer3[23][15:8] = buffer_data_3[1711:1704];
        layer3[23][23:16] = buffer_data_3[1719:1712];
        layer3[23][31:24] = buffer_data_3[1727:1720];
        layer3[23][39:32] = buffer_data_3[1735:1728];
        layer3[23][47:40] = buffer_data_3[1743:1736];
        layer3[23][55:48] = buffer_data_3[1751:1744];
        layer4[23][7:0] = buffer_data_2[1703:1696];
        layer4[23][15:8] = buffer_data_2[1711:1704];
        layer4[23][23:16] = buffer_data_2[1719:1712];
        layer4[23][31:24] = buffer_data_2[1727:1720];
        layer4[23][39:32] = buffer_data_2[1735:1728];
        layer4[23][47:40] = buffer_data_2[1743:1736];
        layer4[23][55:48] = buffer_data_2[1751:1744];
        layer5[23][7:0] = buffer_data_1[1703:1696];
        layer5[23][15:8] = buffer_data_1[1711:1704];
        layer5[23][23:16] = buffer_data_1[1719:1712];
        layer5[23][31:24] = buffer_data_1[1727:1720];
        layer5[23][39:32] = buffer_data_1[1735:1728];
        layer5[23][47:40] = buffer_data_1[1743:1736];
        layer5[23][55:48] = buffer_data_1[1751:1744];
        layer6[23][7:0] = buffer_data_0[1703:1696];
        layer6[23][15:8] = buffer_data_0[1711:1704];
        layer6[23][23:16] = buffer_data_0[1719:1712];
        layer6[23][31:24] = buffer_data_0[1727:1720];
        layer6[23][39:32] = buffer_data_0[1735:1728];
        layer6[23][47:40] = buffer_data_0[1743:1736];
        layer6[23][55:48] = buffer_data_0[1751:1744];
        layer0[24][7:0] = buffer_data_6[1711:1704];
        layer0[24][15:8] = buffer_data_6[1719:1712];
        layer0[24][23:16] = buffer_data_6[1727:1720];
        layer0[24][31:24] = buffer_data_6[1735:1728];
        layer0[24][39:32] = buffer_data_6[1743:1736];
        layer0[24][47:40] = buffer_data_6[1751:1744];
        layer0[24][55:48] = buffer_data_6[1759:1752];
        layer1[24][7:0] = buffer_data_5[1711:1704];
        layer1[24][15:8] = buffer_data_5[1719:1712];
        layer1[24][23:16] = buffer_data_5[1727:1720];
        layer1[24][31:24] = buffer_data_5[1735:1728];
        layer1[24][39:32] = buffer_data_5[1743:1736];
        layer1[24][47:40] = buffer_data_5[1751:1744];
        layer1[24][55:48] = buffer_data_5[1759:1752];
        layer2[24][7:0] = buffer_data_4[1711:1704];
        layer2[24][15:8] = buffer_data_4[1719:1712];
        layer2[24][23:16] = buffer_data_4[1727:1720];
        layer2[24][31:24] = buffer_data_4[1735:1728];
        layer2[24][39:32] = buffer_data_4[1743:1736];
        layer2[24][47:40] = buffer_data_4[1751:1744];
        layer2[24][55:48] = buffer_data_4[1759:1752];
        layer3[24][7:0] = buffer_data_3[1711:1704];
        layer3[24][15:8] = buffer_data_3[1719:1712];
        layer3[24][23:16] = buffer_data_3[1727:1720];
        layer3[24][31:24] = buffer_data_3[1735:1728];
        layer3[24][39:32] = buffer_data_3[1743:1736];
        layer3[24][47:40] = buffer_data_3[1751:1744];
        layer3[24][55:48] = buffer_data_3[1759:1752];
        layer4[24][7:0] = buffer_data_2[1711:1704];
        layer4[24][15:8] = buffer_data_2[1719:1712];
        layer4[24][23:16] = buffer_data_2[1727:1720];
        layer4[24][31:24] = buffer_data_2[1735:1728];
        layer4[24][39:32] = buffer_data_2[1743:1736];
        layer4[24][47:40] = buffer_data_2[1751:1744];
        layer4[24][55:48] = buffer_data_2[1759:1752];
        layer5[24][7:0] = buffer_data_1[1711:1704];
        layer5[24][15:8] = buffer_data_1[1719:1712];
        layer5[24][23:16] = buffer_data_1[1727:1720];
        layer5[24][31:24] = buffer_data_1[1735:1728];
        layer5[24][39:32] = buffer_data_1[1743:1736];
        layer5[24][47:40] = buffer_data_1[1751:1744];
        layer5[24][55:48] = buffer_data_1[1759:1752];
        layer6[24][7:0] = buffer_data_0[1711:1704];
        layer6[24][15:8] = buffer_data_0[1719:1712];
        layer6[24][23:16] = buffer_data_0[1727:1720];
        layer6[24][31:24] = buffer_data_0[1735:1728];
        layer6[24][39:32] = buffer_data_0[1743:1736];
        layer6[24][47:40] = buffer_data_0[1751:1744];
        layer6[24][55:48] = buffer_data_0[1759:1752];
        layer0[25][7:0] = buffer_data_6[1719:1712];
        layer0[25][15:8] = buffer_data_6[1727:1720];
        layer0[25][23:16] = buffer_data_6[1735:1728];
        layer0[25][31:24] = buffer_data_6[1743:1736];
        layer0[25][39:32] = buffer_data_6[1751:1744];
        layer0[25][47:40] = buffer_data_6[1759:1752];
        layer0[25][55:48] = buffer_data_6[1767:1760];
        layer1[25][7:0] = buffer_data_5[1719:1712];
        layer1[25][15:8] = buffer_data_5[1727:1720];
        layer1[25][23:16] = buffer_data_5[1735:1728];
        layer1[25][31:24] = buffer_data_5[1743:1736];
        layer1[25][39:32] = buffer_data_5[1751:1744];
        layer1[25][47:40] = buffer_data_5[1759:1752];
        layer1[25][55:48] = buffer_data_5[1767:1760];
        layer2[25][7:0] = buffer_data_4[1719:1712];
        layer2[25][15:8] = buffer_data_4[1727:1720];
        layer2[25][23:16] = buffer_data_4[1735:1728];
        layer2[25][31:24] = buffer_data_4[1743:1736];
        layer2[25][39:32] = buffer_data_4[1751:1744];
        layer2[25][47:40] = buffer_data_4[1759:1752];
        layer2[25][55:48] = buffer_data_4[1767:1760];
        layer3[25][7:0] = buffer_data_3[1719:1712];
        layer3[25][15:8] = buffer_data_3[1727:1720];
        layer3[25][23:16] = buffer_data_3[1735:1728];
        layer3[25][31:24] = buffer_data_3[1743:1736];
        layer3[25][39:32] = buffer_data_3[1751:1744];
        layer3[25][47:40] = buffer_data_3[1759:1752];
        layer3[25][55:48] = buffer_data_3[1767:1760];
        layer4[25][7:0] = buffer_data_2[1719:1712];
        layer4[25][15:8] = buffer_data_2[1727:1720];
        layer4[25][23:16] = buffer_data_2[1735:1728];
        layer4[25][31:24] = buffer_data_2[1743:1736];
        layer4[25][39:32] = buffer_data_2[1751:1744];
        layer4[25][47:40] = buffer_data_2[1759:1752];
        layer4[25][55:48] = buffer_data_2[1767:1760];
        layer5[25][7:0] = buffer_data_1[1719:1712];
        layer5[25][15:8] = buffer_data_1[1727:1720];
        layer5[25][23:16] = buffer_data_1[1735:1728];
        layer5[25][31:24] = buffer_data_1[1743:1736];
        layer5[25][39:32] = buffer_data_1[1751:1744];
        layer5[25][47:40] = buffer_data_1[1759:1752];
        layer5[25][55:48] = buffer_data_1[1767:1760];
        layer6[25][7:0] = buffer_data_0[1719:1712];
        layer6[25][15:8] = buffer_data_0[1727:1720];
        layer6[25][23:16] = buffer_data_0[1735:1728];
        layer6[25][31:24] = buffer_data_0[1743:1736];
        layer6[25][39:32] = buffer_data_0[1751:1744];
        layer6[25][47:40] = buffer_data_0[1759:1752];
        layer6[25][55:48] = buffer_data_0[1767:1760];
        layer0[26][7:0] = buffer_data_6[1727:1720];
        layer0[26][15:8] = buffer_data_6[1735:1728];
        layer0[26][23:16] = buffer_data_6[1743:1736];
        layer0[26][31:24] = buffer_data_6[1751:1744];
        layer0[26][39:32] = buffer_data_6[1759:1752];
        layer0[26][47:40] = buffer_data_6[1767:1760];
        layer0[26][55:48] = buffer_data_6[1775:1768];
        layer1[26][7:0] = buffer_data_5[1727:1720];
        layer1[26][15:8] = buffer_data_5[1735:1728];
        layer1[26][23:16] = buffer_data_5[1743:1736];
        layer1[26][31:24] = buffer_data_5[1751:1744];
        layer1[26][39:32] = buffer_data_5[1759:1752];
        layer1[26][47:40] = buffer_data_5[1767:1760];
        layer1[26][55:48] = buffer_data_5[1775:1768];
        layer2[26][7:0] = buffer_data_4[1727:1720];
        layer2[26][15:8] = buffer_data_4[1735:1728];
        layer2[26][23:16] = buffer_data_4[1743:1736];
        layer2[26][31:24] = buffer_data_4[1751:1744];
        layer2[26][39:32] = buffer_data_4[1759:1752];
        layer2[26][47:40] = buffer_data_4[1767:1760];
        layer2[26][55:48] = buffer_data_4[1775:1768];
        layer3[26][7:0] = buffer_data_3[1727:1720];
        layer3[26][15:8] = buffer_data_3[1735:1728];
        layer3[26][23:16] = buffer_data_3[1743:1736];
        layer3[26][31:24] = buffer_data_3[1751:1744];
        layer3[26][39:32] = buffer_data_3[1759:1752];
        layer3[26][47:40] = buffer_data_3[1767:1760];
        layer3[26][55:48] = buffer_data_3[1775:1768];
        layer4[26][7:0] = buffer_data_2[1727:1720];
        layer4[26][15:8] = buffer_data_2[1735:1728];
        layer4[26][23:16] = buffer_data_2[1743:1736];
        layer4[26][31:24] = buffer_data_2[1751:1744];
        layer4[26][39:32] = buffer_data_2[1759:1752];
        layer4[26][47:40] = buffer_data_2[1767:1760];
        layer4[26][55:48] = buffer_data_2[1775:1768];
        layer5[26][7:0] = buffer_data_1[1727:1720];
        layer5[26][15:8] = buffer_data_1[1735:1728];
        layer5[26][23:16] = buffer_data_1[1743:1736];
        layer5[26][31:24] = buffer_data_1[1751:1744];
        layer5[26][39:32] = buffer_data_1[1759:1752];
        layer5[26][47:40] = buffer_data_1[1767:1760];
        layer5[26][55:48] = buffer_data_1[1775:1768];
        layer6[26][7:0] = buffer_data_0[1727:1720];
        layer6[26][15:8] = buffer_data_0[1735:1728];
        layer6[26][23:16] = buffer_data_0[1743:1736];
        layer6[26][31:24] = buffer_data_0[1751:1744];
        layer6[26][39:32] = buffer_data_0[1759:1752];
        layer6[26][47:40] = buffer_data_0[1767:1760];
        layer6[26][55:48] = buffer_data_0[1775:1768];
        layer0[27][7:0] = buffer_data_6[1735:1728];
        layer0[27][15:8] = buffer_data_6[1743:1736];
        layer0[27][23:16] = buffer_data_6[1751:1744];
        layer0[27][31:24] = buffer_data_6[1759:1752];
        layer0[27][39:32] = buffer_data_6[1767:1760];
        layer0[27][47:40] = buffer_data_6[1775:1768];
        layer0[27][55:48] = buffer_data_6[1783:1776];
        layer1[27][7:0] = buffer_data_5[1735:1728];
        layer1[27][15:8] = buffer_data_5[1743:1736];
        layer1[27][23:16] = buffer_data_5[1751:1744];
        layer1[27][31:24] = buffer_data_5[1759:1752];
        layer1[27][39:32] = buffer_data_5[1767:1760];
        layer1[27][47:40] = buffer_data_5[1775:1768];
        layer1[27][55:48] = buffer_data_5[1783:1776];
        layer2[27][7:0] = buffer_data_4[1735:1728];
        layer2[27][15:8] = buffer_data_4[1743:1736];
        layer2[27][23:16] = buffer_data_4[1751:1744];
        layer2[27][31:24] = buffer_data_4[1759:1752];
        layer2[27][39:32] = buffer_data_4[1767:1760];
        layer2[27][47:40] = buffer_data_4[1775:1768];
        layer2[27][55:48] = buffer_data_4[1783:1776];
        layer3[27][7:0] = buffer_data_3[1735:1728];
        layer3[27][15:8] = buffer_data_3[1743:1736];
        layer3[27][23:16] = buffer_data_3[1751:1744];
        layer3[27][31:24] = buffer_data_3[1759:1752];
        layer3[27][39:32] = buffer_data_3[1767:1760];
        layer3[27][47:40] = buffer_data_3[1775:1768];
        layer3[27][55:48] = buffer_data_3[1783:1776];
        layer4[27][7:0] = buffer_data_2[1735:1728];
        layer4[27][15:8] = buffer_data_2[1743:1736];
        layer4[27][23:16] = buffer_data_2[1751:1744];
        layer4[27][31:24] = buffer_data_2[1759:1752];
        layer4[27][39:32] = buffer_data_2[1767:1760];
        layer4[27][47:40] = buffer_data_2[1775:1768];
        layer4[27][55:48] = buffer_data_2[1783:1776];
        layer5[27][7:0] = buffer_data_1[1735:1728];
        layer5[27][15:8] = buffer_data_1[1743:1736];
        layer5[27][23:16] = buffer_data_1[1751:1744];
        layer5[27][31:24] = buffer_data_1[1759:1752];
        layer5[27][39:32] = buffer_data_1[1767:1760];
        layer5[27][47:40] = buffer_data_1[1775:1768];
        layer5[27][55:48] = buffer_data_1[1783:1776];
        layer6[27][7:0] = buffer_data_0[1735:1728];
        layer6[27][15:8] = buffer_data_0[1743:1736];
        layer6[27][23:16] = buffer_data_0[1751:1744];
        layer6[27][31:24] = buffer_data_0[1759:1752];
        layer6[27][39:32] = buffer_data_0[1767:1760];
        layer6[27][47:40] = buffer_data_0[1775:1768];
        layer6[27][55:48] = buffer_data_0[1783:1776];
        layer0[28][7:0] = buffer_data_6[1743:1736];
        layer0[28][15:8] = buffer_data_6[1751:1744];
        layer0[28][23:16] = buffer_data_6[1759:1752];
        layer0[28][31:24] = buffer_data_6[1767:1760];
        layer0[28][39:32] = buffer_data_6[1775:1768];
        layer0[28][47:40] = buffer_data_6[1783:1776];
        layer0[28][55:48] = buffer_data_6[1791:1784];
        layer1[28][7:0] = buffer_data_5[1743:1736];
        layer1[28][15:8] = buffer_data_5[1751:1744];
        layer1[28][23:16] = buffer_data_5[1759:1752];
        layer1[28][31:24] = buffer_data_5[1767:1760];
        layer1[28][39:32] = buffer_data_5[1775:1768];
        layer1[28][47:40] = buffer_data_5[1783:1776];
        layer1[28][55:48] = buffer_data_5[1791:1784];
        layer2[28][7:0] = buffer_data_4[1743:1736];
        layer2[28][15:8] = buffer_data_4[1751:1744];
        layer2[28][23:16] = buffer_data_4[1759:1752];
        layer2[28][31:24] = buffer_data_4[1767:1760];
        layer2[28][39:32] = buffer_data_4[1775:1768];
        layer2[28][47:40] = buffer_data_4[1783:1776];
        layer2[28][55:48] = buffer_data_4[1791:1784];
        layer3[28][7:0] = buffer_data_3[1743:1736];
        layer3[28][15:8] = buffer_data_3[1751:1744];
        layer3[28][23:16] = buffer_data_3[1759:1752];
        layer3[28][31:24] = buffer_data_3[1767:1760];
        layer3[28][39:32] = buffer_data_3[1775:1768];
        layer3[28][47:40] = buffer_data_3[1783:1776];
        layer3[28][55:48] = buffer_data_3[1791:1784];
        layer4[28][7:0] = buffer_data_2[1743:1736];
        layer4[28][15:8] = buffer_data_2[1751:1744];
        layer4[28][23:16] = buffer_data_2[1759:1752];
        layer4[28][31:24] = buffer_data_2[1767:1760];
        layer4[28][39:32] = buffer_data_2[1775:1768];
        layer4[28][47:40] = buffer_data_2[1783:1776];
        layer4[28][55:48] = buffer_data_2[1791:1784];
        layer5[28][7:0] = buffer_data_1[1743:1736];
        layer5[28][15:8] = buffer_data_1[1751:1744];
        layer5[28][23:16] = buffer_data_1[1759:1752];
        layer5[28][31:24] = buffer_data_1[1767:1760];
        layer5[28][39:32] = buffer_data_1[1775:1768];
        layer5[28][47:40] = buffer_data_1[1783:1776];
        layer5[28][55:48] = buffer_data_1[1791:1784];
        layer6[28][7:0] = buffer_data_0[1743:1736];
        layer6[28][15:8] = buffer_data_0[1751:1744];
        layer6[28][23:16] = buffer_data_0[1759:1752];
        layer6[28][31:24] = buffer_data_0[1767:1760];
        layer6[28][39:32] = buffer_data_0[1775:1768];
        layer6[28][47:40] = buffer_data_0[1783:1776];
        layer6[28][55:48] = buffer_data_0[1791:1784];
        layer0[29][7:0] = buffer_data_6[1751:1744];
        layer0[29][15:8] = buffer_data_6[1759:1752];
        layer0[29][23:16] = buffer_data_6[1767:1760];
        layer0[29][31:24] = buffer_data_6[1775:1768];
        layer0[29][39:32] = buffer_data_6[1783:1776];
        layer0[29][47:40] = buffer_data_6[1791:1784];
        layer0[29][55:48] = buffer_data_6[1799:1792];
        layer1[29][7:0] = buffer_data_5[1751:1744];
        layer1[29][15:8] = buffer_data_5[1759:1752];
        layer1[29][23:16] = buffer_data_5[1767:1760];
        layer1[29][31:24] = buffer_data_5[1775:1768];
        layer1[29][39:32] = buffer_data_5[1783:1776];
        layer1[29][47:40] = buffer_data_5[1791:1784];
        layer1[29][55:48] = buffer_data_5[1799:1792];
        layer2[29][7:0] = buffer_data_4[1751:1744];
        layer2[29][15:8] = buffer_data_4[1759:1752];
        layer2[29][23:16] = buffer_data_4[1767:1760];
        layer2[29][31:24] = buffer_data_4[1775:1768];
        layer2[29][39:32] = buffer_data_4[1783:1776];
        layer2[29][47:40] = buffer_data_4[1791:1784];
        layer2[29][55:48] = buffer_data_4[1799:1792];
        layer3[29][7:0] = buffer_data_3[1751:1744];
        layer3[29][15:8] = buffer_data_3[1759:1752];
        layer3[29][23:16] = buffer_data_3[1767:1760];
        layer3[29][31:24] = buffer_data_3[1775:1768];
        layer3[29][39:32] = buffer_data_3[1783:1776];
        layer3[29][47:40] = buffer_data_3[1791:1784];
        layer3[29][55:48] = buffer_data_3[1799:1792];
        layer4[29][7:0] = buffer_data_2[1751:1744];
        layer4[29][15:8] = buffer_data_2[1759:1752];
        layer4[29][23:16] = buffer_data_2[1767:1760];
        layer4[29][31:24] = buffer_data_2[1775:1768];
        layer4[29][39:32] = buffer_data_2[1783:1776];
        layer4[29][47:40] = buffer_data_2[1791:1784];
        layer4[29][55:48] = buffer_data_2[1799:1792];
        layer5[29][7:0] = buffer_data_1[1751:1744];
        layer5[29][15:8] = buffer_data_1[1759:1752];
        layer5[29][23:16] = buffer_data_1[1767:1760];
        layer5[29][31:24] = buffer_data_1[1775:1768];
        layer5[29][39:32] = buffer_data_1[1783:1776];
        layer5[29][47:40] = buffer_data_1[1791:1784];
        layer5[29][55:48] = buffer_data_1[1799:1792];
        layer6[29][7:0] = buffer_data_0[1751:1744];
        layer6[29][15:8] = buffer_data_0[1759:1752];
        layer6[29][23:16] = buffer_data_0[1767:1760];
        layer6[29][31:24] = buffer_data_0[1775:1768];
        layer6[29][39:32] = buffer_data_0[1783:1776];
        layer6[29][47:40] = buffer_data_0[1791:1784];
        layer6[29][55:48] = buffer_data_0[1799:1792];
        layer0[30][7:0] = buffer_data_6[1759:1752];
        layer0[30][15:8] = buffer_data_6[1767:1760];
        layer0[30][23:16] = buffer_data_6[1775:1768];
        layer0[30][31:24] = buffer_data_6[1783:1776];
        layer0[30][39:32] = buffer_data_6[1791:1784];
        layer0[30][47:40] = buffer_data_6[1799:1792];
        layer0[30][55:48] = buffer_data_6[1807:1800];
        layer1[30][7:0] = buffer_data_5[1759:1752];
        layer1[30][15:8] = buffer_data_5[1767:1760];
        layer1[30][23:16] = buffer_data_5[1775:1768];
        layer1[30][31:24] = buffer_data_5[1783:1776];
        layer1[30][39:32] = buffer_data_5[1791:1784];
        layer1[30][47:40] = buffer_data_5[1799:1792];
        layer1[30][55:48] = buffer_data_5[1807:1800];
        layer2[30][7:0] = buffer_data_4[1759:1752];
        layer2[30][15:8] = buffer_data_4[1767:1760];
        layer2[30][23:16] = buffer_data_4[1775:1768];
        layer2[30][31:24] = buffer_data_4[1783:1776];
        layer2[30][39:32] = buffer_data_4[1791:1784];
        layer2[30][47:40] = buffer_data_4[1799:1792];
        layer2[30][55:48] = buffer_data_4[1807:1800];
        layer3[30][7:0] = buffer_data_3[1759:1752];
        layer3[30][15:8] = buffer_data_3[1767:1760];
        layer3[30][23:16] = buffer_data_3[1775:1768];
        layer3[30][31:24] = buffer_data_3[1783:1776];
        layer3[30][39:32] = buffer_data_3[1791:1784];
        layer3[30][47:40] = buffer_data_3[1799:1792];
        layer3[30][55:48] = buffer_data_3[1807:1800];
        layer4[30][7:0] = buffer_data_2[1759:1752];
        layer4[30][15:8] = buffer_data_2[1767:1760];
        layer4[30][23:16] = buffer_data_2[1775:1768];
        layer4[30][31:24] = buffer_data_2[1783:1776];
        layer4[30][39:32] = buffer_data_2[1791:1784];
        layer4[30][47:40] = buffer_data_2[1799:1792];
        layer4[30][55:48] = buffer_data_2[1807:1800];
        layer5[30][7:0] = buffer_data_1[1759:1752];
        layer5[30][15:8] = buffer_data_1[1767:1760];
        layer5[30][23:16] = buffer_data_1[1775:1768];
        layer5[30][31:24] = buffer_data_1[1783:1776];
        layer5[30][39:32] = buffer_data_1[1791:1784];
        layer5[30][47:40] = buffer_data_1[1799:1792];
        layer5[30][55:48] = buffer_data_1[1807:1800];
        layer6[30][7:0] = buffer_data_0[1759:1752];
        layer6[30][15:8] = buffer_data_0[1767:1760];
        layer6[30][23:16] = buffer_data_0[1775:1768];
        layer6[30][31:24] = buffer_data_0[1783:1776];
        layer6[30][39:32] = buffer_data_0[1791:1784];
        layer6[30][47:40] = buffer_data_0[1799:1792];
        layer6[30][55:48] = buffer_data_0[1807:1800];
        layer0[31][7:0] = buffer_data_6[1767:1760];
        layer0[31][15:8] = buffer_data_6[1775:1768];
        layer0[31][23:16] = buffer_data_6[1783:1776];
        layer0[31][31:24] = buffer_data_6[1791:1784];
        layer0[31][39:32] = buffer_data_6[1799:1792];
        layer0[31][47:40] = buffer_data_6[1807:1800];
        layer0[31][55:48] = buffer_data_6[1815:1808];
        layer1[31][7:0] = buffer_data_5[1767:1760];
        layer1[31][15:8] = buffer_data_5[1775:1768];
        layer1[31][23:16] = buffer_data_5[1783:1776];
        layer1[31][31:24] = buffer_data_5[1791:1784];
        layer1[31][39:32] = buffer_data_5[1799:1792];
        layer1[31][47:40] = buffer_data_5[1807:1800];
        layer1[31][55:48] = buffer_data_5[1815:1808];
        layer2[31][7:0] = buffer_data_4[1767:1760];
        layer2[31][15:8] = buffer_data_4[1775:1768];
        layer2[31][23:16] = buffer_data_4[1783:1776];
        layer2[31][31:24] = buffer_data_4[1791:1784];
        layer2[31][39:32] = buffer_data_4[1799:1792];
        layer2[31][47:40] = buffer_data_4[1807:1800];
        layer2[31][55:48] = buffer_data_4[1815:1808];
        layer3[31][7:0] = buffer_data_3[1767:1760];
        layer3[31][15:8] = buffer_data_3[1775:1768];
        layer3[31][23:16] = buffer_data_3[1783:1776];
        layer3[31][31:24] = buffer_data_3[1791:1784];
        layer3[31][39:32] = buffer_data_3[1799:1792];
        layer3[31][47:40] = buffer_data_3[1807:1800];
        layer3[31][55:48] = buffer_data_3[1815:1808];
        layer4[31][7:0] = buffer_data_2[1767:1760];
        layer4[31][15:8] = buffer_data_2[1775:1768];
        layer4[31][23:16] = buffer_data_2[1783:1776];
        layer4[31][31:24] = buffer_data_2[1791:1784];
        layer4[31][39:32] = buffer_data_2[1799:1792];
        layer4[31][47:40] = buffer_data_2[1807:1800];
        layer4[31][55:48] = buffer_data_2[1815:1808];
        layer5[31][7:0] = buffer_data_1[1767:1760];
        layer5[31][15:8] = buffer_data_1[1775:1768];
        layer5[31][23:16] = buffer_data_1[1783:1776];
        layer5[31][31:24] = buffer_data_1[1791:1784];
        layer5[31][39:32] = buffer_data_1[1799:1792];
        layer5[31][47:40] = buffer_data_1[1807:1800];
        layer5[31][55:48] = buffer_data_1[1815:1808];
        layer6[31][7:0] = buffer_data_0[1767:1760];
        layer6[31][15:8] = buffer_data_0[1775:1768];
        layer6[31][23:16] = buffer_data_0[1783:1776];
        layer6[31][31:24] = buffer_data_0[1791:1784];
        layer6[31][39:32] = buffer_data_0[1799:1792];
        layer6[31][47:40] = buffer_data_0[1807:1800];
        layer6[31][55:48] = buffer_data_0[1815:1808];
        layer0[32][7:0] = buffer_data_6[1775:1768];
        layer0[32][15:8] = buffer_data_6[1783:1776];
        layer0[32][23:16] = buffer_data_6[1791:1784];
        layer0[32][31:24] = buffer_data_6[1799:1792];
        layer0[32][39:32] = buffer_data_6[1807:1800];
        layer0[32][47:40] = buffer_data_6[1815:1808];
        layer0[32][55:48] = buffer_data_6[1823:1816];
        layer1[32][7:0] = buffer_data_5[1775:1768];
        layer1[32][15:8] = buffer_data_5[1783:1776];
        layer1[32][23:16] = buffer_data_5[1791:1784];
        layer1[32][31:24] = buffer_data_5[1799:1792];
        layer1[32][39:32] = buffer_data_5[1807:1800];
        layer1[32][47:40] = buffer_data_5[1815:1808];
        layer1[32][55:48] = buffer_data_5[1823:1816];
        layer2[32][7:0] = buffer_data_4[1775:1768];
        layer2[32][15:8] = buffer_data_4[1783:1776];
        layer2[32][23:16] = buffer_data_4[1791:1784];
        layer2[32][31:24] = buffer_data_4[1799:1792];
        layer2[32][39:32] = buffer_data_4[1807:1800];
        layer2[32][47:40] = buffer_data_4[1815:1808];
        layer2[32][55:48] = buffer_data_4[1823:1816];
        layer3[32][7:0] = buffer_data_3[1775:1768];
        layer3[32][15:8] = buffer_data_3[1783:1776];
        layer3[32][23:16] = buffer_data_3[1791:1784];
        layer3[32][31:24] = buffer_data_3[1799:1792];
        layer3[32][39:32] = buffer_data_3[1807:1800];
        layer3[32][47:40] = buffer_data_3[1815:1808];
        layer3[32][55:48] = buffer_data_3[1823:1816];
        layer4[32][7:0] = buffer_data_2[1775:1768];
        layer4[32][15:8] = buffer_data_2[1783:1776];
        layer4[32][23:16] = buffer_data_2[1791:1784];
        layer4[32][31:24] = buffer_data_2[1799:1792];
        layer4[32][39:32] = buffer_data_2[1807:1800];
        layer4[32][47:40] = buffer_data_2[1815:1808];
        layer4[32][55:48] = buffer_data_2[1823:1816];
        layer5[32][7:0] = buffer_data_1[1775:1768];
        layer5[32][15:8] = buffer_data_1[1783:1776];
        layer5[32][23:16] = buffer_data_1[1791:1784];
        layer5[32][31:24] = buffer_data_1[1799:1792];
        layer5[32][39:32] = buffer_data_1[1807:1800];
        layer5[32][47:40] = buffer_data_1[1815:1808];
        layer5[32][55:48] = buffer_data_1[1823:1816];
        layer6[32][7:0] = buffer_data_0[1775:1768];
        layer6[32][15:8] = buffer_data_0[1783:1776];
        layer6[32][23:16] = buffer_data_0[1791:1784];
        layer6[32][31:24] = buffer_data_0[1799:1792];
        layer6[32][39:32] = buffer_data_0[1807:1800];
        layer6[32][47:40] = buffer_data_0[1815:1808];
        layer6[32][55:48] = buffer_data_0[1823:1816];
        layer0[33][7:0] = buffer_data_6[1783:1776];
        layer0[33][15:8] = buffer_data_6[1791:1784];
        layer0[33][23:16] = buffer_data_6[1799:1792];
        layer0[33][31:24] = buffer_data_6[1807:1800];
        layer0[33][39:32] = buffer_data_6[1815:1808];
        layer0[33][47:40] = buffer_data_6[1823:1816];
        layer0[33][55:48] = buffer_data_6[1831:1824];
        layer1[33][7:0] = buffer_data_5[1783:1776];
        layer1[33][15:8] = buffer_data_5[1791:1784];
        layer1[33][23:16] = buffer_data_5[1799:1792];
        layer1[33][31:24] = buffer_data_5[1807:1800];
        layer1[33][39:32] = buffer_data_5[1815:1808];
        layer1[33][47:40] = buffer_data_5[1823:1816];
        layer1[33][55:48] = buffer_data_5[1831:1824];
        layer2[33][7:0] = buffer_data_4[1783:1776];
        layer2[33][15:8] = buffer_data_4[1791:1784];
        layer2[33][23:16] = buffer_data_4[1799:1792];
        layer2[33][31:24] = buffer_data_4[1807:1800];
        layer2[33][39:32] = buffer_data_4[1815:1808];
        layer2[33][47:40] = buffer_data_4[1823:1816];
        layer2[33][55:48] = buffer_data_4[1831:1824];
        layer3[33][7:0] = buffer_data_3[1783:1776];
        layer3[33][15:8] = buffer_data_3[1791:1784];
        layer3[33][23:16] = buffer_data_3[1799:1792];
        layer3[33][31:24] = buffer_data_3[1807:1800];
        layer3[33][39:32] = buffer_data_3[1815:1808];
        layer3[33][47:40] = buffer_data_3[1823:1816];
        layer3[33][55:48] = buffer_data_3[1831:1824];
        layer4[33][7:0] = buffer_data_2[1783:1776];
        layer4[33][15:8] = buffer_data_2[1791:1784];
        layer4[33][23:16] = buffer_data_2[1799:1792];
        layer4[33][31:24] = buffer_data_2[1807:1800];
        layer4[33][39:32] = buffer_data_2[1815:1808];
        layer4[33][47:40] = buffer_data_2[1823:1816];
        layer4[33][55:48] = buffer_data_2[1831:1824];
        layer5[33][7:0] = buffer_data_1[1783:1776];
        layer5[33][15:8] = buffer_data_1[1791:1784];
        layer5[33][23:16] = buffer_data_1[1799:1792];
        layer5[33][31:24] = buffer_data_1[1807:1800];
        layer5[33][39:32] = buffer_data_1[1815:1808];
        layer5[33][47:40] = buffer_data_1[1823:1816];
        layer5[33][55:48] = buffer_data_1[1831:1824];
        layer6[33][7:0] = buffer_data_0[1783:1776];
        layer6[33][15:8] = buffer_data_0[1791:1784];
        layer6[33][23:16] = buffer_data_0[1799:1792];
        layer6[33][31:24] = buffer_data_0[1807:1800];
        layer6[33][39:32] = buffer_data_0[1815:1808];
        layer6[33][47:40] = buffer_data_0[1823:1816];
        layer6[33][55:48] = buffer_data_0[1831:1824];
        layer0[34][7:0] = buffer_data_6[1791:1784];
        layer0[34][15:8] = buffer_data_6[1799:1792];
        layer0[34][23:16] = buffer_data_6[1807:1800];
        layer0[34][31:24] = buffer_data_6[1815:1808];
        layer0[34][39:32] = buffer_data_6[1823:1816];
        layer0[34][47:40] = buffer_data_6[1831:1824];
        layer0[34][55:48] = buffer_data_6[1839:1832];
        layer1[34][7:0] = buffer_data_5[1791:1784];
        layer1[34][15:8] = buffer_data_5[1799:1792];
        layer1[34][23:16] = buffer_data_5[1807:1800];
        layer1[34][31:24] = buffer_data_5[1815:1808];
        layer1[34][39:32] = buffer_data_5[1823:1816];
        layer1[34][47:40] = buffer_data_5[1831:1824];
        layer1[34][55:48] = buffer_data_5[1839:1832];
        layer2[34][7:0] = buffer_data_4[1791:1784];
        layer2[34][15:8] = buffer_data_4[1799:1792];
        layer2[34][23:16] = buffer_data_4[1807:1800];
        layer2[34][31:24] = buffer_data_4[1815:1808];
        layer2[34][39:32] = buffer_data_4[1823:1816];
        layer2[34][47:40] = buffer_data_4[1831:1824];
        layer2[34][55:48] = buffer_data_4[1839:1832];
        layer3[34][7:0] = buffer_data_3[1791:1784];
        layer3[34][15:8] = buffer_data_3[1799:1792];
        layer3[34][23:16] = buffer_data_3[1807:1800];
        layer3[34][31:24] = buffer_data_3[1815:1808];
        layer3[34][39:32] = buffer_data_3[1823:1816];
        layer3[34][47:40] = buffer_data_3[1831:1824];
        layer3[34][55:48] = buffer_data_3[1839:1832];
        layer4[34][7:0] = buffer_data_2[1791:1784];
        layer4[34][15:8] = buffer_data_2[1799:1792];
        layer4[34][23:16] = buffer_data_2[1807:1800];
        layer4[34][31:24] = buffer_data_2[1815:1808];
        layer4[34][39:32] = buffer_data_2[1823:1816];
        layer4[34][47:40] = buffer_data_2[1831:1824];
        layer4[34][55:48] = buffer_data_2[1839:1832];
        layer5[34][7:0] = buffer_data_1[1791:1784];
        layer5[34][15:8] = buffer_data_1[1799:1792];
        layer5[34][23:16] = buffer_data_1[1807:1800];
        layer5[34][31:24] = buffer_data_1[1815:1808];
        layer5[34][39:32] = buffer_data_1[1823:1816];
        layer5[34][47:40] = buffer_data_1[1831:1824];
        layer5[34][55:48] = buffer_data_1[1839:1832];
        layer6[34][7:0] = buffer_data_0[1791:1784];
        layer6[34][15:8] = buffer_data_0[1799:1792];
        layer6[34][23:16] = buffer_data_0[1807:1800];
        layer6[34][31:24] = buffer_data_0[1815:1808];
        layer6[34][39:32] = buffer_data_0[1823:1816];
        layer6[34][47:40] = buffer_data_0[1831:1824];
        layer6[34][55:48] = buffer_data_0[1839:1832];
        layer0[35][7:0] = buffer_data_6[1799:1792];
        layer0[35][15:8] = buffer_data_6[1807:1800];
        layer0[35][23:16] = buffer_data_6[1815:1808];
        layer0[35][31:24] = buffer_data_6[1823:1816];
        layer0[35][39:32] = buffer_data_6[1831:1824];
        layer0[35][47:40] = buffer_data_6[1839:1832];
        layer0[35][55:48] = buffer_data_6[1847:1840];
        layer1[35][7:0] = buffer_data_5[1799:1792];
        layer1[35][15:8] = buffer_data_5[1807:1800];
        layer1[35][23:16] = buffer_data_5[1815:1808];
        layer1[35][31:24] = buffer_data_5[1823:1816];
        layer1[35][39:32] = buffer_data_5[1831:1824];
        layer1[35][47:40] = buffer_data_5[1839:1832];
        layer1[35][55:48] = buffer_data_5[1847:1840];
        layer2[35][7:0] = buffer_data_4[1799:1792];
        layer2[35][15:8] = buffer_data_4[1807:1800];
        layer2[35][23:16] = buffer_data_4[1815:1808];
        layer2[35][31:24] = buffer_data_4[1823:1816];
        layer2[35][39:32] = buffer_data_4[1831:1824];
        layer2[35][47:40] = buffer_data_4[1839:1832];
        layer2[35][55:48] = buffer_data_4[1847:1840];
        layer3[35][7:0] = buffer_data_3[1799:1792];
        layer3[35][15:8] = buffer_data_3[1807:1800];
        layer3[35][23:16] = buffer_data_3[1815:1808];
        layer3[35][31:24] = buffer_data_3[1823:1816];
        layer3[35][39:32] = buffer_data_3[1831:1824];
        layer3[35][47:40] = buffer_data_3[1839:1832];
        layer3[35][55:48] = buffer_data_3[1847:1840];
        layer4[35][7:0] = buffer_data_2[1799:1792];
        layer4[35][15:8] = buffer_data_2[1807:1800];
        layer4[35][23:16] = buffer_data_2[1815:1808];
        layer4[35][31:24] = buffer_data_2[1823:1816];
        layer4[35][39:32] = buffer_data_2[1831:1824];
        layer4[35][47:40] = buffer_data_2[1839:1832];
        layer4[35][55:48] = buffer_data_2[1847:1840];
        layer5[35][7:0] = buffer_data_1[1799:1792];
        layer5[35][15:8] = buffer_data_1[1807:1800];
        layer5[35][23:16] = buffer_data_1[1815:1808];
        layer5[35][31:24] = buffer_data_1[1823:1816];
        layer5[35][39:32] = buffer_data_1[1831:1824];
        layer5[35][47:40] = buffer_data_1[1839:1832];
        layer5[35][55:48] = buffer_data_1[1847:1840];
        layer6[35][7:0] = buffer_data_0[1799:1792];
        layer6[35][15:8] = buffer_data_0[1807:1800];
        layer6[35][23:16] = buffer_data_0[1815:1808];
        layer6[35][31:24] = buffer_data_0[1823:1816];
        layer6[35][39:32] = buffer_data_0[1831:1824];
        layer6[35][47:40] = buffer_data_0[1839:1832];
        layer6[35][55:48] = buffer_data_0[1847:1840];
        layer0[36][7:0] = buffer_data_6[1807:1800];
        layer0[36][15:8] = buffer_data_6[1815:1808];
        layer0[36][23:16] = buffer_data_6[1823:1816];
        layer0[36][31:24] = buffer_data_6[1831:1824];
        layer0[36][39:32] = buffer_data_6[1839:1832];
        layer0[36][47:40] = buffer_data_6[1847:1840];
        layer0[36][55:48] = buffer_data_6[1855:1848];
        layer1[36][7:0] = buffer_data_5[1807:1800];
        layer1[36][15:8] = buffer_data_5[1815:1808];
        layer1[36][23:16] = buffer_data_5[1823:1816];
        layer1[36][31:24] = buffer_data_5[1831:1824];
        layer1[36][39:32] = buffer_data_5[1839:1832];
        layer1[36][47:40] = buffer_data_5[1847:1840];
        layer1[36][55:48] = buffer_data_5[1855:1848];
        layer2[36][7:0] = buffer_data_4[1807:1800];
        layer2[36][15:8] = buffer_data_4[1815:1808];
        layer2[36][23:16] = buffer_data_4[1823:1816];
        layer2[36][31:24] = buffer_data_4[1831:1824];
        layer2[36][39:32] = buffer_data_4[1839:1832];
        layer2[36][47:40] = buffer_data_4[1847:1840];
        layer2[36][55:48] = buffer_data_4[1855:1848];
        layer3[36][7:0] = buffer_data_3[1807:1800];
        layer3[36][15:8] = buffer_data_3[1815:1808];
        layer3[36][23:16] = buffer_data_3[1823:1816];
        layer3[36][31:24] = buffer_data_3[1831:1824];
        layer3[36][39:32] = buffer_data_3[1839:1832];
        layer3[36][47:40] = buffer_data_3[1847:1840];
        layer3[36][55:48] = buffer_data_3[1855:1848];
        layer4[36][7:0] = buffer_data_2[1807:1800];
        layer4[36][15:8] = buffer_data_2[1815:1808];
        layer4[36][23:16] = buffer_data_2[1823:1816];
        layer4[36][31:24] = buffer_data_2[1831:1824];
        layer4[36][39:32] = buffer_data_2[1839:1832];
        layer4[36][47:40] = buffer_data_2[1847:1840];
        layer4[36][55:48] = buffer_data_2[1855:1848];
        layer5[36][7:0] = buffer_data_1[1807:1800];
        layer5[36][15:8] = buffer_data_1[1815:1808];
        layer5[36][23:16] = buffer_data_1[1823:1816];
        layer5[36][31:24] = buffer_data_1[1831:1824];
        layer5[36][39:32] = buffer_data_1[1839:1832];
        layer5[36][47:40] = buffer_data_1[1847:1840];
        layer5[36][55:48] = buffer_data_1[1855:1848];
        layer6[36][7:0] = buffer_data_0[1807:1800];
        layer6[36][15:8] = buffer_data_0[1815:1808];
        layer6[36][23:16] = buffer_data_0[1823:1816];
        layer6[36][31:24] = buffer_data_0[1831:1824];
        layer6[36][39:32] = buffer_data_0[1839:1832];
        layer6[36][47:40] = buffer_data_0[1847:1840];
        layer6[36][55:48] = buffer_data_0[1855:1848];
        layer0[37][7:0] = buffer_data_6[1815:1808];
        layer0[37][15:8] = buffer_data_6[1823:1816];
        layer0[37][23:16] = buffer_data_6[1831:1824];
        layer0[37][31:24] = buffer_data_6[1839:1832];
        layer0[37][39:32] = buffer_data_6[1847:1840];
        layer0[37][47:40] = buffer_data_6[1855:1848];
        layer0[37][55:48] = buffer_data_6[1863:1856];
        layer1[37][7:0] = buffer_data_5[1815:1808];
        layer1[37][15:8] = buffer_data_5[1823:1816];
        layer1[37][23:16] = buffer_data_5[1831:1824];
        layer1[37][31:24] = buffer_data_5[1839:1832];
        layer1[37][39:32] = buffer_data_5[1847:1840];
        layer1[37][47:40] = buffer_data_5[1855:1848];
        layer1[37][55:48] = buffer_data_5[1863:1856];
        layer2[37][7:0] = buffer_data_4[1815:1808];
        layer2[37][15:8] = buffer_data_4[1823:1816];
        layer2[37][23:16] = buffer_data_4[1831:1824];
        layer2[37][31:24] = buffer_data_4[1839:1832];
        layer2[37][39:32] = buffer_data_4[1847:1840];
        layer2[37][47:40] = buffer_data_4[1855:1848];
        layer2[37][55:48] = buffer_data_4[1863:1856];
        layer3[37][7:0] = buffer_data_3[1815:1808];
        layer3[37][15:8] = buffer_data_3[1823:1816];
        layer3[37][23:16] = buffer_data_3[1831:1824];
        layer3[37][31:24] = buffer_data_3[1839:1832];
        layer3[37][39:32] = buffer_data_3[1847:1840];
        layer3[37][47:40] = buffer_data_3[1855:1848];
        layer3[37][55:48] = buffer_data_3[1863:1856];
        layer4[37][7:0] = buffer_data_2[1815:1808];
        layer4[37][15:8] = buffer_data_2[1823:1816];
        layer4[37][23:16] = buffer_data_2[1831:1824];
        layer4[37][31:24] = buffer_data_2[1839:1832];
        layer4[37][39:32] = buffer_data_2[1847:1840];
        layer4[37][47:40] = buffer_data_2[1855:1848];
        layer4[37][55:48] = buffer_data_2[1863:1856];
        layer5[37][7:0] = buffer_data_1[1815:1808];
        layer5[37][15:8] = buffer_data_1[1823:1816];
        layer5[37][23:16] = buffer_data_1[1831:1824];
        layer5[37][31:24] = buffer_data_1[1839:1832];
        layer5[37][39:32] = buffer_data_1[1847:1840];
        layer5[37][47:40] = buffer_data_1[1855:1848];
        layer5[37][55:48] = buffer_data_1[1863:1856];
        layer6[37][7:0] = buffer_data_0[1815:1808];
        layer6[37][15:8] = buffer_data_0[1823:1816];
        layer6[37][23:16] = buffer_data_0[1831:1824];
        layer6[37][31:24] = buffer_data_0[1839:1832];
        layer6[37][39:32] = buffer_data_0[1847:1840];
        layer6[37][47:40] = buffer_data_0[1855:1848];
        layer6[37][55:48] = buffer_data_0[1863:1856];
        layer0[38][7:0] = buffer_data_6[1823:1816];
        layer0[38][15:8] = buffer_data_6[1831:1824];
        layer0[38][23:16] = buffer_data_6[1839:1832];
        layer0[38][31:24] = buffer_data_6[1847:1840];
        layer0[38][39:32] = buffer_data_6[1855:1848];
        layer0[38][47:40] = buffer_data_6[1863:1856];
        layer0[38][55:48] = buffer_data_6[1871:1864];
        layer1[38][7:0] = buffer_data_5[1823:1816];
        layer1[38][15:8] = buffer_data_5[1831:1824];
        layer1[38][23:16] = buffer_data_5[1839:1832];
        layer1[38][31:24] = buffer_data_5[1847:1840];
        layer1[38][39:32] = buffer_data_5[1855:1848];
        layer1[38][47:40] = buffer_data_5[1863:1856];
        layer1[38][55:48] = buffer_data_5[1871:1864];
        layer2[38][7:0] = buffer_data_4[1823:1816];
        layer2[38][15:8] = buffer_data_4[1831:1824];
        layer2[38][23:16] = buffer_data_4[1839:1832];
        layer2[38][31:24] = buffer_data_4[1847:1840];
        layer2[38][39:32] = buffer_data_4[1855:1848];
        layer2[38][47:40] = buffer_data_4[1863:1856];
        layer2[38][55:48] = buffer_data_4[1871:1864];
        layer3[38][7:0] = buffer_data_3[1823:1816];
        layer3[38][15:8] = buffer_data_3[1831:1824];
        layer3[38][23:16] = buffer_data_3[1839:1832];
        layer3[38][31:24] = buffer_data_3[1847:1840];
        layer3[38][39:32] = buffer_data_3[1855:1848];
        layer3[38][47:40] = buffer_data_3[1863:1856];
        layer3[38][55:48] = buffer_data_3[1871:1864];
        layer4[38][7:0] = buffer_data_2[1823:1816];
        layer4[38][15:8] = buffer_data_2[1831:1824];
        layer4[38][23:16] = buffer_data_2[1839:1832];
        layer4[38][31:24] = buffer_data_2[1847:1840];
        layer4[38][39:32] = buffer_data_2[1855:1848];
        layer4[38][47:40] = buffer_data_2[1863:1856];
        layer4[38][55:48] = buffer_data_2[1871:1864];
        layer5[38][7:0] = buffer_data_1[1823:1816];
        layer5[38][15:8] = buffer_data_1[1831:1824];
        layer5[38][23:16] = buffer_data_1[1839:1832];
        layer5[38][31:24] = buffer_data_1[1847:1840];
        layer5[38][39:32] = buffer_data_1[1855:1848];
        layer5[38][47:40] = buffer_data_1[1863:1856];
        layer5[38][55:48] = buffer_data_1[1871:1864];
        layer6[38][7:0] = buffer_data_0[1823:1816];
        layer6[38][15:8] = buffer_data_0[1831:1824];
        layer6[38][23:16] = buffer_data_0[1839:1832];
        layer6[38][31:24] = buffer_data_0[1847:1840];
        layer6[38][39:32] = buffer_data_0[1855:1848];
        layer6[38][47:40] = buffer_data_0[1863:1856];
        layer6[38][55:48] = buffer_data_0[1871:1864];
        layer0[39][7:0] = buffer_data_6[1831:1824];
        layer0[39][15:8] = buffer_data_6[1839:1832];
        layer0[39][23:16] = buffer_data_6[1847:1840];
        layer0[39][31:24] = buffer_data_6[1855:1848];
        layer0[39][39:32] = buffer_data_6[1863:1856];
        layer0[39][47:40] = buffer_data_6[1871:1864];
        layer0[39][55:48] = buffer_data_6[1879:1872];
        layer1[39][7:0] = buffer_data_5[1831:1824];
        layer1[39][15:8] = buffer_data_5[1839:1832];
        layer1[39][23:16] = buffer_data_5[1847:1840];
        layer1[39][31:24] = buffer_data_5[1855:1848];
        layer1[39][39:32] = buffer_data_5[1863:1856];
        layer1[39][47:40] = buffer_data_5[1871:1864];
        layer1[39][55:48] = buffer_data_5[1879:1872];
        layer2[39][7:0] = buffer_data_4[1831:1824];
        layer2[39][15:8] = buffer_data_4[1839:1832];
        layer2[39][23:16] = buffer_data_4[1847:1840];
        layer2[39][31:24] = buffer_data_4[1855:1848];
        layer2[39][39:32] = buffer_data_4[1863:1856];
        layer2[39][47:40] = buffer_data_4[1871:1864];
        layer2[39][55:48] = buffer_data_4[1879:1872];
        layer3[39][7:0] = buffer_data_3[1831:1824];
        layer3[39][15:8] = buffer_data_3[1839:1832];
        layer3[39][23:16] = buffer_data_3[1847:1840];
        layer3[39][31:24] = buffer_data_3[1855:1848];
        layer3[39][39:32] = buffer_data_3[1863:1856];
        layer3[39][47:40] = buffer_data_3[1871:1864];
        layer3[39][55:48] = buffer_data_3[1879:1872];
        layer4[39][7:0] = buffer_data_2[1831:1824];
        layer4[39][15:8] = buffer_data_2[1839:1832];
        layer4[39][23:16] = buffer_data_2[1847:1840];
        layer4[39][31:24] = buffer_data_2[1855:1848];
        layer4[39][39:32] = buffer_data_2[1863:1856];
        layer4[39][47:40] = buffer_data_2[1871:1864];
        layer4[39][55:48] = buffer_data_2[1879:1872];
        layer5[39][7:0] = buffer_data_1[1831:1824];
        layer5[39][15:8] = buffer_data_1[1839:1832];
        layer5[39][23:16] = buffer_data_1[1847:1840];
        layer5[39][31:24] = buffer_data_1[1855:1848];
        layer5[39][39:32] = buffer_data_1[1863:1856];
        layer5[39][47:40] = buffer_data_1[1871:1864];
        layer5[39][55:48] = buffer_data_1[1879:1872];
        layer6[39][7:0] = buffer_data_0[1831:1824];
        layer6[39][15:8] = buffer_data_0[1839:1832];
        layer6[39][23:16] = buffer_data_0[1847:1840];
        layer6[39][31:24] = buffer_data_0[1855:1848];
        layer6[39][39:32] = buffer_data_0[1863:1856];
        layer6[39][47:40] = buffer_data_0[1871:1864];
        layer6[39][55:48] = buffer_data_0[1879:1872];
        layer0[40][7:0] = buffer_data_6[1839:1832];
        layer0[40][15:8] = buffer_data_6[1847:1840];
        layer0[40][23:16] = buffer_data_6[1855:1848];
        layer0[40][31:24] = buffer_data_6[1863:1856];
        layer0[40][39:32] = buffer_data_6[1871:1864];
        layer0[40][47:40] = buffer_data_6[1879:1872];
        layer0[40][55:48] = buffer_data_6[1887:1880];
        layer1[40][7:0] = buffer_data_5[1839:1832];
        layer1[40][15:8] = buffer_data_5[1847:1840];
        layer1[40][23:16] = buffer_data_5[1855:1848];
        layer1[40][31:24] = buffer_data_5[1863:1856];
        layer1[40][39:32] = buffer_data_5[1871:1864];
        layer1[40][47:40] = buffer_data_5[1879:1872];
        layer1[40][55:48] = buffer_data_5[1887:1880];
        layer2[40][7:0] = buffer_data_4[1839:1832];
        layer2[40][15:8] = buffer_data_4[1847:1840];
        layer2[40][23:16] = buffer_data_4[1855:1848];
        layer2[40][31:24] = buffer_data_4[1863:1856];
        layer2[40][39:32] = buffer_data_4[1871:1864];
        layer2[40][47:40] = buffer_data_4[1879:1872];
        layer2[40][55:48] = buffer_data_4[1887:1880];
        layer3[40][7:0] = buffer_data_3[1839:1832];
        layer3[40][15:8] = buffer_data_3[1847:1840];
        layer3[40][23:16] = buffer_data_3[1855:1848];
        layer3[40][31:24] = buffer_data_3[1863:1856];
        layer3[40][39:32] = buffer_data_3[1871:1864];
        layer3[40][47:40] = buffer_data_3[1879:1872];
        layer3[40][55:48] = buffer_data_3[1887:1880];
        layer4[40][7:0] = buffer_data_2[1839:1832];
        layer4[40][15:8] = buffer_data_2[1847:1840];
        layer4[40][23:16] = buffer_data_2[1855:1848];
        layer4[40][31:24] = buffer_data_2[1863:1856];
        layer4[40][39:32] = buffer_data_2[1871:1864];
        layer4[40][47:40] = buffer_data_2[1879:1872];
        layer4[40][55:48] = buffer_data_2[1887:1880];
        layer5[40][7:0] = buffer_data_1[1839:1832];
        layer5[40][15:8] = buffer_data_1[1847:1840];
        layer5[40][23:16] = buffer_data_1[1855:1848];
        layer5[40][31:24] = buffer_data_1[1863:1856];
        layer5[40][39:32] = buffer_data_1[1871:1864];
        layer5[40][47:40] = buffer_data_1[1879:1872];
        layer5[40][55:48] = buffer_data_1[1887:1880];
        layer6[40][7:0] = buffer_data_0[1839:1832];
        layer6[40][15:8] = buffer_data_0[1847:1840];
        layer6[40][23:16] = buffer_data_0[1855:1848];
        layer6[40][31:24] = buffer_data_0[1863:1856];
        layer6[40][39:32] = buffer_data_0[1871:1864];
        layer6[40][47:40] = buffer_data_0[1879:1872];
        layer6[40][55:48] = buffer_data_0[1887:1880];
        layer0[41][7:0] = buffer_data_6[1847:1840];
        layer0[41][15:8] = buffer_data_6[1855:1848];
        layer0[41][23:16] = buffer_data_6[1863:1856];
        layer0[41][31:24] = buffer_data_6[1871:1864];
        layer0[41][39:32] = buffer_data_6[1879:1872];
        layer0[41][47:40] = buffer_data_6[1887:1880];
        layer0[41][55:48] = buffer_data_6[1895:1888];
        layer1[41][7:0] = buffer_data_5[1847:1840];
        layer1[41][15:8] = buffer_data_5[1855:1848];
        layer1[41][23:16] = buffer_data_5[1863:1856];
        layer1[41][31:24] = buffer_data_5[1871:1864];
        layer1[41][39:32] = buffer_data_5[1879:1872];
        layer1[41][47:40] = buffer_data_5[1887:1880];
        layer1[41][55:48] = buffer_data_5[1895:1888];
        layer2[41][7:0] = buffer_data_4[1847:1840];
        layer2[41][15:8] = buffer_data_4[1855:1848];
        layer2[41][23:16] = buffer_data_4[1863:1856];
        layer2[41][31:24] = buffer_data_4[1871:1864];
        layer2[41][39:32] = buffer_data_4[1879:1872];
        layer2[41][47:40] = buffer_data_4[1887:1880];
        layer2[41][55:48] = buffer_data_4[1895:1888];
        layer3[41][7:0] = buffer_data_3[1847:1840];
        layer3[41][15:8] = buffer_data_3[1855:1848];
        layer3[41][23:16] = buffer_data_3[1863:1856];
        layer3[41][31:24] = buffer_data_3[1871:1864];
        layer3[41][39:32] = buffer_data_3[1879:1872];
        layer3[41][47:40] = buffer_data_3[1887:1880];
        layer3[41][55:48] = buffer_data_3[1895:1888];
        layer4[41][7:0] = buffer_data_2[1847:1840];
        layer4[41][15:8] = buffer_data_2[1855:1848];
        layer4[41][23:16] = buffer_data_2[1863:1856];
        layer4[41][31:24] = buffer_data_2[1871:1864];
        layer4[41][39:32] = buffer_data_2[1879:1872];
        layer4[41][47:40] = buffer_data_2[1887:1880];
        layer4[41][55:48] = buffer_data_2[1895:1888];
        layer5[41][7:0] = buffer_data_1[1847:1840];
        layer5[41][15:8] = buffer_data_1[1855:1848];
        layer5[41][23:16] = buffer_data_1[1863:1856];
        layer5[41][31:24] = buffer_data_1[1871:1864];
        layer5[41][39:32] = buffer_data_1[1879:1872];
        layer5[41][47:40] = buffer_data_1[1887:1880];
        layer5[41][55:48] = buffer_data_1[1895:1888];
        layer6[41][7:0] = buffer_data_0[1847:1840];
        layer6[41][15:8] = buffer_data_0[1855:1848];
        layer6[41][23:16] = buffer_data_0[1863:1856];
        layer6[41][31:24] = buffer_data_0[1871:1864];
        layer6[41][39:32] = buffer_data_0[1879:1872];
        layer6[41][47:40] = buffer_data_0[1887:1880];
        layer6[41][55:48] = buffer_data_0[1895:1888];
        layer0[42][7:0] = buffer_data_6[1855:1848];
        layer0[42][15:8] = buffer_data_6[1863:1856];
        layer0[42][23:16] = buffer_data_6[1871:1864];
        layer0[42][31:24] = buffer_data_6[1879:1872];
        layer0[42][39:32] = buffer_data_6[1887:1880];
        layer0[42][47:40] = buffer_data_6[1895:1888];
        layer0[42][55:48] = buffer_data_6[1903:1896];
        layer1[42][7:0] = buffer_data_5[1855:1848];
        layer1[42][15:8] = buffer_data_5[1863:1856];
        layer1[42][23:16] = buffer_data_5[1871:1864];
        layer1[42][31:24] = buffer_data_5[1879:1872];
        layer1[42][39:32] = buffer_data_5[1887:1880];
        layer1[42][47:40] = buffer_data_5[1895:1888];
        layer1[42][55:48] = buffer_data_5[1903:1896];
        layer2[42][7:0] = buffer_data_4[1855:1848];
        layer2[42][15:8] = buffer_data_4[1863:1856];
        layer2[42][23:16] = buffer_data_4[1871:1864];
        layer2[42][31:24] = buffer_data_4[1879:1872];
        layer2[42][39:32] = buffer_data_4[1887:1880];
        layer2[42][47:40] = buffer_data_4[1895:1888];
        layer2[42][55:48] = buffer_data_4[1903:1896];
        layer3[42][7:0] = buffer_data_3[1855:1848];
        layer3[42][15:8] = buffer_data_3[1863:1856];
        layer3[42][23:16] = buffer_data_3[1871:1864];
        layer3[42][31:24] = buffer_data_3[1879:1872];
        layer3[42][39:32] = buffer_data_3[1887:1880];
        layer3[42][47:40] = buffer_data_3[1895:1888];
        layer3[42][55:48] = buffer_data_3[1903:1896];
        layer4[42][7:0] = buffer_data_2[1855:1848];
        layer4[42][15:8] = buffer_data_2[1863:1856];
        layer4[42][23:16] = buffer_data_2[1871:1864];
        layer4[42][31:24] = buffer_data_2[1879:1872];
        layer4[42][39:32] = buffer_data_2[1887:1880];
        layer4[42][47:40] = buffer_data_2[1895:1888];
        layer4[42][55:48] = buffer_data_2[1903:1896];
        layer5[42][7:0] = buffer_data_1[1855:1848];
        layer5[42][15:8] = buffer_data_1[1863:1856];
        layer5[42][23:16] = buffer_data_1[1871:1864];
        layer5[42][31:24] = buffer_data_1[1879:1872];
        layer5[42][39:32] = buffer_data_1[1887:1880];
        layer5[42][47:40] = buffer_data_1[1895:1888];
        layer5[42][55:48] = buffer_data_1[1903:1896];
        layer6[42][7:0] = buffer_data_0[1855:1848];
        layer6[42][15:8] = buffer_data_0[1863:1856];
        layer6[42][23:16] = buffer_data_0[1871:1864];
        layer6[42][31:24] = buffer_data_0[1879:1872];
        layer6[42][39:32] = buffer_data_0[1887:1880];
        layer6[42][47:40] = buffer_data_0[1895:1888];
        layer6[42][55:48] = buffer_data_0[1903:1896];
        layer0[43][7:0] = buffer_data_6[1863:1856];
        layer0[43][15:8] = buffer_data_6[1871:1864];
        layer0[43][23:16] = buffer_data_6[1879:1872];
        layer0[43][31:24] = buffer_data_6[1887:1880];
        layer0[43][39:32] = buffer_data_6[1895:1888];
        layer0[43][47:40] = buffer_data_6[1903:1896];
        layer0[43][55:48] = buffer_data_6[1911:1904];
        layer1[43][7:0] = buffer_data_5[1863:1856];
        layer1[43][15:8] = buffer_data_5[1871:1864];
        layer1[43][23:16] = buffer_data_5[1879:1872];
        layer1[43][31:24] = buffer_data_5[1887:1880];
        layer1[43][39:32] = buffer_data_5[1895:1888];
        layer1[43][47:40] = buffer_data_5[1903:1896];
        layer1[43][55:48] = buffer_data_5[1911:1904];
        layer2[43][7:0] = buffer_data_4[1863:1856];
        layer2[43][15:8] = buffer_data_4[1871:1864];
        layer2[43][23:16] = buffer_data_4[1879:1872];
        layer2[43][31:24] = buffer_data_4[1887:1880];
        layer2[43][39:32] = buffer_data_4[1895:1888];
        layer2[43][47:40] = buffer_data_4[1903:1896];
        layer2[43][55:48] = buffer_data_4[1911:1904];
        layer3[43][7:0] = buffer_data_3[1863:1856];
        layer3[43][15:8] = buffer_data_3[1871:1864];
        layer3[43][23:16] = buffer_data_3[1879:1872];
        layer3[43][31:24] = buffer_data_3[1887:1880];
        layer3[43][39:32] = buffer_data_3[1895:1888];
        layer3[43][47:40] = buffer_data_3[1903:1896];
        layer3[43][55:48] = buffer_data_3[1911:1904];
        layer4[43][7:0] = buffer_data_2[1863:1856];
        layer4[43][15:8] = buffer_data_2[1871:1864];
        layer4[43][23:16] = buffer_data_2[1879:1872];
        layer4[43][31:24] = buffer_data_2[1887:1880];
        layer4[43][39:32] = buffer_data_2[1895:1888];
        layer4[43][47:40] = buffer_data_2[1903:1896];
        layer4[43][55:48] = buffer_data_2[1911:1904];
        layer5[43][7:0] = buffer_data_1[1863:1856];
        layer5[43][15:8] = buffer_data_1[1871:1864];
        layer5[43][23:16] = buffer_data_1[1879:1872];
        layer5[43][31:24] = buffer_data_1[1887:1880];
        layer5[43][39:32] = buffer_data_1[1895:1888];
        layer5[43][47:40] = buffer_data_1[1903:1896];
        layer5[43][55:48] = buffer_data_1[1911:1904];
        layer6[43][7:0] = buffer_data_0[1863:1856];
        layer6[43][15:8] = buffer_data_0[1871:1864];
        layer6[43][23:16] = buffer_data_0[1879:1872];
        layer6[43][31:24] = buffer_data_0[1887:1880];
        layer6[43][39:32] = buffer_data_0[1895:1888];
        layer6[43][47:40] = buffer_data_0[1903:1896];
        layer6[43][55:48] = buffer_data_0[1911:1904];
        layer0[44][7:0] = buffer_data_6[1871:1864];
        layer0[44][15:8] = buffer_data_6[1879:1872];
        layer0[44][23:16] = buffer_data_6[1887:1880];
        layer0[44][31:24] = buffer_data_6[1895:1888];
        layer0[44][39:32] = buffer_data_6[1903:1896];
        layer0[44][47:40] = buffer_data_6[1911:1904];
        layer0[44][55:48] = buffer_data_6[1919:1912];
        layer1[44][7:0] = buffer_data_5[1871:1864];
        layer1[44][15:8] = buffer_data_5[1879:1872];
        layer1[44][23:16] = buffer_data_5[1887:1880];
        layer1[44][31:24] = buffer_data_5[1895:1888];
        layer1[44][39:32] = buffer_data_5[1903:1896];
        layer1[44][47:40] = buffer_data_5[1911:1904];
        layer1[44][55:48] = buffer_data_5[1919:1912];
        layer2[44][7:0] = buffer_data_4[1871:1864];
        layer2[44][15:8] = buffer_data_4[1879:1872];
        layer2[44][23:16] = buffer_data_4[1887:1880];
        layer2[44][31:24] = buffer_data_4[1895:1888];
        layer2[44][39:32] = buffer_data_4[1903:1896];
        layer2[44][47:40] = buffer_data_4[1911:1904];
        layer2[44][55:48] = buffer_data_4[1919:1912];
        layer3[44][7:0] = buffer_data_3[1871:1864];
        layer3[44][15:8] = buffer_data_3[1879:1872];
        layer3[44][23:16] = buffer_data_3[1887:1880];
        layer3[44][31:24] = buffer_data_3[1895:1888];
        layer3[44][39:32] = buffer_data_3[1903:1896];
        layer3[44][47:40] = buffer_data_3[1911:1904];
        layer3[44][55:48] = buffer_data_3[1919:1912];
        layer4[44][7:0] = buffer_data_2[1871:1864];
        layer4[44][15:8] = buffer_data_2[1879:1872];
        layer4[44][23:16] = buffer_data_2[1887:1880];
        layer4[44][31:24] = buffer_data_2[1895:1888];
        layer4[44][39:32] = buffer_data_2[1903:1896];
        layer4[44][47:40] = buffer_data_2[1911:1904];
        layer4[44][55:48] = buffer_data_2[1919:1912];
        layer5[44][7:0] = buffer_data_1[1871:1864];
        layer5[44][15:8] = buffer_data_1[1879:1872];
        layer5[44][23:16] = buffer_data_1[1887:1880];
        layer5[44][31:24] = buffer_data_1[1895:1888];
        layer5[44][39:32] = buffer_data_1[1903:1896];
        layer5[44][47:40] = buffer_data_1[1911:1904];
        layer5[44][55:48] = buffer_data_1[1919:1912];
        layer6[44][7:0] = buffer_data_0[1871:1864];
        layer6[44][15:8] = buffer_data_0[1879:1872];
        layer6[44][23:16] = buffer_data_0[1887:1880];
        layer6[44][31:24] = buffer_data_0[1895:1888];
        layer6[44][39:32] = buffer_data_0[1903:1896];
        layer6[44][47:40] = buffer_data_0[1911:1904];
        layer6[44][55:48] = buffer_data_0[1919:1912];
        layer0[45][7:0] = buffer_data_6[1879:1872];
        layer0[45][15:8] = buffer_data_6[1887:1880];
        layer0[45][23:16] = buffer_data_6[1895:1888];
        layer0[45][31:24] = buffer_data_6[1903:1896];
        layer0[45][39:32] = buffer_data_6[1911:1904];
        layer0[45][47:40] = buffer_data_6[1919:1912];
        layer0[45][55:48] = buffer_data_6[1927:1920];
        layer1[45][7:0] = buffer_data_5[1879:1872];
        layer1[45][15:8] = buffer_data_5[1887:1880];
        layer1[45][23:16] = buffer_data_5[1895:1888];
        layer1[45][31:24] = buffer_data_5[1903:1896];
        layer1[45][39:32] = buffer_data_5[1911:1904];
        layer1[45][47:40] = buffer_data_5[1919:1912];
        layer1[45][55:48] = buffer_data_5[1927:1920];
        layer2[45][7:0] = buffer_data_4[1879:1872];
        layer2[45][15:8] = buffer_data_4[1887:1880];
        layer2[45][23:16] = buffer_data_4[1895:1888];
        layer2[45][31:24] = buffer_data_4[1903:1896];
        layer2[45][39:32] = buffer_data_4[1911:1904];
        layer2[45][47:40] = buffer_data_4[1919:1912];
        layer2[45][55:48] = buffer_data_4[1927:1920];
        layer3[45][7:0] = buffer_data_3[1879:1872];
        layer3[45][15:8] = buffer_data_3[1887:1880];
        layer3[45][23:16] = buffer_data_3[1895:1888];
        layer3[45][31:24] = buffer_data_3[1903:1896];
        layer3[45][39:32] = buffer_data_3[1911:1904];
        layer3[45][47:40] = buffer_data_3[1919:1912];
        layer3[45][55:48] = buffer_data_3[1927:1920];
        layer4[45][7:0] = buffer_data_2[1879:1872];
        layer4[45][15:8] = buffer_data_2[1887:1880];
        layer4[45][23:16] = buffer_data_2[1895:1888];
        layer4[45][31:24] = buffer_data_2[1903:1896];
        layer4[45][39:32] = buffer_data_2[1911:1904];
        layer4[45][47:40] = buffer_data_2[1919:1912];
        layer4[45][55:48] = buffer_data_2[1927:1920];
        layer5[45][7:0] = buffer_data_1[1879:1872];
        layer5[45][15:8] = buffer_data_1[1887:1880];
        layer5[45][23:16] = buffer_data_1[1895:1888];
        layer5[45][31:24] = buffer_data_1[1903:1896];
        layer5[45][39:32] = buffer_data_1[1911:1904];
        layer5[45][47:40] = buffer_data_1[1919:1912];
        layer5[45][55:48] = buffer_data_1[1927:1920];
        layer6[45][7:0] = buffer_data_0[1879:1872];
        layer6[45][15:8] = buffer_data_0[1887:1880];
        layer6[45][23:16] = buffer_data_0[1895:1888];
        layer6[45][31:24] = buffer_data_0[1903:1896];
        layer6[45][39:32] = buffer_data_0[1911:1904];
        layer6[45][47:40] = buffer_data_0[1919:1912];
        layer6[45][55:48] = buffer_data_0[1927:1920];
        layer0[46][7:0] = buffer_data_6[1887:1880];
        layer0[46][15:8] = buffer_data_6[1895:1888];
        layer0[46][23:16] = buffer_data_6[1903:1896];
        layer0[46][31:24] = buffer_data_6[1911:1904];
        layer0[46][39:32] = buffer_data_6[1919:1912];
        layer0[46][47:40] = buffer_data_6[1927:1920];
        layer0[46][55:48] = buffer_data_6[1935:1928];
        layer1[46][7:0] = buffer_data_5[1887:1880];
        layer1[46][15:8] = buffer_data_5[1895:1888];
        layer1[46][23:16] = buffer_data_5[1903:1896];
        layer1[46][31:24] = buffer_data_5[1911:1904];
        layer1[46][39:32] = buffer_data_5[1919:1912];
        layer1[46][47:40] = buffer_data_5[1927:1920];
        layer1[46][55:48] = buffer_data_5[1935:1928];
        layer2[46][7:0] = buffer_data_4[1887:1880];
        layer2[46][15:8] = buffer_data_4[1895:1888];
        layer2[46][23:16] = buffer_data_4[1903:1896];
        layer2[46][31:24] = buffer_data_4[1911:1904];
        layer2[46][39:32] = buffer_data_4[1919:1912];
        layer2[46][47:40] = buffer_data_4[1927:1920];
        layer2[46][55:48] = buffer_data_4[1935:1928];
        layer3[46][7:0] = buffer_data_3[1887:1880];
        layer3[46][15:8] = buffer_data_3[1895:1888];
        layer3[46][23:16] = buffer_data_3[1903:1896];
        layer3[46][31:24] = buffer_data_3[1911:1904];
        layer3[46][39:32] = buffer_data_3[1919:1912];
        layer3[46][47:40] = buffer_data_3[1927:1920];
        layer3[46][55:48] = buffer_data_3[1935:1928];
        layer4[46][7:0] = buffer_data_2[1887:1880];
        layer4[46][15:8] = buffer_data_2[1895:1888];
        layer4[46][23:16] = buffer_data_2[1903:1896];
        layer4[46][31:24] = buffer_data_2[1911:1904];
        layer4[46][39:32] = buffer_data_2[1919:1912];
        layer4[46][47:40] = buffer_data_2[1927:1920];
        layer4[46][55:48] = buffer_data_2[1935:1928];
        layer5[46][7:0] = buffer_data_1[1887:1880];
        layer5[46][15:8] = buffer_data_1[1895:1888];
        layer5[46][23:16] = buffer_data_1[1903:1896];
        layer5[46][31:24] = buffer_data_1[1911:1904];
        layer5[46][39:32] = buffer_data_1[1919:1912];
        layer5[46][47:40] = buffer_data_1[1927:1920];
        layer5[46][55:48] = buffer_data_1[1935:1928];
        layer6[46][7:0] = buffer_data_0[1887:1880];
        layer6[46][15:8] = buffer_data_0[1895:1888];
        layer6[46][23:16] = buffer_data_0[1903:1896];
        layer6[46][31:24] = buffer_data_0[1911:1904];
        layer6[46][39:32] = buffer_data_0[1919:1912];
        layer6[46][47:40] = buffer_data_0[1927:1920];
        layer6[46][55:48] = buffer_data_0[1935:1928];
        layer0[47][7:0] = buffer_data_6[1895:1888];
        layer0[47][15:8] = buffer_data_6[1903:1896];
        layer0[47][23:16] = buffer_data_6[1911:1904];
        layer0[47][31:24] = buffer_data_6[1919:1912];
        layer0[47][39:32] = buffer_data_6[1927:1920];
        layer0[47][47:40] = buffer_data_6[1935:1928];
        layer0[47][55:48] = buffer_data_6[1943:1936];
        layer1[47][7:0] = buffer_data_5[1895:1888];
        layer1[47][15:8] = buffer_data_5[1903:1896];
        layer1[47][23:16] = buffer_data_5[1911:1904];
        layer1[47][31:24] = buffer_data_5[1919:1912];
        layer1[47][39:32] = buffer_data_5[1927:1920];
        layer1[47][47:40] = buffer_data_5[1935:1928];
        layer1[47][55:48] = buffer_data_5[1943:1936];
        layer2[47][7:0] = buffer_data_4[1895:1888];
        layer2[47][15:8] = buffer_data_4[1903:1896];
        layer2[47][23:16] = buffer_data_4[1911:1904];
        layer2[47][31:24] = buffer_data_4[1919:1912];
        layer2[47][39:32] = buffer_data_4[1927:1920];
        layer2[47][47:40] = buffer_data_4[1935:1928];
        layer2[47][55:48] = buffer_data_4[1943:1936];
        layer3[47][7:0] = buffer_data_3[1895:1888];
        layer3[47][15:8] = buffer_data_3[1903:1896];
        layer3[47][23:16] = buffer_data_3[1911:1904];
        layer3[47][31:24] = buffer_data_3[1919:1912];
        layer3[47][39:32] = buffer_data_3[1927:1920];
        layer3[47][47:40] = buffer_data_3[1935:1928];
        layer3[47][55:48] = buffer_data_3[1943:1936];
        layer4[47][7:0] = buffer_data_2[1895:1888];
        layer4[47][15:8] = buffer_data_2[1903:1896];
        layer4[47][23:16] = buffer_data_2[1911:1904];
        layer4[47][31:24] = buffer_data_2[1919:1912];
        layer4[47][39:32] = buffer_data_2[1927:1920];
        layer4[47][47:40] = buffer_data_2[1935:1928];
        layer4[47][55:48] = buffer_data_2[1943:1936];
        layer5[47][7:0] = buffer_data_1[1895:1888];
        layer5[47][15:8] = buffer_data_1[1903:1896];
        layer5[47][23:16] = buffer_data_1[1911:1904];
        layer5[47][31:24] = buffer_data_1[1919:1912];
        layer5[47][39:32] = buffer_data_1[1927:1920];
        layer5[47][47:40] = buffer_data_1[1935:1928];
        layer5[47][55:48] = buffer_data_1[1943:1936];
        layer6[47][7:0] = buffer_data_0[1895:1888];
        layer6[47][15:8] = buffer_data_0[1903:1896];
        layer6[47][23:16] = buffer_data_0[1911:1904];
        layer6[47][31:24] = buffer_data_0[1919:1912];
        layer6[47][39:32] = buffer_data_0[1927:1920];
        layer6[47][47:40] = buffer_data_0[1935:1928];
        layer6[47][55:48] = buffer_data_0[1943:1936];
        layer0[48][7:0] = buffer_data_6[1903:1896];
        layer0[48][15:8] = buffer_data_6[1911:1904];
        layer0[48][23:16] = buffer_data_6[1919:1912];
        layer0[48][31:24] = buffer_data_6[1927:1920];
        layer0[48][39:32] = buffer_data_6[1935:1928];
        layer0[48][47:40] = buffer_data_6[1943:1936];
        layer0[48][55:48] = buffer_data_6[1951:1944];
        layer1[48][7:0] = buffer_data_5[1903:1896];
        layer1[48][15:8] = buffer_data_5[1911:1904];
        layer1[48][23:16] = buffer_data_5[1919:1912];
        layer1[48][31:24] = buffer_data_5[1927:1920];
        layer1[48][39:32] = buffer_data_5[1935:1928];
        layer1[48][47:40] = buffer_data_5[1943:1936];
        layer1[48][55:48] = buffer_data_5[1951:1944];
        layer2[48][7:0] = buffer_data_4[1903:1896];
        layer2[48][15:8] = buffer_data_4[1911:1904];
        layer2[48][23:16] = buffer_data_4[1919:1912];
        layer2[48][31:24] = buffer_data_4[1927:1920];
        layer2[48][39:32] = buffer_data_4[1935:1928];
        layer2[48][47:40] = buffer_data_4[1943:1936];
        layer2[48][55:48] = buffer_data_4[1951:1944];
        layer3[48][7:0] = buffer_data_3[1903:1896];
        layer3[48][15:8] = buffer_data_3[1911:1904];
        layer3[48][23:16] = buffer_data_3[1919:1912];
        layer3[48][31:24] = buffer_data_3[1927:1920];
        layer3[48][39:32] = buffer_data_3[1935:1928];
        layer3[48][47:40] = buffer_data_3[1943:1936];
        layer3[48][55:48] = buffer_data_3[1951:1944];
        layer4[48][7:0] = buffer_data_2[1903:1896];
        layer4[48][15:8] = buffer_data_2[1911:1904];
        layer4[48][23:16] = buffer_data_2[1919:1912];
        layer4[48][31:24] = buffer_data_2[1927:1920];
        layer4[48][39:32] = buffer_data_2[1935:1928];
        layer4[48][47:40] = buffer_data_2[1943:1936];
        layer4[48][55:48] = buffer_data_2[1951:1944];
        layer5[48][7:0] = buffer_data_1[1903:1896];
        layer5[48][15:8] = buffer_data_1[1911:1904];
        layer5[48][23:16] = buffer_data_1[1919:1912];
        layer5[48][31:24] = buffer_data_1[1927:1920];
        layer5[48][39:32] = buffer_data_1[1935:1928];
        layer5[48][47:40] = buffer_data_1[1943:1936];
        layer5[48][55:48] = buffer_data_1[1951:1944];
        layer6[48][7:0] = buffer_data_0[1903:1896];
        layer6[48][15:8] = buffer_data_0[1911:1904];
        layer6[48][23:16] = buffer_data_0[1919:1912];
        layer6[48][31:24] = buffer_data_0[1927:1920];
        layer6[48][39:32] = buffer_data_0[1935:1928];
        layer6[48][47:40] = buffer_data_0[1943:1936];
        layer6[48][55:48] = buffer_data_0[1951:1944];
        layer0[49][7:0] = buffer_data_6[1911:1904];
        layer0[49][15:8] = buffer_data_6[1919:1912];
        layer0[49][23:16] = buffer_data_6[1927:1920];
        layer0[49][31:24] = buffer_data_6[1935:1928];
        layer0[49][39:32] = buffer_data_6[1943:1936];
        layer0[49][47:40] = buffer_data_6[1951:1944];
        layer0[49][55:48] = buffer_data_6[1959:1952];
        layer1[49][7:0] = buffer_data_5[1911:1904];
        layer1[49][15:8] = buffer_data_5[1919:1912];
        layer1[49][23:16] = buffer_data_5[1927:1920];
        layer1[49][31:24] = buffer_data_5[1935:1928];
        layer1[49][39:32] = buffer_data_5[1943:1936];
        layer1[49][47:40] = buffer_data_5[1951:1944];
        layer1[49][55:48] = buffer_data_5[1959:1952];
        layer2[49][7:0] = buffer_data_4[1911:1904];
        layer2[49][15:8] = buffer_data_4[1919:1912];
        layer2[49][23:16] = buffer_data_4[1927:1920];
        layer2[49][31:24] = buffer_data_4[1935:1928];
        layer2[49][39:32] = buffer_data_4[1943:1936];
        layer2[49][47:40] = buffer_data_4[1951:1944];
        layer2[49][55:48] = buffer_data_4[1959:1952];
        layer3[49][7:0] = buffer_data_3[1911:1904];
        layer3[49][15:8] = buffer_data_3[1919:1912];
        layer3[49][23:16] = buffer_data_3[1927:1920];
        layer3[49][31:24] = buffer_data_3[1935:1928];
        layer3[49][39:32] = buffer_data_3[1943:1936];
        layer3[49][47:40] = buffer_data_3[1951:1944];
        layer3[49][55:48] = buffer_data_3[1959:1952];
        layer4[49][7:0] = buffer_data_2[1911:1904];
        layer4[49][15:8] = buffer_data_2[1919:1912];
        layer4[49][23:16] = buffer_data_2[1927:1920];
        layer4[49][31:24] = buffer_data_2[1935:1928];
        layer4[49][39:32] = buffer_data_2[1943:1936];
        layer4[49][47:40] = buffer_data_2[1951:1944];
        layer4[49][55:48] = buffer_data_2[1959:1952];
        layer5[49][7:0] = buffer_data_1[1911:1904];
        layer5[49][15:8] = buffer_data_1[1919:1912];
        layer5[49][23:16] = buffer_data_1[1927:1920];
        layer5[49][31:24] = buffer_data_1[1935:1928];
        layer5[49][39:32] = buffer_data_1[1943:1936];
        layer5[49][47:40] = buffer_data_1[1951:1944];
        layer5[49][55:48] = buffer_data_1[1959:1952];
        layer6[49][7:0] = buffer_data_0[1911:1904];
        layer6[49][15:8] = buffer_data_0[1919:1912];
        layer6[49][23:16] = buffer_data_0[1927:1920];
        layer6[49][31:24] = buffer_data_0[1935:1928];
        layer6[49][39:32] = buffer_data_0[1943:1936];
        layer6[49][47:40] = buffer_data_0[1951:1944];
        layer6[49][55:48] = buffer_data_0[1959:1952];
        layer0[50][7:0] = buffer_data_6[1919:1912];
        layer0[50][15:8] = buffer_data_6[1927:1920];
        layer0[50][23:16] = buffer_data_6[1935:1928];
        layer0[50][31:24] = buffer_data_6[1943:1936];
        layer0[50][39:32] = buffer_data_6[1951:1944];
        layer0[50][47:40] = buffer_data_6[1959:1952];
        layer0[50][55:48] = buffer_data_6[1967:1960];
        layer1[50][7:0] = buffer_data_5[1919:1912];
        layer1[50][15:8] = buffer_data_5[1927:1920];
        layer1[50][23:16] = buffer_data_5[1935:1928];
        layer1[50][31:24] = buffer_data_5[1943:1936];
        layer1[50][39:32] = buffer_data_5[1951:1944];
        layer1[50][47:40] = buffer_data_5[1959:1952];
        layer1[50][55:48] = buffer_data_5[1967:1960];
        layer2[50][7:0] = buffer_data_4[1919:1912];
        layer2[50][15:8] = buffer_data_4[1927:1920];
        layer2[50][23:16] = buffer_data_4[1935:1928];
        layer2[50][31:24] = buffer_data_4[1943:1936];
        layer2[50][39:32] = buffer_data_4[1951:1944];
        layer2[50][47:40] = buffer_data_4[1959:1952];
        layer2[50][55:48] = buffer_data_4[1967:1960];
        layer3[50][7:0] = buffer_data_3[1919:1912];
        layer3[50][15:8] = buffer_data_3[1927:1920];
        layer3[50][23:16] = buffer_data_3[1935:1928];
        layer3[50][31:24] = buffer_data_3[1943:1936];
        layer3[50][39:32] = buffer_data_3[1951:1944];
        layer3[50][47:40] = buffer_data_3[1959:1952];
        layer3[50][55:48] = buffer_data_3[1967:1960];
        layer4[50][7:0] = buffer_data_2[1919:1912];
        layer4[50][15:8] = buffer_data_2[1927:1920];
        layer4[50][23:16] = buffer_data_2[1935:1928];
        layer4[50][31:24] = buffer_data_2[1943:1936];
        layer4[50][39:32] = buffer_data_2[1951:1944];
        layer4[50][47:40] = buffer_data_2[1959:1952];
        layer4[50][55:48] = buffer_data_2[1967:1960];
        layer5[50][7:0] = buffer_data_1[1919:1912];
        layer5[50][15:8] = buffer_data_1[1927:1920];
        layer5[50][23:16] = buffer_data_1[1935:1928];
        layer5[50][31:24] = buffer_data_1[1943:1936];
        layer5[50][39:32] = buffer_data_1[1951:1944];
        layer5[50][47:40] = buffer_data_1[1959:1952];
        layer5[50][55:48] = buffer_data_1[1967:1960];
        layer6[50][7:0] = buffer_data_0[1919:1912];
        layer6[50][15:8] = buffer_data_0[1927:1920];
        layer6[50][23:16] = buffer_data_0[1935:1928];
        layer6[50][31:24] = buffer_data_0[1943:1936];
        layer6[50][39:32] = buffer_data_0[1951:1944];
        layer6[50][47:40] = buffer_data_0[1959:1952];
        layer6[50][55:48] = buffer_data_0[1967:1960];
        layer0[51][7:0] = buffer_data_6[1927:1920];
        layer0[51][15:8] = buffer_data_6[1935:1928];
        layer0[51][23:16] = buffer_data_6[1943:1936];
        layer0[51][31:24] = buffer_data_6[1951:1944];
        layer0[51][39:32] = buffer_data_6[1959:1952];
        layer0[51][47:40] = buffer_data_6[1967:1960];
        layer0[51][55:48] = buffer_data_6[1975:1968];
        layer1[51][7:0] = buffer_data_5[1927:1920];
        layer1[51][15:8] = buffer_data_5[1935:1928];
        layer1[51][23:16] = buffer_data_5[1943:1936];
        layer1[51][31:24] = buffer_data_5[1951:1944];
        layer1[51][39:32] = buffer_data_5[1959:1952];
        layer1[51][47:40] = buffer_data_5[1967:1960];
        layer1[51][55:48] = buffer_data_5[1975:1968];
        layer2[51][7:0] = buffer_data_4[1927:1920];
        layer2[51][15:8] = buffer_data_4[1935:1928];
        layer2[51][23:16] = buffer_data_4[1943:1936];
        layer2[51][31:24] = buffer_data_4[1951:1944];
        layer2[51][39:32] = buffer_data_4[1959:1952];
        layer2[51][47:40] = buffer_data_4[1967:1960];
        layer2[51][55:48] = buffer_data_4[1975:1968];
        layer3[51][7:0] = buffer_data_3[1927:1920];
        layer3[51][15:8] = buffer_data_3[1935:1928];
        layer3[51][23:16] = buffer_data_3[1943:1936];
        layer3[51][31:24] = buffer_data_3[1951:1944];
        layer3[51][39:32] = buffer_data_3[1959:1952];
        layer3[51][47:40] = buffer_data_3[1967:1960];
        layer3[51][55:48] = buffer_data_3[1975:1968];
        layer4[51][7:0] = buffer_data_2[1927:1920];
        layer4[51][15:8] = buffer_data_2[1935:1928];
        layer4[51][23:16] = buffer_data_2[1943:1936];
        layer4[51][31:24] = buffer_data_2[1951:1944];
        layer4[51][39:32] = buffer_data_2[1959:1952];
        layer4[51][47:40] = buffer_data_2[1967:1960];
        layer4[51][55:48] = buffer_data_2[1975:1968];
        layer5[51][7:0] = buffer_data_1[1927:1920];
        layer5[51][15:8] = buffer_data_1[1935:1928];
        layer5[51][23:16] = buffer_data_1[1943:1936];
        layer5[51][31:24] = buffer_data_1[1951:1944];
        layer5[51][39:32] = buffer_data_1[1959:1952];
        layer5[51][47:40] = buffer_data_1[1967:1960];
        layer5[51][55:48] = buffer_data_1[1975:1968];
        layer6[51][7:0] = buffer_data_0[1927:1920];
        layer6[51][15:8] = buffer_data_0[1935:1928];
        layer6[51][23:16] = buffer_data_0[1943:1936];
        layer6[51][31:24] = buffer_data_0[1951:1944];
        layer6[51][39:32] = buffer_data_0[1959:1952];
        layer6[51][47:40] = buffer_data_0[1967:1960];
        layer6[51][55:48] = buffer_data_0[1975:1968];
        layer0[52][7:0] = buffer_data_6[1935:1928];
        layer0[52][15:8] = buffer_data_6[1943:1936];
        layer0[52][23:16] = buffer_data_6[1951:1944];
        layer0[52][31:24] = buffer_data_6[1959:1952];
        layer0[52][39:32] = buffer_data_6[1967:1960];
        layer0[52][47:40] = buffer_data_6[1975:1968];
        layer0[52][55:48] = buffer_data_6[1983:1976];
        layer1[52][7:0] = buffer_data_5[1935:1928];
        layer1[52][15:8] = buffer_data_5[1943:1936];
        layer1[52][23:16] = buffer_data_5[1951:1944];
        layer1[52][31:24] = buffer_data_5[1959:1952];
        layer1[52][39:32] = buffer_data_5[1967:1960];
        layer1[52][47:40] = buffer_data_5[1975:1968];
        layer1[52][55:48] = buffer_data_5[1983:1976];
        layer2[52][7:0] = buffer_data_4[1935:1928];
        layer2[52][15:8] = buffer_data_4[1943:1936];
        layer2[52][23:16] = buffer_data_4[1951:1944];
        layer2[52][31:24] = buffer_data_4[1959:1952];
        layer2[52][39:32] = buffer_data_4[1967:1960];
        layer2[52][47:40] = buffer_data_4[1975:1968];
        layer2[52][55:48] = buffer_data_4[1983:1976];
        layer3[52][7:0] = buffer_data_3[1935:1928];
        layer3[52][15:8] = buffer_data_3[1943:1936];
        layer3[52][23:16] = buffer_data_3[1951:1944];
        layer3[52][31:24] = buffer_data_3[1959:1952];
        layer3[52][39:32] = buffer_data_3[1967:1960];
        layer3[52][47:40] = buffer_data_3[1975:1968];
        layer3[52][55:48] = buffer_data_3[1983:1976];
        layer4[52][7:0] = buffer_data_2[1935:1928];
        layer4[52][15:8] = buffer_data_2[1943:1936];
        layer4[52][23:16] = buffer_data_2[1951:1944];
        layer4[52][31:24] = buffer_data_2[1959:1952];
        layer4[52][39:32] = buffer_data_2[1967:1960];
        layer4[52][47:40] = buffer_data_2[1975:1968];
        layer4[52][55:48] = buffer_data_2[1983:1976];
        layer5[52][7:0] = buffer_data_1[1935:1928];
        layer5[52][15:8] = buffer_data_1[1943:1936];
        layer5[52][23:16] = buffer_data_1[1951:1944];
        layer5[52][31:24] = buffer_data_1[1959:1952];
        layer5[52][39:32] = buffer_data_1[1967:1960];
        layer5[52][47:40] = buffer_data_1[1975:1968];
        layer5[52][55:48] = buffer_data_1[1983:1976];
        layer6[52][7:0] = buffer_data_0[1935:1928];
        layer6[52][15:8] = buffer_data_0[1943:1936];
        layer6[52][23:16] = buffer_data_0[1951:1944];
        layer6[52][31:24] = buffer_data_0[1959:1952];
        layer6[52][39:32] = buffer_data_0[1967:1960];
        layer6[52][47:40] = buffer_data_0[1975:1968];
        layer6[52][55:48] = buffer_data_0[1983:1976];
        layer0[53][7:0] = buffer_data_6[1943:1936];
        layer0[53][15:8] = buffer_data_6[1951:1944];
        layer0[53][23:16] = buffer_data_6[1959:1952];
        layer0[53][31:24] = buffer_data_6[1967:1960];
        layer0[53][39:32] = buffer_data_6[1975:1968];
        layer0[53][47:40] = buffer_data_6[1983:1976];
        layer0[53][55:48] = buffer_data_6[1991:1984];
        layer1[53][7:0] = buffer_data_5[1943:1936];
        layer1[53][15:8] = buffer_data_5[1951:1944];
        layer1[53][23:16] = buffer_data_5[1959:1952];
        layer1[53][31:24] = buffer_data_5[1967:1960];
        layer1[53][39:32] = buffer_data_5[1975:1968];
        layer1[53][47:40] = buffer_data_5[1983:1976];
        layer1[53][55:48] = buffer_data_5[1991:1984];
        layer2[53][7:0] = buffer_data_4[1943:1936];
        layer2[53][15:8] = buffer_data_4[1951:1944];
        layer2[53][23:16] = buffer_data_4[1959:1952];
        layer2[53][31:24] = buffer_data_4[1967:1960];
        layer2[53][39:32] = buffer_data_4[1975:1968];
        layer2[53][47:40] = buffer_data_4[1983:1976];
        layer2[53][55:48] = buffer_data_4[1991:1984];
        layer3[53][7:0] = buffer_data_3[1943:1936];
        layer3[53][15:8] = buffer_data_3[1951:1944];
        layer3[53][23:16] = buffer_data_3[1959:1952];
        layer3[53][31:24] = buffer_data_3[1967:1960];
        layer3[53][39:32] = buffer_data_3[1975:1968];
        layer3[53][47:40] = buffer_data_3[1983:1976];
        layer3[53][55:48] = buffer_data_3[1991:1984];
        layer4[53][7:0] = buffer_data_2[1943:1936];
        layer4[53][15:8] = buffer_data_2[1951:1944];
        layer4[53][23:16] = buffer_data_2[1959:1952];
        layer4[53][31:24] = buffer_data_2[1967:1960];
        layer4[53][39:32] = buffer_data_2[1975:1968];
        layer4[53][47:40] = buffer_data_2[1983:1976];
        layer4[53][55:48] = buffer_data_2[1991:1984];
        layer5[53][7:0] = buffer_data_1[1943:1936];
        layer5[53][15:8] = buffer_data_1[1951:1944];
        layer5[53][23:16] = buffer_data_1[1959:1952];
        layer5[53][31:24] = buffer_data_1[1967:1960];
        layer5[53][39:32] = buffer_data_1[1975:1968];
        layer5[53][47:40] = buffer_data_1[1983:1976];
        layer5[53][55:48] = buffer_data_1[1991:1984];
        layer6[53][7:0] = buffer_data_0[1943:1936];
        layer6[53][15:8] = buffer_data_0[1951:1944];
        layer6[53][23:16] = buffer_data_0[1959:1952];
        layer6[53][31:24] = buffer_data_0[1967:1960];
        layer6[53][39:32] = buffer_data_0[1975:1968];
        layer6[53][47:40] = buffer_data_0[1983:1976];
        layer6[53][55:48] = buffer_data_0[1991:1984];
        layer0[54][7:0] = buffer_data_6[1951:1944];
        layer0[54][15:8] = buffer_data_6[1959:1952];
        layer0[54][23:16] = buffer_data_6[1967:1960];
        layer0[54][31:24] = buffer_data_6[1975:1968];
        layer0[54][39:32] = buffer_data_6[1983:1976];
        layer0[54][47:40] = buffer_data_6[1991:1984];
        layer0[54][55:48] = buffer_data_6[1999:1992];
        layer1[54][7:0] = buffer_data_5[1951:1944];
        layer1[54][15:8] = buffer_data_5[1959:1952];
        layer1[54][23:16] = buffer_data_5[1967:1960];
        layer1[54][31:24] = buffer_data_5[1975:1968];
        layer1[54][39:32] = buffer_data_5[1983:1976];
        layer1[54][47:40] = buffer_data_5[1991:1984];
        layer1[54][55:48] = buffer_data_5[1999:1992];
        layer2[54][7:0] = buffer_data_4[1951:1944];
        layer2[54][15:8] = buffer_data_4[1959:1952];
        layer2[54][23:16] = buffer_data_4[1967:1960];
        layer2[54][31:24] = buffer_data_4[1975:1968];
        layer2[54][39:32] = buffer_data_4[1983:1976];
        layer2[54][47:40] = buffer_data_4[1991:1984];
        layer2[54][55:48] = buffer_data_4[1999:1992];
        layer3[54][7:0] = buffer_data_3[1951:1944];
        layer3[54][15:8] = buffer_data_3[1959:1952];
        layer3[54][23:16] = buffer_data_3[1967:1960];
        layer3[54][31:24] = buffer_data_3[1975:1968];
        layer3[54][39:32] = buffer_data_3[1983:1976];
        layer3[54][47:40] = buffer_data_3[1991:1984];
        layer3[54][55:48] = buffer_data_3[1999:1992];
        layer4[54][7:0] = buffer_data_2[1951:1944];
        layer4[54][15:8] = buffer_data_2[1959:1952];
        layer4[54][23:16] = buffer_data_2[1967:1960];
        layer4[54][31:24] = buffer_data_2[1975:1968];
        layer4[54][39:32] = buffer_data_2[1983:1976];
        layer4[54][47:40] = buffer_data_2[1991:1984];
        layer4[54][55:48] = buffer_data_2[1999:1992];
        layer5[54][7:0] = buffer_data_1[1951:1944];
        layer5[54][15:8] = buffer_data_1[1959:1952];
        layer5[54][23:16] = buffer_data_1[1967:1960];
        layer5[54][31:24] = buffer_data_1[1975:1968];
        layer5[54][39:32] = buffer_data_1[1983:1976];
        layer5[54][47:40] = buffer_data_1[1991:1984];
        layer5[54][55:48] = buffer_data_1[1999:1992];
        layer6[54][7:0] = buffer_data_0[1951:1944];
        layer6[54][15:8] = buffer_data_0[1959:1952];
        layer6[54][23:16] = buffer_data_0[1967:1960];
        layer6[54][31:24] = buffer_data_0[1975:1968];
        layer6[54][39:32] = buffer_data_0[1983:1976];
        layer6[54][47:40] = buffer_data_0[1991:1984];
        layer6[54][55:48] = buffer_data_0[1999:1992];
        layer0[55][7:0] = buffer_data_6[1959:1952];
        layer0[55][15:8] = buffer_data_6[1967:1960];
        layer0[55][23:16] = buffer_data_6[1975:1968];
        layer0[55][31:24] = buffer_data_6[1983:1976];
        layer0[55][39:32] = buffer_data_6[1991:1984];
        layer0[55][47:40] = buffer_data_6[1999:1992];
        layer0[55][55:48] = buffer_data_6[2007:2000];
        layer1[55][7:0] = buffer_data_5[1959:1952];
        layer1[55][15:8] = buffer_data_5[1967:1960];
        layer1[55][23:16] = buffer_data_5[1975:1968];
        layer1[55][31:24] = buffer_data_5[1983:1976];
        layer1[55][39:32] = buffer_data_5[1991:1984];
        layer1[55][47:40] = buffer_data_5[1999:1992];
        layer1[55][55:48] = buffer_data_5[2007:2000];
        layer2[55][7:0] = buffer_data_4[1959:1952];
        layer2[55][15:8] = buffer_data_4[1967:1960];
        layer2[55][23:16] = buffer_data_4[1975:1968];
        layer2[55][31:24] = buffer_data_4[1983:1976];
        layer2[55][39:32] = buffer_data_4[1991:1984];
        layer2[55][47:40] = buffer_data_4[1999:1992];
        layer2[55][55:48] = buffer_data_4[2007:2000];
        layer3[55][7:0] = buffer_data_3[1959:1952];
        layer3[55][15:8] = buffer_data_3[1967:1960];
        layer3[55][23:16] = buffer_data_3[1975:1968];
        layer3[55][31:24] = buffer_data_3[1983:1976];
        layer3[55][39:32] = buffer_data_3[1991:1984];
        layer3[55][47:40] = buffer_data_3[1999:1992];
        layer3[55][55:48] = buffer_data_3[2007:2000];
        layer4[55][7:0] = buffer_data_2[1959:1952];
        layer4[55][15:8] = buffer_data_2[1967:1960];
        layer4[55][23:16] = buffer_data_2[1975:1968];
        layer4[55][31:24] = buffer_data_2[1983:1976];
        layer4[55][39:32] = buffer_data_2[1991:1984];
        layer4[55][47:40] = buffer_data_2[1999:1992];
        layer4[55][55:48] = buffer_data_2[2007:2000];
        layer5[55][7:0] = buffer_data_1[1959:1952];
        layer5[55][15:8] = buffer_data_1[1967:1960];
        layer5[55][23:16] = buffer_data_1[1975:1968];
        layer5[55][31:24] = buffer_data_1[1983:1976];
        layer5[55][39:32] = buffer_data_1[1991:1984];
        layer5[55][47:40] = buffer_data_1[1999:1992];
        layer5[55][55:48] = buffer_data_1[2007:2000];
        layer6[55][7:0] = buffer_data_0[1959:1952];
        layer6[55][15:8] = buffer_data_0[1967:1960];
        layer6[55][23:16] = buffer_data_0[1975:1968];
        layer6[55][31:24] = buffer_data_0[1983:1976];
        layer6[55][39:32] = buffer_data_0[1991:1984];
        layer6[55][47:40] = buffer_data_0[1999:1992];
        layer6[55][55:48] = buffer_data_0[2007:2000];
        layer0[56][7:0] = buffer_data_6[1967:1960];
        layer0[56][15:8] = buffer_data_6[1975:1968];
        layer0[56][23:16] = buffer_data_6[1983:1976];
        layer0[56][31:24] = buffer_data_6[1991:1984];
        layer0[56][39:32] = buffer_data_6[1999:1992];
        layer0[56][47:40] = buffer_data_6[2007:2000];
        layer0[56][55:48] = buffer_data_6[2015:2008];
        layer1[56][7:0] = buffer_data_5[1967:1960];
        layer1[56][15:8] = buffer_data_5[1975:1968];
        layer1[56][23:16] = buffer_data_5[1983:1976];
        layer1[56][31:24] = buffer_data_5[1991:1984];
        layer1[56][39:32] = buffer_data_5[1999:1992];
        layer1[56][47:40] = buffer_data_5[2007:2000];
        layer1[56][55:48] = buffer_data_5[2015:2008];
        layer2[56][7:0] = buffer_data_4[1967:1960];
        layer2[56][15:8] = buffer_data_4[1975:1968];
        layer2[56][23:16] = buffer_data_4[1983:1976];
        layer2[56][31:24] = buffer_data_4[1991:1984];
        layer2[56][39:32] = buffer_data_4[1999:1992];
        layer2[56][47:40] = buffer_data_4[2007:2000];
        layer2[56][55:48] = buffer_data_4[2015:2008];
        layer3[56][7:0] = buffer_data_3[1967:1960];
        layer3[56][15:8] = buffer_data_3[1975:1968];
        layer3[56][23:16] = buffer_data_3[1983:1976];
        layer3[56][31:24] = buffer_data_3[1991:1984];
        layer3[56][39:32] = buffer_data_3[1999:1992];
        layer3[56][47:40] = buffer_data_3[2007:2000];
        layer3[56][55:48] = buffer_data_3[2015:2008];
        layer4[56][7:0] = buffer_data_2[1967:1960];
        layer4[56][15:8] = buffer_data_2[1975:1968];
        layer4[56][23:16] = buffer_data_2[1983:1976];
        layer4[56][31:24] = buffer_data_2[1991:1984];
        layer4[56][39:32] = buffer_data_2[1999:1992];
        layer4[56][47:40] = buffer_data_2[2007:2000];
        layer4[56][55:48] = buffer_data_2[2015:2008];
        layer5[56][7:0] = buffer_data_1[1967:1960];
        layer5[56][15:8] = buffer_data_1[1975:1968];
        layer5[56][23:16] = buffer_data_1[1983:1976];
        layer5[56][31:24] = buffer_data_1[1991:1984];
        layer5[56][39:32] = buffer_data_1[1999:1992];
        layer5[56][47:40] = buffer_data_1[2007:2000];
        layer5[56][55:48] = buffer_data_1[2015:2008];
        layer6[56][7:0] = buffer_data_0[1967:1960];
        layer6[56][15:8] = buffer_data_0[1975:1968];
        layer6[56][23:16] = buffer_data_0[1983:1976];
        layer6[56][31:24] = buffer_data_0[1991:1984];
        layer6[56][39:32] = buffer_data_0[1999:1992];
        layer6[56][47:40] = buffer_data_0[2007:2000];
        layer6[56][55:48] = buffer_data_0[2015:2008];
        layer0[57][7:0] = buffer_data_6[1975:1968];
        layer0[57][15:8] = buffer_data_6[1983:1976];
        layer0[57][23:16] = buffer_data_6[1991:1984];
        layer0[57][31:24] = buffer_data_6[1999:1992];
        layer0[57][39:32] = buffer_data_6[2007:2000];
        layer0[57][47:40] = buffer_data_6[2015:2008];
        layer0[57][55:48] = buffer_data_6[2023:2016];
        layer1[57][7:0] = buffer_data_5[1975:1968];
        layer1[57][15:8] = buffer_data_5[1983:1976];
        layer1[57][23:16] = buffer_data_5[1991:1984];
        layer1[57][31:24] = buffer_data_5[1999:1992];
        layer1[57][39:32] = buffer_data_5[2007:2000];
        layer1[57][47:40] = buffer_data_5[2015:2008];
        layer1[57][55:48] = buffer_data_5[2023:2016];
        layer2[57][7:0] = buffer_data_4[1975:1968];
        layer2[57][15:8] = buffer_data_4[1983:1976];
        layer2[57][23:16] = buffer_data_4[1991:1984];
        layer2[57][31:24] = buffer_data_4[1999:1992];
        layer2[57][39:32] = buffer_data_4[2007:2000];
        layer2[57][47:40] = buffer_data_4[2015:2008];
        layer2[57][55:48] = buffer_data_4[2023:2016];
        layer3[57][7:0] = buffer_data_3[1975:1968];
        layer3[57][15:8] = buffer_data_3[1983:1976];
        layer3[57][23:16] = buffer_data_3[1991:1984];
        layer3[57][31:24] = buffer_data_3[1999:1992];
        layer3[57][39:32] = buffer_data_3[2007:2000];
        layer3[57][47:40] = buffer_data_3[2015:2008];
        layer3[57][55:48] = buffer_data_3[2023:2016];
        layer4[57][7:0] = buffer_data_2[1975:1968];
        layer4[57][15:8] = buffer_data_2[1983:1976];
        layer4[57][23:16] = buffer_data_2[1991:1984];
        layer4[57][31:24] = buffer_data_2[1999:1992];
        layer4[57][39:32] = buffer_data_2[2007:2000];
        layer4[57][47:40] = buffer_data_2[2015:2008];
        layer4[57][55:48] = buffer_data_2[2023:2016];
        layer5[57][7:0] = buffer_data_1[1975:1968];
        layer5[57][15:8] = buffer_data_1[1983:1976];
        layer5[57][23:16] = buffer_data_1[1991:1984];
        layer5[57][31:24] = buffer_data_1[1999:1992];
        layer5[57][39:32] = buffer_data_1[2007:2000];
        layer5[57][47:40] = buffer_data_1[2015:2008];
        layer5[57][55:48] = buffer_data_1[2023:2016];
        layer6[57][7:0] = buffer_data_0[1975:1968];
        layer6[57][15:8] = buffer_data_0[1983:1976];
        layer6[57][23:16] = buffer_data_0[1991:1984];
        layer6[57][31:24] = buffer_data_0[1999:1992];
        layer6[57][39:32] = buffer_data_0[2007:2000];
        layer6[57][47:40] = buffer_data_0[2015:2008];
        layer6[57][55:48] = buffer_data_0[2023:2016];
        layer0[58][7:0] = buffer_data_6[1983:1976];
        layer0[58][15:8] = buffer_data_6[1991:1984];
        layer0[58][23:16] = buffer_data_6[1999:1992];
        layer0[58][31:24] = buffer_data_6[2007:2000];
        layer0[58][39:32] = buffer_data_6[2015:2008];
        layer0[58][47:40] = buffer_data_6[2023:2016];
        layer0[58][55:48] = buffer_data_6[2031:2024];
        layer1[58][7:0] = buffer_data_5[1983:1976];
        layer1[58][15:8] = buffer_data_5[1991:1984];
        layer1[58][23:16] = buffer_data_5[1999:1992];
        layer1[58][31:24] = buffer_data_5[2007:2000];
        layer1[58][39:32] = buffer_data_5[2015:2008];
        layer1[58][47:40] = buffer_data_5[2023:2016];
        layer1[58][55:48] = buffer_data_5[2031:2024];
        layer2[58][7:0] = buffer_data_4[1983:1976];
        layer2[58][15:8] = buffer_data_4[1991:1984];
        layer2[58][23:16] = buffer_data_4[1999:1992];
        layer2[58][31:24] = buffer_data_4[2007:2000];
        layer2[58][39:32] = buffer_data_4[2015:2008];
        layer2[58][47:40] = buffer_data_4[2023:2016];
        layer2[58][55:48] = buffer_data_4[2031:2024];
        layer3[58][7:0] = buffer_data_3[1983:1976];
        layer3[58][15:8] = buffer_data_3[1991:1984];
        layer3[58][23:16] = buffer_data_3[1999:1992];
        layer3[58][31:24] = buffer_data_3[2007:2000];
        layer3[58][39:32] = buffer_data_3[2015:2008];
        layer3[58][47:40] = buffer_data_3[2023:2016];
        layer3[58][55:48] = buffer_data_3[2031:2024];
        layer4[58][7:0] = buffer_data_2[1983:1976];
        layer4[58][15:8] = buffer_data_2[1991:1984];
        layer4[58][23:16] = buffer_data_2[1999:1992];
        layer4[58][31:24] = buffer_data_2[2007:2000];
        layer4[58][39:32] = buffer_data_2[2015:2008];
        layer4[58][47:40] = buffer_data_2[2023:2016];
        layer4[58][55:48] = buffer_data_2[2031:2024];
        layer5[58][7:0] = buffer_data_1[1983:1976];
        layer5[58][15:8] = buffer_data_1[1991:1984];
        layer5[58][23:16] = buffer_data_1[1999:1992];
        layer5[58][31:24] = buffer_data_1[2007:2000];
        layer5[58][39:32] = buffer_data_1[2015:2008];
        layer5[58][47:40] = buffer_data_1[2023:2016];
        layer5[58][55:48] = buffer_data_1[2031:2024];
        layer6[58][7:0] = buffer_data_0[1983:1976];
        layer6[58][15:8] = buffer_data_0[1991:1984];
        layer6[58][23:16] = buffer_data_0[1999:1992];
        layer6[58][31:24] = buffer_data_0[2007:2000];
        layer6[58][39:32] = buffer_data_0[2015:2008];
        layer6[58][47:40] = buffer_data_0[2023:2016];
        layer6[58][55:48] = buffer_data_0[2031:2024];
        layer0[59][7:0] = buffer_data_6[1991:1984];
        layer0[59][15:8] = buffer_data_6[1999:1992];
        layer0[59][23:16] = buffer_data_6[2007:2000];
        layer0[59][31:24] = buffer_data_6[2015:2008];
        layer0[59][39:32] = buffer_data_6[2023:2016];
        layer0[59][47:40] = buffer_data_6[2031:2024];
        layer0[59][55:48] = buffer_data_6[2039:2032];
        layer1[59][7:0] = buffer_data_5[1991:1984];
        layer1[59][15:8] = buffer_data_5[1999:1992];
        layer1[59][23:16] = buffer_data_5[2007:2000];
        layer1[59][31:24] = buffer_data_5[2015:2008];
        layer1[59][39:32] = buffer_data_5[2023:2016];
        layer1[59][47:40] = buffer_data_5[2031:2024];
        layer1[59][55:48] = buffer_data_5[2039:2032];
        layer2[59][7:0] = buffer_data_4[1991:1984];
        layer2[59][15:8] = buffer_data_4[1999:1992];
        layer2[59][23:16] = buffer_data_4[2007:2000];
        layer2[59][31:24] = buffer_data_4[2015:2008];
        layer2[59][39:32] = buffer_data_4[2023:2016];
        layer2[59][47:40] = buffer_data_4[2031:2024];
        layer2[59][55:48] = buffer_data_4[2039:2032];
        layer3[59][7:0] = buffer_data_3[1991:1984];
        layer3[59][15:8] = buffer_data_3[1999:1992];
        layer3[59][23:16] = buffer_data_3[2007:2000];
        layer3[59][31:24] = buffer_data_3[2015:2008];
        layer3[59][39:32] = buffer_data_3[2023:2016];
        layer3[59][47:40] = buffer_data_3[2031:2024];
        layer3[59][55:48] = buffer_data_3[2039:2032];
        layer4[59][7:0] = buffer_data_2[1991:1984];
        layer4[59][15:8] = buffer_data_2[1999:1992];
        layer4[59][23:16] = buffer_data_2[2007:2000];
        layer4[59][31:24] = buffer_data_2[2015:2008];
        layer4[59][39:32] = buffer_data_2[2023:2016];
        layer4[59][47:40] = buffer_data_2[2031:2024];
        layer4[59][55:48] = buffer_data_2[2039:2032];
        layer5[59][7:0] = buffer_data_1[1991:1984];
        layer5[59][15:8] = buffer_data_1[1999:1992];
        layer5[59][23:16] = buffer_data_1[2007:2000];
        layer5[59][31:24] = buffer_data_1[2015:2008];
        layer5[59][39:32] = buffer_data_1[2023:2016];
        layer5[59][47:40] = buffer_data_1[2031:2024];
        layer5[59][55:48] = buffer_data_1[2039:2032];
        layer6[59][7:0] = buffer_data_0[1991:1984];
        layer6[59][15:8] = buffer_data_0[1999:1992];
        layer6[59][23:16] = buffer_data_0[2007:2000];
        layer6[59][31:24] = buffer_data_0[2015:2008];
        layer6[59][39:32] = buffer_data_0[2023:2016];
        layer6[59][47:40] = buffer_data_0[2031:2024];
        layer6[59][55:48] = buffer_data_0[2039:2032];
        layer0[60][7:0] = buffer_data_6[1999:1992];
        layer0[60][15:8] = buffer_data_6[2007:2000];
        layer0[60][23:16] = buffer_data_6[2015:2008];
        layer0[60][31:24] = buffer_data_6[2023:2016];
        layer0[60][39:32] = buffer_data_6[2031:2024];
        layer0[60][47:40] = buffer_data_6[2039:2032];
        layer0[60][55:48] = buffer_data_6[2047:2040];
        layer1[60][7:0] = buffer_data_5[1999:1992];
        layer1[60][15:8] = buffer_data_5[2007:2000];
        layer1[60][23:16] = buffer_data_5[2015:2008];
        layer1[60][31:24] = buffer_data_5[2023:2016];
        layer1[60][39:32] = buffer_data_5[2031:2024];
        layer1[60][47:40] = buffer_data_5[2039:2032];
        layer1[60][55:48] = buffer_data_5[2047:2040];
        layer2[60][7:0] = buffer_data_4[1999:1992];
        layer2[60][15:8] = buffer_data_4[2007:2000];
        layer2[60][23:16] = buffer_data_4[2015:2008];
        layer2[60][31:24] = buffer_data_4[2023:2016];
        layer2[60][39:32] = buffer_data_4[2031:2024];
        layer2[60][47:40] = buffer_data_4[2039:2032];
        layer2[60][55:48] = buffer_data_4[2047:2040];
        layer3[60][7:0] = buffer_data_3[1999:1992];
        layer3[60][15:8] = buffer_data_3[2007:2000];
        layer3[60][23:16] = buffer_data_3[2015:2008];
        layer3[60][31:24] = buffer_data_3[2023:2016];
        layer3[60][39:32] = buffer_data_3[2031:2024];
        layer3[60][47:40] = buffer_data_3[2039:2032];
        layer3[60][55:48] = buffer_data_3[2047:2040];
        layer4[60][7:0] = buffer_data_2[1999:1992];
        layer4[60][15:8] = buffer_data_2[2007:2000];
        layer4[60][23:16] = buffer_data_2[2015:2008];
        layer4[60][31:24] = buffer_data_2[2023:2016];
        layer4[60][39:32] = buffer_data_2[2031:2024];
        layer4[60][47:40] = buffer_data_2[2039:2032];
        layer4[60][55:48] = buffer_data_2[2047:2040];
        layer5[60][7:0] = buffer_data_1[1999:1992];
        layer5[60][15:8] = buffer_data_1[2007:2000];
        layer5[60][23:16] = buffer_data_1[2015:2008];
        layer5[60][31:24] = buffer_data_1[2023:2016];
        layer5[60][39:32] = buffer_data_1[2031:2024];
        layer5[60][47:40] = buffer_data_1[2039:2032];
        layer5[60][55:48] = buffer_data_1[2047:2040];
        layer6[60][7:0] = buffer_data_0[1999:1992];
        layer6[60][15:8] = buffer_data_0[2007:2000];
        layer6[60][23:16] = buffer_data_0[2015:2008];
        layer6[60][31:24] = buffer_data_0[2023:2016];
        layer6[60][39:32] = buffer_data_0[2031:2024];
        layer6[60][47:40] = buffer_data_0[2039:2032];
        layer6[60][55:48] = buffer_data_0[2047:2040];
        layer0[61][7:0] = buffer_data_6[2007:2000];
        layer0[61][15:8] = buffer_data_6[2015:2008];
        layer0[61][23:16] = buffer_data_6[2023:2016];
        layer0[61][31:24] = buffer_data_6[2031:2024];
        layer0[61][39:32] = buffer_data_6[2039:2032];
        layer0[61][47:40] = buffer_data_6[2047:2040];
        layer0[61][55:48] = buffer_data_6[2055:2048];
        layer1[61][7:0] = buffer_data_5[2007:2000];
        layer1[61][15:8] = buffer_data_5[2015:2008];
        layer1[61][23:16] = buffer_data_5[2023:2016];
        layer1[61][31:24] = buffer_data_5[2031:2024];
        layer1[61][39:32] = buffer_data_5[2039:2032];
        layer1[61][47:40] = buffer_data_5[2047:2040];
        layer1[61][55:48] = buffer_data_5[2055:2048];
        layer2[61][7:0] = buffer_data_4[2007:2000];
        layer2[61][15:8] = buffer_data_4[2015:2008];
        layer2[61][23:16] = buffer_data_4[2023:2016];
        layer2[61][31:24] = buffer_data_4[2031:2024];
        layer2[61][39:32] = buffer_data_4[2039:2032];
        layer2[61][47:40] = buffer_data_4[2047:2040];
        layer2[61][55:48] = buffer_data_4[2055:2048];
        layer3[61][7:0] = buffer_data_3[2007:2000];
        layer3[61][15:8] = buffer_data_3[2015:2008];
        layer3[61][23:16] = buffer_data_3[2023:2016];
        layer3[61][31:24] = buffer_data_3[2031:2024];
        layer3[61][39:32] = buffer_data_3[2039:2032];
        layer3[61][47:40] = buffer_data_3[2047:2040];
        layer3[61][55:48] = buffer_data_3[2055:2048];
        layer4[61][7:0] = buffer_data_2[2007:2000];
        layer4[61][15:8] = buffer_data_2[2015:2008];
        layer4[61][23:16] = buffer_data_2[2023:2016];
        layer4[61][31:24] = buffer_data_2[2031:2024];
        layer4[61][39:32] = buffer_data_2[2039:2032];
        layer4[61][47:40] = buffer_data_2[2047:2040];
        layer4[61][55:48] = buffer_data_2[2055:2048];
        layer5[61][7:0] = buffer_data_1[2007:2000];
        layer5[61][15:8] = buffer_data_1[2015:2008];
        layer5[61][23:16] = buffer_data_1[2023:2016];
        layer5[61][31:24] = buffer_data_1[2031:2024];
        layer5[61][39:32] = buffer_data_1[2039:2032];
        layer5[61][47:40] = buffer_data_1[2047:2040];
        layer5[61][55:48] = buffer_data_1[2055:2048];
        layer6[61][7:0] = buffer_data_0[2007:2000];
        layer6[61][15:8] = buffer_data_0[2015:2008];
        layer6[61][23:16] = buffer_data_0[2023:2016];
        layer6[61][31:24] = buffer_data_0[2031:2024];
        layer6[61][39:32] = buffer_data_0[2039:2032];
        layer6[61][47:40] = buffer_data_0[2047:2040];
        layer6[61][55:48] = buffer_data_0[2055:2048];
        layer0[62][7:0] = buffer_data_6[2015:2008];
        layer0[62][15:8] = buffer_data_6[2023:2016];
        layer0[62][23:16] = buffer_data_6[2031:2024];
        layer0[62][31:24] = buffer_data_6[2039:2032];
        layer0[62][39:32] = buffer_data_6[2047:2040];
        layer0[62][47:40] = buffer_data_6[2055:2048];
        layer0[62][55:48] = buffer_data_6[2063:2056];
        layer1[62][7:0] = buffer_data_5[2015:2008];
        layer1[62][15:8] = buffer_data_5[2023:2016];
        layer1[62][23:16] = buffer_data_5[2031:2024];
        layer1[62][31:24] = buffer_data_5[2039:2032];
        layer1[62][39:32] = buffer_data_5[2047:2040];
        layer1[62][47:40] = buffer_data_5[2055:2048];
        layer1[62][55:48] = buffer_data_5[2063:2056];
        layer2[62][7:0] = buffer_data_4[2015:2008];
        layer2[62][15:8] = buffer_data_4[2023:2016];
        layer2[62][23:16] = buffer_data_4[2031:2024];
        layer2[62][31:24] = buffer_data_4[2039:2032];
        layer2[62][39:32] = buffer_data_4[2047:2040];
        layer2[62][47:40] = buffer_data_4[2055:2048];
        layer2[62][55:48] = buffer_data_4[2063:2056];
        layer3[62][7:0] = buffer_data_3[2015:2008];
        layer3[62][15:8] = buffer_data_3[2023:2016];
        layer3[62][23:16] = buffer_data_3[2031:2024];
        layer3[62][31:24] = buffer_data_3[2039:2032];
        layer3[62][39:32] = buffer_data_3[2047:2040];
        layer3[62][47:40] = buffer_data_3[2055:2048];
        layer3[62][55:48] = buffer_data_3[2063:2056];
        layer4[62][7:0] = buffer_data_2[2015:2008];
        layer4[62][15:8] = buffer_data_2[2023:2016];
        layer4[62][23:16] = buffer_data_2[2031:2024];
        layer4[62][31:24] = buffer_data_2[2039:2032];
        layer4[62][39:32] = buffer_data_2[2047:2040];
        layer4[62][47:40] = buffer_data_2[2055:2048];
        layer4[62][55:48] = buffer_data_2[2063:2056];
        layer5[62][7:0] = buffer_data_1[2015:2008];
        layer5[62][15:8] = buffer_data_1[2023:2016];
        layer5[62][23:16] = buffer_data_1[2031:2024];
        layer5[62][31:24] = buffer_data_1[2039:2032];
        layer5[62][39:32] = buffer_data_1[2047:2040];
        layer5[62][47:40] = buffer_data_1[2055:2048];
        layer5[62][55:48] = buffer_data_1[2063:2056];
        layer6[62][7:0] = buffer_data_0[2015:2008];
        layer6[62][15:8] = buffer_data_0[2023:2016];
        layer6[62][23:16] = buffer_data_0[2031:2024];
        layer6[62][31:24] = buffer_data_0[2039:2032];
        layer6[62][39:32] = buffer_data_0[2047:2040];
        layer6[62][47:40] = buffer_data_0[2055:2048];
        layer6[62][55:48] = buffer_data_0[2063:2056];
        layer0[63][7:0] = buffer_data_6[2023:2016];
        layer0[63][15:8] = buffer_data_6[2031:2024];
        layer0[63][23:16] = buffer_data_6[2039:2032];
        layer0[63][31:24] = buffer_data_6[2047:2040];
        layer0[63][39:32] = buffer_data_6[2055:2048];
        layer0[63][47:40] = buffer_data_6[2063:2056];
        layer0[63][55:48] = buffer_data_6[2071:2064];
        layer1[63][7:0] = buffer_data_5[2023:2016];
        layer1[63][15:8] = buffer_data_5[2031:2024];
        layer1[63][23:16] = buffer_data_5[2039:2032];
        layer1[63][31:24] = buffer_data_5[2047:2040];
        layer1[63][39:32] = buffer_data_5[2055:2048];
        layer1[63][47:40] = buffer_data_5[2063:2056];
        layer1[63][55:48] = buffer_data_5[2071:2064];
        layer2[63][7:0] = buffer_data_4[2023:2016];
        layer2[63][15:8] = buffer_data_4[2031:2024];
        layer2[63][23:16] = buffer_data_4[2039:2032];
        layer2[63][31:24] = buffer_data_4[2047:2040];
        layer2[63][39:32] = buffer_data_4[2055:2048];
        layer2[63][47:40] = buffer_data_4[2063:2056];
        layer2[63][55:48] = buffer_data_4[2071:2064];
        layer3[63][7:0] = buffer_data_3[2023:2016];
        layer3[63][15:8] = buffer_data_3[2031:2024];
        layer3[63][23:16] = buffer_data_3[2039:2032];
        layer3[63][31:24] = buffer_data_3[2047:2040];
        layer3[63][39:32] = buffer_data_3[2055:2048];
        layer3[63][47:40] = buffer_data_3[2063:2056];
        layer3[63][55:48] = buffer_data_3[2071:2064];
        layer4[63][7:0] = buffer_data_2[2023:2016];
        layer4[63][15:8] = buffer_data_2[2031:2024];
        layer4[63][23:16] = buffer_data_2[2039:2032];
        layer4[63][31:24] = buffer_data_2[2047:2040];
        layer4[63][39:32] = buffer_data_2[2055:2048];
        layer4[63][47:40] = buffer_data_2[2063:2056];
        layer4[63][55:48] = buffer_data_2[2071:2064];
        layer5[63][7:0] = buffer_data_1[2023:2016];
        layer5[63][15:8] = buffer_data_1[2031:2024];
        layer5[63][23:16] = buffer_data_1[2039:2032];
        layer5[63][31:24] = buffer_data_1[2047:2040];
        layer5[63][39:32] = buffer_data_1[2055:2048];
        layer5[63][47:40] = buffer_data_1[2063:2056];
        layer5[63][55:48] = buffer_data_1[2071:2064];
        layer6[63][7:0] = buffer_data_0[2023:2016];
        layer6[63][15:8] = buffer_data_0[2031:2024];
        layer6[63][23:16] = buffer_data_0[2039:2032];
        layer6[63][31:24] = buffer_data_0[2047:2040];
        layer6[63][39:32] = buffer_data_0[2055:2048];
        layer6[63][47:40] = buffer_data_0[2063:2056];
        layer6[63][55:48] = buffer_data_0[2071:2064];
    end
    ST_GAUSSIAN_4: begin
        layer0[0][7:0] = buffer_data_6[2031:2024];
        layer0[0][15:8] = buffer_data_6[2039:2032];
        layer0[0][23:16] = buffer_data_6[2047:2040];
        layer0[0][31:24] = buffer_data_6[2055:2048];
        layer0[0][39:32] = buffer_data_6[2063:2056];
        layer0[0][47:40] = buffer_data_6[2071:2064];
        layer0[0][55:48] = buffer_data_6[2079:2072];
        layer1[0][7:0] = buffer_data_5[2031:2024];
        layer1[0][15:8] = buffer_data_5[2039:2032];
        layer1[0][23:16] = buffer_data_5[2047:2040];
        layer1[0][31:24] = buffer_data_5[2055:2048];
        layer1[0][39:32] = buffer_data_5[2063:2056];
        layer1[0][47:40] = buffer_data_5[2071:2064];
        layer1[0][55:48] = buffer_data_5[2079:2072];
        layer2[0][7:0] = buffer_data_4[2031:2024];
        layer2[0][15:8] = buffer_data_4[2039:2032];
        layer2[0][23:16] = buffer_data_4[2047:2040];
        layer2[0][31:24] = buffer_data_4[2055:2048];
        layer2[0][39:32] = buffer_data_4[2063:2056];
        layer2[0][47:40] = buffer_data_4[2071:2064];
        layer2[0][55:48] = buffer_data_4[2079:2072];
        layer3[0][7:0] = buffer_data_3[2031:2024];
        layer3[0][15:8] = buffer_data_3[2039:2032];
        layer3[0][23:16] = buffer_data_3[2047:2040];
        layer3[0][31:24] = buffer_data_3[2055:2048];
        layer3[0][39:32] = buffer_data_3[2063:2056];
        layer3[0][47:40] = buffer_data_3[2071:2064];
        layer3[0][55:48] = buffer_data_3[2079:2072];
        layer4[0][7:0] = buffer_data_2[2031:2024];
        layer4[0][15:8] = buffer_data_2[2039:2032];
        layer4[0][23:16] = buffer_data_2[2047:2040];
        layer4[0][31:24] = buffer_data_2[2055:2048];
        layer4[0][39:32] = buffer_data_2[2063:2056];
        layer4[0][47:40] = buffer_data_2[2071:2064];
        layer4[0][55:48] = buffer_data_2[2079:2072];
        layer5[0][7:0] = buffer_data_1[2031:2024];
        layer5[0][15:8] = buffer_data_1[2039:2032];
        layer5[0][23:16] = buffer_data_1[2047:2040];
        layer5[0][31:24] = buffer_data_1[2055:2048];
        layer5[0][39:32] = buffer_data_1[2063:2056];
        layer5[0][47:40] = buffer_data_1[2071:2064];
        layer5[0][55:48] = buffer_data_1[2079:2072];
        layer6[0][7:0] = buffer_data_0[2031:2024];
        layer6[0][15:8] = buffer_data_0[2039:2032];
        layer6[0][23:16] = buffer_data_0[2047:2040];
        layer6[0][31:24] = buffer_data_0[2055:2048];
        layer6[0][39:32] = buffer_data_0[2063:2056];
        layer6[0][47:40] = buffer_data_0[2071:2064];
        layer6[0][55:48] = buffer_data_0[2079:2072];
        layer0[1][7:0] = buffer_data_6[2039:2032];
        layer0[1][15:8] = buffer_data_6[2047:2040];
        layer0[1][23:16] = buffer_data_6[2055:2048];
        layer0[1][31:24] = buffer_data_6[2063:2056];
        layer0[1][39:32] = buffer_data_6[2071:2064];
        layer0[1][47:40] = buffer_data_6[2079:2072];
        layer0[1][55:48] = buffer_data_6[2087:2080];
        layer1[1][7:0] = buffer_data_5[2039:2032];
        layer1[1][15:8] = buffer_data_5[2047:2040];
        layer1[1][23:16] = buffer_data_5[2055:2048];
        layer1[1][31:24] = buffer_data_5[2063:2056];
        layer1[1][39:32] = buffer_data_5[2071:2064];
        layer1[1][47:40] = buffer_data_5[2079:2072];
        layer1[1][55:48] = buffer_data_5[2087:2080];
        layer2[1][7:0] = buffer_data_4[2039:2032];
        layer2[1][15:8] = buffer_data_4[2047:2040];
        layer2[1][23:16] = buffer_data_4[2055:2048];
        layer2[1][31:24] = buffer_data_4[2063:2056];
        layer2[1][39:32] = buffer_data_4[2071:2064];
        layer2[1][47:40] = buffer_data_4[2079:2072];
        layer2[1][55:48] = buffer_data_4[2087:2080];
        layer3[1][7:0] = buffer_data_3[2039:2032];
        layer3[1][15:8] = buffer_data_3[2047:2040];
        layer3[1][23:16] = buffer_data_3[2055:2048];
        layer3[1][31:24] = buffer_data_3[2063:2056];
        layer3[1][39:32] = buffer_data_3[2071:2064];
        layer3[1][47:40] = buffer_data_3[2079:2072];
        layer3[1][55:48] = buffer_data_3[2087:2080];
        layer4[1][7:0] = buffer_data_2[2039:2032];
        layer4[1][15:8] = buffer_data_2[2047:2040];
        layer4[1][23:16] = buffer_data_2[2055:2048];
        layer4[1][31:24] = buffer_data_2[2063:2056];
        layer4[1][39:32] = buffer_data_2[2071:2064];
        layer4[1][47:40] = buffer_data_2[2079:2072];
        layer4[1][55:48] = buffer_data_2[2087:2080];
        layer5[1][7:0] = buffer_data_1[2039:2032];
        layer5[1][15:8] = buffer_data_1[2047:2040];
        layer5[1][23:16] = buffer_data_1[2055:2048];
        layer5[1][31:24] = buffer_data_1[2063:2056];
        layer5[1][39:32] = buffer_data_1[2071:2064];
        layer5[1][47:40] = buffer_data_1[2079:2072];
        layer5[1][55:48] = buffer_data_1[2087:2080];
        layer6[1][7:0] = buffer_data_0[2039:2032];
        layer6[1][15:8] = buffer_data_0[2047:2040];
        layer6[1][23:16] = buffer_data_0[2055:2048];
        layer6[1][31:24] = buffer_data_0[2063:2056];
        layer6[1][39:32] = buffer_data_0[2071:2064];
        layer6[1][47:40] = buffer_data_0[2079:2072];
        layer6[1][55:48] = buffer_data_0[2087:2080];
        layer0[2][7:0] = buffer_data_6[2047:2040];
        layer0[2][15:8] = buffer_data_6[2055:2048];
        layer0[2][23:16] = buffer_data_6[2063:2056];
        layer0[2][31:24] = buffer_data_6[2071:2064];
        layer0[2][39:32] = buffer_data_6[2079:2072];
        layer0[2][47:40] = buffer_data_6[2087:2080];
        layer0[2][55:48] = buffer_data_6[2095:2088];
        layer1[2][7:0] = buffer_data_5[2047:2040];
        layer1[2][15:8] = buffer_data_5[2055:2048];
        layer1[2][23:16] = buffer_data_5[2063:2056];
        layer1[2][31:24] = buffer_data_5[2071:2064];
        layer1[2][39:32] = buffer_data_5[2079:2072];
        layer1[2][47:40] = buffer_data_5[2087:2080];
        layer1[2][55:48] = buffer_data_5[2095:2088];
        layer2[2][7:0] = buffer_data_4[2047:2040];
        layer2[2][15:8] = buffer_data_4[2055:2048];
        layer2[2][23:16] = buffer_data_4[2063:2056];
        layer2[2][31:24] = buffer_data_4[2071:2064];
        layer2[2][39:32] = buffer_data_4[2079:2072];
        layer2[2][47:40] = buffer_data_4[2087:2080];
        layer2[2][55:48] = buffer_data_4[2095:2088];
        layer3[2][7:0] = buffer_data_3[2047:2040];
        layer3[2][15:8] = buffer_data_3[2055:2048];
        layer3[2][23:16] = buffer_data_3[2063:2056];
        layer3[2][31:24] = buffer_data_3[2071:2064];
        layer3[2][39:32] = buffer_data_3[2079:2072];
        layer3[2][47:40] = buffer_data_3[2087:2080];
        layer3[2][55:48] = buffer_data_3[2095:2088];
        layer4[2][7:0] = buffer_data_2[2047:2040];
        layer4[2][15:8] = buffer_data_2[2055:2048];
        layer4[2][23:16] = buffer_data_2[2063:2056];
        layer4[2][31:24] = buffer_data_2[2071:2064];
        layer4[2][39:32] = buffer_data_2[2079:2072];
        layer4[2][47:40] = buffer_data_2[2087:2080];
        layer4[2][55:48] = buffer_data_2[2095:2088];
        layer5[2][7:0] = buffer_data_1[2047:2040];
        layer5[2][15:8] = buffer_data_1[2055:2048];
        layer5[2][23:16] = buffer_data_1[2063:2056];
        layer5[2][31:24] = buffer_data_1[2071:2064];
        layer5[2][39:32] = buffer_data_1[2079:2072];
        layer5[2][47:40] = buffer_data_1[2087:2080];
        layer5[2][55:48] = buffer_data_1[2095:2088];
        layer6[2][7:0] = buffer_data_0[2047:2040];
        layer6[2][15:8] = buffer_data_0[2055:2048];
        layer6[2][23:16] = buffer_data_0[2063:2056];
        layer6[2][31:24] = buffer_data_0[2071:2064];
        layer6[2][39:32] = buffer_data_0[2079:2072];
        layer6[2][47:40] = buffer_data_0[2087:2080];
        layer6[2][55:48] = buffer_data_0[2095:2088];
        layer0[3][7:0] = buffer_data_6[2055:2048];
        layer0[3][15:8] = buffer_data_6[2063:2056];
        layer0[3][23:16] = buffer_data_6[2071:2064];
        layer0[3][31:24] = buffer_data_6[2079:2072];
        layer0[3][39:32] = buffer_data_6[2087:2080];
        layer0[3][47:40] = buffer_data_6[2095:2088];
        layer0[3][55:48] = buffer_data_6[2103:2096];
        layer1[3][7:0] = buffer_data_5[2055:2048];
        layer1[3][15:8] = buffer_data_5[2063:2056];
        layer1[3][23:16] = buffer_data_5[2071:2064];
        layer1[3][31:24] = buffer_data_5[2079:2072];
        layer1[3][39:32] = buffer_data_5[2087:2080];
        layer1[3][47:40] = buffer_data_5[2095:2088];
        layer1[3][55:48] = buffer_data_5[2103:2096];
        layer2[3][7:0] = buffer_data_4[2055:2048];
        layer2[3][15:8] = buffer_data_4[2063:2056];
        layer2[3][23:16] = buffer_data_4[2071:2064];
        layer2[3][31:24] = buffer_data_4[2079:2072];
        layer2[3][39:32] = buffer_data_4[2087:2080];
        layer2[3][47:40] = buffer_data_4[2095:2088];
        layer2[3][55:48] = buffer_data_4[2103:2096];
        layer3[3][7:0] = buffer_data_3[2055:2048];
        layer3[3][15:8] = buffer_data_3[2063:2056];
        layer3[3][23:16] = buffer_data_3[2071:2064];
        layer3[3][31:24] = buffer_data_3[2079:2072];
        layer3[3][39:32] = buffer_data_3[2087:2080];
        layer3[3][47:40] = buffer_data_3[2095:2088];
        layer3[3][55:48] = buffer_data_3[2103:2096];
        layer4[3][7:0] = buffer_data_2[2055:2048];
        layer4[3][15:8] = buffer_data_2[2063:2056];
        layer4[3][23:16] = buffer_data_2[2071:2064];
        layer4[3][31:24] = buffer_data_2[2079:2072];
        layer4[3][39:32] = buffer_data_2[2087:2080];
        layer4[3][47:40] = buffer_data_2[2095:2088];
        layer4[3][55:48] = buffer_data_2[2103:2096];
        layer5[3][7:0] = buffer_data_1[2055:2048];
        layer5[3][15:8] = buffer_data_1[2063:2056];
        layer5[3][23:16] = buffer_data_1[2071:2064];
        layer5[3][31:24] = buffer_data_1[2079:2072];
        layer5[3][39:32] = buffer_data_1[2087:2080];
        layer5[3][47:40] = buffer_data_1[2095:2088];
        layer5[3][55:48] = buffer_data_1[2103:2096];
        layer6[3][7:0] = buffer_data_0[2055:2048];
        layer6[3][15:8] = buffer_data_0[2063:2056];
        layer6[3][23:16] = buffer_data_0[2071:2064];
        layer6[3][31:24] = buffer_data_0[2079:2072];
        layer6[3][39:32] = buffer_data_0[2087:2080];
        layer6[3][47:40] = buffer_data_0[2095:2088];
        layer6[3][55:48] = buffer_data_0[2103:2096];
        layer0[4][7:0] = buffer_data_6[2063:2056];
        layer0[4][15:8] = buffer_data_6[2071:2064];
        layer0[4][23:16] = buffer_data_6[2079:2072];
        layer0[4][31:24] = buffer_data_6[2087:2080];
        layer0[4][39:32] = buffer_data_6[2095:2088];
        layer0[4][47:40] = buffer_data_6[2103:2096];
        layer0[4][55:48] = buffer_data_6[2111:2104];
        layer1[4][7:0] = buffer_data_5[2063:2056];
        layer1[4][15:8] = buffer_data_5[2071:2064];
        layer1[4][23:16] = buffer_data_5[2079:2072];
        layer1[4][31:24] = buffer_data_5[2087:2080];
        layer1[4][39:32] = buffer_data_5[2095:2088];
        layer1[4][47:40] = buffer_data_5[2103:2096];
        layer1[4][55:48] = buffer_data_5[2111:2104];
        layer2[4][7:0] = buffer_data_4[2063:2056];
        layer2[4][15:8] = buffer_data_4[2071:2064];
        layer2[4][23:16] = buffer_data_4[2079:2072];
        layer2[4][31:24] = buffer_data_4[2087:2080];
        layer2[4][39:32] = buffer_data_4[2095:2088];
        layer2[4][47:40] = buffer_data_4[2103:2096];
        layer2[4][55:48] = buffer_data_4[2111:2104];
        layer3[4][7:0] = buffer_data_3[2063:2056];
        layer3[4][15:8] = buffer_data_3[2071:2064];
        layer3[4][23:16] = buffer_data_3[2079:2072];
        layer3[4][31:24] = buffer_data_3[2087:2080];
        layer3[4][39:32] = buffer_data_3[2095:2088];
        layer3[4][47:40] = buffer_data_3[2103:2096];
        layer3[4][55:48] = buffer_data_3[2111:2104];
        layer4[4][7:0] = buffer_data_2[2063:2056];
        layer4[4][15:8] = buffer_data_2[2071:2064];
        layer4[4][23:16] = buffer_data_2[2079:2072];
        layer4[4][31:24] = buffer_data_2[2087:2080];
        layer4[4][39:32] = buffer_data_2[2095:2088];
        layer4[4][47:40] = buffer_data_2[2103:2096];
        layer4[4][55:48] = buffer_data_2[2111:2104];
        layer5[4][7:0] = buffer_data_1[2063:2056];
        layer5[4][15:8] = buffer_data_1[2071:2064];
        layer5[4][23:16] = buffer_data_1[2079:2072];
        layer5[4][31:24] = buffer_data_1[2087:2080];
        layer5[4][39:32] = buffer_data_1[2095:2088];
        layer5[4][47:40] = buffer_data_1[2103:2096];
        layer5[4][55:48] = buffer_data_1[2111:2104];
        layer6[4][7:0] = buffer_data_0[2063:2056];
        layer6[4][15:8] = buffer_data_0[2071:2064];
        layer6[4][23:16] = buffer_data_0[2079:2072];
        layer6[4][31:24] = buffer_data_0[2087:2080];
        layer6[4][39:32] = buffer_data_0[2095:2088];
        layer6[4][47:40] = buffer_data_0[2103:2096];
        layer6[4][55:48] = buffer_data_0[2111:2104];
        layer0[5][7:0] = buffer_data_6[2071:2064];
        layer0[5][15:8] = buffer_data_6[2079:2072];
        layer0[5][23:16] = buffer_data_6[2087:2080];
        layer0[5][31:24] = buffer_data_6[2095:2088];
        layer0[5][39:32] = buffer_data_6[2103:2096];
        layer0[5][47:40] = buffer_data_6[2111:2104];
        layer0[5][55:48] = buffer_data_6[2119:2112];
        layer1[5][7:0] = buffer_data_5[2071:2064];
        layer1[5][15:8] = buffer_data_5[2079:2072];
        layer1[5][23:16] = buffer_data_5[2087:2080];
        layer1[5][31:24] = buffer_data_5[2095:2088];
        layer1[5][39:32] = buffer_data_5[2103:2096];
        layer1[5][47:40] = buffer_data_5[2111:2104];
        layer1[5][55:48] = buffer_data_5[2119:2112];
        layer2[5][7:0] = buffer_data_4[2071:2064];
        layer2[5][15:8] = buffer_data_4[2079:2072];
        layer2[5][23:16] = buffer_data_4[2087:2080];
        layer2[5][31:24] = buffer_data_4[2095:2088];
        layer2[5][39:32] = buffer_data_4[2103:2096];
        layer2[5][47:40] = buffer_data_4[2111:2104];
        layer2[5][55:48] = buffer_data_4[2119:2112];
        layer3[5][7:0] = buffer_data_3[2071:2064];
        layer3[5][15:8] = buffer_data_3[2079:2072];
        layer3[5][23:16] = buffer_data_3[2087:2080];
        layer3[5][31:24] = buffer_data_3[2095:2088];
        layer3[5][39:32] = buffer_data_3[2103:2096];
        layer3[5][47:40] = buffer_data_3[2111:2104];
        layer3[5][55:48] = buffer_data_3[2119:2112];
        layer4[5][7:0] = buffer_data_2[2071:2064];
        layer4[5][15:8] = buffer_data_2[2079:2072];
        layer4[5][23:16] = buffer_data_2[2087:2080];
        layer4[5][31:24] = buffer_data_2[2095:2088];
        layer4[5][39:32] = buffer_data_2[2103:2096];
        layer4[5][47:40] = buffer_data_2[2111:2104];
        layer4[5][55:48] = buffer_data_2[2119:2112];
        layer5[5][7:0] = buffer_data_1[2071:2064];
        layer5[5][15:8] = buffer_data_1[2079:2072];
        layer5[5][23:16] = buffer_data_1[2087:2080];
        layer5[5][31:24] = buffer_data_1[2095:2088];
        layer5[5][39:32] = buffer_data_1[2103:2096];
        layer5[5][47:40] = buffer_data_1[2111:2104];
        layer5[5][55:48] = buffer_data_1[2119:2112];
        layer6[5][7:0] = buffer_data_0[2071:2064];
        layer6[5][15:8] = buffer_data_0[2079:2072];
        layer6[5][23:16] = buffer_data_0[2087:2080];
        layer6[5][31:24] = buffer_data_0[2095:2088];
        layer6[5][39:32] = buffer_data_0[2103:2096];
        layer6[5][47:40] = buffer_data_0[2111:2104];
        layer6[5][55:48] = buffer_data_0[2119:2112];
        layer0[6][7:0] = buffer_data_6[2079:2072];
        layer0[6][15:8] = buffer_data_6[2087:2080];
        layer0[6][23:16] = buffer_data_6[2095:2088];
        layer0[6][31:24] = buffer_data_6[2103:2096];
        layer0[6][39:32] = buffer_data_6[2111:2104];
        layer0[6][47:40] = buffer_data_6[2119:2112];
        layer0[6][55:48] = buffer_data_6[2127:2120];
        layer1[6][7:0] = buffer_data_5[2079:2072];
        layer1[6][15:8] = buffer_data_5[2087:2080];
        layer1[6][23:16] = buffer_data_5[2095:2088];
        layer1[6][31:24] = buffer_data_5[2103:2096];
        layer1[6][39:32] = buffer_data_5[2111:2104];
        layer1[6][47:40] = buffer_data_5[2119:2112];
        layer1[6][55:48] = buffer_data_5[2127:2120];
        layer2[6][7:0] = buffer_data_4[2079:2072];
        layer2[6][15:8] = buffer_data_4[2087:2080];
        layer2[6][23:16] = buffer_data_4[2095:2088];
        layer2[6][31:24] = buffer_data_4[2103:2096];
        layer2[6][39:32] = buffer_data_4[2111:2104];
        layer2[6][47:40] = buffer_data_4[2119:2112];
        layer2[6][55:48] = buffer_data_4[2127:2120];
        layer3[6][7:0] = buffer_data_3[2079:2072];
        layer3[6][15:8] = buffer_data_3[2087:2080];
        layer3[6][23:16] = buffer_data_3[2095:2088];
        layer3[6][31:24] = buffer_data_3[2103:2096];
        layer3[6][39:32] = buffer_data_3[2111:2104];
        layer3[6][47:40] = buffer_data_3[2119:2112];
        layer3[6][55:48] = buffer_data_3[2127:2120];
        layer4[6][7:0] = buffer_data_2[2079:2072];
        layer4[6][15:8] = buffer_data_2[2087:2080];
        layer4[6][23:16] = buffer_data_2[2095:2088];
        layer4[6][31:24] = buffer_data_2[2103:2096];
        layer4[6][39:32] = buffer_data_2[2111:2104];
        layer4[6][47:40] = buffer_data_2[2119:2112];
        layer4[6][55:48] = buffer_data_2[2127:2120];
        layer5[6][7:0] = buffer_data_1[2079:2072];
        layer5[6][15:8] = buffer_data_1[2087:2080];
        layer5[6][23:16] = buffer_data_1[2095:2088];
        layer5[6][31:24] = buffer_data_1[2103:2096];
        layer5[6][39:32] = buffer_data_1[2111:2104];
        layer5[6][47:40] = buffer_data_1[2119:2112];
        layer5[6][55:48] = buffer_data_1[2127:2120];
        layer6[6][7:0] = buffer_data_0[2079:2072];
        layer6[6][15:8] = buffer_data_0[2087:2080];
        layer6[6][23:16] = buffer_data_0[2095:2088];
        layer6[6][31:24] = buffer_data_0[2103:2096];
        layer6[6][39:32] = buffer_data_0[2111:2104];
        layer6[6][47:40] = buffer_data_0[2119:2112];
        layer6[6][55:48] = buffer_data_0[2127:2120];
        layer0[7][7:0] = buffer_data_6[2087:2080];
        layer0[7][15:8] = buffer_data_6[2095:2088];
        layer0[7][23:16] = buffer_data_6[2103:2096];
        layer0[7][31:24] = buffer_data_6[2111:2104];
        layer0[7][39:32] = buffer_data_6[2119:2112];
        layer0[7][47:40] = buffer_data_6[2127:2120];
        layer0[7][55:48] = buffer_data_6[2135:2128];
        layer1[7][7:0] = buffer_data_5[2087:2080];
        layer1[7][15:8] = buffer_data_5[2095:2088];
        layer1[7][23:16] = buffer_data_5[2103:2096];
        layer1[7][31:24] = buffer_data_5[2111:2104];
        layer1[7][39:32] = buffer_data_5[2119:2112];
        layer1[7][47:40] = buffer_data_5[2127:2120];
        layer1[7][55:48] = buffer_data_5[2135:2128];
        layer2[7][7:0] = buffer_data_4[2087:2080];
        layer2[7][15:8] = buffer_data_4[2095:2088];
        layer2[7][23:16] = buffer_data_4[2103:2096];
        layer2[7][31:24] = buffer_data_4[2111:2104];
        layer2[7][39:32] = buffer_data_4[2119:2112];
        layer2[7][47:40] = buffer_data_4[2127:2120];
        layer2[7][55:48] = buffer_data_4[2135:2128];
        layer3[7][7:0] = buffer_data_3[2087:2080];
        layer3[7][15:8] = buffer_data_3[2095:2088];
        layer3[7][23:16] = buffer_data_3[2103:2096];
        layer3[7][31:24] = buffer_data_3[2111:2104];
        layer3[7][39:32] = buffer_data_3[2119:2112];
        layer3[7][47:40] = buffer_data_3[2127:2120];
        layer3[7][55:48] = buffer_data_3[2135:2128];
        layer4[7][7:0] = buffer_data_2[2087:2080];
        layer4[7][15:8] = buffer_data_2[2095:2088];
        layer4[7][23:16] = buffer_data_2[2103:2096];
        layer4[7][31:24] = buffer_data_2[2111:2104];
        layer4[7][39:32] = buffer_data_2[2119:2112];
        layer4[7][47:40] = buffer_data_2[2127:2120];
        layer4[7][55:48] = buffer_data_2[2135:2128];
        layer5[7][7:0] = buffer_data_1[2087:2080];
        layer5[7][15:8] = buffer_data_1[2095:2088];
        layer5[7][23:16] = buffer_data_1[2103:2096];
        layer5[7][31:24] = buffer_data_1[2111:2104];
        layer5[7][39:32] = buffer_data_1[2119:2112];
        layer5[7][47:40] = buffer_data_1[2127:2120];
        layer5[7][55:48] = buffer_data_1[2135:2128];
        layer6[7][7:0] = buffer_data_0[2087:2080];
        layer6[7][15:8] = buffer_data_0[2095:2088];
        layer6[7][23:16] = buffer_data_0[2103:2096];
        layer6[7][31:24] = buffer_data_0[2111:2104];
        layer6[7][39:32] = buffer_data_0[2119:2112];
        layer6[7][47:40] = buffer_data_0[2127:2120];
        layer6[7][55:48] = buffer_data_0[2135:2128];
        layer0[8][7:0] = buffer_data_6[2095:2088];
        layer0[8][15:8] = buffer_data_6[2103:2096];
        layer0[8][23:16] = buffer_data_6[2111:2104];
        layer0[8][31:24] = buffer_data_6[2119:2112];
        layer0[8][39:32] = buffer_data_6[2127:2120];
        layer0[8][47:40] = buffer_data_6[2135:2128];
        layer0[8][55:48] = buffer_data_6[2143:2136];
        layer1[8][7:0] = buffer_data_5[2095:2088];
        layer1[8][15:8] = buffer_data_5[2103:2096];
        layer1[8][23:16] = buffer_data_5[2111:2104];
        layer1[8][31:24] = buffer_data_5[2119:2112];
        layer1[8][39:32] = buffer_data_5[2127:2120];
        layer1[8][47:40] = buffer_data_5[2135:2128];
        layer1[8][55:48] = buffer_data_5[2143:2136];
        layer2[8][7:0] = buffer_data_4[2095:2088];
        layer2[8][15:8] = buffer_data_4[2103:2096];
        layer2[8][23:16] = buffer_data_4[2111:2104];
        layer2[8][31:24] = buffer_data_4[2119:2112];
        layer2[8][39:32] = buffer_data_4[2127:2120];
        layer2[8][47:40] = buffer_data_4[2135:2128];
        layer2[8][55:48] = buffer_data_4[2143:2136];
        layer3[8][7:0] = buffer_data_3[2095:2088];
        layer3[8][15:8] = buffer_data_3[2103:2096];
        layer3[8][23:16] = buffer_data_3[2111:2104];
        layer3[8][31:24] = buffer_data_3[2119:2112];
        layer3[8][39:32] = buffer_data_3[2127:2120];
        layer3[8][47:40] = buffer_data_3[2135:2128];
        layer3[8][55:48] = buffer_data_3[2143:2136];
        layer4[8][7:0] = buffer_data_2[2095:2088];
        layer4[8][15:8] = buffer_data_2[2103:2096];
        layer4[8][23:16] = buffer_data_2[2111:2104];
        layer4[8][31:24] = buffer_data_2[2119:2112];
        layer4[8][39:32] = buffer_data_2[2127:2120];
        layer4[8][47:40] = buffer_data_2[2135:2128];
        layer4[8][55:48] = buffer_data_2[2143:2136];
        layer5[8][7:0] = buffer_data_1[2095:2088];
        layer5[8][15:8] = buffer_data_1[2103:2096];
        layer5[8][23:16] = buffer_data_1[2111:2104];
        layer5[8][31:24] = buffer_data_1[2119:2112];
        layer5[8][39:32] = buffer_data_1[2127:2120];
        layer5[8][47:40] = buffer_data_1[2135:2128];
        layer5[8][55:48] = buffer_data_1[2143:2136];
        layer6[8][7:0] = buffer_data_0[2095:2088];
        layer6[8][15:8] = buffer_data_0[2103:2096];
        layer6[8][23:16] = buffer_data_0[2111:2104];
        layer6[8][31:24] = buffer_data_0[2119:2112];
        layer6[8][39:32] = buffer_data_0[2127:2120];
        layer6[8][47:40] = buffer_data_0[2135:2128];
        layer6[8][55:48] = buffer_data_0[2143:2136];
        layer0[9][7:0] = buffer_data_6[2103:2096];
        layer0[9][15:8] = buffer_data_6[2111:2104];
        layer0[9][23:16] = buffer_data_6[2119:2112];
        layer0[9][31:24] = buffer_data_6[2127:2120];
        layer0[9][39:32] = buffer_data_6[2135:2128];
        layer0[9][47:40] = buffer_data_6[2143:2136];
        layer0[9][55:48] = buffer_data_6[2151:2144];
        layer1[9][7:0] = buffer_data_5[2103:2096];
        layer1[9][15:8] = buffer_data_5[2111:2104];
        layer1[9][23:16] = buffer_data_5[2119:2112];
        layer1[9][31:24] = buffer_data_5[2127:2120];
        layer1[9][39:32] = buffer_data_5[2135:2128];
        layer1[9][47:40] = buffer_data_5[2143:2136];
        layer1[9][55:48] = buffer_data_5[2151:2144];
        layer2[9][7:0] = buffer_data_4[2103:2096];
        layer2[9][15:8] = buffer_data_4[2111:2104];
        layer2[9][23:16] = buffer_data_4[2119:2112];
        layer2[9][31:24] = buffer_data_4[2127:2120];
        layer2[9][39:32] = buffer_data_4[2135:2128];
        layer2[9][47:40] = buffer_data_4[2143:2136];
        layer2[9][55:48] = buffer_data_4[2151:2144];
        layer3[9][7:0] = buffer_data_3[2103:2096];
        layer3[9][15:8] = buffer_data_3[2111:2104];
        layer3[9][23:16] = buffer_data_3[2119:2112];
        layer3[9][31:24] = buffer_data_3[2127:2120];
        layer3[9][39:32] = buffer_data_3[2135:2128];
        layer3[9][47:40] = buffer_data_3[2143:2136];
        layer3[9][55:48] = buffer_data_3[2151:2144];
        layer4[9][7:0] = buffer_data_2[2103:2096];
        layer4[9][15:8] = buffer_data_2[2111:2104];
        layer4[9][23:16] = buffer_data_2[2119:2112];
        layer4[9][31:24] = buffer_data_2[2127:2120];
        layer4[9][39:32] = buffer_data_2[2135:2128];
        layer4[9][47:40] = buffer_data_2[2143:2136];
        layer4[9][55:48] = buffer_data_2[2151:2144];
        layer5[9][7:0] = buffer_data_1[2103:2096];
        layer5[9][15:8] = buffer_data_1[2111:2104];
        layer5[9][23:16] = buffer_data_1[2119:2112];
        layer5[9][31:24] = buffer_data_1[2127:2120];
        layer5[9][39:32] = buffer_data_1[2135:2128];
        layer5[9][47:40] = buffer_data_1[2143:2136];
        layer5[9][55:48] = buffer_data_1[2151:2144];
        layer6[9][7:0] = buffer_data_0[2103:2096];
        layer6[9][15:8] = buffer_data_0[2111:2104];
        layer6[9][23:16] = buffer_data_0[2119:2112];
        layer6[9][31:24] = buffer_data_0[2127:2120];
        layer6[9][39:32] = buffer_data_0[2135:2128];
        layer6[9][47:40] = buffer_data_0[2143:2136];
        layer6[9][55:48] = buffer_data_0[2151:2144];
        layer0[10][7:0] = buffer_data_6[2111:2104];
        layer0[10][15:8] = buffer_data_6[2119:2112];
        layer0[10][23:16] = buffer_data_6[2127:2120];
        layer0[10][31:24] = buffer_data_6[2135:2128];
        layer0[10][39:32] = buffer_data_6[2143:2136];
        layer0[10][47:40] = buffer_data_6[2151:2144];
        layer0[10][55:48] = buffer_data_6[2159:2152];
        layer1[10][7:0] = buffer_data_5[2111:2104];
        layer1[10][15:8] = buffer_data_5[2119:2112];
        layer1[10][23:16] = buffer_data_5[2127:2120];
        layer1[10][31:24] = buffer_data_5[2135:2128];
        layer1[10][39:32] = buffer_data_5[2143:2136];
        layer1[10][47:40] = buffer_data_5[2151:2144];
        layer1[10][55:48] = buffer_data_5[2159:2152];
        layer2[10][7:0] = buffer_data_4[2111:2104];
        layer2[10][15:8] = buffer_data_4[2119:2112];
        layer2[10][23:16] = buffer_data_4[2127:2120];
        layer2[10][31:24] = buffer_data_4[2135:2128];
        layer2[10][39:32] = buffer_data_4[2143:2136];
        layer2[10][47:40] = buffer_data_4[2151:2144];
        layer2[10][55:48] = buffer_data_4[2159:2152];
        layer3[10][7:0] = buffer_data_3[2111:2104];
        layer3[10][15:8] = buffer_data_3[2119:2112];
        layer3[10][23:16] = buffer_data_3[2127:2120];
        layer3[10][31:24] = buffer_data_3[2135:2128];
        layer3[10][39:32] = buffer_data_3[2143:2136];
        layer3[10][47:40] = buffer_data_3[2151:2144];
        layer3[10][55:48] = buffer_data_3[2159:2152];
        layer4[10][7:0] = buffer_data_2[2111:2104];
        layer4[10][15:8] = buffer_data_2[2119:2112];
        layer4[10][23:16] = buffer_data_2[2127:2120];
        layer4[10][31:24] = buffer_data_2[2135:2128];
        layer4[10][39:32] = buffer_data_2[2143:2136];
        layer4[10][47:40] = buffer_data_2[2151:2144];
        layer4[10][55:48] = buffer_data_2[2159:2152];
        layer5[10][7:0] = buffer_data_1[2111:2104];
        layer5[10][15:8] = buffer_data_1[2119:2112];
        layer5[10][23:16] = buffer_data_1[2127:2120];
        layer5[10][31:24] = buffer_data_1[2135:2128];
        layer5[10][39:32] = buffer_data_1[2143:2136];
        layer5[10][47:40] = buffer_data_1[2151:2144];
        layer5[10][55:48] = buffer_data_1[2159:2152];
        layer6[10][7:0] = buffer_data_0[2111:2104];
        layer6[10][15:8] = buffer_data_0[2119:2112];
        layer6[10][23:16] = buffer_data_0[2127:2120];
        layer6[10][31:24] = buffer_data_0[2135:2128];
        layer6[10][39:32] = buffer_data_0[2143:2136];
        layer6[10][47:40] = buffer_data_0[2151:2144];
        layer6[10][55:48] = buffer_data_0[2159:2152];
        layer0[11][7:0] = buffer_data_6[2119:2112];
        layer0[11][15:8] = buffer_data_6[2127:2120];
        layer0[11][23:16] = buffer_data_6[2135:2128];
        layer0[11][31:24] = buffer_data_6[2143:2136];
        layer0[11][39:32] = buffer_data_6[2151:2144];
        layer0[11][47:40] = buffer_data_6[2159:2152];
        layer0[11][55:48] = buffer_data_6[2167:2160];
        layer1[11][7:0] = buffer_data_5[2119:2112];
        layer1[11][15:8] = buffer_data_5[2127:2120];
        layer1[11][23:16] = buffer_data_5[2135:2128];
        layer1[11][31:24] = buffer_data_5[2143:2136];
        layer1[11][39:32] = buffer_data_5[2151:2144];
        layer1[11][47:40] = buffer_data_5[2159:2152];
        layer1[11][55:48] = buffer_data_5[2167:2160];
        layer2[11][7:0] = buffer_data_4[2119:2112];
        layer2[11][15:8] = buffer_data_4[2127:2120];
        layer2[11][23:16] = buffer_data_4[2135:2128];
        layer2[11][31:24] = buffer_data_4[2143:2136];
        layer2[11][39:32] = buffer_data_4[2151:2144];
        layer2[11][47:40] = buffer_data_4[2159:2152];
        layer2[11][55:48] = buffer_data_4[2167:2160];
        layer3[11][7:0] = buffer_data_3[2119:2112];
        layer3[11][15:8] = buffer_data_3[2127:2120];
        layer3[11][23:16] = buffer_data_3[2135:2128];
        layer3[11][31:24] = buffer_data_3[2143:2136];
        layer3[11][39:32] = buffer_data_3[2151:2144];
        layer3[11][47:40] = buffer_data_3[2159:2152];
        layer3[11][55:48] = buffer_data_3[2167:2160];
        layer4[11][7:0] = buffer_data_2[2119:2112];
        layer4[11][15:8] = buffer_data_2[2127:2120];
        layer4[11][23:16] = buffer_data_2[2135:2128];
        layer4[11][31:24] = buffer_data_2[2143:2136];
        layer4[11][39:32] = buffer_data_2[2151:2144];
        layer4[11][47:40] = buffer_data_2[2159:2152];
        layer4[11][55:48] = buffer_data_2[2167:2160];
        layer5[11][7:0] = buffer_data_1[2119:2112];
        layer5[11][15:8] = buffer_data_1[2127:2120];
        layer5[11][23:16] = buffer_data_1[2135:2128];
        layer5[11][31:24] = buffer_data_1[2143:2136];
        layer5[11][39:32] = buffer_data_1[2151:2144];
        layer5[11][47:40] = buffer_data_1[2159:2152];
        layer5[11][55:48] = buffer_data_1[2167:2160];
        layer6[11][7:0] = buffer_data_0[2119:2112];
        layer6[11][15:8] = buffer_data_0[2127:2120];
        layer6[11][23:16] = buffer_data_0[2135:2128];
        layer6[11][31:24] = buffer_data_0[2143:2136];
        layer6[11][39:32] = buffer_data_0[2151:2144];
        layer6[11][47:40] = buffer_data_0[2159:2152];
        layer6[11][55:48] = buffer_data_0[2167:2160];
        layer0[12][7:0] = buffer_data_6[2127:2120];
        layer0[12][15:8] = buffer_data_6[2135:2128];
        layer0[12][23:16] = buffer_data_6[2143:2136];
        layer0[12][31:24] = buffer_data_6[2151:2144];
        layer0[12][39:32] = buffer_data_6[2159:2152];
        layer0[12][47:40] = buffer_data_6[2167:2160];
        layer0[12][55:48] = buffer_data_6[2175:2168];
        layer1[12][7:0] = buffer_data_5[2127:2120];
        layer1[12][15:8] = buffer_data_5[2135:2128];
        layer1[12][23:16] = buffer_data_5[2143:2136];
        layer1[12][31:24] = buffer_data_5[2151:2144];
        layer1[12][39:32] = buffer_data_5[2159:2152];
        layer1[12][47:40] = buffer_data_5[2167:2160];
        layer1[12][55:48] = buffer_data_5[2175:2168];
        layer2[12][7:0] = buffer_data_4[2127:2120];
        layer2[12][15:8] = buffer_data_4[2135:2128];
        layer2[12][23:16] = buffer_data_4[2143:2136];
        layer2[12][31:24] = buffer_data_4[2151:2144];
        layer2[12][39:32] = buffer_data_4[2159:2152];
        layer2[12][47:40] = buffer_data_4[2167:2160];
        layer2[12][55:48] = buffer_data_4[2175:2168];
        layer3[12][7:0] = buffer_data_3[2127:2120];
        layer3[12][15:8] = buffer_data_3[2135:2128];
        layer3[12][23:16] = buffer_data_3[2143:2136];
        layer3[12][31:24] = buffer_data_3[2151:2144];
        layer3[12][39:32] = buffer_data_3[2159:2152];
        layer3[12][47:40] = buffer_data_3[2167:2160];
        layer3[12][55:48] = buffer_data_3[2175:2168];
        layer4[12][7:0] = buffer_data_2[2127:2120];
        layer4[12][15:8] = buffer_data_2[2135:2128];
        layer4[12][23:16] = buffer_data_2[2143:2136];
        layer4[12][31:24] = buffer_data_2[2151:2144];
        layer4[12][39:32] = buffer_data_2[2159:2152];
        layer4[12][47:40] = buffer_data_2[2167:2160];
        layer4[12][55:48] = buffer_data_2[2175:2168];
        layer5[12][7:0] = buffer_data_1[2127:2120];
        layer5[12][15:8] = buffer_data_1[2135:2128];
        layer5[12][23:16] = buffer_data_1[2143:2136];
        layer5[12][31:24] = buffer_data_1[2151:2144];
        layer5[12][39:32] = buffer_data_1[2159:2152];
        layer5[12][47:40] = buffer_data_1[2167:2160];
        layer5[12][55:48] = buffer_data_1[2175:2168];
        layer6[12][7:0] = buffer_data_0[2127:2120];
        layer6[12][15:8] = buffer_data_0[2135:2128];
        layer6[12][23:16] = buffer_data_0[2143:2136];
        layer6[12][31:24] = buffer_data_0[2151:2144];
        layer6[12][39:32] = buffer_data_0[2159:2152];
        layer6[12][47:40] = buffer_data_0[2167:2160];
        layer6[12][55:48] = buffer_data_0[2175:2168];
        layer0[13][7:0] = buffer_data_6[2135:2128];
        layer0[13][15:8] = buffer_data_6[2143:2136];
        layer0[13][23:16] = buffer_data_6[2151:2144];
        layer0[13][31:24] = buffer_data_6[2159:2152];
        layer0[13][39:32] = buffer_data_6[2167:2160];
        layer0[13][47:40] = buffer_data_6[2175:2168];
        layer0[13][55:48] = buffer_data_6[2183:2176];
        layer1[13][7:0] = buffer_data_5[2135:2128];
        layer1[13][15:8] = buffer_data_5[2143:2136];
        layer1[13][23:16] = buffer_data_5[2151:2144];
        layer1[13][31:24] = buffer_data_5[2159:2152];
        layer1[13][39:32] = buffer_data_5[2167:2160];
        layer1[13][47:40] = buffer_data_5[2175:2168];
        layer1[13][55:48] = buffer_data_5[2183:2176];
        layer2[13][7:0] = buffer_data_4[2135:2128];
        layer2[13][15:8] = buffer_data_4[2143:2136];
        layer2[13][23:16] = buffer_data_4[2151:2144];
        layer2[13][31:24] = buffer_data_4[2159:2152];
        layer2[13][39:32] = buffer_data_4[2167:2160];
        layer2[13][47:40] = buffer_data_4[2175:2168];
        layer2[13][55:48] = buffer_data_4[2183:2176];
        layer3[13][7:0] = buffer_data_3[2135:2128];
        layer3[13][15:8] = buffer_data_3[2143:2136];
        layer3[13][23:16] = buffer_data_3[2151:2144];
        layer3[13][31:24] = buffer_data_3[2159:2152];
        layer3[13][39:32] = buffer_data_3[2167:2160];
        layer3[13][47:40] = buffer_data_3[2175:2168];
        layer3[13][55:48] = buffer_data_3[2183:2176];
        layer4[13][7:0] = buffer_data_2[2135:2128];
        layer4[13][15:8] = buffer_data_2[2143:2136];
        layer4[13][23:16] = buffer_data_2[2151:2144];
        layer4[13][31:24] = buffer_data_2[2159:2152];
        layer4[13][39:32] = buffer_data_2[2167:2160];
        layer4[13][47:40] = buffer_data_2[2175:2168];
        layer4[13][55:48] = buffer_data_2[2183:2176];
        layer5[13][7:0] = buffer_data_1[2135:2128];
        layer5[13][15:8] = buffer_data_1[2143:2136];
        layer5[13][23:16] = buffer_data_1[2151:2144];
        layer5[13][31:24] = buffer_data_1[2159:2152];
        layer5[13][39:32] = buffer_data_1[2167:2160];
        layer5[13][47:40] = buffer_data_1[2175:2168];
        layer5[13][55:48] = buffer_data_1[2183:2176];
        layer6[13][7:0] = buffer_data_0[2135:2128];
        layer6[13][15:8] = buffer_data_0[2143:2136];
        layer6[13][23:16] = buffer_data_0[2151:2144];
        layer6[13][31:24] = buffer_data_0[2159:2152];
        layer6[13][39:32] = buffer_data_0[2167:2160];
        layer6[13][47:40] = buffer_data_0[2175:2168];
        layer6[13][55:48] = buffer_data_0[2183:2176];
        layer0[14][7:0] = buffer_data_6[2143:2136];
        layer0[14][15:8] = buffer_data_6[2151:2144];
        layer0[14][23:16] = buffer_data_6[2159:2152];
        layer0[14][31:24] = buffer_data_6[2167:2160];
        layer0[14][39:32] = buffer_data_6[2175:2168];
        layer0[14][47:40] = buffer_data_6[2183:2176];
        layer0[14][55:48] = buffer_data_6[2191:2184];
        layer1[14][7:0] = buffer_data_5[2143:2136];
        layer1[14][15:8] = buffer_data_5[2151:2144];
        layer1[14][23:16] = buffer_data_5[2159:2152];
        layer1[14][31:24] = buffer_data_5[2167:2160];
        layer1[14][39:32] = buffer_data_5[2175:2168];
        layer1[14][47:40] = buffer_data_5[2183:2176];
        layer1[14][55:48] = buffer_data_5[2191:2184];
        layer2[14][7:0] = buffer_data_4[2143:2136];
        layer2[14][15:8] = buffer_data_4[2151:2144];
        layer2[14][23:16] = buffer_data_4[2159:2152];
        layer2[14][31:24] = buffer_data_4[2167:2160];
        layer2[14][39:32] = buffer_data_4[2175:2168];
        layer2[14][47:40] = buffer_data_4[2183:2176];
        layer2[14][55:48] = buffer_data_4[2191:2184];
        layer3[14][7:0] = buffer_data_3[2143:2136];
        layer3[14][15:8] = buffer_data_3[2151:2144];
        layer3[14][23:16] = buffer_data_3[2159:2152];
        layer3[14][31:24] = buffer_data_3[2167:2160];
        layer3[14][39:32] = buffer_data_3[2175:2168];
        layer3[14][47:40] = buffer_data_3[2183:2176];
        layer3[14][55:48] = buffer_data_3[2191:2184];
        layer4[14][7:0] = buffer_data_2[2143:2136];
        layer4[14][15:8] = buffer_data_2[2151:2144];
        layer4[14][23:16] = buffer_data_2[2159:2152];
        layer4[14][31:24] = buffer_data_2[2167:2160];
        layer4[14][39:32] = buffer_data_2[2175:2168];
        layer4[14][47:40] = buffer_data_2[2183:2176];
        layer4[14][55:48] = buffer_data_2[2191:2184];
        layer5[14][7:0] = buffer_data_1[2143:2136];
        layer5[14][15:8] = buffer_data_1[2151:2144];
        layer5[14][23:16] = buffer_data_1[2159:2152];
        layer5[14][31:24] = buffer_data_1[2167:2160];
        layer5[14][39:32] = buffer_data_1[2175:2168];
        layer5[14][47:40] = buffer_data_1[2183:2176];
        layer5[14][55:48] = buffer_data_1[2191:2184];
        layer6[14][7:0] = buffer_data_0[2143:2136];
        layer6[14][15:8] = buffer_data_0[2151:2144];
        layer6[14][23:16] = buffer_data_0[2159:2152];
        layer6[14][31:24] = buffer_data_0[2167:2160];
        layer6[14][39:32] = buffer_data_0[2175:2168];
        layer6[14][47:40] = buffer_data_0[2183:2176];
        layer6[14][55:48] = buffer_data_0[2191:2184];
        layer0[15][7:0] = buffer_data_6[2151:2144];
        layer0[15][15:8] = buffer_data_6[2159:2152];
        layer0[15][23:16] = buffer_data_6[2167:2160];
        layer0[15][31:24] = buffer_data_6[2175:2168];
        layer0[15][39:32] = buffer_data_6[2183:2176];
        layer0[15][47:40] = buffer_data_6[2191:2184];
        layer0[15][55:48] = buffer_data_6[2199:2192];
        layer1[15][7:0] = buffer_data_5[2151:2144];
        layer1[15][15:8] = buffer_data_5[2159:2152];
        layer1[15][23:16] = buffer_data_5[2167:2160];
        layer1[15][31:24] = buffer_data_5[2175:2168];
        layer1[15][39:32] = buffer_data_5[2183:2176];
        layer1[15][47:40] = buffer_data_5[2191:2184];
        layer1[15][55:48] = buffer_data_5[2199:2192];
        layer2[15][7:0] = buffer_data_4[2151:2144];
        layer2[15][15:8] = buffer_data_4[2159:2152];
        layer2[15][23:16] = buffer_data_4[2167:2160];
        layer2[15][31:24] = buffer_data_4[2175:2168];
        layer2[15][39:32] = buffer_data_4[2183:2176];
        layer2[15][47:40] = buffer_data_4[2191:2184];
        layer2[15][55:48] = buffer_data_4[2199:2192];
        layer3[15][7:0] = buffer_data_3[2151:2144];
        layer3[15][15:8] = buffer_data_3[2159:2152];
        layer3[15][23:16] = buffer_data_3[2167:2160];
        layer3[15][31:24] = buffer_data_3[2175:2168];
        layer3[15][39:32] = buffer_data_3[2183:2176];
        layer3[15][47:40] = buffer_data_3[2191:2184];
        layer3[15][55:48] = buffer_data_3[2199:2192];
        layer4[15][7:0] = buffer_data_2[2151:2144];
        layer4[15][15:8] = buffer_data_2[2159:2152];
        layer4[15][23:16] = buffer_data_2[2167:2160];
        layer4[15][31:24] = buffer_data_2[2175:2168];
        layer4[15][39:32] = buffer_data_2[2183:2176];
        layer4[15][47:40] = buffer_data_2[2191:2184];
        layer4[15][55:48] = buffer_data_2[2199:2192];
        layer5[15][7:0] = buffer_data_1[2151:2144];
        layer5[15][15:8] = buffer_data_1[2159:2152];
        layer5[15][23:16] = buffer_data_1[2167:2160];
        layer5[15][31:24] = buffer_data_1[2175:2168];
        layer5[15][39:32] = buffer_data_1[2183:2176];
        layer5[15][47:40] = buffer_data_1[2191:2184];
        layer5[15][55:48] = buffer_data_1[2199:2192];
        layer6[15][7:0] = buffer_data_0[2151:2144];
        layer6[15][15:8] = buffer_data_0[2159:2152];
        layer6[15][23:16] = buffer_data_0[2167:2160];
        layer6[15][31:24] = buffer_data_0[2175:2168];
        layer6[15][39:32] = buffer_data_0[2183:2176];
        layer6[15][47:40] = buffer_data_0[2191:2184];
        layer6[15][55:48] = buffer_data_0[2199:2192];
        layer0[16][7:0] = buffer_data_6[2159:2152];
        layer0[16][15:8] = buffer_data_6[2167:2160];
        layer0[16][23:16] = buffer_data_6[2175:2168];
        layer0[16][31:24] = buffer_data_6[2183:2176];
        layer0[16][39:32] = buffer_data_6[2191:2184];
        layer0[16][47:40] = buffer_data_6[2199:2192];
        layer0[16][55:48] = buffer_data_6[2207:2200];
        layer1[16][7:0] = buffer_data_5[2159:2152];
        layer1[16][15:8] = buffer_data_5[2167:2160];
        layer1[16][23:16] = buffer_data_5[2175:2168];
        layer1[16][31:24] = buffer_data_5[2183:2176];
        layer1[16][39:32] = buffer_data_5[2191:2184];
        layer1[16][47:40] = buffer_data_5[2199:2192];
        layer1[16][55:48] = buffer_data_5[2207:2200];
        layer2[16][7:0] = buffer_data_4[2159:2152];
        layer2[16][15:8] = buffer_data_4[2167:2160];
        layer2[16][23:16] = buffer_data_4[2175:2168];
        layer2[16][31:24] = buffer_data_4[2183:2176];
        layer2[16][39:32] = buffer_data_4[2191:2184];
        layer2[16][47:40] = buffer_data_4[2199:2192];
        layer2[16][55:48] = buffer_data_4[2207:2200];
        layer3[16][7:0] = buffer_data_3[2159:2152];
        layer3[16][15:8] = buffer_data_3[2167:2160];
        layer3[16][23:16] = buffer_data_3[2175:2168];
        layer3[16][31:24] = buffer_data_3[2183:2176];
        layer3[16][39:32] = buffer_data_3[2191:2184];
        layer3[16][47:40] = buffer_data_3[2199:2192];
        layer3[16][55:48] = buffer_data_3[2207:2200];
        layer4[16][7:0] = buffer_data_2[2159:2152];
        layer4[16][15:8] = buffer_data_2[2167:2160];
        layer4[16][23:16] = buffer_data_2[2175:2168];
        layer4[16][31:24] = buffer_data_2[2183:2176];
        layer4[16][39:32] = buffer_data_2[2191:2184];
        layer4[16][47:40] = buffer_data_2[2199:2192];
        layer4[16][55:48] = buffer_data_2[2207:2200];
        layer5[16][7:0] = buffer_data_1[2159:2152];
        layer5[16][15:8] = buffer_data_1[2167:2160];
        layer5[16][23:16] = buffer_data_1[2175:2168];
        layer5[16][31:24] = buffer_data_1[2183:2176];
        layer5[16][39:32] = buffer_data_1[2191:2184];
        layer5[16][47:40] = buffer_data_1[2199:2192];
        layer5[16][55:48] = buffer_data_1[2207:2200];
        layer6[16][7:0] = buffer_data_0[2159:2152];
        layer6[16][15:8] = buffer_data_0[2167:2160];
        layer6[16][23:16] = buffer_data_0[2175:2168];
        layer6[16][31:24] = buffer_data_0[2183:2176];
        layer6[16][39:32] = buffer_data_0[2191:2184];
        layer6[16][47:40] = buffer_data_0[2199:2192];
        layer6[16][55:48] = buffer_data_0[2207:2200];
        layer0[17][7:0] = buffer_data_6[2167:2160];
        layer0[17][15:8] = buffer_data_6[2175:2168];
        layer0[17][23:16] = buffer_data_6[2183:2176];
        layer0[17][31:24] = buffer_data_6[2191:2184];
        layer0[17][39:32] = buffer_data_6[2199:2192];
        layer0[17][47:40] = buffer_data_6[2207:2200];
        layer0[17][55:48] = buffer_data_6[2215:2208];
        layer1[17][7:0] = buffer_data_5[2167:2160];
        layer1[17][15:8] = buffer_data_5[2175:2168];
        layer1[17][23:16] = buffer_data_5[2183:2176];
        layer1[17][31:24] = buffer_data_5[2191:2184];
        layer1[17][39:32] = buffer_data_5[2199:2192];
        layer1[17][47:40] = buffer_data_5[2207:2200];
        layer1[17][55:48] = buffer_data_5[2215:2208];
        layer2[17][7:0] = buffer_data_4[2167:2160];
        layer2[17][15:8] = buffer_data_4[2175:2168];
        layer2[17][23:16] = buffer_data_4[2183:2176];
        layer2[17][31:24] = buffer_data_4[2191:2184];
        layer2[17][39:32] = buffer_data_4[2199:2192];
        layer2[17][47:40] = buffer_data_4[2207:2200];
        layer2[17][55:48] = buffer_data_4[2215:2208];
        layer3[17][7:0] = buffer_data_3[2167:2160];
        layer3[17][15:8] = buffer_data_3[2175:2168];
        layer3[17][23:16] = buffer_data_3[2183:2176];
        layer3[17][31:24] = buffer_data_3[2191:2184];
        layer3[17][39:32] = buffer_data_3[2199:2192];
        layer3[17][47:40] = buffer_data_3[2207:2200];
        layer3[17][55:48] = buffer_data_3[2215:2208];
        layer4[17][7:0] = buffer_data_2[2167:2160];
        layer4[17][15:8] = buffer_data_2[2175:2168];
        layer4[17][23:16] = buffer_data_2[2183:2176];
        layer4[17][31:24] = buffer_data_2[2191:2184];
        layer4[17][39:32] = buffer_data_2[2199:2192];
        layer4[17][47:40] = buffer_data_2[2207:2200];
        layer4[17][55:48] = buffer_data_2[2215:2208];
        layer5[17][7:0] = buffer_data_1[2167:2160];
        layer5[17][15:8] = buffer_data_1[2175:2168];
        layer5[17][23:16] = buffer_data_1[2183:2176];
        layer5[17][31:24] = buffer_data_1[2191:2184];
        layer5[17][39:32] = buffer_data_1[2199:2192];
        layer5[17][47:40] = buffer_data_1[2207:2200];
        layer5[17][55:48] = buffer_data_1[2215:2208];
        layer6[17][7:0] = buffer_data_0[2167:2160];
        layer6[17][15:8] = buffer_data_0[2175:2168];
        layer6[17][23:16] = buffer_data_0[2183:2176];
        layer6[17][31:24] = buffer_data_0[2191:2184];
        layer6[17][39:32] = buffer_data_0[2199:2192];
        layer6[17][47:40] = buffer_data_0[2207:2200];
        layer6[17][55:48] = buffer_data_0[2215:2208];
        layer0[18][7:0] = buffer_data_6[2175:2168];
        layer0[18][15:8] = buffer_data_6[2183:2176];
        layer0[18][23:16] = buffer_data_6[2191:2184];
        layer0[18][31:24] = buffer_data_6[2199:2192];
        layer0[18][39:32] = buffer_data_6[2207:2200];
        layer0[18][47:40] = buffer_data_6[2215:2208];
        layer0[18][55:48] = buffer_data_6[2223:2216];
        layer1[18][7:0] = buffer_data_5[2175:2168];
        layer1[18][15:8] = buffer_data_5[2183:2176];
        layer1[18][23:16] = buffer_data_5[2191:2184];
        layer1[18][31:24] = buffer_data_5[2199:2192];
        layer1[18][39:32] = buffer_data_5[2207:2200];
        layer1[18][47:40] = buffer_data_5[2215:2208];
        layer1[18][55:48] = buffer_data_5[2223:2216];
        layer2[18][7:0] = buffer_data_4[2175:2168];
        layer2[18][15:8] = buffer_data_4[2183:2176];
        layer2[18][23:16] = buffer_data_4[2191:2184];
        layer2[18][31:24] = buffer_data_4[2199:2192];
        layer2[18][39:32] = buffer_data_4[2207:2200];
        layer2[18][47:40] = buffer_data_4[2215:2208];
        layer2[18][55:48] = buffer_data_4[2223:2216];
        layer3[18][7:0] = buffer_data_3[2175:2168];
        layer3[18][15:8] = buffer_data_3[2183:2176];
        layer3[18][23:16] = buffer_data_3[2191:2184];
        layer3[18][31:24] = buffer_data_3[2199:2192];
        layer3[18][39:32] = buffer_data_3[2207:2200];
        layer3[18][47:40] = buffer_data_3[2215:2208];
        layer3[18][55:48] = buffer_data_3[2223:2216];
        layer4[18][7:0] = buffer_data_2[2175:2168];
        layer4[18][15:8] = buffer_data_2[2183:2176];
        layer4[18][23:16] = buffer_data_2[2191:2184];
        layer4[18][31:24] = buffer_data_2[2199:2192];
        layer4[18][39:32] = buffer_data_2[2207:2200];
        layer4[18][47:40] = buffer_data_2[2215:2208];
        layer4[18][55:48] = buffer_data_2[2223:2216];
        layer5[18][7:0] = buffer_data_1[2175:2168];
        layer5[18][15:8] = buffer_data_1[2183:2176];
        layer5[18][23:16] = buffer_data_1[2191:2184];
        layer5[18][31:24] = buffer_data_1[2199:2192];
        layer5[18][39:32] = buffer_data_1[2207:2200];
        layer5[18][47:40] = buffer_data_1[2215:2208];
        layer5[18][55:48] = buffer_data_1[2223:2216];
        layer6[18][7:0] = buffer_data_0[2175:2168];
        layer6[18][15:8] = buffer_data_0[2183:2176];
        layer6[18][23:16] = buffer_data_0[2191:2184];
        layer6[18][31:24] = buffer_data_0[2199:2192];
        layer6[18][39:32] = buffer_data_0[2207:2200];
        layer6[18][47:40] = buffer_data_0[2215:2208];
        layer6[18][55:48] = buffer_data_0[2223:2216];
        layer0[19][7:0] = buffer_data_6[2183:2176];
        layer0[19][15:8] = buffer_data_6[2191:2184];
        layer0[19][23:16] = buffer_data_6[2199:2192];
        layer0[19][31:24] = buffer_data_6[2207:2200];
        layer0[19][39:32] = buffer_data_6[2215:2208];
        layer0[19][47:40] = buffer_data_6[2223:2216];
        layer0[19][55:48] = buffer_data_6[2231:2224];
        layer1[19][7:0] = buffer_data_5[2183:2176];
        layer1[19][15:8] = buffer_data_5[2191:2184];
        layer1[19][23:16] = buffer_data_5[2199:2192];
        layer1[19][31:24] = buffer_data_5[2207:2200];
        layer1[19][39:32] = buffer_data_5[2215:2208];
        layer1[19][47:40] = buffer_data_5[2223:2216];
        layer1[19][55:48] = buffer_data_5[2231:2224];
        layer2[19][7:0] = buffer_data_4[2183:2176];
        layer2[19][15:8] = buffer_data_4[2191:2184];
        layer2[19][23:16] = buffer_data_4[2199:2192];
        layer2[19][31:24] = buffer_data_4[2207:2200];
        layer2[19][39:32] = buffer_data_4[2215:2208];
        layer2[19][47:40] = buffer_data_4[2223:2216];
        layer2[19][55:48] = buffer_data_4[2231:2224];
        layer3[19][7:0] = buffer_data_3[2183:2176];
        layer3[19][15:8] = buffer_data_3[2191:2184];
        layer3[19][23:16] = buffer_data_3[2199:2192];
        layer3[19][31:24] = buffer_data_3[2207:2200];
        layer3[19][39:32] = buffer_data_3[2215:2208];
        layer3[19][47:40] = buffer_data_3[2223:2216];
        layer3[19][55:48] = buffer_data_3[2231:2224];
        layer4[19][7:0] = buffer_data_2[2183:2176];
        layer4[19][15:8] = buffer_data_2[2191:2184];
        layer4[19][23:16] = buffer_data_2[2199:2192];
        layer4[19][31:24] = buffer_data_2[2207:2200];
        layer4[19][39:32] = buffer_data_2[2215:2208];
        layer4[19][47:40] = buffer_data_2[2223:2216];
        layer4[19][55:48] = buffer_data_2[2231:2224];
        layer5[19][7:0] = buffer_data_1[2183:2176];
        layer5[19][15:8] = buffer_data_1[2191:2184];
        layer5[19][23:16] = buffer_data_1[2199:2192];
        layer5[19][31:24] = buffer_data_1[2207:2200];
        layer5[19][39:32] = buffer_data_1[2215:2208];
        layer5[19][47:40] = buffer_data_1[2223:2216];
        layer5[19][55:48] = buffer_data_1[2231:2224];
        layer6[19][7:0] = buffer_data_0[2183:2176];
        layer6[19][15:8] = buffer_data_0[2191:2184];
        layer6[19][23:16] = buffer_data_0[2199:2192];
        layer6[19][31:24] = buffer_data_0[2207:2200];
        layer6[19][39:32] = buffer_data_0[2215:2208];
        layer6[19][47:40] = buffer_data_0[2223:2216];
        layer6[19][55:48] = buffer_data_0[2231:2224];
        layer0[20][7:0] = buffer_data_6[2191:2184];
        layer0[20][15:8] = buffer_data_6[2199:2192];
        layer0[20][23:16] = buffer_data_6[2207:2200];
        layer0[20][31:24] = buffer_data_6[2215:2208];
        layer0[20][39:32] = buffer_data_6[2223:2216];
        layer0[20][47:40] = buffer_data_6[2231:2224];
        layer0[20][55:48] = buffer_data_6[2239:2232];
        layer1[20][7:0] = buffer_data_5[2191:2184];
        layer1[20][15:8] = buffer_data_5[2199:2192];
        layer1[20][23:16] = buffer_data_5[2207:2200];
        layer1[20][31:24] = buffer_data_5[2215:2208];
        layer1[20][39:32] = buffer_data_5[2223:2216];
        layer1[20][47:40] = buffer_data_5[2231:2224];
        layer1[20][55:48] = buffer_data_5[2239:2232];
        layer2[20][7:0] = buffer_data_4[2191:2184];
        layer2[20][15:8] = buffer_data_4[2199:2192];
        layer2[20][23:16] = buffer_data_4[2207:2200];
        layer2[20][31:24] = buffer_data_4[2215:2208];
        layer2[20][39:32] = buffer_data_4[2223:2216];
        layer2[20][47:40] = buffer_data_4[2231:2224];
        layer2[20][55:48] = buffer_data_4[2239:2232];
        layer3[20][7:0] = buffer_data_3[2191:2184];
        layer3[20][15:8] = buffer_data_3[2199:2192];
        layer3[20][23:16] = buffer_data_3[2207:2200];
        layer3[20][31:24] = buffer_data_3[2215:2208];
        layer3[20][39:32] = buffer_data_3[2223:2216];
        layer3[20][47:40] = buffer_data_3[2231:2224];
        layer3[20][55:48] = buffer_data_3[2239:2232];
        layer4[20][7:0] = buffer_data_2[2191:2184];
        layer4[20][15:8] = buffer_data_2[2199:2192];
        layer4[20][23:16] = buffer_data_2[2207:2200];
        layer4[20][31:24] = buffer_data_2[2215:2208];
        layer4[20][39:32] = buffer_data_2[2223:2216];
        layer4[20][47:40] = buffer_data_2[2231:2224];
        layer4[20][55:48] = buffer_data_2[2239:2232];
        layer5[20][7:0] = buffer_data_1[2191:2184];
        layer5[20][15:8] = buffer_data_1[2199:2192];
        layer5[20][23:16] = buffer_data_1[2207:2200];
        layer5[20][31:24] = buffer_data_1[2215:2208];
        layer5[20][39:32] = buffer_data_1[2223:2216];
        layer5[20][47:40] = buffer_data_1[2231:2224];
        layer5[20][55:48] = buffer_data_1[2239:2232];
        layer6[20][7:0] = buffer_data_0[2191:2184];
        layer6[20][15:8] = buffer_data_0[2199:2192];
        layer6[20][23:16] = buffer_data_0[2207:2200];
        layer6[20][31:24] = buffer_data_0[2215:2208];
        layer6[20][39:32] = buffer_data_0[2223:2216];
        layer6[20][47:40] = buffer_data_0[2231:2224];
        layer6[20][55:48] = buffer_data_0[2239:2232];
        layer0[21][7:0] = buffer_data_6[2199:2192];
        layer0[21][15:8] = buffer_data_6[2207:2200];
        layer0[21][23:16] = buffer_data_6[2215:2208];
        layer0[21][31:24] = buffer_data_6[2223:2216];
        layer0[21][39:32] = buffer_data_6[2231:2224];
        layer0[21][47:40] = buffer_data_6[2239:2232];
        layer0[21][55:48] = buffer_data_6[2247:2240];
        layer1[21][7:0] = buffer_data_5[2199:2192];
        layer1[21][15:8] = buffer_data_5[2207:2200];
        layer1[21][23:16] = buffer_data_5[2215:2208];
        layer1[21][31:24] = buffer_data_5[2223:2216];
        layer1[21][39:32] = buffer_data_5[2231:2224];
        layer1[21][47:40] = buffer_data_5[2239:2232];
        layer1[21][55:48] = buffer_data_5[2247:2240];
        layer2[21][7:0] = buffer_data_4[2199:2192];
        layer2[21][15:8] = buffer_data_4[2207:2200];
        layer2[21][23:16] = buffer_data_4[2215:2208];
        layer2[21][31:24] = buffer_data_4[2223:2216];
        layer2[21][39:32] = buffer_data_4[2231:2224];
        layer2[21][47:40] = buffer_data_4[2239:2232];
        layer2[21][55:48] = buffer_data_4[2247:2240];
        layer3[21][7:0] = buffer_data_3[2199:2192];
        layer3[21][15:8] = buffer_data_3[2207:2200];
        layer3[21][23:16] = buffer_data_3[2215:2208];
        layer3[21][31:24] = buffer_data_3[2223:2216];
        layer3[21][39:32] = buffer_data_3[2231:2224];
        layer3[21][47:40] = buffer_data_3[2239:2232];
        layer3[21][55:48] = buffer_data_3[2247:2240];
        layer4[21][7:0] = buffer_data_2[2199:2192];
        layer4[21][15:8] = buffer_data_2[2207:2200];
        layer4[21][23:16] = buffer_data_2[2215:2208];
        layer4[21][31:24] = buffer_data_2[2223:2216];
        layer4[21][39:32] = buffer_data_2[2231:2224];
        layer4[21][47:40] = buffer_data_2[2239:2232];
        layer4[21][55:48] = buffer_data_2[2247:2240];
        layer5[21][7:0] = buffer_data_1[2199:2192];
        layer5[21][15:8] = buffer_data_1[2207:2200];
        layer5[21][23:16] = buffer_data_1[2215:2208];
        layer5[21][31:24] = buffer_data_1[2223:2216];
        layer5[21][39:32] = buffer_data_1[2231:2224];
        layer5[21][47:40] = buffer_data_1[2239:2232];
        layer5[21][55:48] = buffer_data_1[2247:2240];
        layer6[21][7:0] = buffer_data_0[2199:2192];
        layer6[21][15:8] = buffer_data_0[2207:2200];
        layer6[21][23:16] = buffer_data_0[2215:2208];
        layer6[21][31:24] = buffer_data_0[2223:2216];
        layer6[21][39:32] = buffer_data_0[2231:2224];
        layer6[21][47:40] = buffer_data_0[2239:2232];
        layer6[21][55:48] = buffer_data_0[2247:2240];
        layer0[22][7:0] = buffer_data_6[2207:2200];
        layer0[22][15:8] = buffer_data_6[2215:2208];
        layer0[22][23:16] = buffer_data_6[2223:2216];
        layer0[22][31:24] = buffer_data_6[2231:2224];
        layer0[22][39:32] = buffer_data_6[2239:2232];
        layer0[22][47:40] = buffer_data_6[2247:2240];
        layer0[22][55:48] = buffer_data_6[2255:2248];
        layer1[22][7:0] = buffer_data_5[2207:2200];
        layer1[22][15:8] = buffer_data_5[2215:2208];
        layer1[22][23:16] = buffer_data_5[2223:2216];
        layer1[22][31:24] = buffer_data_5[2231:2224];
        layer1[22][39:32] = buffer_data_5[2239:2232];
        layer1[22][47:40] = buffer_data_5[2247:2240];
        layer1[22][55:48] = buffer_data_5[2255:2248];
        layer2[22][7:0] = buffer_data_4[2207:2200];
        layer2[22][15:8] = buffer_data_4[2215:2208];
        layer2[22][23:16] = buffer_data_4[2223:2216];
        layer2[22][31:24] = buffer_data_4[2231:2224];
        layer2[22][39:32] = buffer_data_4[2239:2232];
        layer2[22][47:40] = buffer_data_4[2247:2240];
        layer2[22][55:48] = buffer_data_4[2255:2248];
        layer3[22][7:0] = buffer_data_3[2207:2200];
        layer3[22][15:8] = buffer_data_3[2215:2208];
        layer3[22][23:16] = buffer_data_3[2223:2216];
        layer3[22][31:24] = buffer_data_3[2231:2224];
        layer3[22][39:32] = buffer_data_3[2239:2232];
        layer3[22][47:40] = buffer_data_3[2247:2240];
        layer3[22][55:48] = buffer_data_3[2255:2248];
        layer4[22][7:0] = buffer_data_2[2207:2200];
        layer4[22][15:8] = buffer_data_2[2215:2208];
        layer4[22][23:16] = buffer_data_2[2223:2216];
        layer4[22][31:24] = buffer_data_2[2231:2224];
        layer4[22][39:32] = buffer_data_2[2239:2232];
        layer4[22][47:40] = buffer_data_2[2247:2240];
        layer4[22][55:48] = buffer_data_2[2255:2248];
        layer5[22][7:0] = buffer_data_1[2207:2200];
        layer5[22][15:8] = buffer_data_1[2215:2208];
        layer5[22][23:16] = buffer_data_1[2223:2216];
        layer5[22][31:24] = buffer_data_1[2231:2224];
        layer5[22][39:32] = buffer_data_1[2239:2232];
        layer5[22][47:40] = buffer_data_1[2247:2240];
        layer5[22][55:48] = buffer_data_1[2255:2248];
        layer6[22][7:0] = buffer_data_0[2207:2200];
        layer6[22][15:8] = buffer_data_0[2215:2208];
        layer6[22][23:16] = buffer_data_0[2223:2216];
        layer6[22][31:24] = buffer_data_0[2231:2224];
        layer6[22][39:32] = buffer_data_0[2239:2232];
        layer6[22][47:40] = buffer_data_0[2247:2240];
        layer6[22][55:48] = buffer_data_0[2255:2248];
        layer0[23][7:0] = buffer_data_6[2215:2208];
        layer0[23][15:8] = buffer_data_6[2223:2216];
        layer0[23][23:16] = buffer_data_6[2231:2224];
        layer0[23][31:24] = buffer_data_6[2239:2232];
        layer0[23][39:32] = buffer_data_6[2247:2240];
        layer0[23][47:40] = buffer_data_6[2255:2248];
        layer0[23][55:48] = buffer_data_6[2263:2256];
        layer1[23][7:0] = buffer_data_5[2215:2208];
        layer1[23][15:8] = buffer_data_5[2223:2216];
        layer1[23][23:16] = buffer_data_5[2231:2224];
        layer1[23][31:24] = buffer_data_5[2239:2232];
        layer1[23][39:32] = buffer_data_5[2247:2240];
        layer1[23][47:40] = buffer_data_5[2255:2248];
        layer1[23][55:48] = buffer_data_5[2263:2256];
        layer2[23][7:0] = buffer_data_4[2215:2208];
        layer2[23][15:8] = buffer_data_4[2223:2216];
        layer2[23][23:16] = buffer_data_4[2231:2224];
        layer2[23][31:24] = buffer_data_4[2239:2232];
        layer2[23][39:32] = buffer_data_4[2247:2240];
        layer2[23][47:40] = buffer_data_4[2255:2248];
        layer2[23][55:48] = buffer_data_4[2263:2256];
        layer3[23][7:0] = buffer_data_3[2215:2208];
        layer3[23][15:8] = buffer_data_3[2223:2216];
        layer3[23][23:16] = buffer_data_3[2231:2224];
        layer3[23][31:24] = buffer_data_3[2239:2232];
        layer3[23][39:32] = buffer_data_3[2247:2240];
        layer3[23][47:40] = buffer_data_3[2255:2248];
        layer3[23][55:48] = buffer_data_3[2263:2256];
        layer4[23][7:0] = buffer_data_2[2215:2208];
        layer4[23][15:8] = buffer_data_2[2223:2216];
        layer4[23][23:16] = buffer_data_2[2231:2224];
        layer4[23][31:24] = buffer_data_2[2239:2232];
        layer4[23][39:32] = buffer_data_2[2247:2240];
        layer4[23][47:40] = buffer_data_2[2255:2248];
        layer4[23][55:48] = buffer_data_2[2263:2256];
        layer5[23][7:0] = buffer_data_1[2215:2208];
        layer5[23][15:8] = buffer_data_1[2223:2216];
        layer5[23][23:16] = buffer_data_1[2231:2224];
        layer5[23][31:24] = buffer_data_1[2239:2232];
        layer5[23][39:32] = buffer_data_1[2247:2240];
        layer5[23][47:40] = buffer_data_1[2255:2248];
        layer5[23][55:48] = buffer_data_1[2263:2256];
        layer6[23][7:0] = buffer_data_0[2215:2208];
        layer6[23][15:8] = buffer_data_0[2223:2216];
        layer6[23][23:16] = buffer_data_0[2231:2224];
        layer6[23][31:24] = buffer_data_0[2239:2232];
        layer6[23][39:32] = buffer_data_0[2247:2240];
        layer6[23][47:40] = buffer_data_0[2255:2248];
        layer6[23][55:48] = buffer_data_0[2263:2256];
        layer0[24][7:0] = buffer_data_6[2223:2216];
        layer0[24][15:8] = buffer_data_6[2231:2224];
        layer0[24][23:16] = buffer_data_6[2239:2232];
        layer0[24][31:24] = buffer_data_6[2247:2240];
        layer0[24][39:32] = buffer_data_6[2255:2248];
        layer0[24][47:40] = buffer_data_6[2263:2256];
        layer0[24][55:48] = buffer_data_6[2271:2264];
        layer1[24][7:0] = buffer_data_5[2223:2216];
        layer1[24][15:8] = buffer_data_5[2231:2224];
        layer1[24][23:16] = buffer_data_5[2239:2232];
        layer1[24][31:24] = buffer_data_5[2247:2240];
        layer1[24][39:32] = buffer_data_5[2255:2248];
        layer1[24][47:40] = buffer_data_5[2263:2256];
        layer1[24][55:48] = buffer_data_5[2271:2264];
        layer2[24][7:0] = buffer_data_4[2223:2216];
        layer2[24][15:8] = buffer_data_4[2231:2224];
        layer2[24][23:16] = buffer_data_4[2239:2232];
        layer2[24][31:24] = buffer_data_4[2247:2240];
        layer2[24][39:32] = buffer_data_4[2255:2248];
        layer2[24][47:40] = buffer_data_4[2263:2256];
        layer2[24][55:48] = buffer_data_4[2271:2264];
        layer3[24][7:0] = buffer_data_3[2223:2216];
        layer3[24][15:8] = buffer_data_3[2231:2224];
        layer3[24][23:16] = buffer_data_3[2239:2232];
        layer3[24][31:24] = buffer_data_3[2247:2240];
        layer3[24][39:32] = buffer_data_3[2255:2248];
        layer3[24][47:40] = buffer_data_3[2263:2256];
        layer3[24][55:48] = buffer_data_3[2271:2264];
        layer4[24][7:0] = buffer_data_2[2223:2216];
        layer4[24][15:8] = buffer_data_2[2231:2224];
        layer4[24][23:16] = buffer_data_2[2239:2232];
        layer4[24][31:24] = buffer_data_2[2247:2240];
        layer4[24][39:32] = buffer_data_2[2255:2248];
        layer4[24][47:40] = buffer_data_2[2263:2256];
        layer4[24][55:48] = buffer_data_2[2271:2264];
        layer5[24][7:0] = buffer_data_1[2223:2216];
        layer5[24][15:8] = buffer_data_1[2231:2224];
        layer5[24][23:16] = buffer_data_1[2239:2232];
        layer5[24][31:24] = buffer_data_1[2247:2240];
        layer5[24][39:32] = buffer_data_1[2255:2248];
        layer5[24][47:40] = buffer_data_1[2263:2256];
        layer5[24][55:48] = buffer_data_1[2271:2264];
        layer6[24][7:0] = buffer_data_0[2223:2216];
        layer6[24][15:8] = buffer_data_0[2231:2224];
        layer6[24][23:16] = buffer_data_0[2239:2232];
        layer6[24][31:24] = buffer_data_0[2247:2240];
        layer6[24][39:32] = buffer_data_0[2255:2248];
        layer6[24][47:40] = buffer_data_0[2263:2256];
        layer6[24][55:48] = buffer_data_0[2271:2264];
        layer0[25][7:0] = buffer_data_6[2231:2224];
        layer0[25][15:8] = buffer_data_6[2239:2232];
        layer0[25][23:16] = buffer_data_6[2247:2240];
        layer0[25][31:24] = buffer_data_6[2255:2248];
        layer0[25][39:32] = buffer_data_6[2263:2256];
        layer0[25][47:40] = buffer_data_6[2271:2264];
        layer0[25][55:48] = buffer_data_6[2279:2272];
        layer1[25][7:0] = buffer_data_5[2231:2224];
        layer1[25][15:8] = buffer_data_5[2239:2232];
        layer1[25][23:16] = buffer_data_5[2247:2240];
        layer1[25][31:24] = buffer_data_5[2255:2248];
        layer1[25][39:32] = buffer_data_5[2263:2256];
        layer1[25][47:40] = buffer_data_5[2271:2264];
        layer1[25][55:48] = buffer_data_5[2279:2272];
        layer2[25][7:0] = buffer_data_4[2231:2224];
        layer2[25][15:8] = buffer_data_4[2239:2232];
        layer2[25][23:16] = buffer_data_4[2247:2240];
        layer2[25][31:24] = buffer_data_4[2255:2248];
        layer2[25][39:32] = buffer_data_4[2263:2256];
        layer2[25][47:40] = buffer_data_4[2271:2264];
        layer2[25][55:48] = buffer_data_4[2279:2272];
        layer3[25][7:0] = buffer_data_3[2231:2224];
        layer3[25][15:8] = buffer_data_3[2239:2232];
        layer3[25][23:16] = buffer_data_3[2247:2240];
        layer3[25][31:24] = buffer_data_3[2255:2248];
        layer3[25][39:32] = buffer_data_3[2263:2256];
        layer3[25][47:40] = buffer_data_3[2271:2264];
        layer3[25][55:48] = buffer_data_3[2279:2272];
        layer4[25][7:0] = buffer_data_2[2231:2224];
        layer4[25][15:8] = buffer_data_2[2239:2232];
        layer4[25][23:16] = buffer_data_2[2247:2240];
        layer4[25][31:24] = buffer_data_2[2255:2248];
        layer4[25][39:32] = buffer_data_2[2263:2256];
        layer4[25][47:40] = buffer_data_2[2271:2264];
        layer4[25][55:48] = buffer_data_2[2279:2272];
        layer5[25][7:0] = buffer_data_1[2231:2224];
        layer5[25][15:8] = buffer_data_1[2239:2232];
        layer5[25][23:16] = buffer_data_1[2247:2240];
        layer5[25][31:24] = buffer_data_1[2255:2248];
        layer5[25][39:32] = buffer_data_1[2263:2256];
        layer5[25][47:40] = buffer_data_1[2271:2264];
        layer5[25][55:48] = buffer_data_1[2279:2272];
        layer6[25][7:0] = buffer_data_0[2231:2224];
        layer6[25][15:8] = buffer_data_0[2239:2232];
        layer6[25][23:16] = buffer_data_0[2247:2240];
        layer6[25][31:24] = buffer_data_0[2255:2248];
        layer6[25][39:32] = buffer_data_0[2263:2256];
        layer6[25][47:40] = buffer_data_0[2271:2264];
        layer6[25][55:48] = buffer_data_0[2279:2272];
        layer0[26][7:0] = buffer_data_6[2239:2232];
        layer0[26][15:8] = buffer_data_6[2247:2240];
        layer0[26][23:16] = buffer_data_6[2255:2248];
        layer0[26][31:24] = buffer_data_6[2263:2256];
        layer0[26][39:32] = buffer_data_6[2271:2264];
        layer0[26][47:40] = buffer_data_6[2279:2272];
        layer0[26][55:48] = buffer_data_6[2287:2280];
        layer1[26][7:0] = buffer_data_5[2239:2232];
        layer1[26][15:8] = buffer_data_5[2247:2240];
        layer1[26][23:16] = buffer_data_5[2255:2248];
        layer1[26][31:24] = buffer_data_5[2263:2256];
        layer1[26][39:32] = buffer_data_5[2271:2264];
        layer1[26][47:40] = buffer_data_5[2279:2272];
        layer1[26][55:48] = buffer_data_5[2287:2280];
        layer2[26][7:0] = buffer_data_4[2239:2232];
        layer2[26][15:8] = buffer_data_4[2247:2240];
        layer2[26][23:16] = buffer_data_4[2255:2248];
        layer2[26][31:24] = buffer_data_4[2263:2256];
        layer2[26][39:32] = buffer_data_4[2271:2264];
        layer2[26][47:40] = buffer_data_4[2279:2272];
        layer2[26][55:48] = buffer_data_4[2287:2280];
        layer3[26][7:0] = buffer_data_3[2239:2232];
        layer3[26][15:8] = buffer_data_3[2247:2240];
        layer3[26][23:16] = buffer_data_3[2255:2248];
        layer3[26][31:24] = buffer_data_3[2263:2256];
        layer3[26][39:32] = buffer_data_3[2271:2264];
        layer3[26][47:40] = buffer_data_3[2279:2272];
        layer3[26][55:48] = buffer_data_3[2287:2280];
        layer4[26][7:0] = buffer_data_2[2239:2232];
        layer4[26][15:8] = buffer_data_2[2247:2240];
        layer4[26][23:16] = buffer_data_2[2255:2248];
        layer4[26][31:24] = buffer_data_2[2263:2256];
        layer4[26][39:32] = buffer_data_2[2271:2264];
        layer4[26][47:40] = buffer_data_2[2279:2272];
        layer4[26][55:48] = buffer_data_2[2287:2280];
        layer5[26][7:0] = buffer_data_1[2239:2232];
        layer5[26][15:8] = buffer_data_1[2247:2240];
        layer5[26][23:16] = buffer_data_1[2255:2248];
        layer5[26][31:24] = buffer_data_1[2263:2256];
        layer5[26][39:32] = buffer_data_1[2271:2264];
        layer5[26][47:40] = buffer_data_1[2279:2272];
        layer5[26][55:48] = buffer_data_1[2287:2280];
        layer6[26][7:0] = buffer_data_0[2239:2232];
        layer6[26][15:8] = buffer_data_0[2247:2240];
        layer6[26][23:16] = buffer_data_0[2255:2248];
        layer6[26][31:24] = buffer_data_0[2263:2256];
        layer6[26][39:32] = buffer_data_0[2271:2264];
        layer6[26][47:40] = buffer_data_0[2279:2272];
        layer6[26][55:48] = buffer_data_0[2287:2280];
        layer0[27][7:0] = buffer_data_6[2247:2240];
        layer0[27][15:8] = buffer_data_6[2255:2248];
        layer0[27][23:16] = buffer_data_6[2263:2256];
        layer0[27][31:24] = buffer_data_6[2271:2264];
        layer0[27][39:32] = buffer_data_6[2279:2272];
        layer0[27][47:40] = buffer_data_6[2287:2280];
        layer0[27][55:48] = buffer_data_6[2295:2288];
        layer1[27][7:0] = buffer_data_5[2247:2240];
        layer1[27][15:8] = buffer_data_5[2255:2248];
        layer1[27][23:16] = buffer_data_5[2263:2256];
        layer1[27][31:24] = buffer_data_5[2271:2264];
        layer1[27][39:32] = buffer_data_5[2279:2272];
        layer1[27][47:40] = buffer_data_5[2287:2280];
        layer1[27][55:48] = buffer_data_5[2295:2288];
        layer2[27][7:0] = buffer_data_4[2247:2240];
        layer2[27][15:8] = buffer_data_4[2255:2248];
        layer2[27][23:16] = buffer_data_4[2263:2256];
        layer2[27][31:24] = buffer_data_4[2271:2264];
        layer2[27][39:32] = buffer_data_4[2279:2272];
        layer2[27][47:40] = buffer_data_4[2287:2280];
        layer2[27][55:48] = buffer_data_4[2295:2288];
        layer3[27][7:0] = buffer_data_3[2247:2240];
        layer3[27][15:8] = buffer_data_3[2255:2248];
        layer3[27][23:16] = buffer_data_3[2263:2256];
        layer3[27][31:24] = buffer_data_3[2271:2264];
        layer3[27][39:32] = buffer_data_3[2279:2272];
        layer3[27][47:40] = buffer_data_3[2287:2280];
        layer3[27][55:48] = buffer_data_3[2295:2288];
        layer4[27][7:0] = buffer_data_2[2247:2240];
        layer4[27][15:8] = buffer_data_2[2255:2248];
        layer4[27][23:16] = buffer_data_2[2263:2256];
        layer4[27][31:24] = buffer_data_2[2271:2264];
        layer4[27][39:32] = buffer_data_2[2279:2272];
        layer4[27][47:40] = buffer_data_2[2287:2280];
        layer4[27][55:48] = buffer_data_2[2295:2288];
        layer5[27][7:0] = buffer_data_1[2247:2240];
        layer5[27][15:8] = buffer_data_1[2255:2248];
        layer5[27][23:16] = buffer_data_1[2263:2256];
        layer5[27][31:24] = buffer_data_1[2271:2264];
        layer5[27][39:32] = buffer_data_1[2279:2272];
        layer5[27][47:40] = buffer_data_1[2287:2280];
        layer5[27][55:48] = buffer_data_1[2295:2288];
        layer6[27][7:0] = buffer_data_0[2247:2240];
        layer6[27][15:8] = buffer_data_0[2255:2248];
        layer6[27][23:16] = buffer_data_0[2263:2256];
        layer6[27][31:24] = buffer_data_0[2271:2264];
        layer6[27][39:32] = buffer_data_0[2279:2272];
        layer6[27][47:40] = buffer_data_0[2287:2280];
        layer6[27][55:48] = buffer_data_0[2295:2288];
        layer0[28][7:0] = buffer_data_6[2255:2248];
        layer0[28][15:8] = buffer_data_6[2263:2256];
        layer0[28][23:16] = buffer_data_6[2271:2264];
        layer0[28][31:24] = buffer_data_6[2279:2272];
        layer0[28][39:32] = buffer_data_6[2287:2280];
        layer0[28][47:40] = buffer_data_6[2295:2288];
        layer0[28][55:48] = buffer_data_6[2303:2296];
        layer1[28][7:0] = buffer_data_5[2255:2248];
        layer1[28][15:8] = buffer_data_5[2263:2256];
        layer1[28][23:16] = buffer_data_5[2271:2264];
        layer1[28][31:24] = buffer_data_5[2279:2272];
        layer1[28][39:32] = buffer_data_5[2287:2280];
        layer1[28][47:40] = buffer_data_5[2295:2288];
        layer1[28][55:48] = buffer_data_5[2303:2296];
        layer2[28][7:0] = buffer_data_4[2255:2248];
        layer2[28][15:8] = buffer_data_4[2263:2256];
        layer2[28][23:16] = buffer_data_4[2271:2264];
        layer2[28][31:24] = buffer_data_4[2279:2272];
        layer2[28][39:32] = buffer_data_4[2287:2280];
        layer2[28][47:40] = buffer_data_4[2295:2288];
        layer2[28][55:48] = buffer_data_4[2303:2296];
        layer3[28][7:0] = buffer_data_3[2255:2248];
        layer3[28][15:8] = buffer_data_3[2263:2256];
        layer3[28][23:16] = buffer_data_3[2271:2264];
        layer3[28][31:24] = buffer_data_3[2279:2272];
        layer3[28][39:32] = buffer_data_3[2287:2280];
        layer3[28][47:40] = buffer_data_3[2295:2288];
        layer3[28][55:48] = buffer_data_3[2303:2296];
        layer4[28][7:0] = buffer_data_2[2255:2248];
        layer4[28][15:8] = buffer_data_2[2263:2256];
        layer4[28][23:16] = buffer_data_2[2271:2264];
        layer4[28][31:24] = buffer_data_2[2279:2272];
        layer4[28][39:32] = buffer_data_2[2287:2280];
        layer4[28][47:40] = buffer_data_2[2295:2288];
        layer4[28][55:48] = buffer_data_2[2303:2296];
        layer5[28][7:0] = buffer_data_1[2255:2248];
        layer5[28][15:8] = buffer_data_1[2263:2256];
        layer5[28][23:16] = buffer_data_1[2271:2264];
        layer5[28][31:24] = buffer_data_1[2279:2272];
        layer5[28][39:32] = buffer_data_1[2287:2280];
        layer5[28][47:40] = buffer_data_1[2295:2288];
        layer5[28][55:48] = buffer_data_1[2303:2296];
        layer6[28][7:0] = buffer_data_0[2255:2248];
        layer6[28][15:8] = buffer_data_0[2263:2256];
        layer6[28][23:16] = buffer_data_0[2271:2264];
        layer6[28][31:24] = buffer_data_0[2279:2272];
        layer6[28][39:32] = buffer_data_0[2287:2280];
        layer6[28][47:40] = buffer_data_0[2295:2288];
        layer6[28][55:48] = buffer_data_0[2303:2296];
        layer0[29][7:0] = buffer_data_6[2263:2256];
        layer0[29][15:8] = buffer_data_6[2271:2264];
        layer0[29][23:16] = buffer_data_6[2279:2272];
        layer0[29][31:24] = buffer_data_6[2287:2280];
        layer0[29][39:32] = buffer_data_6[2295:2288];
        layer0[29][47:40] = buffer_data_6[2303:2296];
        layer0[29][55:48] = buffer_data_6[2311:2304];
        layer1[29][7:0] = buffer_data_5[2263:2256];
        layer1[29][15:8] = buffer_data_5[2271:2264];
        layer1[29][23:16] = buffer_data_5[2279:2272];
        layer1[29][31:24] = buffer_data_5[2287:2280];
        layer1[29][39:32] = buffer_data_5[2295:2288];
        layer1[29][47:40] = buffer_data_5[2303:2296];
        layer1[29][55:48] = buffer_data_5[2311:2304];
        layer2[29][7:0] = buffer_data_4[2263:2256];
        layer2[29][15:8] = buffer_data_4[2271:2264];
        layer2[29][23:16] = buffer_data_4[2279:2272];
        layer2[29][31:24] = buffer_data_4[2287:2280];
        layer2[29][39:32] = buffer_data_4[2295:2288];
        layer2[29][47:40] = buffer_data_4[2303:2296];
        layer2[29][55:48] = buffer_data_4[2311:2304];
        layer3[29][7:0] = buffer_data_3[2263:2256];
        layer3[29][15:8] = buffer_data_3[2271:2264];
        layer3[29][23:16] = buffer_data_3[2279:2272];
        layer3[29][31:24] = buffer_data_3[2287:2280];
        layer3[29][39:32] = buffer_data_3[2295:2288];
        layer3[29][47:40] = buffer_data_3[2303:2296];
        layer3[29][55:48] = buffer_data_3[2311:2304];
        layer4[29][7:0] = buffer_data_2[2263:2256];
        layer4[29][15:8] = buffer_data_2[2271:2264];
        layer4[29][23:16] = buffer_data_2[2279:2272];
        layer4[29][31:24] = buffer_data_2[2287:2280];
        layer4[29][39:32] = buffer_data_2[2295:2288];
        layer4[29][47:40] = buffer_data_2[2303:2296];
        layer4[29][55:48] = buffer_data_2[2311:2304];
        layer5[29][7:0] = buffer_data_1[2263:2256];
        layer5[29][15:8] = buffer_data_1[2271:2264];
        layer5[29][23:16] = buffer_data_1[2279:2272];
        layer5[29][31:24] = buffer_data_1[2287:2280];
        layer5[29][39:32] = buffer_data_1[2295:2288];
        layer5[29][47:40] = buffer_data_1[2303:2296];
        layer5[29][55:48] = buffer_data_1[2311:2304];
        layer6[29][7:0] = buffer_data_0[2263:2256];
        layer6[29][15:8] = buffer_data_0[2271:2264];
        layer6[29][23:16] = buffer_data_0[2279:2272];
        layer6[29][31:24] = buffer_data_0[2287:2280];
        layer6[29][39:32] = buffer_data_0[2295:2288];
        layer6[29][47:40] = buffer_data_0[2303:2296];
        layer6[29][55:48] = buffer_data_0[2311:2304];
        layer0[30][7:0] = buffer_data_6[2271:2264];
        layer0[30][15:8] = buffer_data_6[2279:2272];
        layer0[30][23:16] = buffer_data_6[2287:2280];
        layer0[30][31:24] = buffer_data_6[2295:2288];
        layer0[30][39:32] = buffer_data_6[2303:2296];
        layer0[30][47:40] = buffer_data_6[2311:2304];
        layer0[30][55:48] = buffer_data_6[2319:2312];
        layer1[30][7:0] = buffer_data_5[2271:2264];
        layer1[30][15:8] = buffer_data_5[2279:2272];
        layer1[30][23:16] = buffer_data_5[2287:2280];
        layer1[30][31:24] = buffer_data_5[2295:2288];
        layer1[30][39:32] = buffer_data_5[2303:2296];
        layer1[30][47:40] = buffer_data_5[2311:2304];
        layer1[30][55:48] = buffer_data_5[2319:2312];
        layer2[30][7:0] = buffer_data_4[2271:2264];
        layer2[30][15:8] = buffer_data_4[2279:2272];
        layer2[30][23:16] = buffer_data_4[2287:2280];
        layer2[30][31:24] = buffer_data_4[2295:2288];
        layer2[30][39:32] = buffer_data_4[2303:2296];
        layer2[30][47:40] = buffer_data_4[2311:2304];
        layer2[30][55:48] = buffer_data_4[2319:2312];
        layer3[30][7:0] = buffer_data_3[2271:2264];
        layer3[30][15:8] = buffer_data_3[2279:2272];
        layer3[30][23:16] = buffer_data_3[2287:2280];
        layer3[30][31:24] = buffer_data_3[2295:2288];
        layer3[30][39:32] = buffer_data_3[2303:2296];
        layer3[30][47:40] = buffer_data_3[2311:2304];
        layer3[30][55:48] = buffer_data_3[2319:2312];
        layer4[30][7:0] = buffer_data_2[2271:2264];
        layer4[30][15:8] = buffer_data_2[2279:2272];
        layer4[30][23:16] = buffer_data_2[2287:2280];
        layer4[30][31:24] = buffer_data_2[2295:2288];
        layer4[30][39:32] = buffer_data_2[2303:2296];
        layer4[30][47:40] = buffer_data_2[2311:2304];
        layer4[30][55:48] = buffer_data_2[2319:2312];
        layer5[30][7:0] = buffer_data_1[2271:2264];
        layer5[30][15:8] = buffer_data_1[2279:2272];
        layer5[30][23:16] = buffer_data_1[2287:2280];
        layer5[30][31:24] = buffer_data_1[2295:2288];
        layer5[30][39:32] = buffer_data_1[2303:2296];
        layer5[30][47:40] = buffer_data_1[2311:2304];
        layer5[30][55:48] = buffer_data_1[2319:2312];
        layer6[30][7:0] = buffer_data_0[2271:2264];
        layer6[30][15:8] = buffer_data_0[2279:2272];
        layer6[30][23:16] = buffer_data_0[2287:2280];
        layer6[30][31:24] = buffer_data_0[2295:2288];
        layer6[30][39:32] = buffer_data_0[2303:2296];
        layer6[30][47:40] = buffer_data_0[2311:2304];
        layer6[30][55:48] = buffer_data_0[2319:2312];
        layer0[31][7:0] = buffer_data_6[2279:2272];
        layer0[31][15:8] = buffer_data_6[2287:2280];
        layer0[31][23:16] = buffer_data_6[2295:2288];
        layer0[31][31:24] = buffer_data_6[2303:2296];
        layer0[31][39:32] = buffer_data_6[2311:2304];
        layer0[31][47:40] = buffer_data_6[2319:2312];
        layer0[31][55:48] = buffer_data_6[2327:2320];
        layer1[31][7:0] = buffer_data_5[2279:2272];
        layer1[31][15:8] = buffer_data_5[2287:2280];
        layer1[31][23:16] = buffer_data_5[2295:2288];
        layer1[31][31:24] = buffer_data_5[2303:2296];
        layer1[31][39:32] = buffer_data_5[2311:2304];
        layer1[31][47:40] = buffer_data_5[2319:2312];
        layer1[31][55:48] = buffer_data_5[2327:2320];
        layer2[31][7:0] = buffer_data_4[2279:2272];
        layer2[31][15:8] = buffer_data_4[2287:2280];
        layer2[31][23:16] = buffer_data_4[2295:2288];
        layer2[31][31:24] = buffer_data_4[2303:2296];
        layer2[31][39:32] = buffer_data_4[2311:2304];
        layer2[31][47:40] = buffer_data_4[2319:2312];
        layer2[31][55:48] = buffer_data_4[2327:2320];
        layer3[31][7:0] = buffer_data_3[2279:2272];
        layer3[31][15:8] = buffer_data_3[2287:2280];
        layer3[31][23:16] = buffer_data_3[2295:2288];
        layer3[31][31:24] = buffer_data_3[2303:2296];
        layer3[31][39:32] = buffer_data_3[2311:2304];
        layer3[31][47:40] = buffer_data_3[2319:2312];
        layer3[31][55:48] = buffer_data_3[2327:2320];
        layer4[31][7:0] = buffer_data_2[2279:2272];
        layer4[31][15:8] = buffer_data_2[2287:2280];
        layer4[31][23:16] = buffer_data_2[2295:2288];
        layer4[31][31:24] = buffer_data_2[2303:2296];
        layer4[31][39:32] = buffer_data_2[2311:2304];
        layer4[31][47:40] = buffer_data_2[2319:2312];
        layer4[31][55:48] = buffer_data_2[2327:2320];
        layer5[31][7:0] = buffer_data_1[2279:2272];
        layer5[31][15:8] = buffer_data_1[2287:2280];
        layer5[31][23:16] = buffer_data_1[2295:2288];
        layer5[31][31:24] = buffer_data_1[2303:2296];
        layer5[31][39:32] = buffer_data_1[2311:2304];
        layer5[31][47:40] = buffer_data_1[2319:2312];
        layer5[31][55:48] = buffer_data_1[2327:2320];
        layer6[31][7:0] = buffer_data_0[2279:2272];
        layer6[31][15:8] = buffer_data_0[2287:2280];
        layer6[31][23:16] = buffer_data_0[2295:2288];
        layer6[31][31:24] = buffer_data_0[2303:2296];
        layer6[31][39:32] = buffer_data_0[2311:2304];
        layer6[31][47:40] = buffer_data_0[2319:2312];
        layer6[31][55:48] = buffer_data_0[2327:2320];
        layer0[32][7:0] = buffer_data_6[2287:2280];
        layer0[32][15:8] = buffer_data_6[2295:2288];
        layer0[32][23:16] = buffer_data_6[2303:2296];
        layer0[32][31:24] = buffer_data_6[2311:2304];
        layer0[32][39:32] = buffer_data_6[2319:2312];
        layer0[32][47:40] = buffer_data_6[2327:2320];
        layer0[32][55:48] = buffer_data_6[2335:2328];
        layer1[32][7:0] = buffer_data_5[2287:2280];
        layer1[32][15:8] = buffer_data_5[2295:2288];
        layer1[32][23:16] = buffer_data_5[2303:2296];
        layer1[32][31:24] = buffer_data_5[2311:2304];
        layer1[32][39:32] = buffer_data_5[2319:2312];
        layer1[32][47:40] = buffer_data_5[2327:2320];
        layer1[32][55:48] = buffer_data_5[2335:2328];
        layer2[32][7:0] = buffer_data_4[2287:2280];
        layer2[32][15:8] = buffer_data_4[2295:2288];
        layer2[32][23:16] = buffer_data_4[2303:2296];
        layer2[32][31:24] = buffer_data_4[2311:2304];
        layer2[32][39:32] = buffer_data_4[2319:2312];
        layer2[32][47:40] = buffer_data_4[2327:2320];
        layer2[32][55:48] = buffer_data_4[2335:2328];
        layer3[32][7:0] = buffer_data_3[2287:2280];
        layer3[32][15:8] = buffer_data_3[2295:2288];
        layer3[32][23:16] = buffer_data_3[2303:2296];
        layer3[32][31:24] = buffer_data_3[2311:2304];
        layer3[32][39:32] = buffer_data_3[2319:2312];
        layer3[32][47:40] = buffer_data_3[2327:2320];
        layer3[32][55:48] = buffer_data_3[2335:2328];
        layer4[32][7:0] = buffer_data_2[2287:2280];
        layer4[32][15:8] = buffer_data_2[2295:2288];
        layer4[32][23:16] = buffer_data_2[2303:2296];
        layer4[32][31:24] = buffer_data_2[2311:2304];
        layer4[32][39:32] = buffer_data_2[2319:2312];
        layer4[32][47:40] = buffer_data_2[2327:2320];
        layer4[32][55:48] = buffer_data_2[2335:2328];
        layer5[32][7:0] = buffer_data_1[2287:2280];
        layer5[32][15:8] = buffer_data_1[2295:2288];
        layer5[32][23:16] = buffer_data_1[2303:2296];
        layer5[32][31:24] = buffer_data_1[2311:2304];
        layer5[32][39:32] = buffer_data_1[2319:2312];
        layer5[32][47:40] = buffer_data_1[2327:2320];
        layer5[32][55:48] = buffer_data_1[2335:2328];
        layer6[32][7:0] = buffer_data_0[2287:2280];
        layer6[32][15:8] = buffer_data_0[2295:2288];
        layer6[32][23:16] = buffer_data_0[2303:2296];
        layer6[32][31:24] = buffer_data_0[2311:2304];
        layer6[32][39:32] = buffer_data_0[2319:2312];
        layer6[32][47:40] = buffer_data_0[2327:2320];
        layer6[32][55:48] = buffer_data_0[2335:2328];
        layer0[33][7:0] = buffer_data_6[2295:2288];
        layer0[33][15:8] = buffer_data_6[2303:2296];
        layer0[33][23:16] = buffer_data_6[2311:2304];
        layer0[33][31:24] = buffer_data_6[2319:2312];
        layer0[33][39:32] = buffer_data_6[2327:2320];
        layer0[33][47:40] = buffer_data_6[2335:2328];
        layer0[33][55:48] = buffer_data_6[2343:2336];
        layer1[33][7:0] = buffer_data_5[2295:2288];
        layer1[33][15:8] = buffer_data_5[2303:2296];
        layer1[33][23:16] = buffer_data_5[2311:2304];
        layer1[33][31:24] = buffer_data_5[2319:2312];
        layer1[33][39:32] = buffer_data_5[2327:2320];
        layer1[33][47:40] = buffer_data_5[2335:2328];
        layer1[33][55:48] = buffer_data_5[2343:2336];
        layer2[33][7:0] = buffer_data_4[2295:2288];
        layer2[33][15:8] = buffer_data_4[2303:2296];
        layer2[33][23:16] = buffer_data_4[2311:2304];
        layer2[33][31:24] = buffer_data_4[2319:2312];
        layer2[33][39:32] = buffer_data_4[2327:2320];
        layer2[33][47:40] = buffer_data_4[2335:2328];
        layer2[33][55:48] = buffer_data_4[2343:2336];
        layer3[33][7:0] = buffer_data_3[2295:2288];
        layer3[33][15:8] = buffer_data_3[2303:2296];
        layer3[33][23:16] = buffer_data_3[2311:2304];
        layer3[33][31:24] = buffer_data_3[2319:2312];
        layer3[33][39:32] = buffer_data_3[2327:2320];
        layer3[33][47:40] = buffer_data_3[2335:2328];
        layer3[33][55:48] = buffer_data_3[2343:2336];
        layer4[33][7:0] = buffer_data_2[2295:2288];
        layer4[33][15:8] = buffer_data_2[2303:2296];
        layer4[33][23:16] = buffer_data_2[2311:2304];
        layer4[33][31:24] = buffer_data_2[2319:2312];
        layer4[33][39:32] = buffer_data_2[2327:2320];
        layer4[33][47:40] = buffer_data_2[2335:2328];
        layer4[33][55:48] = buffer_data_2[2343:2336];
        layer5[33][7:0] = buffer_data_1[2295:2288];
        layer5[33][15:8] = buffer_data_1[2303:2296];
        layer5[33][23:16] = buffer_data_1[2311:2304];
        layer5[33][31:24] = buffer_data_1[2319:2312];
        layer5[33][39:32] = buffer_data_1[2327:2320];
        layer5[33][47:40] = buffer_data_1[2335:2328];
        layer5[33][55:48] = buffer_data_1[2343:2336];
        layer6[33][7:0] = buffer_data_0[2295:2288];
        layer6[33][15:8] = buffer_data_0[2303:2296];
        layer6[33][23:16] = buffer_data_0[2311:2304];
        layer6[33][31:24] = buffer_data_0[2319:2312];
        layer6[33][39:32] = buffer_data_0[2327:2320];
        layer6[33][47:40] = buffer_data_0[2335:2328];
        layer6[33][55:48] = buffer_data_0[2343:2336];
        layer0[34][7:0] = buffer_data_6[2303:2296];
        layer0[34][15:8] = buffer_data_6[2311:2304];
        layer0[34][23:16] = buffer_data_6[2319:2312];
        layer0[34][31:24] = buffer_data_6[2327:2320];
        layer0[34][39:32] = buffer_data_6[2335:2328];
        layer0[34][47:40] = buffer_data_6[2343:2336];
        layer0[34][55:48] = buffer_data_6[2351:2344];
        layer1[34][7:0] = buffer_data_5[2303:2296];
        layer1[34][15:8] = buffer_data_5[2311:2304];
        layer1[34][23:16] = buffer_data_5[2319:2312];
        layer1[34][31:24] = buffer_data_5[2327:2320];
        layer1[34][39:32] = buffer_data_5[2335:2328];
        layer1[34][47:40] = buffer_data_5[2343:2336];
        layer1[34][55:48] = buffer_data_5[2351:2344];
        layer2[34][7:0] = buffer_data_4[2303:2296];
        layer2[34][15:8] = buffer_data_4[2311:2304];
        layer2[34][23:16] = buffer_data_4[2319:2312];
        layer2[34][31:24] = buffer_data_4[2327:2320];
        layer2[34][39:32] = buffer_data_4[2335:2328];
        layer2[34][47:40] = buffer_data_4[2343:2336];
        layer2[34][55:48] = buffer_data_4[2351:2344];
        layer3[34][7:0] = buffer_data_3[2303:2296];
        layer3[34][15:8] = buffer_data_3[2311:2304];
        layer3[34][23:16] = buffer_data_3[2319:2312];
        layer3[34][31:24] = buffer_data_3[2327:2320];
        layer3[34][39:32] = buffer_data_3[2335:2328];
        layer3[34][47:40] = buffer_data_3[2343:2336];
        layer3[34][55:48] = buffer_data_3[2351:2344];
        layer4[34][7:0] = buffer_data_2[2303:2296];
        layer4[34][15:8] = buffer_data_2[2311:2304];
        layer4[34][23:16] = buffer_data_2[2319:2312];
        layer4[34][31:24] = buffer_data_2[2327:2320];
        layer4[34][39:32] = buffer_data_2[2335:2328];
        layer4[34][47:40] = buffer_data_2[2343:2336];
        layer4[34][55:48] = buffer_data_2[2351:2344];
        layer5[34][7:0] = buffer_data_1[2303:2296];
        layer5[34][15:8] = buffer_data_1[2311:2304];
        layer5[34][23:16] = buffer_data_1[2319:2312];
        layer5[34][31:24] = buffer_data_1[2327:2320];
        layer5[34][39:32] = buffer_data_1[2335:2328];
        layer5[34][47:40] = buffer_data_1[2343:2336];
        layer5[34][55:48] = buffer_data_1[2351:2344];
        layer6[34][7:0] = buffer_data_0[2303:2296];
        layer6[34][15:8] = buffer_data_0[2311:2304];
        layer6[34][23:16] = buffer_data_0[2319:2312];
        layer6[34][31:24] = buffer_data_0[2327:2320];
        layer6[34][39:32] = buffer_data_0[2335:2328];
        layer6[34][47:40] = buffer_data_0[2343:2336];
        layer6[34][55:48] = buffer_data_0[2351:2344];
        layer0[35][7:0] = buffer_data_6[2311:2304];
        layer0[35][15:8] = buffer_data_6[2319:2312];
        layer0[35][23:16] = buffer_data_6[2327:2320];
        layer0[35][31:24] = buffer_data_6[2335:2328];
        layer0[35][39:32] = buffer_data_6[2343:2336];
        layer0[35][47:40] = buffer_data_6[2351:2344];
        layer0[35][55:48] = buffer_data_6[2359:2352];
        layer1[35][7:0] = buffer_data_5[2311:2304];
        layer1[35][15:8] = buffer_data_5[2319:2312];
        layer1[35][23:16] = buffer_data_5[2327:2320];
        layer1[35][31:24] = buffer_data_5[2335:2328];
        layer1[35][39:32] = buffer_data_5[2343:2336];
        layer1[35][47:40] = buffer_data_5[2351:2344];
        layer1[35][55:48] = buffer_data_5[2359:2352];
        layer2[35][7:0] = buffer_data_4[2311:2304];
        layer2[35][15:8] = buffer_data_4[2319:2312];
        layer2[35][23:16] = buffer_data_4[2327:2320];
        layer2[35][31:24] = buffer_data_4[2335:2328];
        layer2[35][39:32] = buffer_data_4[2343:2336];
        layer2[35][47:40] = buffer_data_4[2351:2344];
        layer2[35][55:48] = buffer_data_4[2359:2352];
        layer3[35][7:0] = buffer_data_3[2311:2304];
        layer3[35][15:8] = buffer_data_3[2319:2312];
        layer3[35][23:16] = buffer_data_3[2327:2320];
        layer3[35][31:24] = buffer_data_3[2335:2328];
        layer3[35][39:32] = buffer_data_3[2343:2336];
        layer3[35][47:40] = buffer_data_3[2351:2344];
        layer3[35][55:48] = buffer_data_3[2359:2352];
        layer4[35][7:0] = buffer_data_2[2311:2304];
        layer4[35][15:8] = buffer_data_2[2319:2312];
        layer4[35][23:16] = buffer_data_2[2327:2320];
        layer4[35][31:24] = buffer_data_2[2335:2328];
        layer4[35][39:32] = buffer_data_2[2343:2336];
        layer4[35][47:40] = buffer_data_2[2351:2344];
        layer4[35][55:48] = buffer_data_2[2359:2352];
        layer5[35][7:0] = buffer_data_1[2311:2304];
        layer5[35][15:8] = buffer_data_1[2319:2312];
        layer5[35][23:16] = buffer_data_1[2327:2320];
        layer5[35][31:24] = buffer_data_1[2335:2328];
        layer5[35][39:32] = buffer_data_1[2343:2336];
        layer5[35][47:40] = buffer_data_1[2351:2344];
        layer5[35][55:48] = buffer_data_1[2359:2352];
        layer6[35][7:0] = buffer_data_0[2311:2304];
        layer6[35][15:8] = buffer_data_0[2319:2312];
        layer6[35][23:16] = buffer_data_0[2327:2320];
        layer6[35][31:24] = buffer_data_0[2335:2328];
        layer6[35][39:32] = buffer_data_0[2343:2336];
        layer6[35][47:40] = buffer_data_0[2351:2344];
        layer6[35][55:48] = buffer_data_0[2359:2352];
        layer0[36][7:0] = buffer_data_6[2319:2312];
        layer0[36][15:8] = buffer_data_6[2327:2320];
        layer0[36][23:16] = buffer_data_6[2335:2328];
        layer0[36][31:24] = buffer_data_6[2343:2336];
        layer0[36][39:32] = buffer_data_6[2351:2344];
        layer0[36][47:40] = buffer_data_6[2359:2352];
        layer0[36][55:48] = buffer_data_6[2367:2360];
        layer1[36][7:0] = buffer_data_5[2319:2312];
        layer1[36][15:8] = buffer_data_5[2327:2320];
        layer1[36][23:16] = buffer_data_5[2335:2328];
        layer1[36][31:24] = buffer_data_5[2343:2336];
        layer1[36][39:32] = buffer_data_5[2351:2344];
        layer1[36][47:40] = buffer_data_5[2359:2352];
        layer1[36][55:48] = buffer_data_5[2367:2360];
        layer2[36][7:0] = buffer_data_4[2319:2312];
        layer2[36][15:8] = buffer_data_4[2327:2320];
        layer2[36][23:16] = buffer_data_4[2335:2328];
        layer2[36][31:24] = buffer_data_4[2343:2336];
        layer2[36][39:32] = buffer_data_4[2351:2344];
        layer2[36][47:40] = buffer_data_4[2359:2352];
        layer2[36][55:48] = buffer_data_4[2367:2360];
        layer3[36][7:0] = buffer_data_3[2319:2312];
        layer3[36][15:8] = buffer_data_3[2327:2320];
        layer3[36][23:16] = buffer_data_3[2335:2328];
        layer3[36][31:24] = buffer_data_3[2343:2336];
        layer3[36][39:32] = buffer_data_3[2351:2344];
        layer3[36][47:40] = buffer_data_3[2359:2352];
        layer3[36][55:48] = buffer_data_3[2367:2360];
        layer4[36][7:0] = buffer_data_2[2319:2312];
        layer4[36][15:8] = buffer_data_2[2327:2320];
        layer4[36][23:16] = buffer_data_2[2335:2328];
        layer4[36][31:24] = buffer_data_2[2343:2336];
        layer4[36][39:32] = buffer_data_2[2351:2344];
        layer4[36][47:40] = buffer_data_2[2359:2352];
        layer4[36][55:48] = buffer_data_2[2367:2360];
        layer5[36][7:0] = buffer_data_1[2319:2312];
        layer5[36][15:8] = buffer_data_1[2327:2320];
        layer5[36][23:16] = buffer_data_1[2335:2328];
        layer5[36][31:24] = buffer_data_1[2343:2336];
        layer5[36][39:32] = buffer_data_1[2351:2344];
        layer5[36][47:40] = buffer_data_1[2359:2352];
        layer5[36][55:48] = buffer_data_1[2367:2360];
        layer6[36][7:0] = buffer_data_0[2319:2312];
        layer6[36][15:8] = buffer_data_0[2327:2320];
        layer6[36][23:16] = buffer_data_0[2335:2328];
        layer6[36][31:24] = buffer_data_0[2343:2336];
        layer6[36][39:32] = buffer_data_0[2351:2344];
        layer6[36][47:40] = buffer_data_0[2359:2352];
        layer6[36][55:48] = buffer_data_0[2367:2360];
        layer0[37][7:0] = buffer_data_6[2327:2320];
        layer0[37][15:8] = buffer_data_6[2335:2328];
        layer0[37][23:16] = buffer_data_6[2343:2336];
        layer0[37][31:24] = buffer_data_6[2351:2344];
        layer0[37][39:32] = buffer_data_6[2359:2352];
        layer0[37][47:40] = buffer_data_6[2367:2360];
        layer0[37][55:48] = buffer_data_6[2375:2368];
        layer1[37][7:0] = buffer_data_5[2327:2320];
        layer1[37][15:8] = buffer_data_5[2335:2328];
        layer1[37][23:16] = buffer_data_5[2343:2336];
        layer1[37][31:24] = buffer_data_5[2351:2344];
        layer1[37][39:32] = buffer_data_5[2359:2352];
        layer1[37][47:40] = buffer_data_5[2367:2360];
        layer1[37][55:48] = buffer_data_5[2375:2368];
        layer2[37][7:0] = buffer_data_4[2327:2320];
        layer2[37][15:8] = buffer_data_4[2335:2328];
        layer2[37][23:16] = buffer_data_4[2343:2336];
        layer2[37][31:24] = buffer_data_4[2351:2344];
        layer2[37][39:32] = buffer_data_4[2359:2352];
        layer2[37][47:40] = buffer_data_4[2367:2360];
        layer2[37][55:48] = buffer_data_4[2375:2368];
        layer3[37][7:0] = buffer_data_3[2327:2320];
        layer3[37][15:8] = buffer_data_3[2335:2328];
        layer3[37][23:16] = buffer_data_3[2343:2336];
        layer3[37][31:24] = buffer_data_3[2351:2344];
        layer3[37][39:32] = buffer_data_3[2359:2352];
        layer3[37][47:40] = buffer_data_3[2367:2360];
        layer3[37][55:48] = buffer_data_3[2375:2368];
        layer4[37][7:0] = buffer_data_2[2327:2320];
        layer4[37][15:8] = buffer_data_2[2335:2328];
        layer4[37][23:16] = buffer_data_2[2343:2336];
        layer4[37][31:24] = buffer_data_2[2351:2344];
        layer4[37][39:32] = buffer_data_2[2359:2352];
        layer4[37][47:40] = buffer_data_2[2367:2360];
        layer4[37][55:48] = buffer_data_2[2375:2368];
        layer5[37][7:0] = buffer_data_1[2327:2320];
        layer5[37][15:8] = buffer_data_1[2335:2328];
        layer5[37][23:16] = buffer_data_1[2343:2336];
        layer5[37][31:24] = buffer_data_1[2351:2344];
        layer5[37][39:32] = buffer_data_1[2359:2352];
        layer5[37][47:40] = buffer_data_1[2367:2360];
        layer5[37][55:48] = buffer_data_1[2375:2368];
        layer6[37][7:0] = buffer_data_0[2327:2320];
        layer6[37][15:8] = buffer_data_0[2335:2328];
        layer6[37][23:16] = buffer_data_0[2343:2336];
        layer6[37][31:24] = buffer_data_0[2351:2344];
        layer6[37][39:32] = buffer_data_0[2359:2352];
        layer6[37][47:40] = buffer_data_0[2367:2360];
        layer6[37][55:48] = buffer_data_0[2375:2368];
        layer0[38][7:0] = buffer_data_6[2335:2328];
        layer0[38][15:8] = buffer_data_6[2343:2336];
        layer0[38][23:16] = buffer_data_6[2351:2344];
        layer0[38][31:24] = buffer_data_6[2359:2352];
        layer0[38][39:32] = buffer_data_6[2367:2360];
        layer0[38][47:40] = buffer_data_6[2375:2368];
        layer0[38][55:48] = buffer_data_6[2383:2376];
        layer1[38][7:0] = buffer_data_5[2335:2328];
        layer1[38][15:8] = buffer_data_5[2343:2336];
        layer1[38][23:16] = buffer_data_5[2351:2344];
        layer1[38][31:24] = buffer_data_5[2359:2352];
        layer1[38][39:32] = buffer_data_5[2367:2360];
        layer1[38][47:40] = buffer_data_5[2375:2368];
        layer1[38][55:48] = buffer_data_5[2383:2376];
        layer2[38][7:0] = buffer_data_4[2335:2328];
        layer2[38][15:8] = buffer_data_4[2343:2336];
        layer2[38][23:16] = buffer_data_4[2351:2344];
        layer2[38][31:24] = buffer_data_4[2359:2352];
        layer2[38][39:32] = buffer_data_4[2367:2360];
        layer2[38][47:40] = buffer_data_4[2375:2368];
        layer2[38][55:48] = buffer_data_4[2383:2376];
        layer3[38][7:0] = buffer_data_3[2335:2328];
        layer3[38][15:8] = buffer_data_3[2343:2336];
        layer3[38][23:16] = buffer_data_3[2351:2344];
        layer3[38][31:24] = buffer_data_3[2359:2352];
        layer3[38][39:32] = buffer_data_3[2367:2360];
        layer3[38][47:40] = buffer_data_3[2375:2368];
        layer3[38][55:48] = buffer_data_3[2383:2376];
        layer4[38][7:0] = buffer_data_2[2335:2328];
        layer4[38][15:8] = buffer_data_2[2343:2336];
        layer4[38][23:16] = buffer_data_2[2351:2344];
        layer4[38][31:24] = buffer_data_2[2359:2352];
        layer4[38][39:32] = buffer_data_2[2367:2360];
        layer4[38][47:40] = buffer_data_2[2375:2368];
        layer4[38][55:48] = buffer_data_2[2383:2376];
        layer5[38][7:0] = buffer_data_1[2335:2328];
        layer5[38][15:8] = buffer_data_1[2343:2336];
        layer5[38][23:16] = buffer_data_1[2351:2344];
        layer5[38][31:24] = buffer_data_1[2359:2352];
        layer5[38][39:32] = buffer_data_1[2367:2360];
        layer5[38][47:40] = buffer_data_1[2375:2368];
        layer5[38][55:48] = buffer_data_1[2383:2376];
        layer6[38][7:0] = buffer_data_0[2335:2328];
        layer6[38][15:8] = buffer_data_0[2343:2336];
        layer6[38][23:16] = buffer_data_0[2351:2344];
        layer6[38][31:24] = buffer_data_0[2359:2352];
        layer6[38][39:32] = buffer_data_0[2367:2360];
        layer6[38][47:40] = buffer_data_0[2375:2368];
        layer6[38][55:48] = buffer_data_0[2383:2376];
        layer0[39][7:0] = buffer_data_6[2343:2336];
        layer0[39][15:8] = buffer_data_6[2351:2344];
        layer0[39][23:16] = buffer_data_6[2359:2352];
        layer0[39][31:24] = buffer_data_6[2367:2360];
        layer0[39][39:32] = buffer_data_6[2375:2368];
        layer0[39][47:40] = buffer_data_6[2383:2376];
        layer0[39][55:48] = buffer_data_6[2391:2384];
        layer1[39][7:0] = buffer_data_5[2343:2336];
        layer1[39][15:8] = buffer_data_5[2351:2344];
        layer1[39][23:16] = buffer_data_5[2359:2352];
        layer1[39][31:24] = buffer_data_5[2367:2360];
        layer1[39][39:32] = buffer_data_5[2375:2368];
        layer1[39][47:40] = buffer_data_5[2383:2376];
        layer1[39][55:48] = buffer_data_5[2391:2384];
        layer2[39][7:0] = buffer_data_4[2343:2336];
        layer2[39][15:8] = buffer_data_4[2351:2344];
        layer2[39][23:16] = buffer_data_4[2359:2352];
        layer2[39][31:24] = buffer_data_4[2367:2360];
        layer2[39][39:32] = buffer_data_4[2375:2368];
        layer2[39][47:40] = buffer_data_4[2383:2376];
        layer2[39][55:48] = buffer_data_4[2391:2384];
        layer3[39][7:0] = buffer_data_3[2343:2336];
        layer3[39][15:8] = buffer_data_3[2351:2344];
        layer3[39][23:16] = buffer_data_3[2359:2352];
        layer3[39][31:24] = buffer_data_3[2367:2360];
        layer3[39][39:32] = buffer_data_3[2375:2368];
        layer3[39][47:40] = buffer_data_3[2383:2376];
        layer3[39][55:48] = buffer_data_3[2391:2384];
        layer4[39][7:0] = buffer_data_2[2343:2336];
        layer4[39][15:8] = buffer_data_2[2351:2344];
        layer4[39][23:16] = buffer_data_2[2359:2352];
        layer4[39][31:24] = buffer_data_2[2367:2360];
        layer4[39][39:32] = buffer_data_2[2375:2368];
        layer4[39][47:40] = buffer_data_2[2383:2376];
        layer4[39][55:48] = buffer_data_2[2391:2384];
        layer5[39][7:0] = buffer_data_1[2343:2336];
        layer5[39][15:8] = buffer_data_1[2351:2344];
        layer5[39][23:16] = buffer_data_1[2359:2352];
        layer5[39][31:24] = buffer_data_1[2367:2360];
        layer5[39][39:32] = buffer_data_1[2375:2368];
        layer5[39][47:40] = buffer_data_1[2383:2376];
        layer5[39][55:48] = buffer_data_1[2391:2384];
        layer6[39][7:0] = buffer_data_0[2343:2336];
        layer6[39][15:8] = buffer_data_0[2351:2344];
        layer6[39][23:16] = buffer_data_0[2359:2352];
        layer6[39][31:24] = buffer_data_0[2367:2360];
        layer6[39][39:32] = buffer_data_0[2375:2368];
        layer6[39][47:40] = buffer_data_0[2383:2376];
        layer6[39][55:48] = buffer_data_0[2391:2384];
        layer0[40][7:0] = buffer_data_6[2351:2344];
        layer0[40][15:8] = buffer_data_6[2359:2352];
        layer0[40][23:16] = buffer_data_6[2367:2360];
        layer0[40][31:24] = buffer_data_6[2375:2368];
        layer0[40][39:32] = buffer_data_6[2383:2376];
        layer0[40][47:40] = buffer_data_6[2391:2384];
        layer0[40][55:48] = buffer_data_6[2399:2392];
        layer1[40][7:0] = buffer_data_5[2351:2344];
        layer1[40][15:8] = buffer_data_5[2359:2352];
        layer1[40][23:16] = buffer_data_5[2367:2360];
        layer1[40][31:24] = buffer_data_5[2375:2368];
        layer1[40][39:32] = buffer_data_5[2383:2376];
        layer1[40][47:40] = buffer_data_5[2391:2384];
        layer1[40][55:48] = buffer_data_5[2399:2392];
        layer2[40][7:0] = buffer_data_4[2351:2344];
        layer2[40][15:8] = buffer_data_4[2359:2352];
        layer2[40][23:16] = buffer_data_4[2367:2360];
        layer2[40][31:24] = buffer_data_4[2375:2368];
        layer2[40][39:32] = buffer_data_4[2383:2376];
        layer2[40][47:40] = buffer_data_4[2391:2384];
        layer2[40][55:48] = buffer_data_4[2399:2392];
        layer3[40][7:0] = buffer_data_3[2351:2344];
        layer3[40][15:8] = buffer_data_3[2359:2352];
        layer3[40][23:16] = buffer_data_3[2367:2360];
        layer3[40][31:24] = buffer_data_3[2375:2368];
        layer3[40][39:32] = buffer_data_3[2383:2376];
        layer3[40][47:40] = buffer_data_3[2391:2384];
        layer3[40][55:48] = buffer_data_3[2399:2392];
        layer4[40][7:0] = buffer_data_2[2351:2344];
        layer4[40][15:8] = buffer_data_2[2359:2352];
        layer4[40][23:16] = buffer_data_2[2367:2360];
        layer4[40][31:24] = buffer_data_2[2375:2368];
        layer4[40][39:32] = buffer_data_2[2383:2376];
        layer4[40][47:40] = buffer_data_2[2391:2384];
        layer4[40][55:48] = buffer_data_2[2399:2392];
        layer5[40][7:0] = buffer_data_1[2351:2344];
        layer5[40][15:8] = buffer_data_1[2359:2352];
        layer5[40][23:16] = buffer_data_1[2367:2360];
        layer5[40][31:24] = buffer_data_1[2375:2368];
        layer5[40][39:32] = buffer_data_1[2383:2376];
        layer5[40][47:40] = buffer_data_1[2391:2384];
        layer5[40][55:48] = buffer_data_1[2399:2392];
        layer6[40][7:0] = buffer_data_0[2351:2344];
        layer6[40][15:8] = buffer_data_0[2359:2352];
        layer6[40][23:16] = buffer_data_0[2367:2360];
        layer6[40][31:24] = buffer_data_0[2375:2368];
        layer6[40][39:32] = buffer_data_0[2383:2376];
        layer6[40][47:40] = buffer_data_0[2391:2384];
        layer6[40][55:48] = buffer_data_0[2399:2392];
        layer0[41][7:0] = buffer_data_6[2359:2352];
        layer0[41][15:8] = buffer_data_6[2367:2360];
        layer0[41][23:16] = buffer_data_6[2375:2368];
        layer0[41][31:24] = buffer_data_6[2383:2376];
        layer0[41][39:32] = buffer_data_6[2391:2384];
        layer0[41][47:40] = buffer_data_6[2399:2392];
        layer0[41][55:48] = buffer_data_6[2407:2400];
        layer1[41][7:0] = buffer_data_5[2359:2352];
        layer1[41][15:8] = buffer_data_5[2367:2360];
        layer1[41][23:16] = buffer_data_5[2375:2368];
        layer1[41][31:24] = buffer_data_5[2383:2376];
        layer1[41][39:32] = buffer_data_5[2391:2384];
        layer1[41][47:40] = buffer_data_5[2399:2392];
        layer1[41][55:48] = buffer_data_5[2407:2400];
        layer2[41][7:0] = buffer_data_4[2359:2352];
        layer2[41][15:8] = buffer_data_4[2367:2360];
        layer2[41][23:16] = buffer_data_4[2375:2368];
        layer2[41][31:24] = buffer_data_4[2383:2376];
        layer2[41][39:32] = buffer_data_4[2391:2384];
        layer2[41][47:40] = buffer_data_4[2399:2392];
        layer2[41][55:48] = buffer_data_4[2407:2400];
        layer3[41][7:0] = buffer_data_3[2359:2352];
        layer3[41][15:8] = buffer_data_3[2367:2360];
        layer3[41][23:16] = buffer_data_3[2375:2368];
        layer3[41][31:24] = buffer_data_3[2383:2376];
        layer3[41][39:32] = buffer_data_3[2391:2384];
        layer3[41][47:40] = buffer_data_3[2399:2392];
        layer3[41][55:48] = buffer_data_3[2407:2400];
        layer4[41][7:0] = buffer_data_2[2359:2352];
        layer4[41][15:8] = buffer_data_2[2367:2360];
        layer4[41][23:16] = buffer_data_2[2375:2368];
        layer4[41][31:24] = buffer_data_2[2383:2376];
        layer4[41][39:32] = buffer_data_2[2391:2384];
        layer4[41][47:40] = buffer_data_2[2399:2392];
        layer4[41][55:48] = buffer_data_2[2407:2400];
        layer5[41][7:0] = buffer_data_1[2359:2352];
        layer5[41][15:8] = buffer_data_1[2367:2360];
        layer5[41][23:16] = buffer_data_1[2375:2368];
        layer5[41][31:24] = buffer_data_1[2383:2376];
        layer5[41][39:32] = buffer_data_1[2391:2384];
        layer5[41][47:40] = buffer_data_1[2399:2392];
        layer5[41][55:48] = buffer_data_1[2407:2400];
        layer6[41][7:0] = buffer_data_0[2359:2352];
        layer6[41][15:8] = buffer_data_0[2367:2360];
        layer6[41][23:16] = buffer_data_0[2375:2368];
        layer6[41][31:24] = buffer_data_0[2383:2376];
        layer6[41][39:32] = buffer_data_0[2391:2384];
        layer6[41][47:40] = buffer_data_0[2399:2392];
        layer6[41][55:48] = buffer_data_0[2407:2400];
        layer0[42][7:0] = buffer_data_6[2367:2360];
        layer0[42][15:8] = buffer_data_6[2375:2368];
        layer0[42][23:16] = buffer_data_6[2383:2376];
        layer0[42][31:24] = buffer_data_6[2391:2384];
        layer0[42][39:32] = buffer_data_6[2399:2392];
        layer0[42][47:40] = buffer_data_6[2407:2400];
        layer0[42][55:48] = buffer_data_6[2415:2408];
        layer1[42][7:0] = buffer_data_5[2367:2360];
        layer1[42][15:8] = buffer_data_5[2375:2368];
        layer1[42][23:16] = buffer_data_5[2383:2376];
        layer1[42][31:24] = buffer_data_5[2391:2384];
        layer1[42][39:32] = buffer_data_5[2399:2392];
        layer1[42][47:40] = buffer_data_5[2407:2400];
        layer1[42][55:48] = buffer_data_5[2415:2408];
        layer2[42][7:0] = buffer_data_4[2367:2360];
        layer2[42][15:8] = buffer_data_4[2375:2368];
        layer2[42][23:16] = buffer_data_4[2383:2376];
        layer2[42][31:24] = buffer_data_4[2391:2384];
        layer2[42][39:32] = buffer_data_4[2399:2392];
        layer2[42][47:40] = buffer_data_4[2407:2400];
        layer2[42][55:48] = buffer_data_4[2415:2408];
        layer3[42][7:0] = buffer_data_3[2367:2360];
        layer3[42][15:8] = buffer_data_3[2375:2368];
        layer3[42][23:16] = buffer_data_3[2383:2376];
        layer3[42][31:24] = buffer_data_3[2391:2384];
        layer3[42][39:32] = buffer_data_3[2399:2392];
        layer3[42][47:40] = buffer_data_3[2407:2400];
        layer3[42][55:48] = buffer_data_3[2415:2408];
        layer4[42][7:0] = buffer_data_2[2367:2360];
        layer4[42][15:8] = buffer_data_2[2375:2368];
        layer4[42][23:16] = buffer_data_2[2383:2376];
        layer4[42][31:24] = buffer_data_2[2391:2384];
        layer4[42][39:32] = buffer_data_2[2399:2392];
        layer4[42][47:40] = buffer_data_2[2407:2400];
        layer4[42][55:48] = buffer_data_2[2415:2408];
        layer5[42][7:0] = buffer_data_1[2367:2360];
        layer5[42][15:8] = buffer_data_1[2375:2368];
        layer5[42][23:16] = buffer_data_1[2383:2376];
        layer5[42][31:24] = buffer_data_1[2391:2384];
        layer5[42][39:32] = buffer_data_1[2399:2392];
        layer5[42][47:40] = buffer_data_1[2407:2400];
        layer5[42][55:48] = buffer_data_1[2415:2408];
        layer6[42][7:0] = buffer_data_0[2367:2360];
        layer6[42][15:8] = buffer_data_0[2375:2368];
        layer6[42][23:16] = buffer_data_0[2383:2376];
        layer6[42][31:24] = buffer_data_0[2391:2384];
        layer6[42][39:32] = buffer_data_0[2399:2392];
        layer6[42][47:40] = buffer_data_0[2407:2400];
        layer6[42][55:48] = buffer_data_0[2415:2408];
        layer0[43][7:0] = buffer_data_6[2375:2368];
        layer0[43][15:8] = buffer_data_6[2383:2376];
        layer0[43][23:16] = buffer_data_6[2391:2384];
        layer0[43][31:24] = buffer_data_6[2399:2392];
        layer0[43][39:32] = buffer_data_6[2407:2400];
        layer0[43][47:40] = buffer_data_6[2415:2408];
        layer0[43][55:48] = buffer_data_6[2423:2416];
        layer1[43][7:0] = buffer_data_5[2375:2368];
        layer1[43][15:8] = buffer_data_5[2383:2376];
        layer1[43][23:16] = buffer_data_5[2391:2384];
        layer1[43][31:24] = buffer_data_5[2399:2392];
        layer1[43][39:32] = buffer_data_5[2407:2400];
        layer1[43][47:40] = buffer_data_5[2415:2408];
        layer1[43][55:48] = buffer_data_5[2423:2416];
        layer2[43][7:0] = buffer_data_4[2375:2368];
        layer2[43][15:8] = buffer_data_4[2383:2376];
        layer2[43][23:16] = buffer_data_4[2391:2384];
        layer2[43][31:24] = buffer_data_4[2399:2392];
        layer2[43][39:32] = buffer_data_4[2407:2400];
        layer2[43][47:40] = buffer_data_4[2415:2408];
        layer2[43][55:48] = buffer_data_4[2423:2416];
        layer3[43][7:0] = buffer_data_3[2375:2368];
        layer3[43][15:8] = buffer_data_3[2383:2376];
        layer3[43][23:16] = buffer_data_3[2391:2384];
        layer3[43][31:24] = buffer_data_3[2399:2392];
        layer3[43][39:32] = buffer_data_3[2407:2400];
        layer3[43][47:40] = buffer_data_3[2415:2408];
        layer3[43][55:48] = buffer_data_3[2423:2416];
        layer4[43][7:0] = buffer_data_2[2375:2368];
        layer4[43][15:8] = buffer_data_2[2383:2376];
        layer4[43][23:16] = buffer_data_2[2391:2384];
        layer4[43][31:24] = buffer_data_2[2399:2392];
        layer4[43][39:32] = buffer_data_2[2407:2400];
        layer4[43][47:40] = buffer_data_2[2415:2408];
        layer4[43][55:48] = buffer_data_2[2423:2416];
        layer5[43][7:0] = buffer_data_1[2375:2368];
        layer5[43][15:8] = buffer_data_1[2383:2376];
        layer5[43][23:16] = buffer_data_1[2391:2384];
        layer5[43][31:24] = buffer_data_1[2399:2392];
        layer5[43][39:32] = buffer_data_1[2407:2400];
        layer5[43][47:40] = buffer_data_1[2415:2408];
        layer5[43][55:48] = buffer_data_1[2423:2416];
        layer6[43][7:0] = buffer_data_0[2375:2368];
        layer6[43][15:8] = buffer_data_0[2383:2376];
        layer6[43][23:16] = buffer_data_0[2391:2384];
        layer6[43][31:24] = buffer_data_0[2399:2392];
        layer6[43][39:32] = buffer_data_0[2407:2400];
        layer6[43][47:40] = buffer_data_0[2415:2408];
        layer6[43][55:48] = buffer_data_0[2423:2416];
        layer0[44][7:0] = buffer_data_6[2383:2376];
        layer0[44][15:8] = buffer_data_6[2391:2384];
        layer0[44][23:16] = buffer_data_6[2399:2392];
        layer0[44][31:24] = buffer_data_6[2407:2400];
        layer0[44][39:32] = buffer_data_6[2415:2408];
        layer0[44][47:40] = buffer_data_6[2423:2416];
        layer0[44][55:48] = buffer_data_6[2431:2424];
        layer1[44][7:0] = buffer_data_5[2383:2376];
        layer1[44][15:8] = buffer_data_5[2391:2384];
        layer1[44][23:16] = buffer_data_5[2399:2392];
        layer1[44][31:24] = buffer_data_5[2407:2400];
        layer1[44][39:32] = buffer_data_5[2415:2408];
        layer1[44][47:40] = buffer_data_5[2423:2416];
        layer1[44][55:48] = buffer_data_5[2431:2424];
        layer2[44][7:0] = buffer_data_4[2383:2376];
        layer2[44][15:8] = buffer_data_4[2391:2384];
        layer2[44][23:16] = buffer_data_4[2399:2392];
        layer2[44][31:24] = buffer_data_4[2407:2400];
        layer2[44][39:32] = buffer_data_4[2415:2408];
        layer2[44][47:40] = buffer_data_4[2423:2416];
        layer2[44][55:48] = buffer_data_4[2431:2424];
        layer3[44][7:0] = buffer_data_3[2383:2376];
        layer3[44][15:8] = buffer_data_3[2391:2384];
        layer3[44][23:16] = buffer_data_3[2399:2392];
        layer3[44][31:24] = buffer_data_3[2407:2400];
        layer3[44][39:32] = buffer_data_3[2415:2408];
        layer3[44][47:40] = buffer_data_3[2423:2416];
        layer3[44][55:48] = buffer_data_3[2431:2424];
        layer4[44][7:0] = buffer_data_2[2383:2376];
        layer4[44][15:8] = buffer_data_2[2391:2384];
        layer4[44][23:16] = buffer_data_2[2399:2392];
        layer4[44][31:24] = buffer_data_2[2407:2400];
        layer4[44][39:32] = buffer_data_2[2415:2408];
        layer4[44][47:40] = buffer_data_2[2423:2416];
        layer4[44][55:48] = buffer_data_2[2431:2424];
        layer5[44][7:0] = buffer_data_1[2383:2376];
        layer5[44][15:8] = buffer_data_1[2391:2384];
        layer5[44][23:16] = buffer_data_1[2399:2392];
        layer5[44][31:24] = buffer_data_1[2407:2400];
        layer5[44][39:32] = buffer_data_1[2415:2408];
        layer5[44][47:40] = buffer_data_1[2423:2416];
        layer5[44][55:48] = buffer_data_1[2431:2424];
        layer6[44][7:0] = buffer_data_0[2383:2376];
        layer6[44][15:8] = buffer_data_0[2391:2384];
        layer6[44][23:16] = buffer_data_0[2399:2392];
        layer6[44][31:24] = buffer_data_0[2407:2400];
        layer6[44][39:32] = buffer_data_0[2415:2408];
        layer6[44][47:40] = buffer_data_0[2423:2416];
        layer6[44][55:48] = buffer_data_0[2431:2424];
        layer0[45][7:0] = buffer_data_6[2391:2384];
        layer0[45][15:8] = buffer_data_6[2399:2392];
        layer0[45][23:16] = buffer_data_6[2407:2400];
        layer0[45][31:24] = buffer_data_6[2415:2408];
        layer0[45][39:32] = buffer_data_6[2423:2416];
        layer0[45][47:40] = buffer_data_6[2431:2424];
        layer0[45][55:48] = buffer_data_6[2439:2432];
        layer1[45][7:0] = buffer_data_5[2391:2384];
        layer1[45][15:8] = buffer_data_5[2399:2392];
        layer1[45][23:16] = buffer_data_5[2407:2400];
        layer1[45][31:24] = buffer_data_5[2415:2408];
        layer1[45][39:32] = buffer_data_5[2423:2416];
        layer1[45][47:40] = buffer_data_5[2431:2424];
        layer1[45][55:48] = buffer_data_5[2439:2432];
        layer2[45][7:0] = buffer_data_4[2391:2384];
        layer2[45][15:8] = buffer_data_4[2399:2392];
        layer2[45][23:16] = buffer_data_4[2407:2400];
        layer2[45][31:24] = buffer_data_4[2415:2408];
        layer2[45][39:32] = buffer_data_4[2423:2416];
        layer2[45][47:40] = buffer_data_4[2431:2424];
        layer2[45][55:48] = buffer_data_4[2439:2432];
        layer3[45][7:0] = buffer_data_3[2391:2384];
        layer3[45][15:8] = buffer_data_3[2399:2392];
        layer3[45][23:16] = buffer_data_3[2407:2400];
        layer3[45][31:24] = buffer_data_3[2415:2408];
        layer3[45][39:32] = buffer_data_3[2423:2416];
        layer3[45][47:40] = buffer_data_3[2431:2424];
        layer3[45][55:48] = buffer_data_3[2439:2432];
        layer4[45][7:0] = buffer_data_2[2391:2384];
        layer4[45][15:8] = buffer_data_2[2399:2392];
        layer4[45][23:16] = buffer_data_2[2407:2400];
        layer4[45][31:24] = buffer_data_2[2415:2408];
        layer4[45][39:32] = buffer_data_2[2423:2416];
        layer4[45][47:40] = buffer_data_2[2431:2424];
        layer4[45][55:48] = buffer_data_2[2439:2432];
        layer5[45][7:0] = buffer_data_1[2391:2384];
        layer5[45][15:8] = buffer_data_1[2399:2392];
        layer5[45][23:16] = buffer_data_1[2407:2400];
        layer5[45][31:24] = buffer_data_1[2415:2408];
        layer5[45][39:32] = buffer_data_1[2423:2416];
        layer5[45][47:40] = buffer_data_1[2431:2424];
        layer5[45][55:48] = buffer_data_1[2439:2432];
        layer6[45][7:0] = buffer_data_0[2391:2384];
        layer6[45][15:8] = buffer_data_0[2399:2392];
        layer6[45][23:16] = buffer_data_0[2407:2400];
        layer6[45][31:24] = buffer_data_0[2415:2408];
        layer6[45][39:32] = buffer_data_0[2423:2416];
        layer6[45][47:40] = buffer_data_0[2431:2424];
        layer6[45][55:48] = buffer_data_0[2439:2432];
        layer0[46][7:0] = buffer_data_6[2399:2392];
        layer0[46][15:8] = buffer_data_6[2407:2400];
        layer0[46][23:16] = buffer_data_6[2415:2408];
        layer0[46][31:24] = buffer_data_6[2423:2416];
        layer0[46][39:32] = buffer_data_6[2431:2424];
        layer0[46][47:40] = buffer_data_6[2439:2432];
        layer0[46][55:48] = buffer_data_6[2447:2440];
        layer1[46][7:0] = buffer_data_5[2399:2392];
        layer1[46][15:8] = buffer_data_5[2407:2400];
        layer1[46][23:16] = buffer_data_5[2415:2408];
        layer1[46][31:24] = buffer_data_5[2423:2416];
        layer1[46][39:32] = buffer_data_5[2431:2424];
        layer1[46][47:40] = buffer_data_5[2439:2432];
        layer1[46][55:48] = buffer_data_5[2447:2440];
        layer2[46][7:0] = buffer_data_4[2399:2392];
        layer2[46][15:8] = buffer_data_4[2407:2400];
        layer2[46][23:16] = buffer_data_4[2415:2408];
        layer2[46][31:24] = buffer_data_4[2423:2416];
        layer2[46][39:32] = buffer_data_4[2431:2424];
        layer2[46][47:40] = buffer_data_4[2439:2432];
        layer2[46][55:48] = buffer_data_4[2447:2440];
        layer3[46][7:0] = buffer_data_3[2399:2392];
        layer3[46][15:8] = buffer_data_3[2407:2400];
        layer3[46][23:16] = buffer_data_3[2415:2408];
        layer3[46][31:24] = buffer_data_3[2423:2416];
        layer3[46][39:32] = buffer_data_3[2431:2424];
        layer3[46][47:40] = buffer_data_3[2439:2432];
        layer3[46][55:48] = buffer_data_3[2447:2440];
        layer4[46][7:0] = buffer_data_2[2399:2392];
        layer4[46][15:8] = buffer_data_2[2407:2400];
        layer4[46][23:16] = buffer_data_2[2415:2408];
        layer4[46][31:24] = buffer_data_2[2423:2416];
        layer4[46][39:32] = buffer_data_2[2431:2424];
        layer4[46][47:40] = buffer_data_2[2439:2432];
        layer4[46][55:48] = buffer_data_2[2447:2440];
        layer5[46][7:0] = buffer_data_1[2399:2392];
        layer5[46][15:8] = buffer_data_1[2407:2400];
        layer5[46][23:16] = buffer_data_1[2415:2408];
        layer5[46][31:24] = buffer_data_1[2423:2416];
        layer5[46][39:32] = buffer_data_1[2431:2424];
        layer5[46][47:40] = buffer_data_1[2439:2432];
        layer5[46][55:48] = buffer_data_1[2447:2440];
        layer6[46][7:0] = buffer_data_0[2399:2392];
        layer6[46][15:8] = buffer_data_0[2407:2400];
        layer6[46][23:16] = buffer_data_0[2415:2408];
        layer6[46][31:24] = buffer_data_0[2423:2416];
        layer6[46][39:32] = buffer_data_0[2431:2424];
        layer6[46][47:40] = buffer_data_0[2439:2432];
        layer6[46][55:48] = buffer_data_0[2447:2440];
        layer0[47][7:0] = buffer_data_6[2407:2400];
        layer0[47][15:8] = buffer_data_6[2415:2408];
        layer0[47][23:16] = buffer_data_6[2423:2416];
        layer0[47][31:24] = buffer_data_6[2431:2424];
        layer0[47][39:32] = buffer_data_6[2439:2432];
        layer0[47][47:40] = buffer_data_6[2447:2440];
        layer0[47][55:48] = buffer_data_6[2455:2448];
        layer1[47][7:0] = buffer_data_5[2407:2400];
        layer1[47][15:8] = buffer_data_5[2415:2408];
        layer1[47][23:16] = buffer_data_5[2423:2416];
        layer1[47][31:24] = buffer_data_5[2431:2424];
        layer1[47][39:32] = buffer_data_5[2439:2432];
        layer1[47][47:40] = buffer_data_5[2447:2440];
        layer1[47][55:48] = buffer_data_5[2455:2448];
        layer2[47][7:0] = buffer_data_4[2407:2400];
        layer2[47][15:8] = buffer_data_4[2415:2408];
        layer2[47][23:16] = buffer_data_4[2423:2416];
        layer2[47][31:24] = buffer_data_4[2431:2424];
        layer2[47][39:32] = buffer_data_4[2439:2432];
        layer2[47][47:40] = buffer_data_4[2447:2440];
        layer2[47][55:48] = buffer_data_4[2455:2448];
        layer3[47][7:0] = buffer_data_3[2407:2400];
        layer3[47][15:8] = buffer_data_3[2415:2408];
        layer3[47][23:16] = buffer_data_3[2423:2416];
        layer3[47][31:24] = buffer_data_3[2431:2424];
        layer3[47][39:32] = buffer_data_3[2439:2432];
        layer3[47][47:40] = buffer_data_3[2447:2440];
        layer3[47][55:48] = buffer_data_3[2455:2448];
        layer4[47][7:0] = buffer_data_2[2407:2400];
        layer4[47][15:8] = buffer_data_2[2415:2408];
        layer4[47][23:16] = buffer_data_2[2423:2416];
        layer4[47][31:24] = buffer_data_2[2431:2424];
        layer4[47][39:32] = buffer_data_2[2439:2432];
        layer4[47][47:40] = buffer_data_2[2447:2440];
        layer4[47][55:48] = buffer_data_2[2455:2448];
        layer5[47][7:0] = buffer_data_1[2407:2400];
        layer5[47][15:8] = buffer_data_1[2415:2408];
        layer5[47][23:16] = buffer_data_1[2423:2416];
        layer5[47][31:24] = buffer_data_1[2431:2424];
        layer5[47][39:32] = buffer_data_1[2439:2432];
        layer5[47][47:40] = buffer_data_1[2447:2440];
        layer5[47][55:48] = buffer_data_1[2455:2448];
        layer6[47][7:0] = buffer_data_0[2407:2400];
        layer6[47][15:8] = buffer_data_0[2415:2408];
        layer6[47][23:16] = buffer_data_0[2423:2416];
        layer6[47][31:24] = buffer_data_0[2431:2424];
        layer6[47][39:32] = buffer_data_0[2439:2432];
        layer6[47][47:40] = buffer_data_0[2447:2440];
        layer6[47][55:48] = buffer_data_0[2455:2448];
        layer0[48][7:0] = buffer_data_6[2415:2408];
        layer0[48][15:8] = buffer_data_6[2423:2416];
        layer0[48][23:16] = buffer_data_6[2431:2424];
        layer0[48][31:24] = buffer_data_6[2439:2432];
        layer0[48][39:32] = buffer_data_6[2447:2440];
        layer0[48][47:40] = buffer_data_6[2455:2448];
        layer0[48][55:48] = buffer_data_6[2463:2456];
        layer1[48][7:0] = buffer_data_5[2415:2408];
        layer1[48][15:8] = buffer_data_5[2423:2416];
        layer1[48][23:16] = buffer_data_5[2431:2424];
        layer1[48][31:24] = buffer_data_5[2439:2432];
        layer1[48][39:32] = buffer_data_5[2447:2440];
        layer1[48][47:40] = buffer_data_5[2455:2448];
        layer1[48][55:48] = buffer_data_5[2463:2456];
        layer2[48][7:0] = buffer_data_4[2415:2408];
        layer2[48][15:8] = buffer_data_4[2423:2416];
        layer2[48][23:16] = buffer_data_4[2431:2424];
        layer2[48][31:24] = buffer_data_4[2439:2432];
        layer2[48][39:32] = buffer_data_4[2447:2440];
        layer2[48][47:40] = buffer_data_4[2455:2448];
        layer2[48][55:48] = buffer_data_4[2463:2456];
        layer3[48][7:0] = buffer_data_3[2415:2408];
        layer3[48][15:8] = buffer_data_3[2423:2416];
        layer3[48][23:16] = buffer_data_3[2431:2424];
        layer3[48][31:24] = buffer_data_3[2439:2432];
        layer3[48][39:32] = buffer_data_3[2447:2440];
        layer3[48][47:40] = buffer_data_3[2455:2448];
        layer3[48][55:48] = buffer_data_3[2463:2456];
        layer4[48][7:0] = buffer_data_2[2415:2408];
        layer4[48][15:8] = buffer_data_2[2423:2416];
        layer4[48][23:16] = buffer_data_2[2431:2424];
        layer4[48][31:24] = buffer_data_2[2439:2432];
        layer4[48][39:32] = buffer_data_2[2447:2440];
        layer4[48][47:40] = buffer_data_2[2455:2448];
        layer4[48][55:48] = buffer_data_2[2463:2456];
        layer5[48][7:0] = buffer_data_1[2415:2408];
        layer5[48][15:8] = buffer_data_1[2423:2416];
        layer5[48][23:16] = buffer_data_1[2431:2424];
        layer5[48][31:24] = buffer_data_1[2439:2432];
        layer5[48][39:32] = buffer_data_1[2447:2440];
        layer5[48][47:40] = buffer_data_1[2455:2448];
        layer5[48][55:48] = buffer_data_1[2463:2456];
        layer6[48][7:0] = buffer_data_0[2415:2408];
        layer6[48][15:8] = buffer_data_0[2423:2416];
        layer6[48][23:16] = buffer_data_0[2431:2424];
        layer6[48][31:24] = buffer_data_0[2439:2432];
        layer6[48][39:32] = buffer_data_0[2447:2440];
        layer6[48][47:40] = buffer_data_0[2455:2448];
        layer6[48][55:48] = buffer_data_0[2463:2456];
        layer0[49][7:0] = buffer_data_6[2423:2416];
        layer0[49][15:8] = buffer_data_6[2431:2424];
        layer0[49][23:16] = buffer_data_6[2439:2432];
        layer0[49][31:24] = buffer_data_6[2447:2440];
        layer0[49][39:32] = buffer_data_6[2455:2448];
        layer0[49][47:40] = buffer_data_6[2463:2456];
        layer0[49][55:48] = buffer_data_6[2471:2464];
        layer1[49][7:0] = buffer_data_5[2423:2416];
        layer1[49][15:8] = buffer_data_5[2431:2424];
        layer1[49][23:16] = buffer_data_5[2439:2432];
        layer1[49][31:24] = buffer_data_5[2447:2440];
        layer1[49][39:32] = buffer_data_5[2455:2448];
        layer1[49][47:40] = buffer_data_5[2463:2456];
        layer1[49][55:48] = buffer_data_5[2471:2464];
        layer2[49][7:0] = buffer_data_4[2423:2416];
        layer2[49][15:8] = buffer_data_4[2431:2424];
        layer2[49][23:16] = buffer_data_4[2439:2432];
        layer2[49][31:24] = buffer_data_4[2447:2440];
        layer2[49][39:32] = buffer_data_4[2455:2448];
        layer2[49][47:40] = buffer_data_4[2463:2456];
        layer2[49][55:48] = buffer_data_4[2471:2464];
        layer3[49][7:0] = buffer_data_3[2423:2416];
        layer3[49][15:8] = buffer_data_3[2431:2424];
        layer3[49][23:16] = buffer_data_3[2439:2432];
        layer3[49][31:24] = buffer_data_3[2447:2440];
        layer3[49][39:32] = buffer_data_3[2455:2448];
        layer3[49][47:40] = buffer_data_3[2463:2456];
        layer3[49][55:48] = buffer_data_3[2471:2464];
        layer4[49][7:0] = buffer_data_2[2423:2416];
        layer4[49][15:8] = buffer_data_2[2431:2424];
        layer4[49][23:16] = buffer_data_2[2439:2432];
        layer4[49][31:24] = buffer_data_2[2447:2440];
        layer4[49][39:32] = buffer_data_2[2455:2448];
        layer4[49][47:40] = buffer_data_2[2463:2456];
        layer4[49][55:48] = buffer_data_2[2471:2464];
        layer5[49][7:0] = buffer_data_1[2423:2416];
        layer5[49][15:8] = buffer_data_1[2431:2424];
        layer5[49][23:16] = buffer_data_1[2439:2432];
        layer5[49][31:24] = buffer_data_1[2447:2440];
        layer5[49][39:32] = buffer_data_1[2455:2448];
        layer5[49][47:40] = buffer_data_1[2463:2456];
        layer5[49][55:48] = buffer_data_1[2471:2464];
        layer6[49][7:0] = buffer_data_0[2423:2416];
        layer6[49][15:8] = buffer_data_0[2431:2424];
        layer6[49][23:16] = buffer_data_0[2439:2432];
        layer6[49][31:24] = buffer_data_0[2447:2440];
        layer6[49][39:32] = buffer_data_0[2455:2448];
        layer6[49][47:40] = buffer_data_0[2463:2456];
        layer6[49][55:48] = buffer_data_0[2471:2464];
        layer0[50][7:0] = buffer_data_6[2431:2424];
        layer0[50][15:8] = buffer_data_6[2439:2432];
        layer0[50][23:16] = buffer_data_6[2447:2440];
        layer0[50][31:24] = buffer_data_6[2455:2448];
        layer0[50][39:32] = buffer_data_6[2463:2456];
        layer0[50][47:40] = buffer_data_6[2471:2464];
        layer0[50][55:48] = buffer_data_6[2479:2472];
        layer1[50][7:0] = buffer_data_5[2431:2424];
        layer1[50][15:8] = buffer_data_5[2439:2432];
        layer1[50][23:16] = buffer_data_5[2447:2440];
        layer1[50][31:24] = buffer_data_5[2455:2448];
        layer1[50][39:32] = buffer_data_5[2463:2456];
        layer1[50][47:40] = buffer_data_5[2471:2464];
        layer1[50][55:48] = buffer_data_5[2479:2472];
        layer2[50][7:0] = buffer_data_4[2431:2424];
        layer2[50][15:8] = buffer_data_4[2439:2432];
        layer2[50][23:16] = buffer_data_4[2447:2440];
        layer2[50][31:24] = buffer_data_4[2455:2448];
        layer2[50][39:32] = buffer_data_4[2463:2456];
        layer2[50][47:40] = buffer_data_4[2471:2464];
        layer2[50][55:48] = buffer_data_4[2479:2472];
        layer3[50][7:0] = buffer_data_3[2431:2424];
        layer3[50][15:8] = buffer_data_3[2439:2432];
        layer3[50][23:16] = buffer_data_3[2447:2440];
        layer3[50][31:24] = buffer_data_3[2455:2448];
        layer3[50][39:32] = buffer_data_3[2463:2456];
        layer3[50][47:40] = buffer_data_3[2471:2464];
        layer3[50][55:48] = buffer_data_3[2479:2472];
        layer4[50][7:0] = buffer_data_2[2431:2424];
        layer4[50][15:8] = buffer_data_2[2439:2432];
        layer4[50][23:16] = buffer_data_2[2447:2440];
        layer4[50][31:24] = buffer_data_2[2455:2448];
        layer4[50][39:32] = buffer_data_2[2463:2456];
        layer4[50][47:40] = buffer_data_2[2471:2464];
        layer4[50][55:48] = buffer_data_2[2479:2472];
        layer5[50][7:0] = buffer_data_1[2431:2424];
        layer5[50][15:8] = buffer_data_1[2439:2432];
        layer5[50][23:16] = buffer_data_1[2447:2440];
        layer5[50][31:24] = buffer_data_1[2455:2448];
        layer5[50][39:32] = buffer_data_1[2463:2456];
        layer5[50][47:40] = buffer_data_1[2471:2464];
        layer5[50][55:48] = buffer_data_1[2479:2472];
        layer6[50][7:0] = buffer_data_0[2431:2424];
        layer6[50][15:8] = buffer_data_0[2439:2432];
        layer6[50][23:16] = buffer_data_0[2447:2440];
        layer6[50][31:24] = buffer_data_0[2455:2448];
        layer6[50][39:32] = buffer_data_0[2463:2456];
        layer6[50][47:40] = buffer_data_0[2471:2464];
        layer6[50][55:48] = buffer_data_0[2479:2472];
        layer0[51][7:0] = buffer_data_6[2439:2432];
        layer0[51][15:8] = buffer_data_6[2447:2440];
        layer0[51][23:16] = buffer_data_6[2455:2448];
        layer0[51][31:24] = buffer_data_6[2463:2456];
        layer0[51][39:32] = buffer_data_6[2471:2464];
        layer0[51][47:40] = buffer_data_6[2479:2472];
        layer0[51][55:48] = buffer_data_6[2487:2480];
        layer1[51][7:0] = buffer_data_5[2439:2432];
        layer1[51][15:8] = buffer_data_5[2447:2440];
        layer1[51][23:16] = buffer_data_5[2455:2448];
        layer1[51][31:24] = buffer_data_5[2463:2456];
        layer1[51][39:32] = buffer_data_5[2471:2464];
        layer1[51][47:40] = buffer_data_5[2479:2472];
        layer1[51][55:48] = buffer_data_5[2487:2480];
        layer2[51][7:0] = buffer_data_4[2439:2432];
        layer2[51][15:8] = buffer_data_4[2447:2440];
        layer2[51][23:16] = buffer_data_4[2455:2448];
        layer2[51][31:24] = buffer_data_4[2463:2456];
        layer2[51][39:32] = buffer_data_4[2471:2464];
        layer2[51][47:40] = buffer_data_4[2479:2472];
        layer2[51][55:48] = buffer_data_4[2487:2480];
        layer3[51][7:0] = buffer_data_3[2439:2432];
        layer3[51][15:8] = buffer_data_3[2447:2440];
        layer3[51][23:16] = buffer_data_3[2455:2448];
        layer3[51][31:24] = buffer_data_3[2463:2456];
        layer3[51][39:32] = buffer_data_3[2471:2464];
        layer3[51][47:40] = buffer_data_3[2479:2472];
        layer3[51][55:48] = buffer_data_3[2487:2480];
        layer4[51][7:0] = buffer_data_2[2439:2432];
        layer4[51][15:8] = buffer_data_2[2447:2440];
        layer4[51][23:16] = buffer_data_2[2455:2448];
        layer4[51][31:24] = buffer_data_2[2463:2456];
        layer4[51][39:32] = buffer_data_2[2471:2464];
        layer4[51][47:40] = buffer_data_2[2479:2472];
        layer4[51][55:48] = buffer_data_2[2487:2480];
        layer5[51][7:0] = buffer_data_1[2439:2432];
        layer5[51][15:8] = buffer_data_1[2447:2440];
        layer5[51][23:16] = buffer_data_1[2455:2448];
        layer5[51][31:24] = buffer_data_1[2463:2456];
        layer5[51][39:32] = buffer_data_1[2471:2464];
        layer5[51][47:40] = buffer_data_1[2479:2472];
        layer5[51][55:48] = buffer_data_1[2487:2480];
        layer6[51][7:0] = buffer_data_0[2439:2432];
        layer6[51][15:8] = buffer_data_0[2447:2440];
        layer6[51][23:16] = buffer_data_0[2455:2448];
        layer6[51][31:24] = buffer_data_0[2463:2456];
        layer6[51][39:32] = buffer_data_0[2471:2464];
        layer6[51][47:40] = buffer_data_0[2479:2472];
        layer6[51][55:48] = buffer_data_0[2487:2480];
        layer0[52][7:0] = buffer_data_6[2447:2440];
        layer0[52][15:8] = buffer_data_6[2455:2448];
        layer0[52][23:16] = buffer_data_6[2463:2456];
        layer0[52][31:24] = buffer_data_6[2471:2464];
        layer0[52][39:32] = buffer_data_6[2479:2472];
        layer0[52][47:40] = buffer_data_6[2487:2480];
        layer0[52][55:48] = buffer_data_6[2495:2488];
        layer1[52][7:0] = buffer_data_5[2447:2440];
        layer1[52][15:8] = buffer_data_5[2455:2448];
        layer1[52][23:16] = buffer_data_5[2463:2456];
        layer1[52][31:24] = buffer_data_5[2471:2464];
        layer1[52][39:32] = buffer_data_5[2479:2472];
        layer1[52][47:40] = buffer_data_5[2487:2480];
        layer1[52][55:48] = buffer_data_5[2495:2488];
        layer2[52][7:0] = buffer_data_4[2447:2440];
        layer2[52][15:8] = buffer_data_4[2455:2448];
        layer2[52][23:16] = buffer_data_4[2463:2456];
        layer2[52][31:24] = buffer_data_4[2471:2464];
        layer2[52][39:32] = buffer_data_4[2479:2472];
        layer2[52][47:40] = buffer_data_4[2487:2480];
        layer2[52][55:48] = buffer_data_4[2495:2488];
        layer3[52][7:0] = buffer_data_3[2447:2440];
        layer3[52][15:8] = buffer_data_3[2455:2448];
        layer3[52][23:16] = buffer_data_3[2463:2456];
        layer3[52][31:24] = buffer_data_3[2471:2464];
        layer3[52][39:32] = buffer_data_3[2479:2472];
        layer3[52][47:40] = buffer_data_3[2487:2480];
        layer3[52][55:48] = buffer_data_3[2495:2488];
        layer4[52][7:0] = buffer_data_2[2447:2440];
        layer4[52][15:8] = buffer_data_2[2455:2448];
        layer4[52][23:16] = buffer_data_2[2463:2456];
        layer4[52][31:24] = buffer_data_2[2471:2464];
        layer4[52][39:32] = buffer_data_2[2479:2472];
        layer4[52][47:40] = buffer_data_2[2487:2480];
        layer4[52][55:48] = buffer_data_2[2495:2488];
        layer5[52][7:0] = buffer_data_1[2447:2440];
        layer5[52][15:8] = buffer_data_1[2455:2448];
        layer5[52][23:16] = buffer_data_1[2463:2456];
        layer5[52][31:24] = buffer_data_1[2471:2464];
        layer5[52][39:32] = buffer_data_1[2479:2472];
        layer5[52][47:40] = buffer_data_1[2487:2480];
        layer5[52][55:48] = buffer_data_1[2495:2488];
        layer6[52][7:0] = buffer_data_0[2447:2440];
        layer6[52][15:8] = buffer_data_0[2455:2448];
        layer6[52][23:16] = buffer_data_0[2463:2456];
        layer6[52][31:24] = buffer_data_0[2471:2464];
        layer6[52][39:32] = buffer_data_0[2479:2472];
        layer6[52][47:40] = buffer_data_0[2487:2480];
        layer6[52][55:48] = buffer_data_0[2495:2488];
        layer0[53][7:0] = buffer_data_6[2455:2448];
        layer0[53][15:8] = buffer_data_6[2463:2456];
        layer0[53][23:16] = buffer_data_6[2471:2464];
        layer0[53][31:24] = buffer_data_6[2479:2472];
        layer0[53][39:32] = buffer_data_6[2487:2480];
        layer0[53][47:40] = buffer_data_6[2495:2488];
        layer0[53][55:48] = buffer_data_6[2503:2496];
        layer1[53][7:0] = buffer_data_5[2455:2448];
        layer1[53][15:8] = buffer_data_5[2463:2456];
        layer1[53][23:16] = buffer_data_5[2471:2464];
        layer1[53][31:24] = buffer_data_5[2479:2472];
        layer1[53][39:32] = buffer_data_5[2487:2480];
        layer1[53][47:40] = buffer_data_5[2495:2488];
        layer1[53][55:48] = buffer_data_5[2503:2496];
        layer2[53][7:0] = buffer_data_4[2455:2448];
        layer2[53][15:8] = buffer_data_4[2463:2456];
        layer2[53][23:16] = buffer_data_4[2471:2464];
        layer2[53][31:24] = buffer_data_4[2479:2472];
        layer2[53][39:32] = buffer_data_4[2487:2480];
        layer2[53][47:40] = buffer_data_4[2495:2488];
        layer2[53][55:48] = buffer_data_4[2503:2496];
        layer3[53][7:0] = buffer_data_3[2455:2448];
        layer3[53][15:8] = buffer_data_3[2463:2456];
        layer3[53][23:16] = buffer_data_3[2471:2464];
        layer3[53][31:24] = buffer_data_3[2479:2472];
        layer3[53][39:32] = buffer_data_3[2487:2480];
        layer3[53][47:40] = buffer_data_3[2495:2488];
        layer3[53][55:48] = buffer_data_3[2503:2496];
        layer4[53][7:0] = buffer_data_2[2455:2448];
        layer4[53][15:8] = buffer_data_2[2463:2456];
        layer4[53][23:16] = buffer_data_2[2471:2464];
        layer4[53][31:24] = buffer_data_2[2479:2472];
        layer4[53][39:32] = buffer_data_2[2487:2480];
        layer4[53][47:40] = buffer_data_2[2495:2488];
        layer4[53][55:48] = buffer_data_2[2503:2496];
        layer5[53][7:0] = buffer_data_1[2455:2448];
        layer5[53][15:8] = buffer_data_1[2463:2456];
        layer5[53][23:16] = buffer_data_1[2471:2464];
        layer5[53][31:24] = buffer_data_1[2479:2472];
        layer5[53][39:32] = buffer_data_1[2487:2480];
        layer5[53][47:40] = buffer_data_1[2495:2488];
        layer5[53][55:48] = buffer_data_1[2503:2496];
        layer6[53][7:0] = buffer_data_0[2455:2448];
        layer6[53][15:8] = buffer_data_0[2463:2456];
        layer6[53][23:16] = buffer_data_0[2471:2464];
        layer6[53][31:24] = buffer_data_0[2479:2472];
        layer6[53][39:32] = buffer_data_0[2487:2480];
        layer6[53][47:40] = buffer_data_0[2495:2488];
        layer6[53][55:48] = buffer_data_0[2503:2496];
        layer0[54][7:0] = buffer_data_6[2463:2456];
        layer0[54][15:8] = buffer_data_6[2471:2464];
        layer0[54][23:16] = buffer_data_6[2479:2472];
        layer0[54][31:24] = buffer_data_6[2487:2480];
        layer0[54][39:32] = buffer_data_6[2495:2488];
        layer0[54][47:40] = buffer_data_6[2503:2496];
        layer0[54][55:48] = buffer_data_6[2511:2504];
        layer1[54][7:0] = buffer_data_5[2463:2456];
        layer1[54][15:8] = buffer_data_5[2471:2464];
        layer1[54][23:16] = buffer_data_5[2479:2472];
        layer1[54][31:24] = buffer_data_5[2487:2480];
        layer1[54][39:32] = buffer_data_5[2495:2488];
        layer1[54][47:40] = buffer_data_5[2503:2496];
        layer1[54][55:48] = buffer_data_5[2511:2504];
        layer2[54][7:0] = buffer_data_4[2463:2456];
        layer2[54][15:8] = buffer_data_4[2471:2464];
        layer2[54][23:16] = buffer_data_4[2479:2472];
        layer2[54][31:24] = buffer_data_4[2487:2480];
        layer2[54][39:32] = buffer_data_4[2495:2488];
        layer2[54][47:40] = buffer_data_4[2503:2496];
        layer2[54][55:48] = buffer_data_4[2511:2504];
        layer3[54][7:0] = buffer_data_3[2463:2456];
        layer3[54][15:8] = buffer_data_3[2471:2464];
        layer3[54][23:16] = buffer_data_3[2479:2472];
        layer3[54][31:24] = buffer_data_3[2487:2480];
        layer3[54][39:32] = buffer_data_3[2495:2488];
        layer3[54][47:40] = buffer_data_3[2503:2496];
        layer3[54][55:48] = buffer_data_3[2511:2504];
        layer4[54][7:0] = buffer_data_2[2463:2456];
        layer4[54][15:8] = buffer_data_2[2471:2464];
        layer4[54][23:16] = buffer_data_2[2479:2472];
        layer4[54][31:24] = buffer_data_2[2487:2480];
        layer4[54][39:32] = buffer_data_2[2495:2488];
        layer4[54][47:40] = buffer_data_2[2503:2496];
        layer4[54][55:48] = buffer_data_2[2511:2504];
        layer5[54][7:0] = buffer_data_1[2463:2456];
        layer5[54][15:8] = buffer_data_1[2471:2464];
        layer5[54][23:16] = buffer_data_1[2479:2472];
        layer5[54][31:24] = buffer_data_1[2487:2480];
        layer5[54][39:32] = buffer_data_1[2495:2488];
        layer5[54][47:40] = buffer_data_1[2503:2496];
        layer5[54][55:48] = buffer_data_1[2511:2504];
        layer6[54][7:0] = buffer_data_0[2463:2456];
        layer6[54][15:8] = buffer_data_0[2471:2464];
        layer6[54][23:16] = buffer_data_0[2479:2472];
        layer6[54][31:24] = buffer_data_0[2487:2480];
        layer6[54][39:32] = buffer_data_0[2495:2488];
        layer6[54][47:40] = buffer_data_0[2503:2496];
        layer6[54][55:48] = buffer_data_0[2511:2504];
        layer0[55][7:0] = buffer_data_6[2471:2464];
        layer0[55][15:8] = buffer_data_6[2479:2472];
        layer0[55][23:16] = buffer_data_6[2487:2480];
        layer0[55][31:24] = buffer_data_6[2495:2488];
        layer0[55][39:32] = buffer_data_6[2503:2496];
        layer0[55][47:40] = buffer_data_6[2511:2504];
        layer0[55][55:48] = buffer_data_6[2519:2512];
        layer1[55][7:0] = buffer_data_5[2471:2464];
        layer1[55][15:8] = buffer_data_5[2479:2472];
        layer1[55][23:16] = buffer_data_5[2487:2480];
        layer1[55][31:24] = buffer_data_5[2495:2488];
        layer1[55][39:32] = buffer_data_5[2503:2496];
        layer1[55][47:40] = buffer_data_5[2511:2504];
        layer1[55][55:48] = buffer_data_5[2519:2512];
        layer2[55][7:0] = buffer_data_4[2471:2464];
        layer2[55][15:8] = buffer_data_4[2479:2472];
        layer2[55][23:16] = buffer_data_4[2487:2480];
        layer2[55][31:24] = buffer_data_4[2495:2488];
        layer2[55][39:32] = buffer_data_4[2503:2496];
        layer2[55][47:40] = buffer_data_4[2511:2504];
        layer2[55][55:48] = buffer_data_4[2519:2512];
        layer3[55][7:0] = buffer_data_3[2471:2464];
        layer3[55][15:8] = buffer_data_3[2479:2472];
        layer3[55][23:16] = buffer_data_3[2487:2480];
        layer3[55][31:24] = buffer_data_3[2495:2488];
        layer3[55][39:32] = buffer_data_3[2503:2496];
        layer3[55][47:40] = buffer_data_3[2511:2504];
        layer3[55][55:48] = buffer_data_3[2519:2512];
        layer4[55][7:0] = buffer_data_2[2471:2464];
        layer4[55][15:8] = buffer_data_2[2479:2472];
        layer4[55][23:16] = buffer_data_2[2487:2480];
        layer4[55][31:24] = buffer_data_2[2495:2488];
        layer4[55][39:32] = buffer_data_2[2503:2496];
        layer4[55][47:40] = buffer_data_2[2511:2504];
        layer4[55][55:48] = buffer_data_2[2519:2512];
        layer5[55][7:0] = buffer_data_1[2471:2464];
        layer5[55][15:8] = buffer_data_1[2479:2472];
        layer5[55][23:16] = buffer_data_1[2487:2480];
        layer5[55][31:24] = buffer_data_1[2495:2488];
        layer5[55][39:32] = buffer_data_1[2503:2496];
        layer5[55][47:40] = buffer_data_1[2511:2504];
        layer5[55][55:48] = buffer_data_1[2519:2512];
        layer6[55][7:0] = buffer_data_0[2471:2464];
        layer6[55][15:8] = buffer_data_0[2479:2472];
        layer6[55][23:16] = buffer_data_0[2487:2480];
        layer6[55][31:24] = buffer_data_0[2495:2488];
        layer6[55][39:32] = buffer_data_0[2503:2496];
        layer6[55][47:40] = buffer_data_0[2511:2504];
        layer6[55][55:48] = buffer_data_0[2519:2512];
        layer0[56][7:0] = buffer_data_6[2479:2472];
        layer0[56][15:8] = buffer_data_6[2487:2480];
        layer0[56][23:16] = buffer_data_6[2495:2488];
        layer0[56][31:24] = buffer_data_6[2503:2496];
        layer0[56][39:32] = buffer_data_6[2511:2504];
        layer0[56][47:40] = buffer_data_6[2519:2512];
        layer0[56][55:48] = buffer_data_6[2527:2520];
        layer1[56][7:0] = buffer_data_5[2479:2472];
        layer1[56][15:8] = buffer_data_5[2487:2480];
        layer1[56][23:16] = buffer_data_5[2495:2488];
        layer1[56][31:24] = buffer_data_5[2503:2496];
        layer1[56][39:32] = buffer_data_5[2511:2504];
        layer1[56][47:40] = buffer_data_5[2519:2512];
        layer1[56][55:48] = buffer_data_5[2527:2520];
        layer2[56][7:0] = buffer_data_4[2479:2472];
        layer2[56][15:8] = buffer_data_4[2487:2480];
        layer2[56][23:16] = buffer_data_4[2495:2488];
        layer2[56][31:24] = buffer_data_4[2503:2496];
        layer2[56][39:32] = buffer_data_4[2511:2504];
        layer2[56][47:40] = buffer_data_4[2519:2512];
        layer2[56][55:48] = buffer_data_4[2527:2520];
        layer3[56][7:0] = buffer_data_3[2479:2472];
        layer3[56][15:8] = buffer_data_3[2487:2480];
        layer3[56][23:16] = buffer_data_3[2495:2488];
        layer3[56][31:24] = buffer_data_3[2503:2496];
        layer3[56][39:32] = buffer_data_3[2511:2504];
        layer3[56][47:40] = buffer_data_3[2519:2512];
        layer3[56][55:48] = buffer_data_3[2527:2520];
        layer4[56][7:0] = buffer_data_2[2479:2472];
        layer4[56][15:8] = buffer_data_2[2487:2480];
        layer4[56][23:16] = buffer_data_2[2495:2488];
        layer4[56][31:24] = buffer_data_2[2503:2496];
        layer4[56][39:32] = buffer_data_2[2511:2504];
        layer4[56][47:40] = buffer_data_2[2519:2512];
        layer4[56][55:48] = buffer_data_2[2527:2520];
        layer5[56][7:0] = buffer_data_1[2479:2472];
        layer5[56][15:8] = buffer_data_1[2487:2480];
        layer5[56][23:16] = buffer_data_1[2495:2488];
        layer5[56][31:24] = buffer_data_1[2503:2496];
        layer5[56][39:32] = buffer_data_1[2511:2504];
        layer5[56][47:40] = buffer_data_1[2519:2512];
        layer5[56][55:48] = buffer_data_1[2527:2520];
        layer6[56][7:0] = buffer_data_0[2479:2472];
        layer6[56][15:8] = buffer_data_0[2487:2480];
        layer6[56][23:16] = buffer_data_0[2495:2488];
        layer6[56][31:24] = buffer_data_0[2503:2496];
        layer6[56][39:32] = buffer_data_0[2511:2504];
        layer6[56][47:40] = buffer_data_0[2519:2512];
        layer6[56][55:48] = buffer_data_0[2527:2520];
        layer0[57][7:0] = buffer_data_6[2487:2480];
        layer0[57][15:8] = buffer_data_6[2495:2488];
        layer0[57][23:16] = buffer_data_6[2503:2496];
        layer0[57][31:24] = buffer_data_6[2511:2504];
        layer0[57][39:32] = buffer_data_6[2519:2512];
        layer0[57][47:40] = buffer_data_6[2527:2520];
        layer0[57][55:48] = buffer_data_6[2535:2528];
        layer1[57][7:0] = buffer_data_5[2487:2480];
        layer1[57][15:8] = buffer_data_5[2495:2488];
        layer1[57][23:16] = buffer_data_5[2503:2496];
        layer1[57][31:24] = buffer_data_5[2511:2504];
        layer1[57][39:32] = buffer_data_5[2519:2512];
        layer1[57][47:40] = buffer_data_5[2527:2520];
        layer1[57][55:48] = buffer_data_5[2535:2528];
        layer2[57][7:0] = buffer_data_4[2487:2480];
        layer2[57][15:8] = buffer_data_4[2495:2488];
        layer2[57][23:16] = buffer_data_4[2503:2496];
        layer2[57][31:24] = buffer_data_4[2511:2504];
        layer2[57][39:32] = buffer_data_4[2519:2512];
        layer2[57][47:40] = buffer_data_4[2527:2520];
        layer2[57][55:48] = buffer_data_4[2535:2528];
        layer3[57][7:0] = buffer_data_3[2487:2480];
        layer3[57][15:8] = buffer_data_3[2495:2488];
        layer3[57][23:16] = buffer_data_3[2503:2496];
        layer3[57][31:24] = buffer_data_3[2511:2504];
        layer3[57][39:32] = buffer_data_3[2519:2512];
        layer3[57][47:40] = buffer_data_3[2527:2520];
        layer3[57][55:48] = buffer_data_3[2535:2528];
        layer4[57][7:0] = buffer_data_2[2487:2480];
        layer4[57][15:8] = buffer_data_2[2495:2488];
        layer4[57][23:16] = buffer_data_2[2503:2496];
        layer4[57][31:24] = buffer_data_2[2511:2504];
        layer4[57][39:32] = buffer_data_2[2519:2512];
        layer4[57][47:40] = buffer_data_2[2527:2520];
        layer4[57][55:48] = buffer_data_2[2535:2528];
        layer5[57][7:0] = buffer_data_1[2487:2480];
        layer5[57][15:8] = buffer_data_1[2495:2488];
        layer5[57][23:16] = buffer_data_1[2503:2496];
        layer5[57][31:24] = buffer_data_1[2511:2504];
        layer5[57][39:32] = buffer_data_1[2519:2512];
        layer5[57][47:40] = buffer_data_1[2527:2520];
        layer5[57][55:48] = buffer_data_1[2535:2528];
        layer6[57][7:0] = buffer_data_0[2487:2480];
        layer6[57][15:8] = buffer_data_0[2495:2488];
        layer6[57][23:16] = buffer_data_0[2503:2496];
        layer6[57][31:24] = buffer_data_0[2511:2504];
        layer6[57][39:32] = buffer_data_0[2519:2512];
        layer6[57][47:40] = buffer_data_0[2527:2520];
        layer6[57][55:48] = buffer_data_0[2535:2528];
        layer0[58][7:0] = buffer_data_6[2495:2488];
        layer0[58][15:8] = buffer_data_6[2503:2496];
        layer0[58][23:16] = buffer_data_6[2511:2504];
        layer0[58][31:24] = buffer_data_6[2519:2512];
        layer0[58][39:32] = buffer_data_6[2527:2520];
        layer0[58][47:40] = buffer_data_6[2535:2528];
        layer0[58][55:48] = buffer_data_6[2543:2536];
        layer1[58][7:0] = buffer_data_5[2495:2488];
        layer1[58][15:8] = buffer_data_5[2503:2496];
        layer1[58][23:16] = buffer_data_5[2511:2504];
        layer1[58][31:24] = buffer_data_5[2519:2512];
        layer1[58][39:32] = buffer_data_5[2527:2520];
        layer1[58][47:40] = buffer_data_5[2535:2528];
        layer1[58][55:48] = buffer_data_5[2543:2536];
        layer2[58][7:0] = buffer_data_4[2495:2488];
        layer2[58][15:8] = buffer_data_4[2503:2496];
        layer2[58][23:16] = buffer_data_4[2511:2504];
        layer2[58][31:24] = buffer_data_4[2519:2512];
        layer2[58][39:32] = buffer_data_4[2527:2520];
        layer2[58][47:40] = buffer_data_4[2535:2528];
        layer2[58][55:48] = buffer_data_4[2543:2536];
        layer3[58][7:0] = buffer_data_3[2495:2488];
        layer3[58][15:8] = buffer_data_3[2503:2496];
        layer3[58][23:16] = buffer_data_3[2511:2504];
        layer3[58][31:24] = buffer_data_3[2519:2512];
        layer3[58][39:32] = buffer_data_3[2527:2520];
        layer3[58][47:40] = buffer_data_3[2535:2528];
        layer3[58][55:48] = buffer_data_3[2543:2536];
        layer4[58][7:0] = buffer_data_2[2495:2488];
        layer4[58][15:8] = buffer_data_2[2503:2496];
        layer4[58][23:16] = buffer_data_2[2511:2504];
        layer4[58][31:24] = buffer_data_2[2519:2512];
        layer4[58][39:32] = buffer_data_2[2527:2520];
        layer4[58][47:40] = buffer_data_2[2535:2528];
        layer4[58][55:48] = buffer_data_2[2543:2536];
        layer5[58][7:0] = buffer_data_1[2495:2488];
        layer5[58][15:8] = buffer_data_1[2503:2496];
        layer5[58][23:16] = buffer_data_1[2511:2504];
        layer5[58][31:24] = buffer_data_1[2519:2512];
        layer5[58][39:32] = buffer_data_1[2527:2520];
        layer5[58][47:40] = buffer_data_1[2535:2528];
        layer5[58][55:48] = buffer_data_1[2543:2536];
        layer6[58][7:0] = buffer_data_0[2495:2488];
        layer6[58][15:8] = buffer_data_0[2503:2496];
        layer6[58][23:16] = buffer_data_0[2511:2504];
        layer6[58][31:24] = buffer_data_0[2519:2512];
        layer6[58][39:32] = buffer_data_0[2527:2520];
        layer6[58][47:40] = buffer_data_0[2535:2528];
        layer6[58][55:48] = buffer_data_0[2543:2536];
        layer0[59][7:0] = buffer_data_6[2503:2496];
        layer0[59][15:8] = buffer_data_6[2511:2504];
        layer0[59][23:16] = buffer_data_6[2519:2512];
        layer0[59][31:24] = buffer_data_6[2527:2520];
        layer0[59][39:32] = buffer_data_6[2535:2528];
        layer0[59][47:40] = buffer_data_6[2543:2536];
        layer0[59][55:48] = buffer_data_6[2551:2544];
        layer1[59][7:0] = buffer_data_5[2503:2496];
        layer1[59][15:8] = buffer_data_5[2511:2504];
        layer1[59][23:16] = buffer_data_5[2519:2512];
        layer1[59][31:24] = buffer_data_5[2527:2520];
        layer1[59][39:32] = buffer_data_5[2535:2528];
        layer1[59][47:40] = buffer_data_5[2543:2536];
        layer1[59][55:48] = buffer_data_5[2551:2544];
        layer2[59][7:0] = buffer_data_4[2503:2496];
        layer2[59][15:8] = buffer_data_4[2511:2504];
        layer2[59][23:16] = buffer_data_4[2519:2512];
        layer2[59][31:24] = buffer_data_4[2527:2520];
        layer2[59][39:32] = buffer_data_4[2535:2528];
        layer2[59][47:40] = buffer_data_4[2543:2536];
        layer2[59][55:48] = buffer_data_4[2551:2544];
        layer3[59][7:0] = buffer_data_3[2503:2496];
        layer3[59][15:8] = buffer_data_3[2511:2504];
        layer3[59][23:16] = buffer_data_3[2519:2512];
        layer3[59][31:24] = buffer_data_3[2527:2520];
        layer3[59][39:32] = buffer_data_3[2535:2528];
        layer3[59][47:40] = buffer_data_3[2543:2536];
        layer3[59][55:48] = buffer_data_3[2551:2544];
        layer4[59][7:0] = buffer_data_2[2503:2496];
        layer4[59][15:8] = buffer_data_2[2511:2504];
        layer4[59][23:16] = buffer_data_2[2519:2512];
        layer4[59][31:24] = buffer_data_2[2527:2520];
        layer4[59][39:32] = buffer_data_2[2535:2528];
        layer4[59][47:40] = buffer_data_2[2543:2536];
        layer4[59][55:48] = buffer_data_2[2551:2544];
        layer5[59][7:0] = buffer_data_1[2503:2496];
        layer5[59][15:8] = buffer_data_1[2511:2504];
        layer5[59][23:16] = buffer_data_1[2519:2512];
        layer5[59][31:24] = buffer_data_1[2527:2520];
        layer5[59][39:32] = buffer_data_1[2535:2528];
        layer5[59][47:40] = buffer_data_1[2543:2536];
        layer5[59][55:48] = buffer_data_1[2551:2544];
        layer6[59][7:0] = buffer_data_0[2503:2496];
        layer6[59][15:8] = buffer_data_0[2511:2504];
        layer6[59][23:16] = buffer_data_0[2519:2512];
        layer6[59][31:24] = buffer_data_0[2527:2520];
        layer6[59][39:32] = buffer_data_0[2535:2528];
        layer6[59][47:40] = buffer_data_0[2543:2536];
        layer6[59][55:48] = buffer_data_0[2551:2544];
        layer0[60][7:0] = buffer_data_6[2511:2504];
        layer0[60][15:8] = buffer_data_6[2519:2512];
        layer0[60][23:16] = buffer_data_6[2527:2520];
        layer0[60][31:24] = buffer_data_6[2535:2528];
        layer0[60][39:32] = buffer_data_6[2543:2536];
        layer0[60][47:40] = buffer_data_6[2551:2544];
        layer0[60][55:48] = buffer_data_6[2559:2552];
        layer1[60][7:0] = buffer_data_5[2511:2504];
        layer1[60][15:8] = buffer_data_5[2519:2512];
        layer1[60][23:16] = buffer_data_5[2527:2520];
        layer1[60][31:24] = buffer_data_5[2535:2528];
        layer1[60][39:32] = buffer_data_5[2543:2536];
        layer1[60][47:40] = buffer_data_5[2551:2544];
        layer1[60][55:48] = buffer_data_5[2559:2552];
        layer2[60][7:0] = buffer_data_4[2511:2504];
        layer2[60][15:8] = buffer_data_4[2519:2512];
        layer2[60][23:16] = buffer_data_4[2527:2520];
        layer2[60][31:24] = buffer_data_4[2535:2528];
        layer2[60][39:32] = buffer_data_4[2543:2536];
        layer2[60][47:40] = buffer_data_4[2551:2544];
        layer2[60][55:48] = buffer_data_4[2559:2552];
        layer3[60][7:0] = buffer_data_3[2511:2504];
        layer3[60][15:8] = buffer_data_3[2519:2512];
        layer3[60][23:16] = buffer_data_3[2527:2520];
        layer3[60][31:24] = buffer_data_3[2535:2528];
        layer3[60][39:32] = buffer_data_3[2543:2536];
        layer3[60][47:40] = buffer_data_3[2551:2544];
        layer3[60][55:48] = buffer_data_3[2559:2552];
        layer4[60][7:0] = buffer_data_2[2511:2504];
        layer4[60][15:8] = buffer_data_2[2519:2512];
        layer4[60][23:16] = buffer_data_2[2527:2520];
        layer4[60][31:24] = buffer_data_2[2535:2528];
        layer4[60][39:32] = buffer_data_2[2543:2536];
        layer4[60][47:40] = buffer_data_2[2551:2544];
        layer4[60][55:48] = buffer_data_2[2559:2552];
        layer5[60][7:0] = buffer_data_1[2511:2504];
        layer5[60][15:8] = buffer_data_1[2519:2512];
        layer5[60][23:16] = buffer_data_1[2527:2520];
        layer5[60][31:24] = buffer_data_1[2535:2528];
        layer5[60][39:32] = buffer_data_1[2543:2536];
        layer5[60][47:40] = buffer_data_1[2551:2544];
        layer5[60][55:48] = buffer_data_1[2559:2552];
        layer6[60][7:0] = buffer_data_0[2511:2504];
        layer6[60][15:8] = buffer_data_0[2519:2512];
        layer6[60][23:16] = buffer_data_0[2527:2520];
        layer6[60][31:24] = buffer_data_0[2535:2528];
        layer6[60][39:32] = buffer_data_0[2543:2536];
        layer6[60][47:40] = buffer_data_0[2551:2544];
        layer6[60][55:48] = buffer_data_0[2559:2552];
        layer0[61][7:0] = buffer_data_6[2519:2512];
        layer0[61][15:8] = buffer_data_6[2527:2520];
        layer0[61][23:16] = buffer_data_6[2535:2528];
        layer0[61][31:24] = buffer_data_6[2543:2536];
        layer0[61][39:32] = buffer_data_6[2551:2544];
        layer0[61][47:40] = buffer_data_6[2559:2552];
        layer0[61][55:48] = buffer_data_6[2567:2560];
        layer1[61][7:0] = buffer_data_5[2519:2512];
        layer1[61][15:8] = buffer_data_5[2527:2520];
        layer1[61][23:16] = buffer_data_5[2535:2528];
        layer1[61][31:24] = buffer_data_5[2543:2536];
        layer1[61][39:32] = buffer_data_5[2551:2544];
        layer1[61][47:40] = buffer_data_5[2559:2552];
        layer1[61][55:48] = buffer_data_5[2567:2560];
        layer2[61][7:0] = buffer_data_4[2519:2512];
        layer2[61][15:8] = buffer_data_4[2527:2520];
        layer2[61][23:16] = buffer_data_4[2535:2528];
        layer2[61][31:24] = buffer_data_4[2543:2536];
        layer2[61][39:32] = buffer_data_4[2551:2544];
        layer2[61][47:40] = buffer_data_4[2559:2552];
        layer2[61][55:48] = buffer_data_4[2567:2560];
        layer3[61][7:0] = buffer_data_3[2519:2512];
        layer3[61][15:8] = buffer_data_3[2527:2520];
        layer3[61][23:16] = buffer_data_3[2535:2528];
        layer3[61][31:24] = buffer_data_3[2543:2536];
        layer3[61][39:32] = buffer_data_3[2551:2544];
        layer3[61][47:40] = buffer_data_3[2559:2552];
        layer3[61][55:48] = buffer_data_3[2567:2560];
        layer4[61][7:0] = buffer_data_2[2519:2512];
        layer4[61][15:8] = buffer_data_2[2527:2520];
        layer4[61][23:16] = buffer_data_2[2535:2528];
        layer4[61][31:24] = buffer_data_2[2543:2536];
        layer4[61][39:32] = buffer_data_2[2551:2544];
        layer4[61][47:40] = buffer_data_2[2559:2552];
        layer4[61][55:48] = buffer_data_2[2567:2560];
        layer5[61][7:0] = buffer_data_1[2519:2512];
        layer5[61][15:8] = buffer_data_1[2527:2520];
        layer5[61][23:16] = buffer_data_1[2535:2528];
        layer5[61][31:24] = buffer_data_1[2543:2536];
        layer5[61][39:32] = buffer_data_1[2551:2544];
        layer5[61][47:40] = buffer_data_1[2559:2552];
        layer5[61][55:48] = buffer_data_1[2567:2560];
        layer6[61][7:0] = buffer_data_0[2519:2512];
        layer6[61][15:8] = buffer_data_0[2527:2520];
        layer6[61][23:16] = buffer_data_0[2535:2528];
        layer6[61][31:24] = buffer_data_0[2543:2536];
        layer6[61][39:32] = buffer_data_0[2551:2544];
        layer6[61][47:40] = buffer_data_0[2559:2552];
        layer6[61][55:48] = buffer_data_0[2567:2560];
        layer0[62][7:0] = buffer_data_6[2527:2520];
        layer0[62][15:8] = buffer_data_6[2535:2528];
        layer0[62][23:16] = buffer_data_6[2543:2536];
        layer0[62][31:24] = buffer_data_6[2551:2544];
        layer0[62][39:32] = buffer_data_6[2559:2552];
        layer0[62][47:40] = buffer_data_6[2567:2560];
        layer0[62][55:48] = buffer_data_6[2575:2568];
        layer1[62][7:0] = buffer_data_5[2527:2520];
        layer1[62][15:8] = buffer_data_5[2535:2528];
        layer1[62][23:16] = buffer_data_5[2543:2536];
        layer1[62][31:24] = buffer_data_5[2551:2544];
        layer1[62][39:32] = buffer_data_5[2559:2552];
        layer1[62][47:40] = buffer_data_5[2567:2560];
        layer1[62][55:48] = buffer_data_5[2575:2568];
        layer2[62][7:0] = buffer_data_4[2527:2520];
        layer2[62][15:8] = buffer_data_4[2535:2528];
        layer2[62][23:16] = buffer_data_4[2543:2536];
        layer2[62][31:24] = buffer_data_4[2551:2544];
        layer2[62][39:32] = buffer_data_4[2559:2552];
        layer2[62][47:40] = buffer_data_4[2567:2560];
        layer2[62][55:48] = buffer_data_4[2575:2568];
        layer3[62][7:0] = buffer_data_3[2527:2520];
        layer3[62][15:8] = buffer_data_3[2535:2528];
        layer3[62][23:16] = buffer_data_3[2543:2536];
        layer3[62][31:24] = buffer_data_3[2551:2544];
        layer3[62][39:32] = buffer_data_3[2559:2552];
        layer3[62][47:40] = buffer_data_3[2567:2560];
        layer3[62][55:48] = buffer_data_3[2575:2568];
        layer4[62][7:0] = buffer_data_2[2527:2520];
        layer4[62][15:8] = buffer_data_2[2535:2528];
        layer4[62][23:16] = buffer_data_2[2543:2536];
        layer4[62][31:24] = buffer_data_2[2551:2544];
        layer4[62][39:32] = buffer_data_2[2559:2552];
        layer4[62][47:40] = buffer_data_2[2567:2560];
        layer4[62][55:48] = buffer_data_2[2575:2568];
        layer5[62][7:0] = buffer_data_1[2527:2520];
        layer5[62][15:8] = buffer_data_1[2535:2528];
        layer5[62][23:16] = buffer_data_1[2543:2536];
        layer5[62][31:24] = buffer_data_1[2551:2544];
        layer5[62][39:32] = buffer_data_1[2559:2552];
        layer5[62][47:40] = buffer_data_1[2567:2560];
        layer5[62][55:48] = buffer_data_1[2575:2568];
        layer6[62][7:0] = buffer_data_0[2527:2520];
        layer6[62][15:8] = buffer_data_0[2535:2528];
        layer6[62][23:16] = buffer_data_0[2543:2536];
        layer6[62][31:24] = buffer_data_0[2551:2544];
        layer6[62][39:32] = buffer_data_0[2559:2552];
        layer6[62][47:40] = buffer_data_0[2567:2560];
        layer6[62][55:48] = buffer_data_0[2575:2568];
        layer0[63][7:0] = buffer_data_6[2535:2528];
        layer0[63][15:8] = buffer_data_6[2543:2536];
        layer0[63][23:16] = buffer_data_6[2551:2544];
        layer0[63][31:24] = buffer_data_6[2559:2552];
        layer0[63][39:32] = buffer_data_6[2567:2560];
        layer0[63][47:40] = buffer_data_6[2575:2568];
        layer0[63][55:48] = buffer_data_6[2583:2576];
        layer1[63][7:0] = buffer_data_5[2535:2528];
        layer1[63][15:8] = buffer_data_5[2543:2536];
        layer1[63][23:16] = buffer_data_5[2551:2544];
        layer1[63][31:24] = buffer_data_5[2559:2552];
        layer1[63][39:32] = buffer_data_5[2567:2560];
        layer1[63][47:40] = buffer_data_5[2575:2568];
        layer1[63][55:48] = buffer_data_5[2583:2576];
        layer2[63][7:0] = buffer_data_4[2535:2528];
        layer2[63][15:8] = buffer_data_4[2543:2536];
        layer2[63][23:16] = buffer_data_4[2551:2544];
        layer2[63][31:24] = buffer_data_4[2559:2552];
        layer2[63][39:32] = buffer_data_4[2567:2560];
        layer2[63][47:40] = buffer_data_4[2575:2568];
        layer2[63][55:48] = buffer_data_4[2583:2576];
        layer3[63][7:0] = buffer_data_3[2535:2528];
        layer3[63][15:8] = buffer_data_3[2543:2536];
        layer3[63][23:16] = buffer_data_3[2551:2544];
        layer3[63][31:24] = buffer_data_3[2559:2552];
        layer3[63][39:32] = buffer_data_3[2567:2560];
        layer3[63][47:40] = buffer_data_3[2575:2568];
        layer3[63][55:48] = buffer_data_3[2583:2576];
        layer4[63][7:0] = buffer_data_2[2535:2528];
        layer4[63][15:8] = buffer_data_2[2543:2536];
        layer4[63][23:16] = buffer_data_2[2551:2544];
        layer4[63][31:24] = buffer_data_2[2559:2552];
        layer4[63][39:32] = buffer_data_2[2567:2560];
        layer4[63][47:40] = buffer_data_2[2575:2568];
        layer4[63][55:48] = buffer_data_2[2583:2576];
        layer5[63][7:0] = buffer_data_1[2535:2528];
        layer5[63][15:8] = buffer_data_1[2543:2536];
        layer5[63][23:16] = buffer_data_1[2551:2544];
        layer5[63][31:24] = buffer_data_1[2559:2552];
        layer5[63][39:32] = buffer_data_1[2567:2560];
        layer5[63][47:40] = buffer_data_1[2575:2568];
        layer5[63][55:48] = buffer_data_1[2583:2576];
        layer6[63][7:0] = buffer_data_0[2535:2528];
        layer6[63][15:8] = buffer_data_0[2543:2536];
        layer6[63][23:16] = buffer_data_0[2551:2544];
        layer6[63][31:24] = buffer_data_0[2559:2552];
        layer6[63][39:32] = buffer_data_0[2567:2560];
        layer6[63][47:40] = buffer_data_0[2575:2568];
        layer6[63][55:48] = buffer_data_0[2583:2576];
    end
    ST_GAUSSIAN_5: begin
        layer0[0][7:0] = buffer_data_6[2543:2536];
        layer0[0][15:8] = buffer_data_6[2551:2544];
        layer0[0][23:16] = buffer_data_6[2559:2552];
        layer0[0][31:24] = buffer_data_6[2567:2560];
        layer0[0][39:32] = buffer_data_6[2575:2568];
        layer0[0][47:40] = buffer_data_6[2583:2576];
        layer0[0][55:48] = buffer_data_6[2591:2584];
        layer1[0][7:0] = buffer_data_5[2543:2536];
        layer1[0][15:8] = buffer_data_5[2551:2544];
        layer1[0][23:16] = buffer_data_5[2559:2552];
        layer1[0][31:24] = buffer_data_5[2567:2560];
        layer1[0][39:32] = buffer_data_5[2575:2568];
        layer1[0][47:40] = buffer_data_5[2583:2576];
        layer1[0][55:48] = buffer_data_5[2591:2584];
        layer2[0][7:0] = buffer_data_4[2543:2536];
        layer2[0][15:8] = buffer_data_4[2551:2544];
        layer2[0][23:16] = buffer_data_4[2559:2552];
        layer2[0][31:24] = buffer_data_4[2567:2560];
        layer2[0][39:32] = buffer_data_4[2575:2568];
        layer2[0][47:40] = buffer_data_4[2583:2576];
        layer2[0][55:48] = buffer_data_4[2591:2584];
        layer3[0][7:0] = buffer_data_3[2543:2536];
        layer3[0][15:8] = buffer_data_3[2551:2544];
        layer3[0][23:16] = buffer_data_3[2559:2552];
        layer3[0][31:24] = buffer_data_3[2567:2560];
        layer3[0][39:32] = buffer_data_3[2575:2568];
        layer3[0][47:40] = buffer_data_3[2583:2576];
        layer3[0][55:48] = buffer_data_3[2591:2584];
        layer4[0][7:0] = buffer_data_2[2543:2536];
        layer4[0][15:8] = buffer_data_2[2551:2544];
        layer4[0][23:16] = buffer_data_2[2559:2552];
        layer4[0][31:24] = buffer_data_2[2567:2560];
        layer4[0][39:32] = buffer_data_2[2575:2568];
        layer4[0][47:40] = buffer_data_2[2583:2576];
        layer4[0][55:48] = buffer_data_2[2591:2584];
        layer5[0][7:0] = buffer_data_1[2543:2536];
        layer5[0][15:8] = buffer_data_1[2551:2544];
        layer5[0][23:16] = buffer_data_1[2559:2552];
        layer5[0][31:24] = buffer_data_1[2567:2560];
        layer5[0][39:32] = buffer_data_1[2575:2568];
        layer5[0][47:40] = buffer_data_1[2583:2576];
        layer5[0][55:48] = buffer_data_1[2591:2584];
        layer6[0][7:0] = buffer_data_0[2543:2536];
        layer6[0][15:8] = buffer_data_0[2551:2544];
        layer6[0][23:16] = buffer_data_0[2559:2552];
        layer6[0][31:24] = buffer_data_0[2567:2560];
        layer6[0][39:32] = buffer_data_0[2575:2568];
        layer6[0][47:40] = buffer_data_0[2583:2576];
        layer6[0][55:48] = buffer_data_0[2591:2584];
        layer0[1][7:0] = buffer_data_6[2551:2544];
        layer0[1][15:8] = buffer_data_6[2559:2552];
        layer0[1][23:16] = buffer_data_6[2567:2560];
        layer0[1][31:24] = buffer_data_6[2575:2568];
        layer0[1][39:32] = buffer_data_6[2583:2576];
        layer0[1][47:40] = buffer_data_6[2591:2584];
        layer0[1][55:48] = buffer_data_6[2599:2592];
        layer1[1][7:0] = buffer_data_5[2551:2544];
        layer1[1][15:8] = buffer_data_5[2559:2552];
        layer1[1][23:16] = buffer_data_5[2567:2560];
        layer1[1][31:24] = buffer_data_5[2575:2568];
        layer1[1][39:32] = buffer_data_5[2583:2576];
        layer1[1][47:40] = buffer_data_5[2591:2584];
        layer1[1][55:48] = buffer_data_5[2599:2592];
        layer2[1][7:0] = buffer_data_4[2551:2544];
        layer2[1][15:8] = buffer_data_4[2559:2552];
        layer2[1][23:16] = buffer_data_4[2567:2560];
        layer2[1][31:24] = buffer_data_4[2575:2568];
        layer2[1][39:32] = buffer_data_4[2583:2576];
        layer2[1][47:40] = buffer_data_4[2591:2584];
        layer2[1][55:48] = buffer_data_4[2599:2592];
        layer3[1][7:0] = buffer_data_3[2551:2544];
        layer3[1][15:8] = buffer_data_3[2559:2552];
        layer3[1][23:16] = buffer_data_3[2567:2560];
        layer3[1][31:24] = buffer_data_3[2575:2568];
        layer3[1][39:32] = buffer_data_3[2583:2576];
        layer3[1][47:40] = buffer_data_3[2591:2584];
        layer3[1][55:48] = buffer_data_3[2599:2592];
        layer4[1][7:0] = buffer_data_2[2551:2544];
        layer4[1][15:8] = buffer_data_2[2559:2552];
        layer4[1][23:16] = buffer_data_2[2567:2560];
        layer4[1][31:24] = buffer_data_2[2575:2568];
        layer4[1][39:32] = buffer_data_2[2583:2576];
        layer4[1][47:40] = buffer_data_2[2591:2584];
        layer4[1][55:48] = buffer_data_2[2599:2592];
        layer5[1][7:0] = buffer_data_1[2551:2544];
        layer5[1][15:8] = buffer_data_1[2559:2552];
        layer5[1][23:16] = buffer_data_1[2567:2560];
        layer5[1][31:24] = buffer_data_1[2575:2568];
        layer5[1][39:32] = buffer_data_1[2583:2576];
        layer5[1][47:40] = buffer_data_1[2591:2584];
        layer5[1][55:48] = buffer_data_1[2599:2592];
        layer6[1][7:0] = buffer_data_0[2551:2544];
        layer6[1][15:8] = buffer_data_0[2559:2552];
        layer6[1][23:16] = buffer_data_0[2567:2560];
        layer6[1][31:24] = buffer_data_0[2575:2568];
        layer6[1][39:32] = buffer_data_0[2583:2576];
        layer6[1][47:40] = buffer_data_0[2591:2584];
        layer6[1][55:48] = buffer_data_0[2599:2592];
        layer0[2][7:0] = buffer_data_6[2559:2552];
        layer0[2][15:8] = buffer_data_6[2567:2560];
        layer0[2][23:16] = buffer_data_6[2575:2568];
        layer0[2][31:24] = buffer_data_6[2583:2576];
        layer0[2][39:32] = buffer_data_6[2591:2584];
        layer0[2][47:40] = buffer_data_6[2599:2592];
        layer0[2][55:48] = buffer_data_6[2607:2600];
        layer1[2][7:0] = buffer_data_5[2559:2552];
        layer1[2][15:8] = buffer_data_5[2567:2560];
        layer1[2][23:16] = buffer_data_5[2575:2568];
        layer1[2][31:24] = buffer_data_5[2583:2576];
        layer1[2][39:32] = buffer_data_5[2591:2584];
        layer1[2][47:40] = buffer_data_5[2599:2592];
        layer1[2][55:48] = buffer_data_5[2607:2600];
        layer2[2][7:0] = buffer_data_4[2559:2552];
        layer2[2][15:8] = buffer_data_4[2567:2560];
        layer2[2][23:16] = buffer_data_4[2575:2568];
        layer2[2][31:24] = buffer_data_4[2583:2576];
        layer2[2][39:32] = buffer_data_4[2591:2584];
        layer2[2][47:40] = buffer_data_4[2599:2592];
        layer2[2][55:48] = buffer_data_4[2607:2600];
        layer3[2][7:0] = buffer_data_3[2559:2552];
        layer3[2][15:8] = buffer_data_3[2567:2560];
        layer3[2][23:16] = buffer_data_3[2575:2568];
        layer3[2][31:24] = buffer_data_3[2583:2576];
        layer3[2][39:32] = buffer_data_3[2591:2584];
        layer3[2][47:40] = buffer_data_3[2599:2592];
        layer3[2][55:48] = buffer_data_3[2607:2600];
        layer4[2][7:0] = buffer_data_2[2559:2552];
        layer4[2][15:8] = buffer_data_2[2567:2560];
        layer4[2][23:16] = buffer_data_2[2575:2568];
        layer4[2][31:24] = buffer_data_2[2583:2576];
        layer4[2][39:32] = buffer_data_2[2591:2584];
        layer4[2][47:40] = buffer_data_2[2599:2592];
        layer4[2][55:48] = buffer_data_2[2607:2600];
        layer5[2][7:0] = buffer_data_1[2559:2552];
        layer5[2][15:8] = buffer_data_1[2567:2560];
        layer5[2][23:16] = buffer_data_1[2575:2568];
        layer5[2][31:24] = buffer_data_1[2583:2576];
        layer5[2][39:32] = buffer_data_1[2591:2584];
        layer5[2][47:40] = buffer_data_1[2599:2592];
        layer5[2][55:48] = buffer_data_1[2607:2600];
        layer6[2][7:0] = buffer_data_0[2559:2552];
        layer6[2][15:8] = buffer_data_0[2567:2560];
        layer6[2][23:16] = buffer_data_0[2575:2568];
        layer6[2][31:24] = buffer_data_0[2583:2576];
        layer6[2][39:32] = buffer_data_0[2591:2584];
        layer6[2][47:40] = buffer_data_0[2599:2592];
        layer6[2][55:48] = buffer_data_0[2607:2600];
        layer0[3][7:0] = buffer_data_6[2567:2560];
        layer0[3][15:8] = buffer_data_6[2575:2568];
        layer0[3][23:16] = buffer_data_6[2583:2576];
        layer0[3][31:24] = buffer_data_6[2591:2584];
        layer0[3][39:32] = buffer_data_6[2599:2592];
        layer0[3][47:40] = buffer_data_6[2607:2600];
        layer0[3][55:48] = buffer_data_6[2615:2608];
        layer1[3][7:0] = buffer_data_5[2567:2560];
        layer1[3][15:8] = buffer_data_5[2575:2568];
        layer1[3][23:16] = buffer_data_5[2583:2576];
        layer1[3][31:24] = buffer_data_5[2591:2584];
        layer1[3][39:32] = buffer_data_5[2599:2592];
        layer1[3][47:40] = buffer_data_5[2607:2600];
        layer1[3][55:48] = buffer_data_5[2615:2608];
        layer2[3][7:0] = buffer_data_4[2567:2560];
        layer2[3][15:8] = buffer_data_4[2575:2568];
        layer2[3][23:16] = buffer_data_4[2583:2576];
        layer2[3][31:24] = buffer_data_4[2591:2584];
        layer2[3][39:32] = buffer_data_4[2599:2592];
        layer2[3][47:40] = buffer_data_4[2607:2600];
        layer2[3][55:48] = buffer_data_4[2615:2608];
        layer3[3][7:0] = buffer_data_3[2567:2560];
        layer3[3][15:8] = buffer_data_3[2575:2568];
        layer3[3][23:16] = buffer_data_3[2583:2576];
        layer3[3][31:24] = buffer_data_3[2591:2584];
        layer3[3][39:32] = buffer_data_3[2599:2592];
        layer3[3][47:40] = buffer_data_3[2607:2600];
        layer3[3][55:48] = buffer_data_3[2615:2608];
        layer4[3][7:0] = buffer_data_2[2567:2560];
        layer4[3][15:8] = buffer_data_2[2575:2568];
        layer4[3][23:16] = buffer_data_2[2583:2576];
        layer4[3][31:24] = buffer_data_2[2591:2584];
        layer4[3][39:32] = buffer_data_2[2599:2592];
        layer4[3][47:40] = buffer_data_2[2607:2600];
        layer4[3][55:48] = buffer_data_2[2615:2608];
        layer5[3][7:0] = buffer_data_1[2567:2560];
        layer5[3][15:8] = buffer_data_1[2575:2568];
        layer5[3][23:16] = buffer_data_1[2583:2576];
        layer5[3][31:24] = buffer_data_1[2591:2584];
        layer5[3][39:32] = buffer_data_1[2599:2592];
        layer5[3][47:40] = buffer_data_1[2607:2600];
        layer5[3][55:48] = buffer_data_1[2615:2608];
        layer6[3][7:0] = buffer_data_0[2567:2560];
        layer6[3][15:8] = buffer_data_0[2575:2568];
        layer6[3][23:16] = buffer_data_0[2583:2576];
        layer6[3][31:24] = buffer_data_0[2591:2584];
        layer6[3][39:32] = buffer_data_0[2599:2592];
        layer6[3][47:40] = buffer_data_0[2607:2600];
        layer6[3][55:48] = buffer_data_0[2615:2608];
        layer0[4][7:0] = buffer_data_6[2575:2568];
        layer0[4][15:8] = buffer_data_6[2583:2576];
        layer0[4][23:16] = buffer_data_6[2591:2584];
        layer0[4][31:24] = buffer_data_6[2599:2592];
        layer0[4][39:32] = buffer_data_6[2607:2600];
        layer0[4][47:40] = buffer_data_6[2615:2608];
        layer0[4][55:48] = buffer_data_6[2623:2616];
        layer1[4][7:0] = buffer_data_5[2575:2568];
        layer1[4][15:8] = buffer_data_5[2583:2576];
        layer1[4][23:16] = buffer_data_5[2591:2584];
        layer1[4][31:24] = buffer_data_5[2599:2592];
        layer1[4][39:32] = buffer_data_5[2607:2600];
        layer1[4][47:40] = buffer_data_5[2615:2608];
        layer1[4][55:48] = buffer_data_5[2623:2616];
        layer2[4][7:0] = buffer_data_4[2575:2568];
        layer2[4][15:8] = buffer_data_4[2583:2576];
        layer2[4][23:16] = buffer_data_4[2591:2584];
        layer2[4][31:24] = buffer_data_4[2599:2592];
        layer2[4][39:32] = buffer_data_4[2607:2600];
        layer2[4][47:40] = buffer_data_4[2615:2608];
        layer2[4][55:48] = buffer_data_4[2623:2616];
        layer3[4][7:0] = buffer_data_3[2575:2568];
        layer3[4][15:8] = buffer_data_3[2583:2576];
        layer3[4][23:16] = buffer_data_3[2591:2584];
        layer3[4][31:24] = buffer_data_3[2599:2592];
        layer3[4][39:32] = buffer_data_3[2607:2600];
        layer3[4][47:40] = buffer_data_3[2615:2608];
        layer3[4][55:48] = buffer_data_3[2623:2616];
        layer4[4][7:0] = buffer_data_2[2575:2568];
        layer4[4][15:8] = buffer_data_2[2583:2576];
        layer4[4][23:16] = buffer_data_2[2591:2584];
        layer4[4][31:24] = buffer_data_2[2599:2592];
        layer4[4][39:32] = buffer_data_2[2607:2600];
        layer4[4][47:40] = buffer_data_2[2615:2608];
        layer4[4][55:48] = buffer_data_2[2623:2616];
        layer5[4][7:0] = buffer_data_1[2575:2568];
        layer5[4][15:8] = buffer_data_1[2583:2576];
        layer5[4][23:16] = buffer_data_1[2591:2584];
        layer5[4][31:24] = buffer_data_1[2599:2592];
        layer5[4][39:32] = buffer_data_1[2607:2600];
        layer5[4][47:40] = buffer_data_1[2615:2608];
        layer5[4][55:48] = buffer_data_1[2623:2616];
        layer6[4][7:0] = buffer_data_0[2575:2568];
        layer6[4][15:8] = buffer_data_0[2583:2576];
        layer6[4][23:16] = buffer_data_0[2591:2584];
        layer6[4][31:24] = buffer_data_0[2599:2592];
        layer6[4][39:32] = buffer_data_0[2607:2600];
        layer6[4][47:40] = buffer_data_0[2615:2608];
        layer6[4][55:48] = buffer_data_0[2623:2616];
        layer0[5][7:0] = buffer_data_6[2583:2576];
        layer0[5][15:8] = buffer_data_6[2591:2584];
        layer0[5][23:16] = buffer_data_6[2599:2592];
        layer0[5][31:24] = buffer_data_6[2607:2600];
        layer0[5][39:32] = buffer_data_6[2615:2608];
        layer0[5][47:40] = buffer_data_6[2623:2616];
        layer0[5][55:48] = buffer_data_6[2631:2624];
        layer1[5][7:0] = buffer_data_5[2583:2576];
        layer1[5][15:8] = buffer_data_5[2591:2584];
        layer1[5][23:16] = buffer_data_5[2599:2592];
        layer1[5][31:24] = buffer_data_5[2607:2600];
        layer1[5][39:32] = buffer_data_5[2615:2608];
        layer1[5][47:40] = buffer_data_5[2623:2616];
        layer1[5][55:48] = buffer_data_5[2631:2624];
        layer2[5][7:0] = buffer_data_4[2583:2576];
        layer2[5][15:8] = buffer_data_4[2591:2584];
        layer2[5][23:16] = buffer_data_4[2599:2592];
        layer2[5][31:24] = buffer_data_4[2607:2600];
        layer2[5][39:32] = buffer_data_4[2615:2608];
        layer2[5][47:40] = buffer_data_4[2623:2616];
        layer2[5][55:48] = buffer_data_4[2631:2624];
        layer3[5][7:0] = buffer_data_3[2583:2576];
        layer3[5][15:8] = buffer_data_3[2591:2584];
        layer3[5][23:16] = buffer_data_3[2599:2592];
        layer3[5][31:24] = buffer_data_3[2607:2600];
        layer3[5][39:32] = buffer_data_3[2615:2608];
        layer3[5][47:40] = buffer_data_3[2623:2616];
        layer3[5][55:48] = buffer_data_3[2631:2624];
        layer4[5][7:0] = buffer_data_2[2583:2576];
        layer4[5][15:8] = buffer_data_2[2591:2584];
        layer4[5][23:16] = buffer_data_2[2599:2592];
        layer4[5][31:24] = buffer_data_2[2607:2600];
        layer4[5][39:32] = buffer_data_2[2615:2608];
        layer4[5][47:40] = buffer_data_2[2623:2616];
        layer4[5][55:48] = buffer_data_2[2631:2624];
        layer5[5][7:0] = buffer_data_1[2583:2576];
        layer5[5][15:8] = buffer_data_1[2591:2584];
        layer5[5][23:16] = buffer_data_1[2599:2592];
        layer5[5][31:24] = buffer_data_1[2607:2600];
        layer5[5][39:32] = buffer_data_1[2615:2608];
        layer5[5][47:40] = buffer_data_1[2623:2616];
        layer5[5][55:48] = buffer_data_1[2631:2624];
        layer6[5][7:0] = buffer_data_0[2583:2576];
        layer6[5][15:8] = buffer_data_0[2591:2584];
        layer6[5][23:16] = buffer_data_0[2599:2592];
        layer6[5][31:24] = buffer_data_0[2607:2600];
        layer6[5][39:32] = buffer_data_0[2615:2608];
        layer6[5][47:40] = buffer_data_0[2623:2616];
        layer6[5][55:48] = buffer_data_0[2631:2624];
        layer0[6][7:0] = buffer_data_6[2591:2584];
        layer0[6][15:8] = buffer_data_6[2599:2592];
        layer0[6][23:16] = buffer_data_6[2607:2600];
        layer0[6][31:24] = buffer_data_6[2615:2608];
        layer0[6][39:32] = buffer_data_6[2623:2616];
        layer0[6][47:40] = buffer_data_6[2631:2624];
        layer0[6][55:48] = buffer_data_6[2639:2632];
        layer1[6][7:0] = buffer_data_5[2591:2584];
        layer1[6][15:8] = buffer_data_5[2599:2592];
        layer1[6][23:16] = buffer_data_5[2607:2600];
        layer1[6][31:24] = buffer_data_5[2615:2608];
        layer1[6][39:32] = buffer_data_5[2623:2616];
        layer1[6][47:40] = buffer_data_5[2631:2624];
        layer1[6][55:48] = buffer_data_5[2639:2632];
        layer2[6][7:0] = buffer_data_4[2591:2584];
        layer2[6][15:8] = buffer_data_4[2599:2592];
        layer2[6][23:16] = buffer_data_4[2607:2600];
        layer2[6][31:24] = buffer_data_4[2615:2608];
        layer2[6][39:32] = buffer_data_4[2623:2616];
        layer2[6][47:40] = buffer_data_4[2631:2624];
        layer2[6][55:48] = buffer_data_4[2639:2632];
        layer3[6][7:0] = buffer_data_3[2591:2584];
        layer3[6][15:8] = buffer_data_3[2599:2592];
        layer3[6][23:16] = buffer_data_3[2607:2600];
        layer3[6][31:24] = buffer_data_3[2615:2608];
        layer3[6][39:32] = buffer_data_3[2623:2616];
        layer3[6][47:40] = buffer_data_3[2631:2624];
        layer3[6][55:48] = buffer_data_3[2639:2632];
        layer4[6][7:0] = buffer_data_2[2591:2584];
        layer4[6][15:8] = buffer_data_2[2599:2592];
        layer4[6][23:16] = buffer_data_2[2607:2600];
        layer4[6][31:24] = buffer_data_2[2615:2608];
        layer4[6][39:32] = buffer_data_2[2623:2616];
        layer4[6][47:40] = buffer_data_2[2631:2624];
        layer4[6][55:48] = buffer_data_2[2639:2632];
        layer5[6][7:0] = buffer_data_1[2591:2584];
        layer5[6][15:8] = buffer_data_1[2599:2592];
        layer5[6][23:16] = buffer_data_1[2607:2600];
        layer5[6][31:24] = buffer_data_1[2615:2608];
        layer5[6][39:32] = buffer_data_1[2623:2616];
        layer5[6][47:40] = buffer_data_1[2631:2624];
        layer5[6][55:48] = buffer_data_1[2639:2632];
        layer6[6][7:0] = buffer_data_0[2591:2584];
        layer6[6][15:8] = buffer_data_0[2599:2592];
        layer6[6][23:16] = buffer_data_0[2607:2600];
        layer6[6][31:24] = buffer_data_0[2615:2608];
        layer6[6][39:32] = buffer_data_0[2623:2616];
        layer6[6][47:40] = buffer_data_0[2631:2624];
        layer6[6][55:48] = buffer_data_0[2639:2632];
        layer0[7][7:0] = buffer_data_6[2599:2592];
        layer0[7][15:8] = buffer_data_6[2607:2600];
        layer0[7][23:16] = buffer_data_6[2615:2608];
        layer0[7][31:24] = buffer_data_6[2623:2616];
        layer0[7][39:32] = buffer_data_6[2631:2624];
        layer0[7][47:40] = buffer_data_6[2639:2632];
        layer0[7][55:48] = buffer_data_6[2647:2640];
        layer1[7][7:0] = buffer_data_5[2599:2592];
        layer1[7][15:8] = buffer_data_5[2607:2600];
        layer1[7][23:16] = buffer_data_5[2615:2608];
        layer1[7][31:24] = buffer_data_5[2623:2616];
        layer1[7][39:32] = buffer_data_5[2631:2624];
        layer1[7][47:40] = buffer_data_5[2639:2632];
        layer1[7][55:48] = buffer_data_5[2647:2640];
        layer2[7][7:0] = buffer_data_4[2599:2592];
        layer2[7][15:8] = buffer_data_4[2607:2600];
        layer2[7][23:16] = buffer_data_4[2615:2608];
        layer2[7][31:24] = buffer_data_4[2623:2616];
        layer2[7][39:32] = buffer_data_4[2631:2624];
        layer2[7][47:40] = buffer_data_4[2639:2632];
        layer2[7][55:48] = buffer_data_4[2647:2640];
        layer3[7][7:0] = buffer_data_3[2599:2592];
        layer3[7][15:8] = buffer_data_3[2607:2600];
        layer3[7][23:16] = buffer_data_3[2615:2608];
        layer3[7][31:24] = buffer_data_3[2623:2616];
        layer3[7][39:32] = buffer_data_3[2631:2624];
        layer3[7][47:40] = buffer_data_3[2639:2632];
        layer3[7][55:48] = buffer_data_3[2647:2640];
        layer4[7][7:0] = buffer_data_2[2599:2592];
        layer4[7][15:8] = buffer_data_2[2607:2600];
        layer4[7][23:16] = buffer_data_2[2615:2608];
        layer4[7][31:24] = buffer_data_2[2623:2616];
        layer4[7][39:32] = buffer_data_2[2631:2624];
        layer4[7][47:40] = buffer_data_2[2639:2632];
        layer4[7][55:48] = buffer_data_2[2647:2640];
        layer5[7][7:0] = buffer_data_1[2599:2592];
        layer5[7][15:8] = buffer_data_1[2607:2600];
        layer5[7][23:16] = buffer_data_1[2615:2608];
        layer5[7][31:24] = buffer_data_1[2623:2616];
        layer5[7][39:32] = buffer_data_1[2631:2624];
        layer5[7][47:40] = buffer_data_1[2639:2632];
        layer5[7][55:48] = buffer_data_1[2647:2640];
        layer6[7][7:0] = buffer_data_0[2599:2592];
        layer6[7][15:8] = buffer_data_0[2607:2600];
        layer6[7][23:16] = buffer_data_0[2615:2608];
        layer6[7][31:24] = buffer_data_0[2623:2616];
        layer6[7][39:32] = buffer_data_0[2631:2624];
        layer6[7][47:40] = buffer_data_0[2639:2632];
        layer6[7][55:48] = buffer_data_0[2647:2640];
        layer0[8][7:0] = buffer_data_6[2607:2600];
        layer0[8][15:8] = buffer_data_6[2615:2608];
        layer0[8][23:16] = buffer_data_6[2623:2616];
        layer0[8][31:24] = buffer_data_6[2631:2624];
        layer0[8][39:32] = buffer_data_6[2639:2632];
        layer0[8][47:40] = buffer_data_6[2647:2640];
        layer0[8][55:48] = buffer_data_6[2655:2648];
        layer1[8][7:0] = buffer_data_5[2607:2600];
        layer1[8][15:8] = buffer_data_5[2615:2608];
        layer1[8][23:16] = buffer_data_5[2623:2616];
        layer1[8][31:24] = buffer_data_5[2631:2624];
        layer1[8][39:32] = buffer_data_5[2639:2632];
        layer1[8][47:40] = buffer_data_5[2647:2640];
        layer1[8][55:48] = buffer_data_5[2655:2648];
        layer2[8][7:0] = buffer_data_4[2607:2600];
        layer2[8][15:8] = buffer_data_4[2615:2608];
        layer2[8][23:16] = buffer_data_4[2623:2616];
        layer2[8][31:24] = buffer_data_4[2631:2624];
        layer2[8][39:32] = buffer_data_4[2639:2632];
        layer2[8][47:40] = buffer_data_4[2647:2640];
        layer2[8][55:48] = buffer_data_4[2655:2648];
        layer3[8][7:0] = buffer_data_3[2607:2600];
        layer3[8][15:8] = buffer_data_3[2615:2608];
        layer3[8][23:16] = buffer_data_3[2623:2616];
        layer3[8][31:24] = buffer_data_3[2631:2624];
        layer3[8][39:32] = buffer_data_3[2639:2632];
        layer3[8][47:40] = buffer_data_3[2647:2640];
        layer3[8][55:48] = buffer_data_3[2655:2648];
        layer4[8][7:0] = buffer_data_2[2607:2600];
        layer4[8][15:8] = buffer_data_2[2615:2608];
        layer4[8][23:16] = buffer_data_2[2623:2616];
        layer4[8][31:24] = buffer_data_2[2631:2624];
        layer4[8][39:32] = buffer_data_2[2639:2632];
        layer4[8][47:40] = buffer_data_2[2647:2640];
        layer4[8][55:48] = buffer_data_2[2655:2648];
        layer5[8][7:0] = buffer_data_1[2607:2600];
        layer5[8][15:8] = buffer_data_1[2615:2608];
        layer5[8][23:16] = buffer_data_1[2623:2616];
        layer5[8][31:24] = buffer_data_1[2631:2624];
        layer5[8][39:32] = buffer_data_1[2639:2632];
        layer5[8][47:40] = buffer_data_1[2647:2640];
        layer5[8][55:48] = buffer_data_1[2655:2648];
        layer6[8][7:0] = buffer_data_0[2607:2600];
        layer6[8][15:8] = buffer_data_0[2615:2608];
        layer6[8][23:16] = buffer_data_0[2623:2616];
        layer6[8][31:24] = buffer_data_0[2631:2624];
        layer6[8][39:32] = buffer_data_0[2639:2632];
        layer6[8][47:40] = buffer_data_0[2647:2640];
        layer6[8][55:48] = buffer_data_0[2655:2648];
        layer0[9][7:0] = buffer_data_6[2615:2608];
        layer0[9][15:8] = buffer_data_6[2623:2616];
        layer0[9][23:16] = buffer_data_6[2631:2624];
        layer0[9][31:24] = buffer_data_6[2639:2632];
        layer0[9][39:32] = buffer_data_6[2647:2640];
        layer0[9][47:40] = buffer_data_6[2655:2648];
        layer0[9][55:48] = buffer_data_6[2663:2656];
        layer1[9][7:0] = buffer_data_5[2615:2608];
        layer1[9][15:8] = buffer_data_5[2623:2616];
        layer1[9][23:16] = buffer_data_5[2631:2624];
        layer1[9][31:24] = buffer_data_5[2639:2632];
        layer1[9][39:32] = buffer_data_5[2647:2640];
        layer1[9][47:40] = buffer_data_5[2655:2648];
        layer1[9][55:48] = buffer_data_5[2663:2656];
        layer2[9][7:0] = buffer_data_4[2615:2608];
        layer2[9][15:8] = buffer_data_4[2623:2616];
        layer2[9][23:16] = buffer_data_4[2631:2624];
        layer2[9][31:24] = buffer_data_4[2639:2632];
        layer2[9][39:32] = buffer_data_4[2647:2640];
        layer2[9][47:40] = buffer_data_4[2655:2648];
        layer2[9][55:48] = buffer_data_4[2663:2656];
        layer3[9][7:0] = buffer_data_3[2615:2608];
        layer3[9][15:8] = buffer_data_3[2623:2616];
        layer3[9][23:16] = buffer_data_3[2631:2624];
        layer3[9][31:24] = buffer_data_3[2639:2632];
        layer3[9][39:32] = buffer_data_3[2647:2640];
        layer3[9][47:40] = buffer_data_3[2655:2648];
        layer3[9][55:48] = buffer_data_3[2663:2656];
        layer4[9][7:0] = buffer_data_2[2615:2608];
        layer4[9][15:8] = buffer_data_2[2623:2616];
        layer4[9][23:16] = buffer_data_2[2631:2624];
        layer4[9][31:24] = buffer_data_2[2639:2632];
        layer4[9][39:32] = buffer_data_2[2647:2640];
        layer4[9][47:40] = buffer_data_2[2655:2648];
        layer4[9][55:48] = buffer_data_2[2663:2656];
        layer5[9][7:0] = buffer_data_1[2615:2608];
        layer5[9][15:8] = buffer_data_1[2623:2616];
        layer5[9][23:16] = buffer_data_1[2631:2624];
        layer5[9][31:24] = buffer_data_1[2639:2632];
        layer5[9][39:32] = buffer_data_1[2647:2640];
        layer5[9][47:40] = buffer_data_1[2655:2648];
        layer5[9][55:48] = buffer_data_1[2663:2656];
        layer6[9][7:0] = buffer_data_0[2615:2608];
        layer6[9][15:8] = buffer_data_0[2623:2616];
        layer6[9][23:16] = buffer_data_0[2631:2624];
        layer6[9][31:24] = buffer_data_0[2639:2632];
        layer6[9][39:32] = buffer_data_0[2647:2640];
        layer6[9][47:40] = buffer_data_0[2655:2648];
        layer6[9][55:48] = buffer_data_0[2663:2656];
        layer0[10][7:0] = buffer_data_6[2623:2616];
        layer0[10][15:8] = buffer_data_6[2631:2624];
        layer0[10][23:16] = buffer_data_6[2639:2632];
        layer0[10][31:24] = buffer_data_6[2647:2640];
        layer0[10][39:32] = buffer_data_6[2655:2648];
        layer0[10][47:40] = buffer_data_6[2663:2656];
        layer0[10][55:48] = buffer_data_6[2671:2664];
        layer1[10][7:0] = buffer_data_5[2623:2616];
        layer1[10][15:8] = buffer_data_5[2631:2624];
        layer1[10][23:16] = buffer_data_5[2639:2632];
        layer1[10][31:24] = buffer_data_5[2647:2640];
        layer1[10][39:32] = buffer_data_5[2655:2648];
        layer1[10][47:40] = buffer_data_5[2663:2656];
        layer1[10][55:48] = buffer_data_5[2671:2664];
        layer2[10][7:0] = buffer_data_4[2623:2616];
        layer2[10][15:8] = buffer_data_4[2631:2624];
        layer2[10][23:16] = buffer_data_4[2639:2632];
        layer2[10][31:24] = buffer_data_4[2647:2640];
        layer2[10][39:32] = buffer_data_4[2655:2648];
        layer2[10][47:40] = buffer_data_4[2663:2656];
        layer2[10][55:48] = buffer_data_4[2671:2664];
        layer3[10][7:0] = buffer_data_3[2623:2616];
        layer3[10][15:8] = buffer_data_3[2631:2624];
        layer3[10][23:16] = buffer_data_3[2639:2632];
        layer3[10][31:24] = buffer_data_3[2647:2640];
        layer3[10][39:32] = buffer_data_3[2655:2648];
        layer3[10][47:40] = buffer_data_3[2663:2656];
        layer3[10][55:48] = buffer_data_3[2671:2664];
        layer4[10][7:0] = buffer_data_2[2623:2616];
        layer4[10][15:8] = buffer_data_2[2631:2624];
        layer4[10][23:16] = buffer_data_2[2639:2632];
        layer4[10][31:24] = buffer_data_2[2647:2640];
        layer4[10][39:32] = buffer_data_2[2655:2648];
        layer4[10][47:40] = buffer_data_2[2663:2656];
        layer4[10][55:48] = buffer_data_2[2671:2664];
        layer5[10][7:0] = buffer_data_1[2623:2616];
        layer5[10][15:8] = buffer_data_1[2631:2624];
        layer5[10][23:16] = buffer_data_1[2639:2632];
        layer5[10][31:24] = buffer_data_1[2647:2640];
        layer5[10][39:32] = buffer_data_1[2655:2648];
        layer5[10][47:40] = buffer_data_1[2663:2656];
        layer5[10][55:48] = buffer_data_1[2671:2664];
        layer6[10][7:0] = buffer_data_0[2623:2616];
        layer6[10][15:8] = buffer_data_0[2631:2624];
        layer6[10][23:16] = buffer_data_0[2639:2632];
        layer6[10][31:24] = buffer_data_0[2647:2640];
        layer6[10][39:32] = buffer_data_0[2655:2648];
        layer6[10][47:40] = buffer_data_0[2663:2656];
        layer6[10][55:48] = buffer_data_0[2671:2664];
        layer0[11][7:0] = buffer_data_6[2631:2624];
        layer0[11][15:8] = buffer_data_6[2639:2632];
        layer0[11][23:16] = buffer_data_6[2647:2640];
        layer0[11][31:24] = buffer_data_6[2655:2648];
        layer0[11][39:32] = buffer_data_6[2663:2656];
        layer0[11][47:40] = buffer_data_6[2671:2664];
        layer0[11][55:48] = buffer_data_6[2679:2672];
        layer1[11][7:0] = buffer_data_5[2631:2624];
        layer1[11][15:8] = buffer_data_5[2639:2632];
        layer1[11][23:16] = buffer_data_5[2647:2640];
        layer1[11][31:24] = buffer_data_5[2655:2648];
        layer1[11][39:32] = buffer_data_5[2663:2656];
        layer1[11][47:40] = buffer_data_5[2671:2664];
        layer1[11][55:48] = buffer_data_5[2679:2672];
        layer2[11][7:0] = buffer_data_4[2631:2624];
        layer2[11][15:8] = buffer_data_4[2639:2632];
        layer2[11][23:16] = buffer_data_4[2647:2640];
        layer2[11][31:24] = buffer_data_4[2655:2648];
        layer2[11][39:32] = buffer_data_4[2663:2656];
        layer2[11][47:40] = buffer_data_4[2671:2664];
        layer2[11][55:48] = buffer_data_4[2679:2672];
        layer3[11][7:0] = buffer_data_3[2631:2624];
        layer3[11][15:8] = buffer_data_3[2639:2632];
        layer3[11][23:16] = buffer_data_3[2647:2640];
        layer3[11][31:24] = buffer_data_3[2655:2648];
        layer3[11][39:32] = buffer_data_3[2663:2656];
        layer3[11][47:40] = buffer_data_3[2671:2664];
        layer3[11][55:48] = buffer_data_3[2679:2672];
        layer4[11][7:0] = buffer_data_2[2631:2624];
        layer4[11][15:8] = buffer_data_2[2639:2632];
        layer4[11][23:16] = buffer_data_2[2647:2640];
        layer4[11][31:24] = buffer_data_2[2655:2648];
        layer4[11][39:32] = buffer_data_2[2663:2656];
        layer4[11][47:40] = buffer_data_2[2671:2664];
        layer4[11][55:48] = buffer_data_2[2679:2672];
        layer5[11][7:0] = buffer_data_1[2631:2624];
        layer5[11][15:8] = buffer_data_1[2639:2632];
        layer5[11][23:16] = buffer_data_1[2647:2640];
        layer5[11][31:24] = buffer_data_1[2655:2648];
        layer5[11][39:32] = buffer_data_1[2663:2656];
        layer5[11][47:40] = buffer_data_1[2671:2664];
        layer5[11][55:48] = buffer_data_1[2679:2672];
        layer6[11][7:0] = buffer_data_0[2631:2624];
        layer6[11][15:8] = buffer_data_0[2639:2632];
        layer6[11][23:16] = buffer_data_0[2647:2640];
        layer6[11][31:24] = buffer_data_0[2655:2648];
        layer6[11][39:32] = buffer_data_0[2663:2656];
        layer6[11][47:40] = buffer_data_0[2671:2664];
        layer6[11][55:48] = buffer_data_0[2679:2672];
        layer0[12][7:0] = buffer_data_6[2639:2632];
        layer0[12][15:8] = buffer_data_6[2647:2640];
        layer0[12][23:16] = buffer_data_6[2655:2648];
        layer0[12][31:24] = buffer_data_6[2663:2656];
        layer0[12][39:32] = buffer_data_6[2671:2664];
        layer0[12][47:40] = buffer_data_6[2679:2672];
        layer0[12][55:48] = buffer_data_6[2687:2680];
        layer1[12][7:0] = buffer_data_5[2639:2632];
        layer1[12][15:8] = buffer_data_5[2647:2640];
        layer1[12][23:16] = buffer_data_5[2655:2648];
        layer1[12][31:24] = buffer_data_5[2663:2656];
        layer1[12][39:32] = buffer_data_5[2671:2664];
        layer1[12][47:40] = buffer_data_5[2679:2672];
        layer1[12][55:48] = buffer_data_5[2687:2680];
        layer2[12][7:0] = buffer_data_4[2639:2632];
        layer2[12][15:8] = buffer_data_4[2647:2640];
        layer2[12][23:16] = buffer_data_4[2655:2648];
        layer2[12][31:24] = buffer_data_4[2663:2656];
        layer2[12][39:32] = buffer_data_4[2671:2664];
        layer2[12][47:40] = buffer_data_4[2679:2672];
        layer2[12][55:48] = buffer_data_4[2687:2680];
        layer3[12][7:0] = buffer_data_3[2639:2632];
        layer3[12][15:8] = buffer_data_3[2647:2640];
        layer3[12][23:16] = buffer_data_3[2655:2648];
        layer3[12][31:24] = buffer_data_3[2663:2656];
        layer3[12][39:32] = buffer_data_3[2671:2664];
        layer3[12][47:40] = buffer_data_3[2679:2672];
        layer3[12][55:48] = buffer_data_3[2687:2680];
        layer4[12][7:0] = buffer_data_2[2639:2632];
        layer4[12][15:8] = buffer_data_2[2647:2640];
        layer4[12][23:16] = buffer_data_2[2655:2648];
        layer4[12][31:24] = buffer_data_2[2663:2656];
        layer4[12][39:32] = buffer_data_2[2671:2664];
        layer4[12][47:40] = buffer_data_2[2679:2672];
        layer4[12][55:48] = buffer_data_2[2687:2680];
        layer5[12][7:0] = buffer_data_1[2639:2632];
        layer5[12][15:8] = buffer_data_1[2647:2640];
        layer5[12][23:16] = buffer_data_1[2655:2648];
        layer5[12][31:24] = buffer_data_1[2663:2656];
        layer5[12][39:32] = buffer_data_1[2671:2664];
        layer5[12][47:40] = buffer_data_1[2679:2672];
        layer5[12][55:48] = buffer_data_1[2687:2680];
        layer6[12][7:0] = buffer_data_0[2639:2632];
        layer6[12][15:8] = buffer_data_0[2647:2640];
        layer6[12][23:16] = buffer_data_0[2655:2648];
        layer6[12][31:24] = buffer_data_0[2663:2656];
        layer6[12][39:32] = buffer_data_0[2671:2664];
        layer6[12][47:40] = buffer_data_0[2679:2672];
        layer6[12][55:48] = buffer_data_0[2687:2680];
        layer0[13][7:0] = buffer_data_6[2647:2640];
        layer0[13][15:8] = buffer_data_6[2655:2648];
        layer0[13][23:16] = buffer_data_6[2663:2656];
        layer0[13][31:24] = buffer_data_6[2671:2664];
        layer0[13][39:32] = buffer_data_6[2679:2672];
        layer0[13][47:40] = buffer_data_6[2687:2680];
        layer0[13][55:48] = buffer_data_6[2695:2688];
        layer1[13][7:0] = buffer_data_5[2647:2640];
        layer1[13][15:8] = buffer_data_5[2655:2648];
        layer1[13][23:16] = buffer_data_5[2663:2656];
        layer1[13][31:24] = buffer_data_5[2671:2664];
        layer1[13][39:32] = buffer_data_5[2679:2672];
        layer1[13][47:40] = buffer_data_5[2687:2680];
        layer1[13][55:48] = buffer_data_5[2695:2688];
        layer2[13][7:0] = buffer_data_4[2647:2640];
        layer2[13][15:8] = buffer_data_4[2655:2648];
        layer2[13][23:16] = buffer_data_4[2663:2656];
        layer2[13][31:24] = buffer_data_4[2671:2664];
        layer2[13][39:32] = buffer_data_4[2679:2672];
        layer2[13][47:40] = buffer_data_4[2687:2680];
        layer2[13][55:48] = buffer_data_4[2695:2688];
        layer3[13][7:0] = buffer_data_3[2647:2640];
        layer3[13][15:8] = buffer_data_3[2655:2648];
        layer3[13][23:16] = buffer_data_3[2663:2656];
        layer3[13][31:24] = buffer_data_3[2671:2664];
        layer3[13][39:32] = buffer_data_3[2679:2672];
        layer3[13][47:40] = buffer_data_3[2687:2680];
        layer3[13][55:48] = buffer_data_3[2695:2688];
        layer4[13][7:0] = buffer_data_2[2647:2640];
        layer4[13][15:8] = buffer_data_2[2655:2648];
        layer4[13][23:16] = buffer_data_2[2663:2656];
        layer4[13][31:24] = buffer_data_2[2671:2664];
        layer4[13][39:32] = buffer_data_2[2679:2672];
        layer4[13][47:40] = buffer_data_2[2687:2680];
        layer4[13][55:48] = buffer_data_2[2695:2688];
        layer5[13][7:0] = buffer_data_1[2647:2640];
        layer5[13][15:8] = buffer_data_1[2655:2648];
        layer5[13][23:16] = buffer_data_1[2663:2656];
        layer5[13][31:24] = buffer_data_1[2671:2664];
        layer5[13][39:32] = buffer_data_1[2679:2672];
        layer5[13][47:40] = buffer_data_1[2687:2680];
        layer5[13][55:48] = buffer_data_1[2695:2688];
        layer6[13][7:0] = buffer_data_0[2647:2640];
        layer6[13][15:8] = buffer_data_0[2655:2648];
        layer6[13][23:16] = buffer_data_0[2663:2656];
        layer6[13][31:24] = buffer_data_0[2671:2664];
        layer6[13][39:32] = buffer_data_0[2679:2672];
        layer6[13][47:40] = buffer_data_0[2687:2680];
        layer6[13][55:48] = buffer_data_0[2695:2688];
        layer0[14][7:0] = buffer_data_6[2655:2648];
        layer0[14][15:8] = buffer_data_6[2663:2656];
        layer0[14][23:16] = buffer_data_6[2671:2664];
        layer0[14][31:24] = buffer_data_6[2679:2672];
        layer0[14][39:32] = buffer_data_6[2687:2680];
        layer0[14][47:40] = buffer_data_6[2695:2688];
        layer0[14][55:48] = buffer_data_6[2703:2696];
        layer1[14][7:0] = buffer_data_5[2655:2648];
        layer1[14][15:8] = buffer_data_5[2663:2656];
        layer1[14][23:16] = buffer_data_5[2671:2664];
        layer1[14][31:24] = buffer_data_5[2679:2672];
        layer1[14][39:32] = buffer_data_5[2687:2680];
        layer1[14][47:40] = buffer_data_5[2695:2688];
        layer1[14][55:48] = buffer_data_5[2703:2696];
        layer2[14][7:0] = buffer_data_4[2655:2648];
        layer2[14][15:8] = buffer_data_4[2663:2656];
        layer2[14][23:16] = buffer_data_4[2671:2664];
        layer2[14][31:24] = buffer_data_4[2679:2672];
        layer2[14][39:32] = buffer_data_4[2687:2680];
        layer2[14][47:40] = buffer_data_4[2695:2688];
        layer2[14][55:48] = buffer_data_4[2703:2696];
        layer3[14][7:0] = buffer_data_3[2655:2648];
        layer3[14][15:8] = buffer_data_3[2663:2656];
        layer3[14][23:16] = buffer_data_3[2671:2664];
        layer3[14][31:24] = buffer_data_3[2679:2672];
        layer3[14][39:32] = buffer_data_3[2687:2680];
        layer3[14][47:40] = buffer_data_3[2695:2688];
        layer3[14][55:48] = buffer_data_3[2703:2696];
        layer4[14][7:0] = buffer_data_2[2655:2648];
        layer4[14][15:8] = buffer_data_2[2663:2656];
        layer4[14][23:16] = buffer_data_2[2671:2664];
        layer4[14][31:24] = buffer_data_2[2679:2672];
        layer4[14][39:32] = buffer_data_2[2687:2680];
        layer4[14][47:40] = buffer_data_2[2695:2688];
        layer4[14][55:48] = buffer_data_2[2703:2696];
        layer5[14][7:0] = buffer_data_1[2655:2648];
        layer5[14][15:8] = buffer_data_1[2663:2656];
        layer5[14][23:16] = buffer_data_1[2671:2664];
        layer5[14][31:24] = buffer_data_1[2679:2672];
        layer5[14][39:32] = buffer_data_1[2687:2680];
        layer5[14][47:40] = buffer_data_1[2695:2688];
        layer5[14][55:48] = buffer_data_1[2703:2696];
        layer6[14][7:0] = buffer_data_0[2655:2648];
        layer6[14][15:8] = buffer_data_0[2663:2656];
        layer6[14][23:16] = buffer_data_0[2671:2664];
        layer6[14][31:24] = buffer_data_0[2679:2672];
        layer6[14][39:32] = buffer_data_0[2687:2680];
        layer6[14][47:40] = buffer_data_0[2695:2688];
        layer6[14][55:48] = buffer_data_0[2703:2696];
        layer0[15][7:0] = buffer_data_6[2663:2656];
        layer0[15][15:8] = buffer_data_6[2671:2664];
        layer0[15][23:16] = buffer_data_6[2679:2672];
        layer0[15][31:24] = buffer_data_6[2687:2680];
        layer0[15][39:32] = buffer_data_6[2695:2688];
        layer0[15][47:40] = buffer_data_6[2703:2696];
        layer0[15][55:48] = buffer_data_6[2711:2704];
        layer1[15][7:0] = buffer_data_5[2663:2656];
        layer1[15][15:8] = buffer_data_5[2671:2664];
        layer1[15][23:16] = buffer_data_5[2679:2672];
        layer1[15][31:24] = buffer_data_5[2687:2680];
        layer1[15][39:32] = buffer_data_5[2695:2688];
        layer1[15][47:40] = buffer_data_5[2703:2696];
        layer1[15][55:48] = buffer_data_5[2711:2704];
        layer2[15][7:0] = buffer_data_4[2663:2656];
        layer2[15][15:8] = buffer_data_4[2671:2664];
        layer2[15][23:16] = buffer_data_4[2679:2672];
        layer2[15][31:24] = buffer_data_4[2687:2680];
        layer2[15][39:32] = buffer_data_4[2695:2688];
        layer2[15][47:40] = buffer_data_4[2703:2696];
        layer2[15][55:48] = buffer_data_4[2711:2704];
        layer3[15][7:0] = buffer_data_3[2663:2656];
        layer3[15][15:8] = buffer_data_3[2671:2664];
        layer3[15][23:16] = buffer_data_3[2679:2672];
        layer3[15][31:24] = buffer_data_3[2687:2680];
        layer3[15][39:32] = buffer_data_3[2695:2688];
        layer3[15][47:40] = buffer_data_3[2703:2696];
        layer3[15][55:48] = buffer_data_3[2711:2704];
        layer4[15][7:0] = buffer_data_2[2663:2656];
        layer4[15][15:8] = buffer_data_2[2671:2664];
        layer4[15][23:16] = buffer_data_2[2679:2672];
        layer4[15][31:24] = buffer_data_2[2687:2680];
        layer4[15][39:32] = buffer_data_2[2695:2688];
        layer4[15][47:40] = buffer_data_2[2703:2696];
        layer4[15][55:48] = buffer_data_2[2711:2704];
        layer5[15][7:0] = buffer_data_1[2663:2656];
        layer5[15][15:8] = buffer_data_1[2671:2664];
        layer5[15][23:16] = buffer_data_1[2679:2672];
        layer5[15][31:24] = buffer_data_1[2687:2680];
        layer5[15][39:32] = buffer_data_1[2695:2688];
        layer5[15][47:40] = buffer_data_1[2703:2696];
        layer5[15][55:48] = buffer_data_1[2711:2704];
        layer6[15][7:0] = buffer_data_0[2663:2656];
        layer6[15][15:8] = buffer_data_0[2671:2664];
        layer6[15][23:16] = buffer_data_0[2679:2672];
        layer6[15][31:24] = buffer_data_0[2687:2680];
        layer6[15][39:32] = buffer_data_0[2695:2688];
        layer6[15][47:40] = buffer_data_0[2703:2696];
        layer6[15][55:48] = buffer_data_0[2711:2704];
        layer0[16][7:0] = buffer_data_6[2671:2664];
        layer0[16][15:8] = buffer_data_6[2679:2672];
        layer0[16][23:16] = buffer_data_6[2687:2680];
        layer0[16][31:24] = buffer_data_6[2695:2688];
        layer0[16][39:32] = buffer_data_6[2703:2696];
        layer0[16][47:40] = buffer_data_6[2711:2704];
        layer0[16][55:48] = buffer_data_6[2719:2712];
        layer1[16][7:0] = buffer_data_5[2671:2664];
        layer1[16][15:8] = buffer_data_5[2679:2672];
        layer1[16][23:16] = buffer_data_5[2687:2680];
        layer1[16][31:24] = buffer_data_5[2695:2688];
        layer1[16][39:32] = buffer_data_5[2703:2696];
        layer1[16][47:40] = buffer_data_5[2711:2704];
        layer1[16][55:48] = buffer_data_5[2719:2712];
        layer2[16][7:0] = buffer_data_4[2671:2664];
        layer2[16][15:8] = buffer_data_4[2679:2672];
        layer2[16][23:16] = buffer_data_4[2687:2680];
        layer2[16][31:24] = buffer_data_4[2695:2688];
        layer2[16][39:32] = buffer_data_4[2703:2696];
        layer2[16][47:40] = buffer_data_4[2711:2704];
        layer2[16][55:48] = buffer_data_4[2719:2712];
        layer3[16][7:0] = buffer_data_3[2671:2664];
        layer3[16][15:8] = buffer_data_3[2679:2672];
        layer3[16][23:16] = buffer_data_3[2687:2680];
        layer3[16][31:24] = buffer_data_3[2695:2688];
        layer3[16][39:32] = buffer_data_3[2703:2696];
        layer3[16][47:40] = buffer_data_3[2711:2704];
        layer3[16][55:48] = buffer_data_3[2719:2712];
        layer4[16][7:0] = buffer_data_2[2671:2664];
        layer4[16][15:8] = buffer_data_2[2679:2672];
        layer4[16][23:16] = buffer_data_2[2687:2680];
        layer4[16][31:24] = buffer_data_2[2695:2688];
        layer4[16][39:32] = buffer_data_2[2703:2696];
        layer4[16][47:40] = buffer_data_2[2711:2704];
        layer4[16][55:48] = buffer_data_2[2719:2712];
        layer5[16][7:0] = buffer_data_1[2671:2664];
        layer5[16][15:8] = buffer_data_1[2679:2672];
        layer5[16][23:16] = buffer_data_1[2687:2680];
        layer5[16][31:24] = buffer_data_1[2695:2688];
        layer5[16][39:32] = buffer_data_1[2703:2696];
        layer5[16][47:40] = buffer_data_1[2711:2704];
        layer5[16][55:48] = buffer_data_1[2719:2712];
        layer6[16][7:0] = buffer_data_0[2671:2664];
        layer6[16][15:8] = buffer_data_0[2679:2672];
        layer6[16][23:16] = buffer_data_0[2687:2680];
        layer6[16][31:24] = buffer_data_0[2695:2688];
        layer6[16][39:32] = buffer_data_0[2703:2696];
        layer6[16][47:40] = buffer_data_0[2711:2704];
        layer6[16][55:48] = buffer_data_0[2719:2712];
        layer0[17][7:0] = buffer_data_6[2679:2672];
        layer0[17][15:8] = buffer_data_6[2687:2680];
        layer0[17][23:16] = buffer_data_6[2695:2688];
        layer0[17][31:24] = buffer_data_6[2703:2696];
        layer0[17][39:32] = buffer_data_6[2711:2704];
        layer0[17][47:40] = buffer_data_6[2719:2712];
        layer0[17][55:48] = buffer_data_6[2727:2720];
        layer1[17][7:0] = buffer_data_5[2679:2672];
        layer1[17][15:8] = buffer_data_5[2687:2680];
        layer1[17][23:16] = buffer_data_5[2695:2688];
        layer1[17][31:24] = buffer_data_5[2703:2696];
        layer1[17][39:32] = buffer_data_5[2711:2704];
        layer1[17][47:40] = buffer_data_5[2719:2712];
        layer1[17][55:48] = buffer_data_5[2727:2720];
        layer2[17][7:0] = buffer_data_4[2679:2672];
        layer2[17][15:8] = buffer_data_4[2687:2680];
        layer2[17][23:16] = buffer_data_4[2695:2688];
        layer2[17][31:24] = buffer_data_4[2703:2696];
        layer2[17][39:32] = buffer_data_4[2711:2704];
        layer2[17][47:40] = buffer_data_4[2719:2712];
        layer2[17][55:48] = buffer_data_4[2727:2720];
        layer3[17][7:0] = buffer_data_3[2679:2672];
        layer3[17][15:8] = buffer_data_3[2687:2680];
        layer3[17][23:16] = buffer_data_3[2695:2688];
        layer3[17][31:24] = buffer_data_3[2703:2696];
        layer3[17][39:32] = buffer_data_3[2711:2704];
        layer3[17][47:40] = buffer_data_3[2719:2712];
        layer3[17][55:48] = buffer_data_3[2727:2720];
        layer4[17][7:0] = buffer_data_2[2679:2672];
        layer4[17][15:8] = buffer_data_2[2687:2680];
        layer4[17][23:16] = buffer_data_2[2695:2688];
        layer4[17][31:24] = buffer_data_2[2703:2696];
        layer4[17][39:32] = buffer_data_2[2711:2704];
        layer4[17][47:40] = buffer_data_2[2719:2712];
        layer4[17][55:48] = buffer_data_2[2727:2720];
        layer5[17][7:0] = buffer_data_1[2679:2672];
        layer5[17][15:8] = buffer_data_1[2687:2680];
        layer5[17][23:16] = buffer_data_1[2695:2688];
        layer5[17][31:24] = buffer_data_1[2703:2696];
        layer5[17][39:32] = buffer_data_1[2711:2704];
        layer5[17][47:40] = buffer_data_1[2719:2712];
        layer5[17][55:48] = buffer_data_1[2727:2720];
        layer6[17][7:0] = buffer_data_0[2679:2672];
        layer6[17][15:8] = buffer_data_0[2687:2680];
        layer6[17][23:16] = buffer_data_0[2695:2688];
        layer6[17][31:24] = buffer_data_0[2703:2696];
        layer6[17][39:32] = buffer_data_0[2711:2704];
        layer6[17][47:40] = buffer_data_0[2719:2712];
        layer6[17][55:48] = buffer_data_0[2727:2720];
        layer0[18][7:0] = buffer_data_6[2687:2680];
        layer0[18][15:8] = buffer_data_6[2695:2688];
        layer0[18][23:16] = buffer_data_6[2703:2696];
        layer0[18][31:24] = buffer_data_6[2711:2704];
        layer0[18][39:32] = buffer_data_6[2719:2712];
        layer0[18][47:40] = buffer_data_6[2727:2720];
        layer0[18][55:48] = buffer_data_6[2735:2728];
        layer1[18][7:0] = buffer_data_5[2687:2680];
        layer1[18][15:8] = buffer_data_5[2695:2688];
        layer1[18][23:16] = buffer_data_5[2703:2696];
        layer1[18][31:24] = buffer_data_5[2711:2704];
        layer1[18][39:32] = buffer_data_5[2719:2712];
        layer1[18][47:40] = buffer_data_5[2727:2720];
        layer1[18][55:48] = buffer_data_5[2735:2728];
        layer2[18][7:0] = buffer_data_4[2687:2680];
        layer2[18][15:8] = buffer_data_4[2695:2688];
        layer2[18][23:16] = buffer_data_4[2703:2696];
        layer2[18][31:24] = buffer_data_4[2711:2704];
        layer2[18][39:32] = buffer_data_4[2719:2712];
        layer2[18][47:40] = buffer_data_4[2727:2720];
        layer2[18][55:48] = buffer_data_4[2735:2728];
        layer3[18][7:0] = buffer_data_3[2687:2680];
        layer3[18][15:8] = buffer_data_3[2695:2688];
        layer3[18][23:16] = buffer_data_3[2703:2696];
        layer3[18][31:24] = buffer_data_3[2711:2704];
        layer3[18][39:32] = buffer_data_3[2719:2712];
        layer3[18][47:40] = buffer_data_3[2727:2720];
        layer3[18][55:48] = buffer_data_3[2735:2728];
        layer4[18][7:0] = buffer_data_2[2687:2680];
        layer4[18][15:8] = buffer_data_2[2695:2688];
        layer4[18][23:16] = buffer_data_2[2703:2696];
        layer4[18][31:24] = buffer_data_2[2711:2704];
        layer4[18][39:32] = buffer_data_2[2719:2712];
        layer4[18][47:40] = buffer_data_2[2727:2720];
        layer4[18][55:48] = buffer_data_2[2735:2728];
        layer5[18][7:0] = buffer_data_1[2687:2680];
        layer5[18][15:8] = buffer_data_1[2695:2688];
        layer5[18][23:16] = buffer_data_1[2703:2696];
        layer5[18][31:24] = buffer_data_1[2711:2704];
        layer5[18][39:32] = buffer_data_1[2719:2712];
        layer5[18][47:40] = buffer_data_1[2727:2720];
        layer5[18][55:48] = buffer_data_1[2735:2728];
        layer6[18][7:0] = buffer_data_0[2687:2680];
        layer6[18][15:8] = buffer_data_0[2695:2688];
        layer6[18][23:16] = buffer_data_0[2703:2696];
        layer6[18][31:24] = buffer_data_0[2711:2704];
        layer6[18][39:32] = buffer_data_0[2719:2712];
        layer6[18][47:40] = buffer_data_0[2727:2720];
        layer6[18][55:48] = buffer_data_0[2735:2728];
        layer0[19][7:0] = buffer_data_6[2695:2688];
        layer0[19][15:8] = buffer_data_6[2703:2696];
        layer0[19][23:16] = buffer_data_6[2711:2704];
        layer0[19][31:24] = buffer_data_6[2719:2712];
        layer0[19][39:32] = buffer_data_6[2727:2720];
        layer0[19][47:40] = buffer_data_6[2735:2728];
        layer0[19][55:48] = buffer_data_6[2743:2736];
        layer1[19][7:0] = buffer_data_5[2695:2688];
        layer1[19][15:8] = buffer_data_5[2703:2696];
        layer1[19][23:16] = buffer_data_5[2711:2704];
        layer1[19][31:24] = buffer_data_5[2719:2712];
        layer1[19][39:32] = buffer_data_5[2727:2720];
        layer1[19][47:40] = buffer_data_5[2735:2728];
        layer1[19][55:48] = buffer_data_5[2743:2736];
        layer2[19][7:0] = buffer_data_4[2695:2688];
        layer2[19][15:8] = buffer_data_4[2703:2696];
        layer2[19][23:16] = buffer_data_4[2711:2704];
        layer2[19][31:24] = buffer_data_4[2719:2712];
        layer2[19][39:32] = buffer_data_4[2727:2720];
        layer2[19][47:40] = buffer_data_4[2735:2728];
        layer2[19][55:48] = buffer_data_4[2743:2736];
        layer3[19][7:0] = buffer_data_3[2695:2688];
        layer3[19][15:8] = buffer_data_3[2703:2696];
        layer3[19][23:16] = buffer_data_3[2711:2704];
        layer3[19][31:24] = buffer_data_3[2719:2712];
        layer3[19][39:32] = buffer_data_3[2727:2720];
        layer3[19][47:40] = buffer_data_3[2735:2728];
        layer3[19][55:48] = buffer_data_3[2743:2736];
        layer4[19][7:0] = buffer_data_2[2695:2688];
        layer4[19][15:8] = buffer_data_2[2703:2696];
        layer4[19][23:16] = buffer_data_2[2711:2704];
        layer4[19][31:24] = buffer_data_2[2719:2712];
        layer4[19][39:32] = buffer_data_2[2727:2720];
        layer4[19][47:40] = buffer_data_2[2735:2728];
        layer4[19][55:48] = buffer_data_2[2743:2736];
        layer5[19][7:0] = buffer_data_1[2695:2688];
        layer5[19][15:8] = buffer_data_1[2703:2696];
        layer5[19][23:16] = buffer_data_1[2711:2704];
        layer5[19][31:24] = buffer_data_1[2719:2712];
        layer5[19][39:32] = buffer_data_1[2727:2720];
        layer5[19][47:40] = buffer_data_1[2735:2728];
        layer5[19][55:48] = buffer_data_1[2743:2736];
        layer6[19][7:0] = buffer_data_0[2695:2688];
        layer6[19][15:8] = buffer_data_0[2703:2696];
        layer6[19][23:16] = buffer_data_0[2711:2704];
        layer6[19][31:24] = buffer_data_0[2719:2712];
        layer6[19][39:32] = buffer_data_0[2727:2720];
        layer6[19][47:40] = buffer_data_0[2735:2728];
        layer6[19][55:48] = buffer_data_0[2743:2736];
        layer0[20][7:0] = buffer_data_6[2703:2696];
        layer0[20][15:8] = buffer_data_6[2711:2704];
        layer0[20][23:16] = buffer_data_6[2719:2712];
        layer0[20][31:24] = buffer_data_6[2727:2720];
        layer0[20][39:32] = buffer_data_6[2735:2728];
        layer0[20][47:40] = buffer_data_6[2743:2736];
        layer0[20][55:48] = buffer_data_6[2751:2744];
        layer1[20][7:0] = buffer_data_5[2703:2696];
        layer1[20][15:8] = buffer_data_5[2711:2704];
        layer1[20][23:16] = buffer_data_5[2719:2712];
        layer1[20][31:24] = buffer_data_5[2727:2720];
        layer1[20][39:32] = buffer_data_5[2735:2728];
        layer1[20][47:40] = buffer_data_5[2743:2736];
        layer1[20][55:48] = buffer_data_5[2751:2744];
        layer2[20][7:0] = buffer_data_4[2703:2696];
        layer2[20][15:8] = buffer_data_4[2711:2704];
        layer2[20][23:16] = buffer_data_4[2719:2712];
        layer2[20][31:24] = buffer_data_4[2727:2720];
        layer2[20][39:32] = buffer_data_4[2735:2728];
        layer2[20][47:40] = buffer_data_4[2743:2736];
        layer2[20][55:48] = buffer_data_4[2751:2744];
        layer3[20][7:0] = buffer_data_3[2703:2696];
        layer3[20][15:8] = buffer_data_3[2711:2704];
        layer3[20][23:16] = buffer_data_3[2719:2712];
        layer3[20][31:24] = buffer_data_3[2727:2720];
        layer3[20][39:32] = buffer_data_3[2735:2728];
        layer3[20][47:40] = buffer_data_3[2743:2736];
        layer3[20][55:48] = buffer_data_3[2751:2744];
        layer4[20][7:0] = buffer_data_2[2703:2696];
        layer4[20][15:8] = buffer_data_2[2711:2704];
        layer4[20][23:16] = buffer_data_2[2719:2712];
        layer4[20][31:24] = buffer_data_2[2727:2720];
        layer4[20][39:32] = buffer_data_2[2735:2728];
        layer4[20][47:40] = buffer_data_2[2743:2736];
        layer4[20][55:48] = buffer_data_2[2751:2744];
        layer5[20][7:0] = buffer_data_1[2703:2696];
        layer5[20][15:8] = buffer_data_1[2711:2704];
        layer5[20][23:16] = buffer_data_1[2719:2712];
        layer5[20][31:24] = buffer_data_1[2727:2720];
        layer5[20][39:32] = buffer_data_1[2735:2728];
        layer5[20][47:40] = buffer_data_1[2743:2736];
        layer5[20][55:48] = buffer_data_1[2751:2744];
        layer6[20][7:0] = buffer_data_0[2703:2696];
        layer6[20][15:8] = buffer_data_0[2711:2704];
        layer6[20][23:16] = buffer_data_0[2719:2712];
        layer6[20][31:24] = buffer_data_0[2727:2720];
        layer6[20][39:32] = buffer_data_0[2735:2728];
        layer6[20][47:40] = buffer_data_0[2743:2736];
        layer6[20][55:48] = buffer_data_0[2751:2744];
        layer0[21][7:0] = buffer_data_6[2711:2704];
        layer0[21][15:8] = buffer_data_6[2719:2712];
        layer0[21][23:16] = buffer_data_6[2727:2720];
        layer0[21][31:24] = buffer_data_6[2735:2728];
        layer0[21][39:32] = buffer_data_6[2743:2736];
        layer0[21][47:40] = buffer_data_6[2751:2744];
        layer0[21][55:48] = buffer_data_6[2759:2752];
        layer1[21][7:0] = buffer_data_5[2711:2704];
        layer1[21][15:8] = buffer_data_5[2719:2712];
        layer1[21][23:16] = buffer_data_5[2727:2720];
        layer1[21][31:24] = buffer_data_5[2735:2728];
        layer1[21][39:32] = buffer_data_5[2743:2736];
        layer1[21][47:40] = buffer_data_5[2751:2744];
        layer1[21][55:48] = buffer_data_5[2759:2752];
        layer2[21][7:0] = buffer_data_4[2711:2704];
        layer2[21][15:8] = buffer_data_4[2719:2712];
        layer2[21][23:16] = buffer_data_4[2727:2720];
        layer2[21][31:24] = buffer_data_4[2735:2728];
        layer2[21][39:32] = buffer_data_4[2743:2736];
        layer2[21][47:40] = buffer_data_4[2751:2744];
        layer2[21][55:48] = buffer_data_4[2759:2752];
        layer3[21][7:0] = buffer_data_3[2711:2704];
        layer3[21][15:8] = buffer_data_3[2719:2712];
        layer3[21][23:16] = buffer_data_3[2727:2720];
        layer3[21][31:24] = buffer_data_3[2735:2728];
        layer3[21][39:32] = buffer_data_3[2743:2736];
        layer3[21][47:40] = buffer_data_3[2751:2744];
        layer3[21][55:48] = buffer_data_3[2759:2752];
        layer4[21][7:0] = buffer_data_2[2711:2704];
        layer4[21][15:8] = buffer_data_2[2719:2712];
        layer4[21][23:16] = buffer_data_2[2727:2720];
        layer4[21][31:24] = buffer_data_2[2735:2728];
        layer4[21][39:32] = buffer_data_2[2743:2736];
        layer4[21][47:40] = buffer_data_2[2751:2744];
        layer4[21][55:48] = buffer_data_2[2759:2752];
        layer5[21][7:0] = buffer_data_1[2711:2704];
        layer5[21][15:8] = buffer_data_1[2719:2712];
        layer5[21][23:16] = buffer_data_1[2727:2720];
        layer5[21][31:24] = buffer_data_1[2735:2728];
        layer5[21][39:32] = buffer_data_1[2743:2736];
        layer5[21][47:40] = buffer_data_1[2751:2744];
        layer5[21][55:48] = buffer_data_1[2759:2752];
        layer6[21][7:0] = buffer_data_0[2711:2704];
        layer6[21][15:8] = buffer_data_0[2719:2712];
        layer6[21][23:16] = buffer_data_0[2727:2720];
        layer6[21][31:24] = buffer_data_0[2735:2728];
        layer6[21][39:32] = buffer_data_0[2743:2736];
        layer6[21][47:40] = buffer_data_0[2751:2744];
        layer6[21][55:48] = buffer_data_0[2759:2752];
        layer0[22][7:0] = buffer_data_6[2719:2712];
        layer0[22][15:8] = buffer_data_6[2727:2720];
        layer0[22][23:16] = buffer_data_6[2735:2728];
        layer0[22][31:24] = buffer_data_6[2743:2736];
        layer0[22][39:32] = buffer_data_6[2751:2744];
        layer0[22][47:40] = buffer_data_6[2759:2752];
        layer0[22][55:48] = buffer_data_6[2767:2760];
        layer1[22][7:0] = buffer_data_5[2719:2712];
        layer1[22][15:8] = buffer_data_5[2727:2720];
        layer1[22][23:16] = buffer_data_5[2735:2728];
        layer1[22][31:24] = buffer_data_5[2743:2736];
        layer1[22][39:32] = buffer_data_5[2751:2744];
        layer1[22][47:40] = buffer_data_5[2759:2752];
        layer1[22][55:48] = buffer_data_5[2767:2760];
        layer2[22][7:0] = buffer_data_4[2719:2712];
        layer2[22][15:8] = buffer_data_4[2727:2720];
        layer2[22][23:16] = buffer_data_4[2735:2728];
        layer2[22][31:24] = buffer_data_4[2743:2736];
        layer2[22][39:32] = buffer_data_4[2751:2744];
        layer2[22][47:40] = buffer_data_4[2759:2752];
        layer2[22][55:48] = buffer_data_4[2767:2760];
        layer3[22][7:0] = buffer_data_3[2719:2712];
        layer3[22][15:8] = buffer_data_3[2727:2720];
        layer3[22][23:16] = buffer_data_3[2735:2728];
        layer3[22][31:24] = buffer_data_3[2743:2736];
        layer3[22][39:32] = buffer_data_3[2751:2744];
        layer3[22][47:40] = buffer_data_3[2759:2752];
        layer3[22][55:48] = buffer_data_3[2767:2760];
        layer4[22][7:0] = buffer_data_2[2719:2712];
        layer4[22][15:8] = buffer_data_2[2727:2720];
        layer4[22][23:16] = buffer_data_2[2735:2728];
        layer4[22][31:24] = buffer_data_2[2743:2736];
        layer4[22][39:32] = buffer_data_2[2751:2744];
        layer4[22][47:40] = buffer_data_2[2759:2752];
        layer4[22][55:48] = buffer_data_2[2767:2760];
        layer5[22][7:0] = buffer_data_1[2719:2712];
        layer5[22][15:8] = buffer_data_1[2727:2720];
        layer5[22][23:16] = buffer_data_1[2735:2728];
        layer5[22][31:24] = buffer_data_1[2743:2736];
        layer5[22][39:32] = buffer_data_1[2751:2744];
        layer5[22][47:40] = buffer_data_1[2759:2752];
        layer5[22][55:48] = buffer_data_1[2767:2760];
        layer6[22][7:0] = buffer_data_0[2719:2712];
        layer6[22][15:8] = buffer_data_0[2727:2720];
        layer6[22][23:16] = buffer_data_0[2735:2728];
        layer6[22][31:24] = buffer_data_0[2743:2736];
        layer6[22][39:32] = buffer_data_0[2751:2744];
        layer6[22][47:40] = buffer_data_0[2759:2752];
        layer6[22][55:48] = buffer_data_0[2767:2760];
        layer0[23][7:0] = buffer_data_6[2727:2720];
        layer0[23][15:8] = buffer_data_6[2735:2728];
        layer0[23][23:16] = buffer_data_6[2743:2736];
        layer0[23][31:24] = buffer_data_6[2751:2744];
        layer0[23][39:32] = buffer_data_6[2759:2752];
        layer0[23][47:40] = buffer_data_6[2767:2760];
        layer0[23][55:48] = buffer_data_6[2775:2768];
        layer1[23][7:0] = buffer_data_5[2727:2720];
        layer1[23][15:8] = buffer_data_5[2735:2728];
        layer1[23][23:16] = buffer_data_5[2743:2736];
        layer1[23][31:24] = buffer_data_5[2751:2744];
        layer1[23][39:32] = buffer_data_5[2759:2752];
        layer1[23][47:40] = buffer_data_5[2767:2760];
        layer1[23][55:48] = buffer_data_5[2775:2768];
        layer2[23][7:0] = buffer_data_4[2727:2720];
        layer2[23][15:8] = buffer_data_4[2735:2728];
        layer2[23][23:16] = buffer_data_4[2743:2736];
        layer2[23][31:24] = buffer_data_4[2751:2744];
        layer2[23][39:32] = buffer_data_4[2759:2752];
        layer2[23][47:40] = buffer_data_4[2767:2760];
        layer2[23][55:48] = buffer_data_4[2775:2768];
        layer3[23][7:0] = buffer_data_3[2727:2720];
        layer3[23][15:8] = buffer_data_3[2735:2728];
        layer3[23][23:16] = buffer_data_3[2743:2736];
        layer3[23][31:24] = buffer_data_3[2751:2744];
        layer3[23][39:32] = buffer_data_3[2759:2752];
        layer3[23][47:40] = buffer_data_3[2767:2760];
        layer3[23][55:48] = buffer_data_3[2775:2768];
        layer4[23][7:0] = buffer_data_2[2727:2720];
        layer4[23][15:8] = buffer_data_2[2735:2728];
        layer4[23][23:16] = buffer_data_2[2743:2736];
        layer4[23][31:24] = buffer_data_2[2751:2744];
        layer4[23][39:32] = buffer_data_2[2759:2752];
        layer4[23][47:40] = buffer_data_2[2767:2760];
        layer4[23][55:48] = buffer_data_2[2775:2768];
        layer5[23][7:0] = buffer_data_1[2727:2720];
        layer5[23][15:8] = buffer_data_1[2735:2728];
        layer5[23][23:16] = buffer_data_1[2743:2736];
        layer5[23][31:24] = buffer_data_1[2751:2744];
        layer5[23][39:32] = buffer_data_1[2759:2752];
        layer5[23][47:40] = buffer_data_1[2767:2760];
        layer5[23][55:48] = buffer_data_1[2775:2768];
        layer6[23][7:0] = buffer_data_0[2727:2720];
        layer6[23][15:8] = buffer_data_0[2735:2728];
        layer6[23][23:16] = buffer_data_0[2743:2736];
        layer6[23][31:24] = buffer_data_0[2751:2744];
        layer6[23][39:32] = buffer_data_0[2759:2752];
        layer6[23][47:40] = buffer_data_0[2767:2760];
        layer6[23][55:48] = buffer_data_0[2775:2768];
        layer0[24][7:0] = buffer_data_6[2735:2728];
        layer0[24][15:8] = buffer_data_6[2743:2736];
        layer0[24][23:16] = buffer_data_6[2751:2744];
        layer0[24][31:24] = buffer_data_6[2759:2752];
        layer0[24][39:32] = buffer_data_6[2767:2760];
        layer0[24][47:40] = buffer_data_6[2775:2768];
        layer0[24][55:48] = buffer_data_6[2783:2776];
        layer1[24][7:0] = buffer_data_5[2735:2728];
        layer1[24][15:8] = buffer_data_5[2743:2736];
        layer1[24][23:16] = buffer_data_5[2751:2744];
        layer1[24][31:24] = buffer_data_5[2759:2752];
        layer1[24][39:32] = buffer_data_5[2767:2760];
        layer1[24][47:40] = buffer_data_5[2775:2768];
        layer1[24][55:48] = buffer_data_5[2783:2776];
        layer2[24][7:0] = buffer_data_4[2735:2728];
        layer2[24][15:8] = buffer_data_4[2743:2736];
        layer2[24][23:16] = buffer_data_4[2751:2744];
        layer2[24][31:24] = buffer_data_4[2759:2752];
        layer2[24][39:32] = buffer_data_4[2767:2760];
        layer2[24][47:40] = buffer_data_4[2775:2768];
        layer2[24][55:48] = buffer_data_4[2783:2776];
        layer3[24][7:0] = buffer_data_3[2735:2728];
        layer3[24][15:8] = buffer_data_3[2743:2736];
        layer3[24][23:16] = buffer_data_3[2751:2744];
        layer3[24][31:24] = buffer_data_3[2759:2752];
        layer3[24][39:32] = buffer_data_3[2767:2760];
        layer3[24][47:40] = buffer_data_3[2775:2768];
        layer3[24][55:48] = buffer_data_3[2783:2776];
        layer4[24][7:0] = buffer_data_2[2735:2728];
        layer4[24][15:8] = buffer_data_2[2743:2736];
        layer4[24][23:16] = buffer_data_2[2751:2744];
        layer4[24][31:24] = buffer_data_2[2759:2752];
        layer4[24][39:32] = buffer_data_2[2767:2760];
        layer4[24][47:40] = buffer_data_2[2775:2768];
        layer4[24][55:48] = buffer_data_2[2783:2776];
        layer5[24][7:0] = buffer_data_1[2735:2728];
        layer5[24][15:8] = buffer_data_1[2743:2736];
        layer5[24][23:16] = buffer_data_1[2751:2744];
        layer5[24][31:24] = buffer_data_1[2759:2752];
        layer5[24][39:32] = buffer_data_1[2767:2760];
        layer5[24][47:40] = buffer_data_1[2775:2768];
        layer5[24][55:48] = buffer_data_1[2783:2776];
        layer6[24][7:0] = buffer_data_0[2735:2728];
        layer6[24][15:8] = buffer_data_0[2743:2736];
        layer6[24][23:16] = buffer_data_0[2751:2744];
        layer6[24][31:24] = buffer_data_0[2759:2752];
        layer6[24][39:32] = buffer_data_0[2767:2760];
        layer6[24][47:40] = buffer_data_0[2775:2768];
        layer6[24][55:48] = buffer_data_0[2783:2776];
        layer0[25][7:0] = buffer_data_6[2743:2736];
        layer0[25][15:8] = buffer_data_6[2751:2744];
        layer0[25][23:16] = buffer_data_6[2759:2752];
        layer0[25][31:24] = buffer_data_6[2767:2760];
        layer0[25][39:32] = buffer_data_6[2775:2768];
        layer0[25][47:40] = buffer_data_6[2783:2776];
        layer0[25][55:48] = buffer_data_6[2791:2784];
        layer1[25][7:0] = buffer_data_5[2743:2736];
        layer1[25][15:8] = buffer_data_5[2751:2744];
        layer1[25][23:16] = buffer_data_5[2759:2752];
        layer1[25][31:24] = buffer_data_5[2767:2760];
        layer1[25][39:32] = buffer_data_5[2775:2768];
        layer1[25][47:40] = buffer_data_5[2783:2776];
        layer1[25][55:48] = buffer_data_5[2791:2784];
        layer2[25][7:0] = buffer_data_4[2743:2736];
        layer2[25][15:8] = buffer_data_4[2751:2744];
        layer2[25][23:16] = buffer_data_4[2759:2752];
        layer2[25][31:24] = buffer_data_4[2767:2760];
        layer2[25][39:32] = buffer_data_4[2775:2768];
        layer2[25][47:40] = buffer_data_4[2783:2776];
        layer2[25][55:48] = buffer_data_4[2791:2784];
        layer3[25][7:0] = buffer_data_3[2743:2736];
        layer3[25][15:8] = buffer_data_3[2751:2744];
        layer3[25][23:16] = buffer_data_3[2759:2752];
        layer3[25][31:24] = buffer_data_3[2767:2760];
        layer3[25][39:32] = buffer_data_3[2775:2768];
        layer3[25][47:40] = buffer_data_3[2783:2776];
        layer3[25][55:48] = buffer_data_3[2791:2784];
        layer4[25][7:0] = buffer_data_2[2743:2736];
        layer4[25][15:8] = buffer_data_2[2751:2744];
        layer4[25][23:16] = buffer_data_2[2759:2752];
        layer4[25][31:24] = buffer_data_2[2767:2760];
        layer4[25][39:32] = buffer_data_2[2775:2768];
        layer4[25][47:40] = buffer_data_2[2783:2776];
        layer4[25][55:48] = buffer_data_2[2791:2784];
        layer5[25][7:0] = buffer_data_1[2743:2736];
        layer5[25][15:8] = buffer_data_1[2751:2744];
        layer5[25][23:16] = buffer_data_1[2759:2752];
        layer5[25][31:24] = buffer_data_1[2767:2760];
        layer5[25][39:32] = buffer_data_1[2775:2768];
        layer5[25][47:40] = buffer_data_1[2783:2776];
        layer5[25][55:48] = buffer_data_1[2791:2784];
        layer6[25][7:0] = buffer_data_0[2743:2736];
        layer6[25][15:8] = buffer_data_0[2751:2744];
        layer6[25][23:16] = buffer_data_0[2759:2752];
        layer6[25][31:24] = buffer_data_0[2767:2760];
        layer6[25][39:32] = buffer_data_0[2775:2768];
        layer6[25][47:40] = buffer_data_0[2783:2776];
        layer6[25][55:48] = buffer_data_0[2791:2784];
        layer0[26][7:0] = buffer_data_6[2751:2744];
        layer0[26][15:8] = buffer_data_6[2759:2752];
        layer0[26][23:16] = buffer_data_6[2767:2760];
        layer0[26][31:24] = buffer_data_6[2775:2768];
        layer0[26][39:32] = buffer_data_6[2783:2776];
        layer0[26][47:40] = buffer_data_6[2791:2784];
        layer0[26][55:48] = buffer_data_6[2799:2792];
        layer1[26][7:0] = buffer_data_5[2751:2744];
        layer1[26][15:8] = buffer_data_5[2759:2752];
        layer1[26][23:16] = buffer_data_5[2767:2760];
        layer1[26][31:24] = buffer_data_5[2775:2768];
        layer1[26][39:32] = buffer_data_5[2783:2776];
        layer1[26][47:40] = buffer_data_5[2791:2784];
        layer1[26][55:48] = buffer_data_5[2799:2792];
        layer2[26][7:0] = buffer_data_4[2751:2744];
        layer2[26][15:8] = buffer_data_4[2759:2752];
        layer2[26][23:16] = buffer_data_4[2767:2760];
        layer2[26][31:24] = buffer_data_4[2775:2768];
        layer2[26][39:32] = buffer_data_4[2783:2776];
        layer2[26][47:40] = buffer_data_4[2791:2784];
        layer2[26][55:48] = buffer_data_4[2799:2792];
        layer3[26][7:0] = buffer_data_3[2751:2744];
        layer3[26][15:8] = buffer_data_3[2759:2752];
        layer3[26][23:16] = buffer_data_3[2767:2760];
        layer3[26][31:24] = buffer_data_3[2775:2768];
        layer3[26][39:32] = buffer_data_3[2783:2776];
        layer3[26][47:40] = buffer_data_3[2791:2784];
        layer3[26][55:48] = buffer_data_3[2799:2792];
        layer4[26][7:0] = buffer_data_2[2751:2744];
        layer4[26][15:8] = buffer_data_2[2759:2752];
        layer4[26][23:16] = buffer_data_2[2767:2760];
        layer4[26][31:24] = buffer_data_2[2775:2768];
        layer4[26][39:32] = buffer_data_2[2783:2776];
        layer4[26][47:40] = buffer_data_2[2791:2784];
        layer4[26][55:48] = buffer_data_2[2799:2792];
        layer5[26][7:0] = buffer_data_1[2751:2744];
        layer5[26][15:8] = buffer_data_1[2759:2752];
        layer5[26][23:16] = buffer_data_1[2767:2760];
        layer5[26][31:24] = buffer_data_1[2775:2768];
        layer5[26][39:32] = buffer_data_1[2783:2776];
        layer5[26][47:40] = buffer_data_1[2791:2784];
        layer5[26][55:48] = buffer_data_1[2799:2792];
        layer6[26][7:0] = buffer_data_0[2751:2744];
        layer6[26][15:8] = buffer_data_0[2759:2752];
        layer6[26][23:16] = buffer_data_0[2767:2760];
        layer6[26][31:24] = buffer_data_0[2775:2768];
        layer6[26][39:32] = buffer_data_0[2783:2776];
        layer6[26][47:40] = buffer_data_0[2791:2784];
        layer6[26][55:48] = buffer_data_0[2799:2792];
        layer0[27][7:0] = buffer_data_6[2759:2752];
        layer0[27][15:8] = buffer_data_6[2767:2760];
        layer0[27][23:16] = buffer_data_6[2775:2768];
        layer0[27][31:24] = buffer_data_6[2783:2776];
        layer0[27][39:32] = buffer_data_6[2791:2784];
        layer0[27][47:40] = buffer_data_6[2799:2792];
        layer0[27][55:48] = buffer_data_6[2807:2800];
        layer1[27][7:0] = buffer_data_5[2759:2752];
        layer1[27][15:8] = buffer_data_5[2767:2760];
        layer1[27][23:16] = buffer_data_5[2775:2768];
        layer1[27][31:24] = buffer_data_5[2783:2776];
        layer1[27][39:32] = buffer_data_5[2791:2784];
        layer1[27][47:40] = buffer_data_5[2799:2792];
        layer1[27][55:48] = buffer_data_5[2807:2800];
        layer2[27][7:0] = buffer_data_4[2759:2752];
        layer2[27][15:8] = buffer_data_4[2767:2760];
        layer2[27][23:16] = buffer_data_4[2775:2768];
        layer2[27][31:24] = buffer_data_4[2783:2776];
        layer2[27][39:32] = buffer_data_4[2791:2784];
        layer2[27][47:40] = buffer_data_4[2799:2792];
        layer2[27][55:48] = buffer_data_4[2807:2800];
        layer3[27][7:0] = buffer_data_3[2759:2752];
        layer3[27][15:8] = buffer_data_3[2767:2760];
        layer3[27][23:16] = buffer_data_3[2775:2768];
        layer3[27][31:24] = buffer_data_3[2783:2776];
        layer3[27][39:32] = buffer_data_3[2791:2784];
        layer3[27][47:40] = buffer_data_3[2799:2792];
        layer3[27][55:48] = buffer_data_3[2807:2800];
        layer4[27][7:0] = buffer_data_2[2759:2752];
        layer4[27][15:8] = buffer_data_2[2767:2760];
        layer4[27][23:16] = buffer_data_2[2775:2768];
        layer4[27][31:24] = buffer_data_2[2783:2776];
        layer4[27][39:32] = buffer_data_2[2791:2784];
        layer4[27][47:40] = buffer_data_2[2799:2792];
        layer4[27][55:48] = buffer_data_2[2807:2800];
        layer5[27][7:0] = buffer_data_1[2759:2752];
        layer5[27][15:8] = buffer_data_1[2767:2760];
        layer5[27][23:16] = buffer_data_1[2775:2768];
        layer5[27][31:24] = buffer_data_1[2783:2776];
        layer5[27][39:32] = buffer_data_1[2791:2784];
        layer5[27][47:40] = buffer_data_1[2799:2792];
        layer5[27][55:48] = buffer_data_1[2807:2800];
        layer6[27][7:0] = buffer_data_0[2759:2752];
        layer6[27][15:8] = buffer_data_0[2767:2760];
        layer6[27][23:16] = buffer_data_0[2775:2768];
        layer6[27][31:24] = buffer_data_0[2783:2776];
        layer6[27][39:32] = buffer_data_0[2791:2784];
        layer6[27][47:40] = buffer_data_0[2799:2792];
        layer6[27][55:48] = buffer_data_0[2807:2800];
        layer0[28][7:0] = buffer_data_6[2767:2760];
        layer0[28][15:8] = buffer_data_6[2775:2768];
        layer0[28][23:16] = buffer_data_6[2783:2776];
        layer0[28][31:24] = buffer_data_6[2791:2784];
        layer0[28][39:32] = buffer_data_6[2799:2792];
        layer0[28][47:40] = buffer_data_6[2807:2800];
        layer0[28][55:48] = buffer_data_6[2815:2808];
        layer1[28][7:0] = buffer_data_5[2767:2760];
        layer1[28][15:8] = buffer_data_5[2775:2768];
        layer1[28][23:16] = buffer_data_5[2783:2776];
        layer1[28][31:24] = buffer_data_5[2791:2784];
        layer1[28][39:32] = buffer_data_5[2799:2792];
        layer1[28][47:40] = buffer_data_5[2807:2800];
        layer1[28][55:48] = buffer_data_5[2815:2808];
        layer2[28][7:0] = buffer_data_4[2767:2760];
        layer2[28][15:8] = buffer_data_4[2775:2768];
        layer2[28][23:16] = buffer_data_4[2783:2776];
        layer2[28][31:24] = buffer_data_4[2791:2784];
        layer2[28][39:32] = buffer_data_4[2799:2792];
        layer2[28][47:40] = buffer_data_4[2807:2800];
        layer2[28][55:48] = buffer_data_4[2815:2808];
        layer3[28][7:0] = buffer_data_3[2767:2760];
        layer3[28][15:8] = buffer_data_3[2775:2768];
        layer3[28][23:16] = buffer_data_3[2783:2776];
        layer3[28][31:24] = buffer_data_3[2791:2784];
        layer3[28][39:32] = buffer_data_3[2799:2792];
        layer3[28][47:40] = buffer_data_3[2807:2800];
        layer3[28][55:48] = buffer_data_3[2815:2808];
        layer4[28][7:0] = buffer_data_2[2767:2760];
        layer4[28][15:8] = buffer_data_2[2775:2768];
        layer4[28][23:16] = buffer_data_2[2783:2776];
        layer4[28][31:24] = buffer_data_2[2791:2784];
        layer4[28][39:32] = buffer_data_2[2799:2792];
        layer4[28][47:40] = buffer_data_2[2807:2800];
        layer4[28][55:48] = buffer_data_2[2815:2808];
        layer5[28][7:0] = buffer_data_1[2767:2760];
        layer5[28][15:8] = buffer_data_1[2775:2768];
        layer5[28][23:16] = buffer_data_1[2783:2776];
        layer5[28][31:24] = buffer_data_1[2791:2784];
        layer5[28][39:32] = buffer_data_1[2799:2792];
        layer5[28][47:40] = buffer_data_1[2807:2800];
        layer5[28][55:48] = buffer_data_1[2815:2808];
        layer6[28][7:0] = buffer_data_0[2767:2760];
        layer6[28][15:8] = buffer_data_0[2775:2768];
        layer6[28][23:16] = buffer_data_0[2783:2776];
        layer6[28][31:24] = buffer_data_0[2791:2784];
        layer6[28][39:32] = buffer_data_0[2799:2792];
        layer6[28][47:40] = buffer_data_0[2807:2800];
        layer6[28][55:48] = buffer_data_0[2815:2808];
        layer0[29][7:0] = buffer_data_6[2775:2768];
        layer0[29][15:8] = buffer_data_6[2783:2776];
        layer0[29][23:16] = buffer_data_6[2791:2784];
        layer0[29][31:24] = buffer_data_6[2799:2792];
        layer0[29][39:32] = buffer_data_6[2807:2800];
        layer0[29][47:40] = buffer_data_6[2815:2808];
        layer0[29][55:48] = buffer_data_6[2823:2816];
        layer1[29][7:0] = buffer_data_5[2775:2768];
        layer1[29][15:8] = buffer_data_5[2783:2776];
        layer1[29][23:16] = buffer_data_5[2791:2784];
        layer1[29][31:24] = buffer_data_5[2799:2792];
        layer1[29][39:32] = buffer_data_5[2807:2800];
        layer1[29][47:40] = buffer_data_5[2815:2808];
        layer1[29][55:48] = buffer_data_5[2823:2816];
        layer2[29][7:0] = buffer_data_4[2775:2768];
        layer2[29][15:8] = buffer_data_4[2783:2776];
        layer2[29][23:16] = buffer_data_4[2791:2784];
        layer2[29][31:24] = buffer_data_4[2799:2792];
        layer2[29][39:32] = buffer_data_4[2807:2800];
        layer2[29][47:40] = buffer_data_4[2815:2808];
        layer2[29][55:48] = buffer_data_4[2823:2816];
        layer3[29][7:0] = buffer_data_3[2775:2768];
        layer3[29][15:8] = buffer_data_3[2783:2776];
        layer3[29][23:16] = buffer_data_3[2791:2784];
        layer3[29][31:24] = buffer_data_3[2799:2792];
        layer3[29][39:32] = buffer_data_3[2807:2800];
        layer3[29][47:40] = buffer_data_3[2815:2808];
        layer3[29][55:48] = buffer_data_3[2823:2816];
        layer4[29][7:0] = buffer_data_2[2775:2768];
        layer4[29][15:8] = buffer_data_2[2783:2776];
        layer4[29][23:16] = buffer_data_2[2791:2784];
        layer4[29][31:24] = buffer_data_2[2799:2792];
        layer4[29][39:32] = buffer_data_2[2807:2800];
        layer4[29][47:40] = buffer_data_2[2815:2808];
        layer4[29][55:48] = buffer_data_2[2823:2816];
        layer5[29][7:0] = buffer_data_1[2775:2768];
        layer5[29][15:8] = buffer_data_1[2783:2776];
        layer5[29][23:16] = buffer_data_1[2791:2784];
        layer5[29][31:24] = buffer_data_1[2799:2792];
        layer5[29][39:32] = buffer_data_1[2807:2800];
        layer5[29][47:40] = buffer_data_1[2815:2808];
        layer5[29][55:48] = buffer_data_1[2823:2816];
        layer6[29][7:0] = buffer_data_0[2775:2768];
        layer6[29][15:8] = buffer_data_0[2783:2776];
        layer6[29][23:16] = buffer_data_0[2791:2784];
        layer6[29][31:24] = buffer_data_0[2799:2792];
        layer6[29][39:32] = buffer_data_0[2807:2800];
        layer6[29][47:40] = buffer_data_0[2815:2808];
        layer6[29][55:48] = buffer_data_0[2823:2816];
        layer0[30][7:0] = buffer_data_6[2783:2776];
        layer0[30][15:8] = buffer_data_6[2791:2784];
        layer0[30][23:16] = buffer_data_6[2799:2792];
        layer0[30][31:24] = buffer_data_6[2807:2800];
        layer0[30][39:32] = buffer_data_6[2815:2808];
        layer0[30][47:40] = buffer_data_6[2823:2816];
        layer0[30][55:48] = buffer_data_6[2831:2824];
        layer1[30][7:0] = buffer_data_5[2783:2776];
        layer1[30][15:8] = buffer_data_5[2791:2784];
        layer1[30][23:16] = buffer_data_5[2799:2792];
        layer1[30][31:24] = buffer_data_5[2807:2800];
        layer1[30][39:32] = buffer_data_5[2815:2808];
        layer1[30][47:40] = buffer_data_5[2823:2816];
        layer1[30][55:48] = buffer_data_5[2831:2824];
        layer2[30][7:0] = buffer_data_4[2783:2776];
        layer2[30][15:8] = buffer_data_4[2791:2784];
        layer2[30][23:16] = buffer_data_4[2799:2792];
        layer2[30][31:24] = buffer_data_4[2807:2800];
        layer2[30][39:32] = buffer_data_4[2815:2808];
        layer2[30][47:40] = buffer_data_4[2823:2816];
        layer2[30][55:48] = buffer_data_4[2831:2824];
        layer3[30][7:0] = buffer_data_3[2783:2776];
        layer3[30][15:8] = buffer_data_3[2791:2784];
        layer3[30][23:16] = buffer_data_3[2799:2792];
        layer3[30][31:24] = buffer_data_3[2807:2800];
        layer3[30][39:32] = buffer_data_3[2815:2808];
        layer3[30][47:40] = buffer_data_3[2823:2816];
        layer3[30][55:48] = buffer_data_3[2831:2824];
        layer4[30][7:0] = buffer_data_2[2783:2776];
        layer4[30][15:8] = buffer_data_2[2791:2784];
        layer4[30][23:16] = buffer_data_2[2799:2792];
        layer4[30][31:24] = buffer_data_2[2807:2800];
        layer4[30][39:32] = buffer_data_2[2815:2808];
        layer4[30][47:40] = buffer_data_2[2823:2816];
        layer4[30][55:48] = buffer_data_2[2831:2824];
        layer5[30][7:0] = buffer_data_1[2783:2776];
        layer5[30][15:8] = buffer_data_1[2791:2784];
        layer5[30][23:16] = buffer_data_1[2799:2792];
        layer5[30][31:24] = buffer_data_1[2807:2800];
        layer5[30][39:32] = buffer_data_1[2815:2808];
        layer5[30][47:40] = buffer_data_1[2823:2816];
        layer5[30][55:48] = buffer_data_1[2831:2824];
        layer6[30][7:0] = buffer_data_0[2783:2776];
        layer6[30][15:8] = buffer_data_0[2791:2784];
        layer6[30][23:16] = buffer_data_0[2799:2792];
        layer6[30][31:24] = buffer_data_0[2807:2800];
        layer6[30][39:32] = buffer_data_0[2815:2808];
        layer6[30][47:40] = buffer_data_0[2823:2816];
        layer6[30][55:48] = buffer_data_0[2831:2824];
        layer0[31][7:0] = buffer_data_6[2791:2784];
        layer0[31][15:8] = buffer_data_6[2799:2792];
        layer0[31][23:16] = buffer_data_6[2807:2800];
        layer0[31][31:24] = buffer_data_6[2815:2808];
        layer0[31][39:32] = buffer_data_6[2823:2816];
        layer0[31][47:40] = buffer_data_6[2831:2824];
        layer0[31][55:48] = buffer_data_6[2839:2832];
        layer1[31][7:0] = buffer_data_5[2791:2784];
        layer1[31][15:8] = buffer_data_5[2799:2792];
        layer1[31][23:16] = buffer_data_5[2807:2800];
        layer1[31][31:24] = buffer_data_5[2815:2808];
        layer1[31][39:32] = buffer_data_5[2823:2816];
        layer1[31][47:40] = buffer_data_5[2831:2824];
        layer1[31][55:48] = buffer_data_5[2839:2832];
        layer2[31][7:0] = buffer_data_4[2791:2784];
        layer2[31][15:8] = buffer_data_4[2799:2792];
        layer2[31][23:16] = buffer_data_4[2807:2800];
        layer2[31][31:24] = buffer_data_4[2815:2808];
        layer2[31][39:32] = buffer_data_4[2823:2816];
        layer2[31][47:40] = buffer_data_4[2831:2824];
        layer2[31][55:48] = buffer_data_4[2839:2832];
        layer3[31][7:0] = buffer_data_3[2791:2784];
        layer3[31][15:8] = buffer_data_3[2799:2792];
        layer3[31][23:16] = buffer_data_3[2807:2800];
        layer3[31][31:24] = buffer_data_3[2815:2808];
        layer3[31][39:32] = buffer_data_3[2823:2816];
        layer3[31][47:40] = buffer_data_3[2831:2824];
        layer3[31][55:48] = buffer_data_3[2839:2832];
        layer4[31][7:0] = buffer_data_2[2791:2784];
        layer4[31][15:8] = buffer_data_2[2799:2792];
        layer4[31][23:16] = buffer_data_2[2807:2800];
        layer4[31][31:24] = buffer_data_2[2815:2808];
        layer4[31][39:32] = buffer_data_2[2823:2816];
        layer4[31][47:40] = buffer_data_2[2831:2824];
        layer4[31][55:48] = buffer_data_2[2839:2832];
        layer5[31][7:0] = buffer_data_1[2791:2784];
        layer5[31][15:8] = buffer_data_1[2799:2792];
        layer5[31][23:16] = buffer_data_1[2807:2800];
        layer5[31][31:24] = buffer_data_1[2815:2808];
        layer5[31][39:32] = buffer_data_1[2823:2816];
        layer5[31][47:40] = buffer_data_1[2831:2824];
        layer5[31][55:48] = buffer_data_1[2839:2832];
        layer6[31][7:0] = buffer_data_0[2791:2784];
        layer6[31][15:8] = buffer_data_0[2799:2792];
        layer6[31][23:16] = buffer_data_0[2807:2800];
        layer6[31][31:24] = buffer_data_0[2815:2808];
        layer6[31][39:32] = buffer_data_0[2823:2816];
        layer6[31][47:40] = buffer_data_0[2831:2824];
        layer6[31][55:48] = buffer_data_0[2839:2832];
        layer0[32][7:0] = buffer_data_6[2799:2792];
        layer0[32][15:8] = buffer_data_6[2807:2800];
        layer0[32][23:16] = buffer_data_6[2815:2808];
        layer0[32][31:24] = buffer_data_6[2823:2816];
        layer0[32][39:32] = buffer_data_6[2831:2824];
        layer0[32][47:40] = buffer_data_6[2839:2832];
        layer0[32][55:48] = buffer_data_6[2847:2840];
        layer1[32][7:0] = buffer_data_5[2799:2792];
        layer1[32][15:8] = buffer_data_5[2807:2800];
        layer1[32][23:16] = buffer_data_5[2815:2808];
        layer1[32][31:24] = buffer_data_5[2823:2816];
        layer1[32][39:32] = buffer_data_5[2831:2824];
        layer1[32][47:40] = buffer_data_5[2839:2832];
        layer1[32][55:48] = buffer_data_5[2847:2840];
        layer2[32][7:0] = buffer_data_4[2799:2792];
        layer2[32][15:8] = buffer_data_4[2807:2800];
        layer2[32][23:16] = buffer_data_4[2815:2808];
        layer2[32][31:24] = buffer_data_4[2823:2816];
        layer2[32][39:32] = buffer_data_4[2831:2824];
        layer2[32][47:40] = buffer_data_4[2839:2832];
        layer2[32][55:48] = buffer_data_4[2847:2840];
        layer3[32][7:0] = buffer_data_3[2799:2792];
        layer3[32][15:8] = buffer_data_3[2807:2800];
        layer3[32][23:16] = buffer_data_3[2815:2808];
        layer3[32][31:24] = buffer_data_3[2823:2816];
        layer3[32][39:32] = buffer_data_3[2831:2824];
        layer3[32][47:40] = buffer_data_3[2839:2832];
        layer3[32][55:48] = buffer_data_3[2847:2840];
        layer4[32][7:0] = buffer_data_2[2799:2792];
        layer4[32][15:8] = buffer_data_2[2807:2800];
        layer4[32][23:16] = buffer_data_2[2815:2808];
        layer4[32][31:24] = buffer_data_2[2823:2816];
        layer4[32][39:32] = buffer_data_2[2831:2824];
        layer4[32][47:40] = buffer_data_2[2839:2832];
        layer4[32][55:48] = buffer_data_2[2847:2840];
        layer5[32][7:0] = buffer_data_1[2799:2792];
        layer5[32][15:8] = buffer_data_1[2807:2800];
        layer5[32][23:16] = buffer_data_1[2815:2808];
        layer5[32][31:24] = buffer_data_1[2823:2816];
        layer5[32][39:32] = buffer_data_1[2831:2824];
        layer5[32][47:40] = buffer_data_1[2839:2832];
        layer5[32][55:48] = buffer_data_1[2847:2840];
        layer6[32][7:0] = buffer_data_0[2799:2792];
        layer6[32][15:8] = buffer_data_0[2807:2800];
        layer6[32][23:16] = buffer_data_0[2815:2808];
        layer6[32][31:24] = buffer_data_0[2823:2816];
        layer6[32][39:32] = buffer_data_0[2831:2824];
        layer6[32][47:40] = buffer_data_0[2839:2832];
        layer6[32][55:48] = buffer_data_0[2847:2840];
        layer0[33][7:0] = buffer_data_6[2807:2800];
        layer0[33][15:8] = buffer_data_6[2815:2808];
        layer0[33][23:16] = buffer_data_6[2823:2816];
        layer0[33][31:24] = buffer_data_6[2831:2824];
        layer0[33][39:32] = buffer_data_6[2839:2832];
        layer0[33][47:40] = buffer_data_6[2847:2840];
        layer0[33][55:48] = buffer_data_6[2855:2848];
        layer1[33][7:0] = buffer_data_5[2807:2800];
        layer1[33][15:8] = buffer_data_5[2815:2808];
        layer1[33][23:16] = buffer_data_5[2823:2816];
        layer1[33][31:24] = buffer_data_5[2831:2824];
        layer1[33][39:32] = buffer_data_5[2839:2832];
        layer1[33][47:40] = buffer_data_5[2847:2840];
        layer1[33][55:48] = buffer_data_5[2855:2848];
        layer2[33][7:0] = buffer_data_4[2807:2800];
        layer2[33][15:8] = buffer_data_4[2815:2808];
        layer2[33][23:16] = buffer_data_4[2823:2816];
        layer2[33][31:24] = buffer_data_4[2831:2824];
        layer2[33][39:32] = buffer_data_4[2839:2832];
        layer2[33][47:40] = buffer_data_4[2847:2840];
        layer2[33][55:48] = buffer_data_4[2855:2848];
        layer3[33][7:0] = buffer_data_3[2807:2800];
        layer3[33][15:8] = buffer_data_3[2815:2808];
        layer3[33][23:16] = buffer_data_3[2823:2816];
        layer3[33][31:24] = buffer_data_3[2831:2824];
        layer3[33][39:32] = buffer_data_3[2839:2832];
        layer3[33][47:40] = buffer_data_3[2847:2840];
        layer3[33][55:48] = buffer_data_3[2855:2848];
        layer4[33][7:0] = buffer_data_2[2807:2800];
        layer4[33][15:8] = buffer_data_2[2815:2808];
        layer4[33][23:16] = buffer_data_2[2823:2816];
        layer4[33][31:24] = buffer_data_2[2831:2824];
        layer4[33][39:32] = buffer_data_2[2839:2832];
        layer4[33][47:40] = buffer_data_2[2847:2840];
        layer4[33][55:48] = buffer_data_2[2855:2848];
        layer5[33][7:0] = buffer_data_1[2807:2800];
        layer5[33][15:8] = buffer_data_1[2815:2808];
        layer5[33][23:16] = buffer_data_1[2823:2816];
        layer5[33][31:24] = buffer_data_1[2831:2824];
        layer5[33][39:32] = buffer_data_1[2839:2832];
        layer5[33][47:40] = buffer_data_1[2847:2840];
        layer5[33][55:48] = buffer_data_1[2855:2848];
        layer6[33][7:0] = buffer_data_0[2807:2800];
        layer6[33][15:8] = buffer_data_0[2815:2808];
        layer6[33][23:16] = buffer_data_0[2823:2816];
        layer6[33][31:24] = buffer_data_0[2831:2824];
        layer6[33][39:32] = buffer_data_0[2839:2832];
        layer6[33][47:40] = buffer_data_0[2847:2840];
        layer6[33][55:48] = buffer_data_0[2855:2848];
        layer0[34][7:0] = buffer_data_6[2815:2808];
        layer0[34][15:8] = buffer_data_6[2823:2816];
        layer0[34][23:16] = buffer_data_6[2831:2824];
        layer0[34][31:24] = buffer_data_6[2839:2832];
        layer0[34][39:32] = buffer_data_6[2847:2840];
        layer0[34][47:40] = buffer_data_6[2855:2848];
        layer0[34][55:48] = buffer_data_6[2863:2856];
        layer1[34][7:0] = buffer_data_5[2815:2808];
        layer1[34][15:8] = buffer_data_5[2823:2816];
        layer1[34][23:16] = buffer_data_5[2831:2824];
        layer1[34][31:24] = buffer_data_5[2839:2832];
        layer1[34][39:32] = buffer_data_5[2847:2840];
        layer1[34][47:40] = buffer_data_5[2855:2848];
        layer1[34][55:48] = buffer_data_5[2863:2856];
        layer2[34][7:0] = buffer_data_4[2815:2808];
        layer2[34][15:8] = buffer_data_4[2823:2816];
        layer2[34][23:16] = buffer_data_4[2831:2824];
        layer2[34][31:24] = buffer_data_4[2839:2832];
        layer2[34][39:32] = buffer_data_4[2847:2840];
        layer2[34][47:40] = buffer_data_4[2855:2848];
        layer2[34][55:48] = buffer_data_4[2863:2856];
        layer3[34][7:0] = buffer_data_3[2815:2808];
        layer3[34][15:8] = buffer_data_3[2823:2816];
        layer3[34][23:16] = buffer_data_3[2831:2824];
        layer3[34][31:24] = buffer_data_3[2839:2832];
        layer3[34][39:32] = buffer_data_3[2847:2840];
        layer3[34][47:40] = buffer_data_3[2855:2848];
        layer3[34][55:48] = buffer_data_3[2863:2856];
        layer4[34][7:0] = buffer_data_2[2815:2808];
        layer4[34][15:8] = buffer_data_2[2823:2816];
        layer4[34][23:16] = buffer_data_2[2831:2824];
        layer4[34][31:24] = buffer_data_2[2839:2832];
        layer4[34][39:32] = buffer_data_2[2847:2840];
        layer4[34][47:40] = buffer_data_2[2855:2848];
        layer4[34][55:48] = buffer_data_2[2863:2856];
        layer5[34][7:0] = buffer_data_1[2815:2808];
        layer5[34][15:8] = buffer_data_1[2823:2816];
        layer5[34][23:16] = buffer_data_1[2831:2824];
        layer5[34][31:24] = buffer_data_1[2839:2832];
        layer5[34][39:32] = buffer_data_1[2847:2840];
        layer5[34][47:40] = buffer_data_1[2855:2848];
        layer5[34][55:48] = buffer_data_1[2863:2856];
        layer6[34][7:0] = buffer_data_0[2815:2808];
        layer6[34][15:8] = buffer_data_0[2823:2816];
        layer6[34][23:16] = buffer_data_0[2831:2824];
        layer6[34][31:24] = buffer_data_0[2839:2832];
        layer6[34][39:32] = buffer_data_0[2847:2840];
        layer6[34][47:40] = buffer_data_0[2855:2848];
        layer6[34][55:48] = buffer_data_0[2863:2856];
        layer0[35][7:0] = buffer_data_6[2823:2816];
        layer0[35][15:8] = buffer_data_6[2831:2824];
        layer0[35][23:16] = buffer_data_6[2839:2832];
        layer0[35][31:24] = buffer_data_6[2847:2840];
        layer0[35][39:32] = buffer_data_6[2855:2848];
        layer0[35][47:40] = buffer_data_6[2863:2856];
        layer0[35][55:48] = buffer_data_6[2871:2864];
        layer1[35][7:0] = buffer_data_5[2823:2816];
        layer1[35][15:8] = buffer_data_5[2831:2824];
        layer1[35][23:16] = buffer_data_5[2839:2832];
        layer1[35][31:24] = buffer_data_5[2847:2840];
        layer1[35][39:32] = buffer_data_5[2855:2848];
        layer1[35][47:40] = buffer_data_5[2863:2856];
        layer1[35][55:48] = buffer_data_5[2871:2864];
        layer2[35][7:0] = buffer_data_4[2823:2816];
        layer2[35][15:8] = buffer_data_4[2831:2824];
        layer2[35][23:16] = buffer_data_4[2839:2832];
        layer2[35][31:24] = buffer_data_4[2847:2840];
        layer2[35][39:32] = buffer_data_4[2855:2848];
        layer2[35][47:40] = buffer_data_4[2863:2856];
        layer2[35][55:48] = buffer_data_4[2871:2864];
        layer3[35][7:0] = buffer_data_3[2823:2816];
        layer3[35][15:8] = buffer_data_3[2831:2824];
        layer3[35][23:16] = buffer_data_3[2839:2832];
        layer3[35][31:24] = buffer_data_3[2847:2840];
        layer3[35][39:32] = buffer_data_3[2855:2848];
        layer3[35][47:40] = buffer_data_3[2863:2856];
        layer3[35][55:48] = buffer_data_3[2871:2864];
        layer4[35][7:0] = buffer_data_2[2823:2816];
        layer4[35][15:8] = buffer_data_2[2831:2824];
        layer4[35][23:16] = buffer_data_2[2839:2832];
        layer4[35][31:24] = buffer_data_2[2847:2840];
        layer4[35][39:32] = buffer_data_2[2855:2848];
        layer4[35][47:40] = buffer_data_2[2863:2856];
        layer4[35][55:48] = buffer_data_2[2871:2864];
        layer5[35][7:0] = buffer_data_1[2823:2816];
        layer5[35][15:8] = buffer_data_1[2831:2824];
        layer5[35][23:16] = buffer_data_1[2839:2832];
        layer5[35][31:24] = buffer_data_1[2847:2840];
        layer5[35][39:32] = buffer_data_1[2855:2848];
        layer5[35][47:40] = buffer_data_1[2863:2856];
        layer5[35][55:48] = buffer_data_1[2871:2864];
        layer6[35][7:0] = buffer_data_0[2823:2816];
        layer6[35][15:8] = buffer_data_0[2831:2824];
        layer6[35][23:16] = buffer_data_0[2839:2832];
        layer6[35][31:24] = buffer_data_0[2847:2840];
        layer6[35][39:32] = buffer_data_0[2855:2848];
        layer6[35][47:40] = buffer_data_0[2863:2856];
        layer6[35][55:48] = buffer_data_0[2871:2864];
        layer0[36][7:0] = buffer_data_6[2831:2824];
        layer0[36][15:8] = buffer_data_6[2839:2832];
        layer0[36][23:16] = buffer_data_6[2847:2840];
        layer0[36][31:24] = buffer_data_6[2855:2848];
        layer0[36][39:32] = buffer_data_6[2863:2856];
        layer0[36][47:40] = buffer_data_6[2871:2864];
        layer0[36][55:48] = buffer_data_6[2879:2872];
        layer1[36][7:0] = buffer_data_5[2831:2824];
        layer1[36][15:8] = buffer_data_5[2839:2832];
        layer1[36][23:16] = buffer_data_5[2847:2840];
        layer1[36][31:24] = buffer_data_5[2855:2848];
        layer1[36][39:32] = buffer_data_5[2863:2856];
        layer1[36][47:40] = buffer_data_5[2871:2864];
        layer1[36][55:48] = buffer_data_5[2879:2872];
        layer2[36][7:0] = buffer_data_4[2831:2824];
        layer2[36][15:8] = buffer_data_4[2839:2832];
        layer2[36][23:16] = buffer_data_4[2847:2840];
        layer2[36][31:24] = buffer_data_4[2855:2848];
        layer2[36][39:32] = buffer_data_4[2863:2856];
        layer2[36][47:40] = buffer_data_4[2871:2864];
        layer2[36][55:48] = buffer_data_4[2879:2872];
        layer3[36][7:0] = buffer_data_3[2831:2824];
        layer3[36][15:8] = buffer_data_3[2839:2832];
        layer3[36][23:16] = buffer_data_3[2847:2840];
        layer3[36][31:24] = buffer_data_3[2855:2848];
        layer3[36][39:32] = buffer_data_3[2863:2856];
        layer3[36][47:40] = buffer_data_3[2871:2864];
        layer3[36][55:48] = buffer_data_3[2879:2872];
        layer4[36][7:0] = buffer_data_2[2831:2824];
        layer4[36][15:8] = buffer_data_2[2839:2832];
        layer4[36][23:16] = buffer_data_2[2847:2840];
        layer4[36][31:24] = buffer_data_2[2855:2848];
        layer4[36][39:32] = buffer_data_2[2863:2856];
        layer4[36][47:40] = buffer_data_2[2871:2864];
        layer4[36][55:48] = buffer_data_2[2879:2872];
        layer5[36][7:0] = buffer_data_1[2831:2824];
        layer5[36][15:8] = buffer_data_1[2839:2832];
        layer5[36][23:16] = buffer_data_1[2847:2840];
        layer5[36][31:24] = buffer_data_1[2855:2848];
        layer5[36][39:32] = buffer_data_1[2863:2856];
        layer5[36][47:40] = buffer_data_1[2871:2864];
        layer5[36][55:48] = buffer_data_1[2879:2872];
        layer6[36][7:0] = buffer_data_0[2831:2824];
        layer6[36][15:8] = buffer_data_0[2839:2832];
        layer6[36][23:16] = buffer_data_0[2847:2840];
        layer6[36][31:24] = buffer_data_0[2855:2848];
        layer6[36][39:32] = buffer_data_0[2863:2856];
        layer6[36][47:40] = buffer_data_0[2871:2864];
        layer6[36][55:48] = buffer_data_0[2879:2872];
        layer0[37][7:0] = buffer_data_6[2839:2832];
        layer0[37][15:8] = buffer_data_6[2847:2840];
        layer0[37][23:16] = buffer_data_6[2855:2848];
        layer0[37][31:24] = buffer_data_6[2863:2856];
        layer0[37][39:32] = buffer_data_6[2871:2864];
        layer0[37][47:40] = buffer_data_6[2879:2872];
        layer0[37][55:48] = buffer_data_6[2887:2880];
        layer1[37][7:0] = buffer_data_5[2839:2832];
        layer1[37][15:8] = buffer_data_5[2847:2840];
        layer1[37][23:16] = buffer_data_5[2855:2848];
        layer1[37][31:24] = buffer_data_5[2863:2856];
        layer1[37][39:32] = buffer_data_5[2871:2864];
        layer1[37][47:40] = buffer_data_5[2879:2872];
        layer1[37][55:48] = buffer_data_5[2887:2880];
        layer2[37][7:0] = buffer_data_4[2839:2832];
        layer2[37][15:8] = buffer_data_4[2847:2840];
        layer2[37][23:16] = buffer_data_4[2855:2848];
        layer2[37][31:24] = buffer_data_4[2863:2856];
        layer2[37][39:32] = buffer_data_4[2871:2864];
        layer2[37][47:40] = buffer_data_4[2879:2872];
        layer2[37][55:48] = buffer_data_4[2887:2880];
        layer3[37][7:0] = buffer_data_3[2839:2832];
        layer3[37][15:8] = buffer_data_3[2847:2840];
        layer3[37][23:16] = buffer_data_3[2855:2848];
        layer3[37][31:24] = buffer_data_3[2863:2856];
        layer3[37][39:32] = buffer_data_3[2871:2864];
        layer3[37][47:40] = buffer_data_3[2879:2872];
        layer3[37][55:48] = buffer_data_3[2887:2880];
        layer4[37][7:0] = buffer_data_2[2839:2832];
        layer4[37][15:8] = buffer_data_2[2847:2840];
        layer4[37][23:16] = buffer_data_2[2855:2848];
        layer4[37][31:24] = buffer_data_2[2863:2856];
        layer4[37][39:32] = buffer_data_2[2871:2864];
        layer4[37][47:40] = buffer_data_2[2879:2872];
        layer4[37][55:48] = buffer_data_2[2887:2880];
        layer5[37][7:0] = buffer_data_1[2839:2832];
        layer5[37][15:8] = buffer_data_1[2847:2840];
        layer5[37][23:16] = buffer_data_1[2855:2848];
        layer5[37][31:24] = buffer_data_1[2863:2856];
        layer5[37][39:32] = buffer_data_1[2871:2864];
        layer5[37][47:40] = buffer_data_1[2879:2872];
        layer5[37][55:48] = buffer_data_1[2887:2880];
        layer6[37][7:0] = buffer_data_0[2839:2832];
        layer6[37][15:8] = buffer_data_0[2847:2840];
        layer6[37][23:16] = buffer_data_0[2855:2848];
        layer6[37][31:24] = buffer_data_0[2863:2856];
        layer6[37][39:32] = buffer_data_0[2871:2864];
        layer6[37][47:40] = buffer_data_0[2879:2872];
        layer6[37][55:48] = buffer_data_0[2887:2880];
        layer0[38][7:0] = buffer_data_6[2847:2840];
        layer0[38][15:8] = buffer_data_6[2855:2848];
        layer0[38][23:16] = buffer_data_6[2863:2856];
        layer0[38][31:24] = buffer_data_6[2871:2864];
        layer0[38][39:32] = buffer_data_6[2879:2872];
        layer0[38][47:40] = buffer_data_6[2887:2880];
        layer0[38][55:48] = buffer_data_6[2895:2888];
        layer1[38][7:0] = buffer_data_5[2847:2840];
        layer1[38][15:8] = buffer_data_5[2855:2848];
        layer1[38][23:16] = buffer_data_5[2863:2856];
        layer1[38][31:24] = buffer_data_5[2871:2864];
        layer1[38][39:32] = buffer_data_5[2879:2872];
        layer1[38][47:40] = buffer_data_5[2887:2880];
        layer1[38][55:48] = buffer_data_5[2895:2888];
        layer2[38][7:0] = buffer_data_4[2847:2840];
        layer2[38][15:8] = buffer_data_4[2855:2848];
        layer2[38][23:16] = buffer_data_4[2863:2856];
        layer2[38][31:24] = buffer_data_4[2871:2864];
        layer2[38][39:32] = buffer_data_4[2879:2872];
        layer2[38][47:40] = buffer_data_4[2887:2880];
        layer2[38][55:48] = buffer_data_4[2895:2888];
        layer3[38][7:0] = buffer_data_3[2847:2840];
        layer3[38][15:8] = buffer_data_3[2855:2848];
        layer3[38][23:16] = buffer_data_3[2863:2856];
        layer3[38][31:24] = buffer_data_3[2871:2864];
        layer3[38][39:32] = buffer_data_3[2879:2872];
        layer3[38][47:40] = buffer_data_3[2887:2880];
        layer3[38][55:48] = buffer_data_3[2895:2888];
        layer4[38][7:0] = buffer_data_2[2847:2840];
        layer4[38][15:8] = buffer_data_2[2855:2848];
        layer4[38][23:16] = buffer_data_2[2863:2856];
        layer4[38][31:24] = buffer_data_2[2871:2864];
        layer4[38][39:32] = buffer_data_2[2879:2872];
        layer4[38][47:40] = buffer_data_2[2887:2880];
        layer4[38][55:48] = buffer_data_2[2895:2888];
        layer5[38][7:0] = buffer_data_1[2847:2840];
        layer5[38][15:8] = buffer_data_1[2855:2848];
        layer5[38][23:16] = buffer_data_1[2863:2856];
        layer5[38][31:24] = buffer_data_1[2871:2864];
        layer5[38][39:32] = buffer_data_1[2879:2872];
        layer5[38][47:40] = buffer_data_1[2887:2880];
        layer5[38][55:48] = buffer_data_1[2895:2888];
        layer6[38][7:0] = buffer_data_0[2847:2840];
        layer6[38][15:8] = buffer_data_0[2855:2848];
        layer6[38][23:16] = buffer_data_0[2863:2856];
        layer6[38][31:24] = buffer_data_0[2871:2864];
        layer6[38][39:32] = buffer_data_0[2879:2872];
        layer6[38][47:40] = buffer_data_0[2887:2880];
        layer6[38][55:48] = buffer_data_0[2895:2888];
        layer0[39][7:0] = buffer_data_6[2855:2848];
        layer0[39][15:8] = buffer_data_6[2863:2856];
        layer0[39][23:16] = buffer_data_6[2871:2864];
        layer0[39][31:24] = buffer_data_6[2879:2872];
        layer0[39][39:32] = buffer_data_6[2887:2880];
        layer0[39][47:40] = buffer_data_6[2895:2888];
        layer0[39][55:48] = buffer_data_6[2903:2896];
        layer1[39][7:0] = buffer_data_5[2855:2848];
        layer1[39][15:8] = buffer_data_5[2863:2856];
        layer1[39][23:16] = buffer_data_5[2871:2864];
        layer1[39][31:24] = buffer_data_5[2879:2872];
        layer1[39][39:32] = buffer_data_5[2887:2880];
        layer1[39][47:40] = buffer_data_5[2895:2888];
        layer1[39][55:48] = buffer_data_5[2903:2896];
        layer2[39][7:0] = buffer_data_4[2855:2848];
        layer2[39][15:8] = buffer_data_4[2863:2856];
        layer2[39][23:16] = buffer_data_4[2871:2864];
        layer2[39][31:24] = buffer_data_4[2879:2872];
        layer2[39][39:32] = buffer_data_4[2887:2880];
        layer2[39][47:40] = buffer_data_4[2895:2888];
        layer2[39][55:48] = buffer_data_4[2903:2896];
        layer3[39][7:0] = buffer_data_3[2855:2848];
        layer3[39][15:8] = buffer_data_3[2863:2856];
        layer3[39][23:16] = buffer_data_3[2871:2864];
        layer3[39][31:24] = buffer_data_3[2879:2872];
        layer3[39][39:32] = buffer_data_3[2887:2880];
        layer3[39][47:40] = buffer_data_3[2895:2888];
        layer3[39][55:48] = buffer_data_3[2903:2896];
        layer4[39][7:0] = buffer_data_2[2855:2848];
        layer4[39][15:8] = buffer_data_2[2863:2856];
        layer4[39][23:16] = buffer_data_2[2871:2864];
        layer4[39][31:24] = buffer_data_2[2879:2872];
        layer4[39][39:32] = buffer_data_2[2887:2880];
        layer4[39][47:40] = buffer_data_2[2895:2888];
        layer4[39][55:48] = buffer_data_2[2903:2896];
        layer5[39][7:0] = buffer_data_1[2855:2848];
        layer5[39][15:8] = buffer_data_1[2863:2856];
        layer5[39][23:16] = buffer_data_1[2871:2864];
        layer5[39][31:24] = buffer_data_1[2879:2872];
        layer5[39][39:32] = buffer_data_1[2887:2880];
        layer5[39][47:40] = buffer_data_1[2895:2888];
        layer5[39][55:48] = buffer_data_1[2903:2896];
        layer6[39][7:0] = buffer_data_0[2855:2848];
        layer6[39][15:8] = buffer_data_0[2863:2856];
        layer6[39][23:16] = buffer_data_0[2871:2864];
        layer6[39][31:24] = buffer_data_0[2879:2872];
        layer6[39][39:32] = buffer_data_0[2887:2880];
        layer6[39][47:40] = buffer_data_0[2895:2888];
        layer6[39][55:48] = buffer_data_0[2903:2896];
        layer0[40][7:0] = buffer_data_6[2863:2856];
        layer0[40][15:8] = buffer_data_6[2871:2864];
        layer0[40][23:16] = buffer_data_6[2879:2872];
        layer0[40][31:24] = buffer_data_6[2887:2880];
        layer0[40][39:32] = buffer_data_6[2895:2888];
        layer0[40][47:40] = buffer_data_6[2903:2896];
        layer0[40][55:48] = buffer_data_6[2911:2904];
        layer1[40][7:0] = buffer_data_5[2863:2856];
        layer1[40][15:8] = buffer_data_5[2871:2864];
        layer1[40][23:16] = buffer_data_5[2879:2872];
        layer1[40][31:24] = buffer_data_5[2887:2880];
        layer1[40][39:32] = buffer_data_5[2895:2888];
        layer1[40][47:40] = buffer_data_5[2903:2896];
        layer1[40][55:48] = buffer_data_5[2911:2904];
        layer2[40][7:0] = buffer_data_4[2863:2856];
        layer2[40][15:8] = buffer_data_4[2871:2864];
        layer2[40][23:16] = buffer_data_4[2879:2872];
        layer2[40][31:24] = buffer_data_4[2887:2880];
        layer2[40][39:32] = buffer_data_4[2895:2888];
        layer2[40][47:40] = buffer_data_4[2903:2896];
        layer2[40][55:48] = buffer_data_4[2911:2904];
        layer3[40][7:0] = buffer_data_3[2863:2856];
        layer3[40][15:8] = buffer_data_3[2871:2864];
        layer3[40][23:16] = buffer_data_3[2879:2872];
        layer3[40][31:24] = buffer_data_3[2887:2880];
        layer3[40][39:32] = buffer_data_3[2895:2888];
        layer3[40][47:40] = buffer_data_3[2903:2896];
        layer3[40][55:48] = buffer_data_3[2911:2904];
        layer4[40][7:0] = buffer_data_2[2863:2856];
        layer4[40][15:8] = buffer_data_2[2871:2864];
        layer4[40][23:16] = buffer_data_2[2879:2872];
        layer4[40][31:24] = buffer_data_2[2887:2880];
        layer4[40][39:32] = buffer_data_2[2895:2888];
        layer4[40][47:40] = buffer_data_2[2903:2896];
        layer4[40][55:48] = buffer_data_2[2911:2904];
        layer5[40][7:0] = buffer_data_1[2863:2856];
        layer5[40][15:8] = buffer_data_1[2871:2864];
        layer5[40][23:16] = buffer_data_1[2879:2872];
        layer5[40][31:24] = buffer_data_1[2887:2880];
        layer5[40][39:32] = buffer_data_1[2895:2888];
        layer5[40][47:40] = buffer_data_1[2903:2896];
        layer5[40][55:48] = buffer_data_1[2911:2904];
        layer6[40][7:0] = buffer_data_0[2863:2856];
        layer6[40][15:8] = buffer_data_0[2871:2864];
        layer6[40][23:16] = buffer_data_0[2879:2872];
        layer6[40][31:24] = buffer_data_0[2887:2880];
        layer6[40][39:32] = buffer_data_0[2895:2888];
        layer6[40][47:40] = buffer_data_0[2903:2896];
        layer6[40][55:48] = buffer_data_0[2911:2904];
        layer0[41][7:0] = buffer_data_6[2871:2864];
        layer0[41][15:8] = buffer_data_6[2879:2872];
        layer0[41][23:16] = buffer_data_6[2887:2880];
        layer0[41][31:24] = buffer_data_6[2895:2888];
        layer0[41][39:32] = buffer_data_6[2903:2896];
        layer0[41][47:40] = buffer_data_6[2911:2904];
        layer0[41][55:48] = buffer_data_6[2919:2912];
        layer1[41][7:0] = buffer_data_5[2871:2864];
        layer1[41][15:8] = buffer_data_5[2879:2872];
        layer1[41][23:16] = buffer_data_5[2887:2880];
        layer1[41][31:24] = buffer_data_5[2895:2888];
        layer1[41][39:32] = buffer_data_5[2903:2896];
        layer1[41][47:40] = buffer_data_5[2911:2904];
        layer1[41][55:48] = buffer_data_5[2919:2912];
        layer2[41][7:0] = buffer_data_4[2871:2864];
        layer2[41][15:8] = buffer_data_4[2879:2872];
        layer2[41][23:16] = buffer_data_4[2887:2880];
        layer2[41][31:24] = buffer_data_4[2895:2888];
        layer2[41][39:32] = buffer_data_4[2903:2896];
        layer2[41][47:40] = buffer_data_4[2911:2904];
        layer2[41][55:48] = buffer_data_4[2919:2912];
        layer3[41][7:0] = buffer_data_3[2871:2864];
        layer3[41][15:8] = buffer_data_3[2879:2872];
        layer3[41][23:16] = buffer_data_3[2887:2880];
        layer3[41][31:24] = buffer_data_3[2895:2888];
        layer3[41][39:32] = buffer_data_3[2903:2896];
        layer3[41][47:40] = buffer_data_3[2911:2904];
        layer3[41][55:48] = buffer_data_3[2919:2912];
        layer4[41][7:0] = buffer_data_2[2871:2864];
        layer4[41][15:8] = buffer_data_2[2879:2872];
        layer4[41][23:16] = buffer_data_2[2887:2880];
        layer4[41][31:24] = buffer_data_2[2895:2888];
        layer4[41][39:32] = buffer_data_2[2903:2896];
        layer4[41][47:40] = buffer_data_2[2911:2904];
        layer4[41][55:48] = buffer_data_2[2919:2912];
        layer5[41][7:0] = buffer_data_1[2871:2864];
        layer5[41][15:8] = buffer_data_1[2879:2872];
        layer5[41][23:16] = buffer_data_1[2887:2880];
        layer5[41][31:24] = buffer_data_1[2895:2888];
        layer5[41][39:32] = buffer_data_1[2903:2896];
        layer5[41][47:40] = buffer_data_1[2911:2904];
        layer5[41][55:48] = buffer_data_1[2919:2912];
        layer6[41][7:0] = buffer_data_0[2871:2864];
        layer6[41][15:8] = buffer_data_0[2879:2872];
        layer6[41][23:16] = buffer_data_0[2887:2880];
        layer6[41][31:24] = buffer_data_0[2895:2888];
        layer6[41][39:32] = buffer_data_0[2903:2896];
        layer6[41][47:40] = buffer_data_0[2911:2904];
        layer6[41][55:48] = buffer_data_0[2919:2912];
        layer0[42][7:0] = buffer_data_6[2879:2872];
        layer0[42][15:8] = buffer_data_6[2887:2880];
        layer0[42][23:16] = buffer_data_6[2895:2888];
        layer0[42][31:24] = buffer_data_6[2903:2896];
        layer0[42][39:32] = buffer_data_6[2911:2904];
        layer0[42][47:40] = buffer_data_6[2919:2912];
        layer0[42][55:48] = buffer_data_6[2927:2920];
        layer1[42][7:0] = buffer_data_5[2879:2872];
        layer1[42][15:8] = buffer_data_5[2887:2880];
        layer1[42][23:16] = buffer_data_5[2895:2888];
        layer1[42][31:24] = buffer_data_5[2903:2896];
        layer1[42][39:32] = buffer_data_5[2911:2904];
        layer1[42][47:40] = buffer_data_5[2919:2912];
        layer1[42][55:48] = buffer_data_5[2927:2920];
        layer2[42][7:0] = buffer_data_4[2879:2872];
        layer2[42][15:8] = buffer_data_4[2887:2880];
        layer2[42][23:16] = buffer_data_4[2895:2888];
        layer2[42][31:24] = buffer_data_4[2903:2896];
        layer2[42][39:32] = buffer_data_4[2911:2904];
        layer2[42][47:40] = buffer_data_4[2919:2912];
        layer2[42][55:48] = buffer_data_4[2927:2920];
        layer3[42][7:0] = buffer_data_3[2879:2872];
        layer3[42][15:8] = buffer_data_3[2887:2880];
        layer3[42][23:16] = buffer_data_3[2895:2888];
        layer3[42][31:24] = buffer_data_3[2903:2896];
        layer3[42][39:32] = buffer_data_3[2911:2904];
        layer3[42][47:40] = buffer_data_3[2919:2912];
        layer3[42][55:48] = buffer_data_3[2927:2920];
        layer4[42][7:0] = buffer_data_2[2879:2872];
        layer4[42][15:8] = buffer_data_2[2887:2880];
        layer4[42][23:16] = buffer_data_2[2895:2888];
        layer4[42][31:24] = buffer_data_2[2903:2896];
        layer4[42][39:32] = buffer_data_2[2911:2904];
        layer4[42][47:40] = buffer_data_2[2919:2912];
        layer4[42][55:48] = buffer_data_2[2927:2920];
        layer5[42][7:0] = buffer_data_1[2879:2872];
        layer5[42][15:8] = buffer_data_1[2887:2880];
        layer5[42][23:16] = buffer_data_1[2895:2888];
        layer5[42][31:24] = buffer_data_1[2903:2896];
        layer5[42][39:32] = buffer_data_1[2911:2904];
        layer5[42][47:40] = buffer_data_1[2919:2912];
        layer5[42][55:48] = buffer_data_1[2927:2920];
        layer6[42][7:0] = buffer_data_0[2879:2872];
        layer6[42][15:8] = buffer_data_0[2887:2880];
        layer6[42][23:16] = buffer_data_0[2895:2888];
        layer6[42][31:24] = buffer_data_0[2903:2896];
        layer6[42][39:32] = buffer_data_0[2911:2904];
        layer6[42][47:40] = buffer_data_0[2919:2912];
        layer6[42][55:48] = buffer_data_0[2927:2920];
        layer0[43][7:0] = buffer_data_6[2887:2880];
        layer0[43][15:8] = buffer_data_6[2895:2888];
        layer0[43][23:16] = buffer_data_6[2903:2896];
        layer0[43][31:24] = buffer_data_6[2911:2904];
        layer0[43][39:32] = buffer_data_6[2919:2912];
        layer0[43][47:40] = buffer_data_6[2927:2920];
        layer0[43][55:48] = buffer_data_6[2935:2928];
        layer1[43][7:0] = buffer_data_5[2887:2880];
        layer1[43][15:8] = buffer_data_5[2895:2888];
        layer1[43][23:16] = buffer_data_5[2903:2896];
        layer1[43][31:24] = buffer_data_5[2911:2904];
        layer1[43][39:32] = buffer_data_5[2919:2912];
        layer1[43][47:40] = buffer_data_5[2927:2920];
        layer1[43][55:48] = buffer_data_5[2935:2928];
        layer2[43][7:0] = buffer_data_4[2887:2880];
        layer2[43][15:8] = buffer_data_4[2895:2888];
        layer2[43][23:16] = buffer_data_4[2903:2896];
        layer2[43][31:24] = buffer_data_4[2911:2904];
        layer2[43][39:32] = buffer_data_4[2919:2912];
        layer2[43][47:40] = buffer_data_4[2927:2920];
        layer2[43][55:48] = buffer_data_4[2935:2928];
        layer3[43][7:0] = buffer_data_3[2887:2880];
        layer3[43][15:8] = buffer_data_3[2895:2888];
        layer3[43][23:16] = buffer_data_3[2903:2896];
        layer3[43][31:24] = buffer_data_3[2911:2904];
        layer3[43][39:32] = buffer_data_3[2919:2912];
        layer3[43][47:40] = buffer_data_3[2927:2920];
        layer3[43][55:48] = buffer_data_3[2935:2928];
        layer4[43][7:0] = buffer_data_2[2887:2880];
        layer4[43][15:8] = buffer_data_2[2895:2888];
        layer4[43][23:16] = buffer_data_2[2903:2896];
        layer4[43][31:24] = buffer_data_2[2911:2904];
        layer4[43][39:32] = buffer_data_2[2919:2912];
        layer4[43][47:40] = buffer_data_2[2927:2920];
        layer4[43][55:48] = buffer_data_2[2935:2928];
        layer5[43][7:0] = buffer_data_1[2887:2880];
        layer5[43][15:8] = buffer_data_1[2895:2888];
        layer5[43][23:16] = buffer_data_1[2903:2896];
        layer5[43][31:24] = buffer_data_1[2911:2904];
        layer5[43][39:32] = buffer_data_1[2919:2912];
        layer5[43][47:40] = buffer_data_1[2927:2920];
        layer5[43][55:48] = buffer_data_1[2935:2928];
        layer6[43][7:0] = buffer_data_0[2887:2880];
        layer6[43][15:8] = buffer_data_0[2895:2888];
        layer6[43][23:16] = buffer_data_0[2903:2896];
        layer6[43][31:24] = buffer_data_0[2911:2904];
        layer6[43][39:32] = buffer_data_0[2919:2912];
        layer6[43][47:40] = buffer_data_0[2927:2920];
        layer6[43][55:48] = buffer_data_0[2935:2928];
        layer0[44][7:0] = buffer_data_6[2895:2888];
        layer0[44][15:8] = buffer_data_6[2903:2896];
        layer0[44][23:16] = buffer_data_6[2911:2904];
        layer0[44][31:24] = buffer_data_6[2919:2912];
        layer0[44][39:32] = buffer_data_6[2927:2920];
        layer0[44][47:40] = buffer_data_6[2935:2928];
        layer0[44][55:48] = buffer_data_6[2943:2936];
        layer1[44][7:0] = buffer_data_5[2895:2888];
        layer1[44][15:8] = buffer_data_5[2903:2896];
        layer1[44][23:16] = buffer_data_5[2911:2904];
        layer1[44][31:24] = buffer_data_5[2919:2912];
        layer1[44][39:32] = buffer_data_5[2927:2920];
        layer1[44][47:40] = buffer_data_5[2935:2928];
        layer1[44][55:48] = buffer_data_5[2943:2936];
        layer2[44][7:0] = buffer_data_4[2895:2888];
        layer2[44][15:8] = buffer_data_4[2903:2896];
        layer2[44][23:16] = buffer_data_4[2911:2904];
        layer2[44][31:24] = buffer_data_4[2919:2912];
        layer2[44][39:32] = buffer_data_4[2927:2920];
        layer2[44][47:40] = buffer_data_4[2935:2928];
        layer2[44][55:48] = buffer_data_4[2943:2936];
        layer3[44][7:0] = buffer_data_3[2895:2888];
        layer3[44][15:8] = buffer_data_3[2903:2896];
        layer3[44][23:16] = buffer_data_3[2911:2904];
        layer3[44][31:24] = buffer_data_3[2919:2912];
        layer3[44][39:32] = buffer_data_3[2927:2920];
        layer3[44][47:40] = buffer_data_3[2935:2928];
        layer3[44][55:48] = buffer_data_3[2943:2936];
        layer4[44][7:0] = buffer_data_2[2895:2888];
        layer4[44][15:8] = buffer_data_2[2903:2896];
        layer4[44][23:16] = buffer_data_2[2911:2904];
        layer4[44][31:24] = buffer_data_2[2919:2912];
        layer4[44][39:32] = buffer_data_2[2927:2920];
        layer4[44][47:40] = buffer_data_2[2935:2928];
        layer4[44][55:48] = buffer_data_2[2943:2936];
        layer5[44][7:0] = buffer_data_1[2895:2888];
        layer5[44][15:8] = buffer_data_1[2903:2896];
        layer5[44][23:16] = buffer_data_1[2911:2904];
        layer5[44][31:24] = buffer_data_1[2919:2912];
        layer5[44][39:32] = buffer_data_1[2927:2920];
        layer5[44][47:40] = buffer_data_1[2935:2928];
        layer5[44][55:48] = buffer_data_1[2943:2936];
        layer6[44][7:0] = buffer_data_0[2895:2888];
        layer6[44][15:8] = buffer_data_0[2903:2896];
        layer6[44][23:16] = buffer_data_0[2911:2904];
        layer6[44][31:24] = buffer_data_0[2919:2912];
        layer6[44][39:32] = buffer_data_0[2927:2920];
        layer6[44][47:40] = buffer_data_0[2935:2928];
        layer6[44][55:48] = buffer_data_0[2943:2936];
        layer0[45][7:0] = buffer_data_6[2903:2896];
        layer0[45][15:8] = buffer_data_6[2911:2904];
        layer0[45][23:16] = buffer_data_6[2919:2912];
        layer0[45][31:24] = buffer_data_6[2927:2920];
        layer0[45][39:32] = buffer_data_6[2935:2928];
        layer0[45][47:40] = buffer_data_6[2943:2936];
        layer0[45][55:48] = buffer_data_6[2951:2944];
        layer1[45][7:0] = buffer_data_5[2903:2896];
        layer1[45][15:8] = buffer_data_5[2911:2904];
        layer1[45][23:16] = buffer_data_5[2919:2912];
        layer1[45][31:24] = buffer_data_5[2927:2920];
        layer1[45][39:32] = buffer_data_5[2935:2928];
        layer1[45][47:40] = buffer_data_5[2943:2936];
        layer1[45][55:48] = buffer_data_5[2951:2944];
        layer2[45][7:0] = buffer_data_4[2903:2896];
        layer2[45][15:8] = buffer_data_4[2911:2904];
        layer2[45][23:16] = buffer_data_4[2919:2912];
        layer2[45][31:24] = buffer_data_4[2927:2920];
        layer2[45][39:32] = buffer_data_4[2935:2928];
        layer2[45][47:40] = buffer_data_4[2943:2936];
        layer2[45][55:48] = buffer_data_4[2951:2944];
        layer3[45][7:0] = buffer_data_3[2903:2896];
        layer3[45][15:8] = buffer_data_3[2911:2904];
        layer3[45][23:16] = buffer_data_3[2919:2912];
        layer3[45][31:24] = buffer_data_3[2927:2920];
        layer3[45][39:32] = buffer_data_3[2935:2928];
        layer3[45][47:40] = buffer_data_3[2943:2936];
        layer3[45][55:48] = buffer_data_3[2951:2944];
        layer4[45][7:0] = buffer_data_2[2903:2896];
        layer4[45][15:8] = buffer_data_2[2911:2904];
        layer4[45][23:16] = buffer_data_2[2919:2912];
        layer4[45][31:24] = buffer_data_2[2927:2920];
        layer4[45][39:32] = buffer_data_2[2935:2928];
        layer4[45][47:40] = buffer_data_2[2943:2936];
        layer4[45][55:48] = buffer_data_2[2951:2944];
        layer5[45][7:0] = buffer_data_1[2903:2896];
        layer5[45][15:8] = buffer_data_1[2911:2904];
        layer5[45][23:16] = buffer_data_1[2919:2912];
        layer5[45][31:24] = buffer_data_1[2927:2920];
        layer5[45][39:32] = buffer_data_1[2935:2928];
        layer5[45][47:40] = buffer_data_1[2943:2936];
        layer5[45][55:48] = buffer_data_1[2951:2944];
        layer6[45][7:0] = buffer_data_0[2903:2896];
        layer6[45][15:8] = buffer_data_0[2911:2904];
        layer6[45][23:16] = buffer_data_0[2919:2912];
        layer6[45][31:24] = buffer_data_0[2927:2920];
        layer6[45][39:32] = buffer_data_0[2935:2928];
        layer6[45][47:40] = buffer_data_0[2943:2936];
        layer6[45][55:48] = buffer_data_0[2951:2944];
        layer0[46][7:0] = buffer_data_6[2911:2904];
        layer0[46][15:8] = buffer_data_6[2919:2912];
        layer0[46][23:16] = buffer_data_6[2927:2920];
        layer0[46][31:24] = buffer_data_6[2935:2928];
        layer0[46][39:32] = buffer_data_6[2943:2936];
        layer0[46][47:40] = buffer_data_6[2951:2944];
        layer0[46][55:48] = buffer_data_6[2959:2952];
        layer1[46][7:0] = buffer_data_5[2911:2904];
        layer1[46][15:8] = buffer_data_5[2919:2912];
        layer1[46][23:16] = buffer_data_5[2927:2920];
        layer1[46][31:24] = buffer_data_5[2935:2928];
        layer1[46][39:32] = buffer_data_5[2943:2936];
        layer1[46][47:40] = buffer_data_5[2951:2944];
        layer1[46][55:48] = buffer_data_5[2959:2952];
        layer2[46][7:0] = buffer_data_4[2911:2904];
        layer2[46][15:8] = buffer_data_4[2919:2912];
        layer2[46][23:16] = buffer_data_4[2927:2920];
        layer2[46][31:24] = buffer_data_4[2935:2928];
        layer2[46][39:32] = buffer_data_4[2943:2936];
        layer2[46][47:40] = buffer_data_4[2951:2944];
        layer2[46][55:48] = buffer_data_4[2959:2952];
        layer3[46][7:0] = buffer_data_3[2911:2904];
        layer3[46][15:8] = buffer_data_3[2919:2912];
        layer3[46][23:16] = buffer_data_3[2927:2920];
        layer3[46][31:24] = buffer_data_3[2935:2928];
        layer3[46][39:32] = buffer_data_3[2943:2936];
        layer3[46][47:40] = buffer_data_3[2951:2944];
        layer3[46][55:48] = buffer_data_3[2959:2952];
        layer4[46][7:0] = buffer_data_2[2911:2904];
        layer4[46][15:8] = buffer_data_2[2919:2912];
        layer4[46][23:16] = buffer_data_2[2927:2920];
        layer4[46][31:24] = buffer_data_2[2935:2928];
        layer4[46][39:32] = buffer_data_2[2943:2936];
        layer4[46][47:40] = buffer_data_2[2951:2944];
        layer4[46][55:48] = buffer_data_2[2959:2952];
        layer5[46][7:0] = buffer_data_1[2911:2904];
        layer5[46][15:8] = buffer_data_1[2919:2912];
        layer5[46][23:16] = buffer_data_1[2927:2920];
        layer5[46][31:24] = buffer_data_1[2935:2928];
        layer5[46][39:32] = buffer_data_1[2943:2936];
        layer5[46][47:40] = buffer_data_1[2951:2944];
        layer5[46][55:48] = buffer_data_1[2959:2952];
        layer6[46][7:0] = buffer_data_0[2911:2904];
        layer6[46][15:8] = buffer_data_0[2919:2912];
        layer6[46][23:16] = buffer_data_0[2927:2920];
        layer6[46][31:24] = buffer_data_0[2935:2928];
        layer6[46][39:32] = buffer_data_0[2943:2936];
        layer6[46][47:40] = buffer_data_0[2951:2944];
        layer6[46][55:48] = buffer_data_0[2959:2952];
        layer0[47][7:0] = buffer_data_6[2919:2912];
        layer0[47][15:8] = buffer_data_6[2927:2920];
        layer0[47][23:16] = buffer_data_6[2935:2928];
        layer0[47][31:24] = buffer_data_6[2943:2936];
        layer0[47][39:32] = buffer_data_6[2951:2944];
        layer0[47][47:40] = buffer_data_6[2959:2952];
        layer0[47][55:48] = buffer_data_6[2967:2960];
        layer1[47][7:0] = buffer_data_5[2919:2912];
        layer1[47][15:8] = buffer_data_5[2927:2920];
        layer1[47][23:16] = buffer_data_5[2935:2928];
        layer1[47][31:24] = buffer_data_5[2943:2936];
        layer1[47][39:32] = buffer_data_5[2951:2944];
        layer1[47][47:40] = buffer_data_5[2959:2952];
        layer1[47][55:48] = buffer_data_5[2967:2960];
        layer2[47][7:0] = buffer_data_4[2919:2912];
        layer2[47][15:8] = buffer_data_4[2927:2920];
        layer2[47][23:16] = buffer_data_4[2935:2928];
        layer2[47][31:24] = buffer_data_4[2943:2936];
        layer2[47][39:32] = buffer_data_4[2951:2944];
        layer2[47][47:40] = buffer_data_4[2959:2952];
        layer2[47][55:48] = buffer_data_4[2967:2960];
        layer3[47][7:0] = buffer_data_3[2919:2912];
        layer3[47][15:8] = buffer_data_3[2927:2920];
        layer3[47][23:16] = buffer_data_3[2935:2928];
        layer3[47][31:24] = buffer_data_3[2943:2936];
        layer3[47][39:32] = buffer_data_3[2951:2944];
        layer3[47][47:40] = buffer_data_3[2959:2952];
        layer3[47][55:48] = buffer_data_3[2967:2960];
        layer4[47][7:0] = buffer_data_2[2919:2912];
        layer4[47][15:8] = buffer_data_2[2927:2920];
        layer4[47][23:16] = buffer_data_2[2935:2928];
        layer4[47][31:24] = buffer_data_2[2943:2936];
        layer4[47][39:32] = buffer_data_2[2951:2944];
        layer4[47][47:40] = buffer_data_2[2959:2952];
        layer4[47][55:48] = buffer_data_2[2967:2960];
        layer5[47][7:0] = buffer_data_1[2919:2912];
        layer5[47][15:8] = buffer_data_1[2927:2920];
        layer5[47][23:16] = buffer_data_1[2935:2928];
        layer5[47][31:24] = buffer_data_1[2943:2936];
        layer5[47][39:32] = buffer_data_1[2951:2944];
        layer5[47][47:40] = buffer_data_1[2959:2952];
        layer5[47][55:48] = buffer_data_1[2967:2960];
        layer6[47][7:0] = buffer_data_0[2919:2912];
        layer6[47][15:8] = buffer_data_0[2927:2920];
        layer6[47][23:16] = buffer_data_0[2935:2928];
        layer6[47][31:24] = buffer_data_0[2943:2936];
        layer6[47][39:32] = buffer_data_0[2951:2944];
        layer6[47][47:40] = buffer_data_0[2959:2952];
        layer6[47][55:48] = buffer_data_0[2967:2960];
        layer0[48][7:0] = buffer_data_6[2927:2920];
        layer0[48][15:8] = buffer_data_6[2935:2928];
        layer0[48][23:16] = buffer_data_6[2943:2936];
        layer0[48][31:24] = buffer_data_6[2951:2944];
        layer0[48][39:32] = buffer_data_6[2959:2952];
        layer0[48][47:40] = buffer_data_6[2967:2960];
        layer0[48][55:48] = buffer_data_6[2975:2968];
        layer1[48][7:0] = buffer_data_5[2927:2920];
        layer1[48][15:8] = buffer_data_5[2935:2928];
        layer1[48][23:16] = buffer_data_5[2943:2936];
        layer1[48][31:24] = buffer_data_5[2951:2944];
        layer1[48][39:32] = buffer_data_5[2959:2952];
        layer1[48][47:40] = buffer_data_5[2967:2960];
        layer1[48][55:48] = buffer_data_5[2975:2968];
        layer2[48][7:0] = buffer_data_4[2927:2920];
        layer2[48][15:8] = buffer_data_4[2935:2928];
        layer2[48][23:16] = buffer_data_4[2943:2936];
        layer2[48][31:24] = buffer_data_4[2951:2944];
        layer2[48][39:32] = buffer_data_4[2959:2952];
        layer2[48][47:40] = buffer_data_4[2967:2960];
        layer2[48][55:48] = buffer_data_4[2975:2968];
        layer3[48][7:0] = buffer_data_3[2927:2920];
        layer3[48][15:8] = buffer_data_3[2935:2928];
        layer3[48][23:16] = buffer_data_3[2943:2936];
        layer3[48][31:24] = buffer_data_3[2951:2944];
        layer3[48][39:32] = buffer_data_3[2959:2952];
        layer3[48][47:40] = buffer_data_3[2967:2960];
        layer3[48][55:48] = buffer_data_3[2975:2968];
        layer4[48][7:0] = buffer_data_2[2927:2920];
        layer4[48][15:8] = buffer_data_2[2935:2928];
        layer4[48][23:16] = buffer_data_2[2943:2936];
        layer4[48][31:24] = buffer_data_2[2951:2944];
        layer4[48][39:32] = buffer_data_2[2959:2952];
        layer4[48][47:40] = buffer_data_2[2967:2960];
        layer4[48][55:48] = buffer_data_2[2975:2968];
        layer5[48][7:0] = buffer_data_1[2927:2920];
        layer5[48][15:8] = buffer_data_1[2935:2928];
        layer5[48][23:16] = buffer_data_1[2943:2936];
        layer5[48][31:24] = buffer_data_1[2951:2944];
        layer5[48][39:32] = buffer_data_1[2959:2952];
        layer5[48][47:40] = buffer_data_1[2967:2960];
        layer5[48][55:48] = buffer_data_1[2975:2968];
        layer6[48][7:0] = buffer_data_0[2927:2920];
        layer6[48][15:8] = buffer_data_0[2935:2928];
        layer6[48][23:16] = buffer_data_0[2943:2936];
        layer6[48][31:24] = buffer_data_0[2951:2944];
        layer6[48][39:32] = buffer_data_0[2959:2952];
        layer6[48][47:40] = buffer_data_0[2967:2960];
        layer6[48][55:48] = buffer_data_0[2975:2968];
        layer0[49][7:0] = buffer_data_6[2935:2928];
        layer0[49][15:8] = buffer_data_6[2943:2936];
        layer0[49][23:16] = buffer_data_6[2951:2944];
        layer0[49][31:24] = buffer_data_6[2959:2952];
        layer0[49][39:32] = buffer_data_6[2967:2960];
        layer0[49][47:40] = buffer_data_6[2975:2968];
        layer0[49][55:48] = buffer_data_6[2983:2976];
        layer1[49][7:0] = buffer_data_5[2935:2928];
        layer1[49][15:8] = buffer_data_5[2943:2936];
        layer1[49][23:16] = buffer_data_5[2951:2944];
        layer1[49][31:24] = buffer_data_5[2959:2952];
        layer1[49][39:32] = buffer_data_5[2967:2960];
        layer1[49][47:40] = buffer_data_5[2975:2968];
        layer1[49][55:48] = buffer_data_5[2983:2976];
        layer2[49][7:0] = buffer_data_4[2935:2928];
        layer2[49][15:8] = buffer_data_4[2943:2936];
        layer2[49][23:16] = buffer_data_4[2951:2944];
        layer2[49][31:24] = buffer_data_4[2959:2952];
        layer2[49][39:32] = buffer_data_4[2967:2960];
        layer2[49][47:40] = buffer_data_4[2975:2968];
        layer2[49][55:48] = buffer_data_4[2983:2976];
        layer3[49][7:0] = buffer_data_3[2935:2928];
        layer3[49][15:8] = buffer_data_3[2943:2936];
        layer3[49][23:16] = buffer_data_3[2951:2944];
        layer3[49][31:24] = buffer_data_3[2959:2952];
        layer3[49][39:32] = buffer_data_3[2967:2960];
        layer3[49][47:40] = buffer_data_3[2975:2968];
        layer3[49][55:48] = buffer_data_3[2983:2976];
        layer4[49][7:0] = buffer_data_2[2935:2928];
        layer4[49][15:8] = buffer_data_2[2943:2936];
        layer4[49][23:16] = buffer_data_2[2951:2944];
        layer4[49][31:24] = buffer_data_2[2959:2952];
        layer4[49][39:32] = buffer_data_2[2967:2960];
        layer4[49][47:40] = buffer_data_2[2975:2968];
        layer4[49][55:48] = buffer_data_2[2983:2976];
        layer5[49][7:0] = buffer_data_1[2935:2928];
        layer5[49][15:8] = buffer_data_1[2943:2936];
        layer5[49][23:16] = buffer_data_1[2951:2944];
        layer5[49][31:24] = buffer_data_1[2959:2952];
        layer5[49][39:32] = buffer_data_1[2967:2960];
        layer5[49][47:40] = buffer_data_1[2975:2968];
        layer5[49][55:48] = buffer_data_1[2983:2976];
        layer6[49][7:0] = buffer_data_0[2935:2928];
        layer6[49][15:8] = buffer_data_0[2943:2936];
        layer6[49][23:16] = buffer_data_0[2951:2944];
        layer6[49][31:24] = buffer_data_0[2959:2952];
        layer6[49][39:32] = buffer_data_0[2967:2960];
        layer6[49][47:40] = buffer_data_0[2975:2968];
        layer6[49][55:48] = buffer_data_0[2983:2976];
        layer0[50][7:0] = buffer_data_6[2943:2936];
        layer0[50][15:8] = buffer_data_6[2951:2944];
        layer0[50][23:16] = buffer_data_6[2959:2952];
        layer0[50][31:24] = buffer_data_6[2967:2960];
        layer0[50][39:32] = buffer_data_6[2975:2968];
        layer0[50][47:40] = buffer_data_6[2983:2976];
        layer0[50][55:48] = buffer_data_6[2991:2984];
        layer1[50][7:0] = buffer_data_5[2943:2936];
        layer1[50][15:8] = buffer_data_5[2951:2944];
        layer1[50][23:16] = buffer_data_5[2959:2952];
        layer1[50][31:24] = buffer_data_5[2967:2960];
        layer1[50][39:32] = buffer_data_5[2975:2968];
        layer1[50][47:40] = buffer_data_5[2983:2976];
        layer1[50][55:48] = buffer_data_5[2991:2984];
        layer2[50][7:0] = buffer_data_4[2943:2936];
        layer2[50][15:8] = buffer_data_4[2951:2944];
        layer2[50][23:16] = buffer_data_4[2959:2952];
        layer2[50][31:24] = buffer_data_4[2967:2960];
        layer2[50][39:32] = buffer_data_4[2975:2968];
        layer2[50][47:40] = buffer_data_4[2983:2976];
        layer2[50][55:48] = buffer_data_4[2991:2984];
        layer3[50][7:0] = buffer_data_3[2943:2936];
        layer3[50][15:8] = buffer_data_3[2951:2944];
        layer3[50][23:16] = buffer_data_3[2959:2952];
        layer3[50][31:24] = buffer_data_3[2967:2960];
        layer3[50][39:32] = buffer_data_3[2975:2968];
        layer3[50][47:40] = buffer_data_3[2983:2976];
        layer3[50][55:48] = buffer_data_3[2991:2984];
        layer4[50][7:0] = buffer_data_2[2943:2936];
        layer4[50][15:8] = buffer_data_2[2951:2944];
        layer4[50][23:16] = buffer_data_2[2959:2952];
        layer4[50][31:24] = buffer_data_2[2967:2960];
        layer4[50][39:32] = buffer_data_2[2975:2968];
        layer4[50][47:40] = buffer_data_2[2983:2976];
        layer4[50][55:48] = buffer_data_2[2991:2984];
        layer5[50][7:0] = buffer_data_1[2943:2936];
        layer5[50][15:8] = buffer_data_1[2951:2944];
        layer5[50][23:16] = buffer_data_1[2959:2952];
        layer5[50][31:24] = buffer_data_1[2967:2960];
        layer5[50][39:32] = buffer_data_1[2975:2968];
        layer5[50][47:40] = buffer_data_1[2983:2976];
        layer5[50][55:48] = buffer_data_1[2991:2984];
        layer6[50][7:0] = buffer_data_0[2943:2936];
        layer6[50][15:8] = buffer_data_0[2951:2944];
        layer6[50][23:16] = buffer_data_0[2959:2952];
        layer6[50][31:24] = buffer_data_0[2967:2960];
        layer6[50][39:32] = buffer_data_0[2975:2968];
        layer6[50][47:40] = buffer_data_0[2983:2976];
        layer6[50][55:48] = buffer_data_0[2991:2984];
        layer0[51][7:0] = buffer_data_6[2951:2944];
        layer0[51][15:8] = buffer_data_6[2959:2952];
        layer0[51][23:16] = buffer_data_6[2967:2960];
        layer0[51][31:24] = buffer_data_6[2975:2968];
        layer0[51][39:32] = buffer_data_6[2983:2976];
        layer0[51][47:40] = buffer_data_6[2991:2984];
        layer0[51][55:48] = buffer_data_6[2999:2992];
        layer1[51][7:0] = buffer_data_5[2951:2944];
        layer1[51][15:8] = buffer_data_5[2959:2952];
        layer1[51][23:16] = buffer_data_5[2967:2960];
        layer1[51][31:24] = buffer_data_5[2975:2968];
        layer1[51][39:32] = buffer_data_5[2983:2976];
        layer1[51][47:40] = buffer_data_5[2991:2984];
        layer1[51][55:48] = buffer_data_5[2999:2992];
        layer2[51][7:0] = buffer_data_4[2951:2944];
        layer2[51][15:8] = buffer_data_4[2959:2952];
        layer2[51][23:16] = buffer_data_4[2967:2960];
        layer2[51][31:24] = buffer_data_4[2975:2968];
        layer2[51][39:32] = buffer_data_4[2983:2976];
        layer2[51][47:40] = buffer_data_4[2991:2984];
        layer2[51][55:48] = buffer_data_4[2999:2992];
        layer3[51][7:0] = buffer_data_3[2951:2944];
        layer3[51][15:8] = buffer_data_3[2959:2952];
        layer3[51][23:16] = buffer_data_3[2967:2960];
        layer3[51][31:24] = buffer_data_3[2975:2968];
        layer3[51][39:32] = buffer_data_3[2983:2976];
        layer3[51][47:40] = buffer_data_3[2991:2984];
        layer3[51][55:48] = buffer_data_3[2999:2992];
        layer4[51][7:0] = buffer_data_2[2951:2944];
        layer4[51][15:8] = buffer_data_2[2959:2952];
        layer4[51][23:16] = buffer_data_2[2967:2960];
        layer4[51][31:24] = buffer_data_2[2975:2968];
        layer4[51][39:32] = buffer_data_2[2983:2976];
        layer4[51][47:40] = buffer_data_2[2991:2984];
        layer4[51][55:48] = buffer_data_2[2999:2992];
        layer5[51][7:0] = buffer_data_1[2951:2944];
        layer5[51][15:8] = buffer_data_1[2959:2952];
        layer5[51][23:16] = buffer_data_1[2967:2960];
        layer5[51][31:24] = buffer_data_1[2975:2968];
        layer5[51][39:32] = buffer_data_1[2983:2976];
        layer5[51][47:40] = buffer_data_1[2991:2984];
        layer5[51][55:48] = buffer_data_1[2999:2992];
        layer6[51][7:0] = buffer_data_0[2951:2944];
        layer6[51][15:8] = buffer_data_0[2959:2952];
        layer6[51][23:16] = buffer_data_0[2967:2960];
        layer6[51][31:24] = buffer_data_0[2975:2968];
        layer6[51][39:32] = buffer_data_0[2983:2976];
        layer6[51][47:40] = buffer_data_0[2991:2984];
        layer6[51][55:48] = buffer_data_0[2999:2992];
        layer0[52][7:0] = buffer_data_6[2959:2952];
        layer0[52][15:8] = buffer_data_6[2967:2960];
        layer0[52][23:16] = buffer_data_6[2975:2968];
        layer0[52][31:24] = buffer_data_6[2983:2976];
        layer0[52][39:32] = buffer_data_6[2991:2984];
        layer0[52][47:40] = buffer_data_6[2999:2992];
        layer0[52][55:48] = buffer_data_6[3007:3000];
        layer1[52][7:0] = buffer_data_5[2959:2952];
        layer1[52][15:8] = buffer_data_5[2967:2960];
        layer1[52][23:16] = buffer_data_5[2975:2968];
        layer1[52][31:24] = buffer_data_5[2983:2976];
        layer1[52][39:32] = buffer_data_5[2991:2984];
        layer1[52][47:40] = buffer_data_5[2999:2992];
        layer1[52][55:48] = buffer_data_5[3007:3000];
        layer2[52][7:0] = buffer_data_4[2959:2952];
        layer2[52][15:8] = buffer_data_4[2967:2960];
        layer2[52][23:16] = buffer_data_4[2975:2968];
        layer2[52][31:24] = buffer_data_4[2983:2976];
        layer2[52][39:32] = buffer_data_4[2991:2984];
        layer2[52][47:40] = buffer_data_4[2999:2992];
        layer2[52][55:48] = buffer_data_4[3007:3000];
        layer3[52][7:0] = buffer_data_3[2959:2952];
        layer3[52][15:8] = buffer_data_3[2967:2960];
        layer3[52][23:16] = buffer_data_3[2975:2968];
        layer3[52][31:24] = buffer_data_3[2983:2976];
        layer3[52][39:32] = buffer_data_3[2991:2984];
        layer3[52][47:40] = buffer_data_3[2999:2992];
        layer3[52][55:48] = buffer_data_3[3007:3000];
        layer4[52][7:0] = buffer_data_2[2959:2952];
        layer4[52][15:8] = buffer_data_2[2967:2960];
        layer4[52][23:16] = buffer_data_2[2975:2968];
        layer4[52][31:24] = buffer_data_2[2983:2976];
        layer4[52][39:32] = buffer_data_2[2991:2984];
        layer4[52][47:40] = buffer_data_2[2999:2992];
        layer4[52][55:48] = buffer_data_2[3007:3000];
        layer5[52][7:0] = buffer_data_1[2959:2952];
        layer5[52][15:8] = buffer_data_1[2967:2960];
        layer5[52][23:16] = buffer_data_1[2975:2968];
        layer5[52][31:24] = buffer_data_1[2983:2976];
        layer5[52][39:32] = buffer_data_1[2991:2984];
        layer5[52][47:40] = buffer_data_1[2999:2992];
        layer5[52][55:48] = buffer_data_1[3007:3000];
        layer6[52][7:0] = buffer_data_0[2959:2952];
        layer6[52][15:8] = buffer_data_0[2967:2960];
        layer6[52][23:16] = buffer_data_0[2975:2968];
        layer6[52][31:24] = buffer_data_0[2983:2976];
        layer6[52][39:32] = buffer_data_0[2991:2984];
        layer6[52][47:40] = buffer_data_0[2999:2992];
        layer6[52][55:48] = buffer_data_0[3007:3000];
        layer0[53][7:0] = buffer_data_6[2967:2960];
        layer0[53][15:8] = buffer_data_6[2975:2968];
        layer0[53][23:16] = buffer_data_6[2983:2976];
        layer0[53][31:24] = buffer_data_6[2991:2984];
        layer0[53][39:32] = buffer_data_6[2999:2992];
        layer0[53][47:40] = buffer_data_6[3007:3000];
        layer0[53][55:48] = buffer_data_6[3015:3008];
        layer1[53][7:0] = buffer_data_5[2967:2960];
        layer1[53][15:8] = buffer_data_5[2975:2968];
        layer1[53][23:16] = buffer_data_5[2983:2976];
        layer1[53][31:24] = buffer_data_5[2991:2984];
        layer1[53][39:32] = buffer_data_5[2999:2992];
        layer1[53][47:40] = buffer_data_5[3007:3000];
        layer1[53][55:48] = buffer_data_5[3015:3008];
        layer2[53][7:0] = buffer_data_4[2967:2960];
        layer2[53][15:8] = buffer_data_4[2975:2968];
        layer2[53][23:16] = buffer_data_4[2983:2976];
        layer2[53][31:24] = buffer_data_4[2991:2984];
        layer2[53][39:32] = buffer_data_4[2999:2992];
        layer2[53][47:40] = buffer_data_4[3007:3000];
        layer2[53][55:48] = buffer_data_4[3015:3008];
        layer3[53][7:0] = buffer_data_3[2967:2960];
        layer3[53][15:8] = buffer_data_3[2975:2968];
        layer3[53][23:16] = buffer_data_3[2983:2976];
        layer3[53][31:24] = buffer_data_3[2991:2984];
        layer3[53][39:32] = buffer_data_3[2999:2992];
        layer3[53][47:40] = buffer_data_3[3007:3000];
        layer3[53][55:48] = buffer_data_3[3015:3008];
        layer4[53][7:0] = buffer_data_2[2967:2960];
        layer4[53][15:8] = buffer_data_2[2975:2968];
        layer4[53][23:16] = buffer_data_2[2983:2976];
        layer4[53][31:24] = buffer_data_2[2991:2984];
        layer4[53][39:32] = buffer_data_2[2999:2992];
        layer4[53][47:40] = buffer_data_2[3007:3000];
        layer4[53][55:48] = buffer_data_2[3015:3008];
        layer5[53][7:0] = buffer_data_1[2967:2960];
        layer5[53][15:8] = buffer_data_1[2975:2968];
        layer5[53][23:16] = buffer_data_1[2983:2976];
        layer5[53][31:24] = buffer_data_1[2991:2984];
        layer5[53][39:32] = buffer_data_1[2999:2992];
        layer5[53][47:40] = buffer_data_1[3007:3000];
        layer5[53][55:48] = buffer_data_1[3015:3008];
        layer6[53][7:0] = buffer_data_0[2967:2960];
        layer6[53][15:8] = buffer_data_0[2975:2968];
        layer6[53][23:16] = buffer_data_0[2983:2976];
        layer6[53][31:24] = buffer_data_0[2991:2984];
        layer6[53][39:32] = buffer_data_0[2999:2992];
        layer6[53][47:40] = buffer_data_0[3007:3000];
        layer6[53][55:48] = buffer_data_0[3015:3008];
        layer0[54][7:0] = buffer_data_6[2975:2968];
        layer0[54][15:8] = buffer_data_6[2983:2976];
        layer0[54][23:16] = buffer_data_6[2991:2984];
        layer0[54][31:24] = buffer_data_6[2999:2992];
        layer0[54][39:32] = buffer_data_6[3007:3000];
        layer0[54][47:40] = buffer_data_6[3015:3008];
        layer0[54][55:48] = buffer_data_6[3023:3016];
        layer1[54][7:0] = buffer_data_5[2975:2968];
        layer1[54][15:8] = buffer_data_5[2983:2976];
        layer1[54][23:16] = buffer_data_5[2991:2984];
        layer1[54][31:24] = buffer_data_5[2999:2992];
        layer1[54][39:32] = buffer_data_5[3007:3000];
        layer1[54][47:40] = buffer_data_5[3015:3008];
        layer1[54][55:48] = buffer_data_5[3023:3016];
        layer2[54][7:0] = buffer_data_4[2975:2968];
        layer2[54][15:8] = buffer_data_4[2983:2976];
        layer2[54][23:16] = buffer_data_4[2991:2984];
        layer2[54][31:24] = buffer_data_4[2999:2992];
        layer2[54][39:32] = buffer_data_4[3007:3000];
        layer2[54][47:40] = buffer_data_4[3015:3008];
        layer2[54][55:48] = buffer_data_4[3023:3016];
        layer3[54][7:0] = buffer_data_3[2975:2968];
        layer3[54][15:8] = buffer_data_3[2983:2976];
        layer3[54][23:16] = buffer_data_3[2991:2984];
        layer3[54][31:24] = buffer_data_3[2999:2992];
        layer3[54][39:32] = buffer_data_3[3007:3000];
        layer3[54][47:40] = buffer_data_3[3015:3008];
        layer3[54][55:48] = buffer_data_3[3023:3016];
        layer4[54][7:0] = buffer_data_2[2975:2968];
        layer4[54][15:8] = buffer_data_2[2983:2976];
        layer4[54][23:16] = buffer_data_2[2991:2984];
        layer4[54][31:24] = buffer_data_2[2999:2992];
        layer4[54][39:32] = buffer_data_2[3007:3000];
        layer4[54][47:40] = buffer_data_2[3015:3008];
        layer4[54][55:48] = buffer_data_2[3023:3016];
        layer5[54][7:0] = buffer_data_1[2975:2968];
        layer5[54][15:8] = buffer_data_1[2983:2976];
        layer5[54][23:16] = buffer_data_1[2991:2984];
        layer5[54][31:24] = buffer_data_1[2999:2992];
        layer5[54][39:32] = buffer_data_1[3007:3000];
        layer5[54][47:40] = buffer_data_1[3015:3008];
        layer5[54][55:48] = buffer_data_1[3023:3016];
        layer6[54][7:0] = buffer_data_0[2975:2968];
        layer6[54][15:8] = buffer_data_0[2983:2976];
        layer6[54][23:16] = buffer_data_0[2991:2984];
        layer6[54][31:24] = buffer_data_0[2999:2992];
        layer6[54][39:32] = buffer_data_0[3007:3000];
        layer6[54][47:40] = buffer_data_0[3015:3008];
        layer6[54][55:48] = buffer_data_0[3023:3016];
        layer0[55][7:0] = buffer_data_6[2983:2976];
        layer0[55][15:8] = buffer_data_6[2991:2984];
        layer0[55][23:16] = buffer_data_6[2999:2992];
        layer0[55][31:24] = buffer_data_6[3007:3000];
        layer0[55][39:32] = buffer_data_6[3015:3008];
        layer0[55][47:40] = buffer_data_6[3023:3016];
        layer0[55][55:48] = buffer_data_6[3031:3024];
        layer1[55][7:0] = buffer_data_5[2983:2976];
        layer1[55][15:8] = buffer_data_5[2991:2984];
        layer1[55][23:16] = buffer_data_5[2999:2992];
        layer1[55][31:24] = buffer_data_5[3007:3000];
        layer1[55][39:32] = buffer_data_5[3015:3008];
        layer1[55][47:40] = buffer_data_5[3023:3016];
        layer1[55][55:48] = buffer_data_5[3031:3024];
        layer2[55][7:0] = buffer_data_4[2983:2976];
        layer2[55][15:8] = buffer_data_4[2991:2984];
        layer2[55][23:16] = buffer_data_4[2999:2992];
        layer2[55][31:24] = buffer_data_4[3007:3000];
        layer2[55][39:32] = buffer_data_4[3015:3008];
        layer2[55][47:40] = buffer_data_4[3023:3016];
        layer2[55][55:48] = buffer_data_4[3031:3024];
        layer3[55][7:0] = buffer_data_3[2983:2976];
        layer3[55][15:8] = buffer_data_3[2991:2984];
        layer3[55][23:16] = buffer_data_3[2999:2992];
        layer3[55][31:24] = buffer_data_3[3007:3000];
        layer3[55][39:32] = buffer_data_3[3015:3008];
        layer3[55][47:40] = buffer_data_3[3023:3016];
        layer3[55][55:48] = buffer_data_3[3031:3024];
        layer4[55][7:0] = buffer_data_2[2983:2976];
        layer4[55][15:8] = buffer_data_2[2991:2984];
        layer4[55][23:16] = buffer_data_2[2999:2992];
        layer4[55][31:24] = buffer_data_2[3007:3000];
        layer4[55][39:32] = buffer_data_2[3015:3008];
        layer4[55][47:40] = buffer_data_2[3023:3016];
        layer4[55][55:48] = buffer_data_2[3031:3024];
        layer5[55][7:0] = buffer_data_1[2983:2976];
        layer5[55][15:8] = buffer_data_1[2991:2984];
        layer5[55][23:16] = buffer_data_1[2999:2992];
        layer5[55][31:24] = buffer_data_1[3007:3000];
        layer5[55][39:32] = buffer_data_1[3015:3008];
        layer5[55][47:40] = buffer_data_1[3023:3016];
        layer5[55][55:48] = buffer_data_1[3031:3024];
        layer6[55][7:0] = buffer_data_0[2983:2976];
        layer6[55][15:8] = buffer_data_0[2991:2984];
        layer6[55][23:16] = buffer_data_0[2999:2992];
        layer6[55][31:24] = buffer_data_0[3007:3000];
        layer6[55][39:32] = buffer_data_0[3015:3008];
        layer6[55][47:40] = buffer_data_0[3023:3016];
        layer6[55][55:48] = buffer_data_0[3031:3024];
        layer0[56][7:0] = buffer_data_6[2991:2984];
        layer0[56][15:8] = buffer_data_6[2999:2992];
        layer0[56][23:16] = buffer_data_6[3007:3000];
        layer0[56][31:24] = buffer_data_6[3015:3008];
        layer0[56][39:32] = buffer_data_6[3023:3016];
        layer0[56][47:40] = buffer_data_6[3031:3024];
        layer0[56][55:48] = buffer_data_6[3039:3032];
        layer1[56][7:0] = buffer_data_5[2991:2984];
        layer1[56][15:8] = buffer_data_5[2999:2992];
        layer1[56][23:16] = buffer_data_5[3007:3000];
        layer1[56][31:24] = buffer_data_5[3015:3008];
        layer1[56][39:32] = buffer_data_5[3023:3016];
        layer1[56][47:40] = buffer_data_5[3031:3024];
        layer1[56][55:48] = buffer_data_5[3039:3032];
        layer2[56][7:0] = buffer_data_4[2991:2984];
        layer2[56][15:8] = buffer_data_4[2999:2992];
        layer2[56][23:16] = buffer_data_4[3007:3000];
        layer2[56][31:24] = buffer_data_4[3015:3008];
        layer2[56][39:32] = buffer_data_4[3023:3016];
        layer2[56][47:40] = buffer_data_4[3031:3024];
        layer2[56][55:48] = buffer_data_4[3039:3032];
        layer3[56][7:0] = buffer_data_3[2991:2984];
        layer3[56][15:8] = buffer_data_3[2999:2992];
        layer3[56][23:16] = buffer_data_3[3007:3000];
        layer3[56][31:24] = buffer_data_3[3015:3008];
        layer3[56][39:32] = buffer_data_3[3023:3016];
        layer3[56][47:40] = buffer_data_3[3031:3024];
        layer3[56][55:48] = buffer_data_3[3039:3032];
        layer4[56][7:0] = buffer_data_2[2991:2984];
        layer4[56][15:8] = buffer_data_2[2999:2992];
        layer4[56][23:16] = buffer_data_2[3007:3000];
        layer4[56][31:24] = buffer_data_2[3015:3008];
        layer4[56][39:32] = buffer_data_2[3023:3016];
        layer4[56][47:40] = buffer_data_2[3031:3024];
        layer4[56][55:48] = buffer_data_2[3039:3032];
        layer5[56][7:0] = buffer_data_1[2991:2984];
        layer5[56][15:8] = buffer_data_1[2999:2992];
        layer5[56][23:16] = buffer_data_1[3007:3000];
        layer5[56][31:24] = buffer_data_1[3015:3008];
        layer5[56][39:32] = buffer_data_1[3023:3016];
        layer5[56][47:40] = buffer_data_1[3031:3024];
        layer5[56][55:48] = buffer_data_1[3039:3032];
        layer6[56][7:0] = buffer_data_0[2991:2984];
        layer6[56][15:8] = buffer_data_0[2999:2992];
        layer6[56][23:16] = buffer_data_0[3007:3000];
        layer6[56][31:24] = buffer_data_0[3015:3008];
        layer6[56][39:32] = buffer_data_0[3023:3016];
        layer6[56][47:40] = buffer_data_0[3031:3024];
        layer6[56][55:48] = buffer_data_0[3039:3032];
        layer0[57][7:0] = buffer_data_6[2999:2992];
        layer0[57][15:8] = buffer_data_6[3007:3000];
        layer0[57][23:16] = buffer_data_6[3015:3008];
        layer0[57][31:24] = buffer_data_6[3023:3016];
        layer0[57][39:32] = buffer_data_6[3031:3024];
        layer0[57][47:40] = buffer_data_6[3039:3032];
        layer0[57][55:48] = buffer_data_6[3047:3040];
        layer1[57][7:0] = buffer_data_5[2999:2992];
        layer1[57][15:8] = buffer_data_5[3007:3000];
        layer1[57][23:16] = buffer_data_5[3015:3008];
        layer1[57][31:24] = buffer_data_5[3023:3016];
        layer1[57][39:32] = buffer_data_5[3031:3024];
        layer1[57][47:40] = buffer_data_5[3039:3032];
        layer1[57][55:48] = buffer_data_5[3047:3040];
        layer2[57][7:0] = buffer_data_4[2999:2992];
        layer2[57][15:8] = buffer_data_4[3007:3000];
        layer2[57][23:16] = buffer_data_4[3015:3008];
        layer2[57][31:24] = buffer_data_4[3023:3016];
        layer2[57][39:32] = buffer_data_4[3031:3024];
        layer2[57][47:40] = buffer_data_4[3039:3032];
        layer2[57][55:48] = buffer_data_4[3047:3040];
        layer3[57][7:0] = buffer_data_3[2999:2992];
        layer3[57][15:8] = buffer_data_3[3007:3000];
        layer3[57][23:16] = buffer_data_3[3015:3008];
        layer3[57][31:24] = buffer_data_3[3023:3016];
        layer3[57][39:32] = buffer_data_3[3031:3024];
        layer3[57][47:40] = buffer_data_3[3039:3032];
        layer3[57][55:48] = buffer_data_3[3047:3040];
        layer4[57][7:0] = buffer_data_2[2999:2992];
        layer4[57][15:8] = buffer_data_2[3007:3000];
        layer4[57][23:16] = buffer_data_2[3015:3008];
        layer4[57][31:24] = buffer_data_2[3023:3016];
        layer4[57][39:32] = buffer_data_2[3031:3024];
        layer4[57][47:40] = buffer_data_2[3039:3032];
        layer4[57][55:48] = buffer_data_2[3047:3040];
        layer5[57][7:0] = buffer_data_1[2999:2992];
        layer5[57][15:8] = buffer_data_1[3007:3000];
        layer5[57][23:16] = buffer_data_1[3015:3008];
        layer5[57][31:24] = buffer_data_1[3023:3016];
        layer5[57][39:32] = buffer_data_1[3031:3024];
        layer5[57][47:40] = buffer_data_1[3039:3032];
        layer5[57][55:48] = buffer_data_1[3047:3040];
        layer6[57][7:0] = buffer_data_0[2999:2992];
        layer6[57][15:8] = buffer_data_0[3007:3000];
        layer6[57][23:16] = buffer_data_0[3015:3008];
        layer6[57][31:24] = buffer_data_0[3023:3016];
        layer6[57][39:32] = buffer_data_0[3031:3024];
        layer6[57][47:40] = buffer_data_0[3039:3032];
        layer6[57][55:48] = buffer_data_0[3047:3040];
        layer0[58][7:0] = buffer_data_6[3007:3000];
        layer0[58][15:8] = buffer_data_6[3015:3008];
        layer0[58][23:16] = buffer_data_6[3023:3016];
        layer0[58][31:24] = buffer_data_6[3031:3024];
        layer0[58][39:32] = buffer_data_6[3039:3032];
        layer0[58][47:40] = buffer_data_6[3047:3040];
        layer0[58][55:48] = buffer_data_6[3055:3048];
        layer1[58][7:0] = buffer_data_5[3007:3000];
        layer1[58][15:8] = buffer_data_5[3015:3008];
        layer1[58][23:16] = buffer_data_5[3023:3016];
        layer1[58][31:24] = buffer_data_5[3031:3024];
        layer1[58][39:32] = buffer_data_5[3039:3032];
        layer1[58][47:40] = buffer_data_5[3047:3040];
        layer1[58][55:48] = buffer_data_5[3055:3048];
        layer2[58][7:0] = buffer_data_4[3007:3000];
        layer2[58][15:8] = buffer_data_4[3015:3008];
        layer2[58][23:16] = buffer_data_4[3023:3016];
        layer2[58][31:24] = buffer_data_4[3031:3024];
        layer2[58][39:32] = buffer_data_4[3039:3032];
        layer2[58][47:40] = buffer_data_4[3047:3040];
        layer2[58][55:48] = buffer_data_4[3055:3048];
        layer3[58][7:0] = buffer_data_3[3007:3000];
        layer3[58][15:8] = buffer_data_3[3015:3008];
        layer3[58][23:16] = buffer_data_3[3023:3016];
        layer3[58][31:24] = buffer_data_3[3031:3024];
        layer3[58][39:32] = buffer_data_3[3039:3032];
        layer3[58][47:40] = buffer_data_3[3047:3040];
        layer3[58][55:48] = buffer_data_3[3055:3048];
        layer4[58][7:0] = buffer_data_2[3007:3000];
        layer4[58][15:8] = buffer_data_2[3015:3008];
        layer4[58][23:16] = buffer_data_2[3023:3016];
        layer4[58][31:24] = buffer_data_2[3031:3024];
        layer4[58][39:32] = buffer_data_2[3039:3032];
        layer4[58][47:40] = buffer_data_2[3047:3040];
        layer4[58][55:48] = buffer_data_2[3055:3048];
        layer5[58][7:0] = buffer_data_1[3007:3000];
        layer5[58][15:8] = buffer_data_1[3015:3008];
        layer5[58][23:16] = buffer_data_1[3023:3016];
        layer5[58][31:24] = buffer_data_1[3031:3024];
        layer5[58][39:32] = buffer_data_1[3039:3032];
        layer5[58][47:40] = buffer_data_1[3047:3040];
        layer5[58][55:48] = buffer_data_1[3055:3048];
        layer6[58][7:0] = buffer_data_0[3007:3000];
        layer6[58][15:8] = buffer_data_0[3015:3008];
        layer6[58][23:16] = buffer_data_0[3023:3016];
        layer6[58][31:24] = buffer_data_0[3031:3024];
        layer6[58][39:32] = buffer_data_0[3039:3032];
        layer6[58][47:40] = buffer_data_0[3047:3040];
        layer6[58][55:48] = buffer_data_0[3055:3048];
        layer0[59][7:0] = buffer_data_6[3015:3008];
        layer0[59][15:8] = buffer_data_6[3023:3016];
        layer0[59][23:16] = buffer_data_6[3031:3024];
        layer0[59][31:24] = buffer_data_6[3039:3032];
        layer0[59][39:32] = buffer_data_6[3047:3040];
        layer0[59][47:40] = buffer_data_6[3055:3048];
        layer0[59][55:48] = buffer_data_6[3063:3056];
        layer1[59][7:0] = buffer_data_5[3015:3008];
        layer1[59][15:8] = buffer_data_5[3023:3016];
        layer1[59][23:16] = buffer_data_5[3031:3024];
        layer1[59][31:24] = buffer_data_5[3039:3032];
        layer1[59][39:32] = buffer_data_5[3047:3040];
        layer1[59][47:40] = buffer_data_5[3055:3048];
        layer1[59][55:48] = buffer_data_5[3063:3056];
        layer2[59][7:0] = buffer_data_4[3015:3008];
        layer2[59][15:8] = buffer_data_4[3023:3016];
        layer2[59][23:16] = buffer_data_4[3031:3024];
        layer2[59][31:24] = buffer_data_4[3039:3032];
        layer2[59][39:32] = buffer_data_4[3047:3040];
        layer2[59][47:40] = buffer_data_4[3055:3048];
        layer2[59][55:48] = buffer_data_4[3063:3056];
        layer3[59][7:0] = buffer_data_3[3015:3008];
        layer3[59][15:8] = buffer_data_3[3023:3016];
        layer3[59][23:16] = buffer_data_3[3031:3024];
        layer3[59][31:24] = buffer_data_3[3039:3032];
        layer3[59][39:32] = buffer_data_3[3047:3040];
        layer3[59][47:40] = buffer_data_3[3055:3048];
        layer3[59][55:48] = buffer_data_3[3063:3056];
        layer4[59][7:0] = buffer_data_2[3015:3008];
        layer4[59][15:8] = buffer_data_2[3023:3016];
        layer4[59][23:16] = buffer_data_2[3031:3024];
        layer4[59][31:24] = buffer_data_2[3039:3032];
        layer4[59][39:32] = buffer_data_2[3047:3040];
        layer4[59][47:40] = buffer_data_2[3055:3048];
        layer4[59][55:48] = buffer_data_2[3063:3056];
        layer5[59][7:0] = buffer_data_1[3015:3008];
        layer5[59][15:8] = buffer_data_1[3023:3016];
        layer5[59][23:16] = buffer_data_1[3031:3024];
        layer5[59][31:24] = buffer_data_1[3039:3032];
        layer5[59][39:32] = buffer_data_1[3047:3040];
        layer5[59][47:40] = buffer_data_1[3055:3048];
        layer5[59][55:48] = buffer_data_1[3063:3056];
        layer6[59][7:0] = buffer_data_0[3015:3008];
        layer6[59][15:8] = buffer_data_0[3023:3016];
        layer6[59][23:16] = buffer_data_0[3031:3024];
        layer6[59][31:24] = buffer_data_0[3039:3032];
        layer6[59][39:32] = buffer_data_0[3047:3040];
        layer6[59][47:40] = buffer_data_0[3055:3048];
        layer6[59][55:48] = buffer_data_0[3063:3056];
        layer0[60][7:0] = buffer_data_6[3023:3016];
        layer0[60][15:8] = buffer_data_6[3031:3024];
        layer0[60][23:16] = buffer_data_6[3039:3032];
        layer0[60][31:24] = buffer_data_6[3047:3040];
        layer0[60][39:32] = buffer_data_6[3055:3048];
        layer0[60][47:40] = buffer_data_6[3063:3056];
        layer0[60][55:48] = buffer_data_6[3071:3064];
        layer1[60][7:0] = buffer_data_5[3023:3016];
        layer1[60][15:8] = buffer_data_5[3031:3024];
        layer1[60][23:16] = buffer_data_5[3039:3032];
        layer1[60][31:24] = buffer_data_5[3047:3040];
        layer1[60][39:32] = buffer_data_5[3055:3048];
        layer1[60][47:40] = buffer_data_5[3063:3056];
        layer1[60][55:48] = buffer_data_5[3071:3064];
        layer2[60][7:0] = buffer_data_4[3023:3016];
        layer2[60][15:8] = buffer_data_4[3031:3024];
        layer2[60][23:16] = buffer_data_4[3039:3032];
        layer2[60][31:24] = buffer_data_4[3047:3040];
        layer2[60][39:32] = buffer_data_4[3055:3048];
        layer2[60][47:40] = buffer_data_4[3063:3056];
        layer2[60][55:48] = buffer_data_4[3071:3064];
        layer3[60][7:0] = buffer_data_3[3023:3016];
        layer3[60][15:8] = buffer_data_3[3031:3024];
        layer3[60][23:16] = buffer_data_3[3039:3032];
        layer3[60][31:24] = buffer_data_3[3047:3040];
        layer3[60][39:32] = buffer_data_3[3055:3048];
        layer3[60][47:40] = buffer_data_3[3063:3056];
        layer3[60][55:48] = buffer_data_3[3071:3064];
        layer4[60][7:0] = buffer_data_2[3023:3016];
        layer4[60][15:8] = buffer_data_2[3031:3024];
        layer4[60][23:16] = buffer_data_2[3039:3032];
        layer4[60][31:24] = buffer_data_2[3047:3040];
        layer4[60][39:32] = buffer_data_2[3055:3048];
        layer4[60][47:40] = buffer_data_2[3063:3056];
        layer4[60][55:48] = buffer_data_2[3071:3064];
        layer5[60][7:0] = buffer_data_1[3023:3016];
        layer5[60][15:8] = buffer_data_1[3031:3024];
        layer5[60][23:16] = buffer_data_1[3039:3032];
        layer5[60][31:24] = buffer_data_1[3047:3040];
        layer5[60][39:32] = buffer_data_1[3055:3048];
        layer5[60][47:40] = buffer_data_1[3063:3056];
        layer5[60][55:48] = buffer_data_1[3071:3064];
        layer6[60][7:0] = buffer_data_0[3023:3016];
        layer6[60][15:8] = buffer_data_0[3031:3024];
        layer6[60][23:16] = buffer_data_0[3039:3032];
        layer6[60][31:24] = buffer_data_0[3047:3040];
        layer6[60][39:32] = buffer_data_0[3055:3048];
        layer6[60][47:40] = buffer_data_0[3063:3056];
        layer6[60][55:48] = buffer_data_0[3071:3064];
        layer0[61][7:0] = buffer_data_6[3031:3024];
        layer0[61][15:8] = buffer_data_6[3039:3032];
        layer0[61][23:16] = buffer_data_6[3047:3040];
        layer0[61][31:24] = buffer_data_6[3055:3048];
        layer0[61][39:32] = buffer_data_6[3063:3056];
        layer0[61][47:40] = buffer_data_6[3071:3064];
        layer0[61][55:48] = buffer_data_6[3079:3072];
        layer1[61][7:0] = buffer_data_5[3031:3024];
        layer1[61][15:8] = buffer_data_5[3039:3032];
        layer1[61][23:16] = buffer_data_5[3047:3040];
        layer1[61][31:24] = buffer_data_5[3055:3048];
        layer1[61][39:32] = buffer_data_5[3063:3056];
        layer1[61][47:40] = buffer_data_5[3071:3064];
        layer1[61][55:48] = buffer_data_5[3079:3072];
        layer2[61][7:0] = buffer_data_4[3031:3024];
        layer2[61][15:8] = buffer_data_4[3039:3032];
        layer2[61][23:16] = buffer_data_4[3047:3040];
        layer2[61][31:24] = buffer_data_4[3055:3048];
        layer2[61][39:32] = buffer_data_4[3063:3056];
        layer2[61][47:40] = buffer_data_4[3071:3064];
        layer2[61][55:48] = buffer_data_4[3079:3072];
        layer3[61][7:0] = buffer_data_3[3031:3024];
        layer3[61][15:8] = buffer_data_3[3039:3032];
        layer3[61][23:16] = buffer_data_3[3047:3040];
        layer3[61][31:24] = buffer_data_3[3055:3048];
        layer3[61][39:32] = buffer_data_3[3063:3056];
        layer3[61][47:40] = buffer_data_3[3071:3064];
        layer3[61][55:48] = buffer_data_3[3079:3072];
        layer4[61][7:0] = buffer_data_2[3031:3024];
        layer4[61][15:8] = buffer_data_2[3039:3032];
        layer4[61][23:16] = buffer_data_2[3047:3040];
        layer4[61][31:24] = buffer_data_2[3055:3048];
        layer4[61][39:32] = buffer_data_2[3063:3056];
        layer4[61][47:40] = buffer_data_2[3071:3064];
        layer4[61][55:48] = buffer_data_2[3079:3072];
        layer5[61][7:0] = buffer_data_1[3031:3024];
        layer5[61][15:8] = buffer_data_1[3039:3032];
        layer5[61][23:16] = buffer_data_1[3047:3040];
        layer5[61][31:24] = buffer_data_1[3055:3048];
        layer5[61][39:32] = buffer_data_1[3063:3056];
        layer5[61][47:40] = buffer_data_1[3071:3064];
        layer5[61][55:48] = buffer_data_1[3079:3072];
        layer6[61][7:0] = buffer_data_0[3031:3024];
        layer6[61][15:8] = buffer_data_0[3039:3032];
        layer6[61][23:16] = buffer_data_0[3047:3040];
        layer6[61][31:24] = buffer_data_0[3055:3048];
        layer6[61][39:32] = buffer_data_0[3063:3056];
        layer6[61][47:40] = buffer_data_0[3071:3064];
        layer6[61][55:48] = buffer_data_0[3079:3072];
        layer0[62][7:0] = buffer_data_6[3039:3032];
        layer0[62][15:8] = buffer_data_6[3047:3040];
        layer0[62][23:16] = buffer_data_6[3055:3048];
        layer0[62][31:24] = buffer_data_6[3063:3056];
        layer0[62][39:32] = buffer_data_6[3071:3064];
        layer0[62][47:40] = buffer_data_6[3079:3072];
        layer0[62][55:48] = buffer_data_6[3087:3080];
        layer1[62][7:0] = buffer_data_5[3039:3032];
        layer1[62][15:8] = buffer_data_5[3047:3040];
        layer1[62][23:16] = buffer_data_5[3055:3048];
        layer1[62][31:24] = buffer_data_5[3063:3056];
        layer1[62][39:32] = buffer_data_5[3071:3064];
        layer1[62][47:40] = buffer_data_5[3079:3072];
        layer1[62][55:48] = buffer_data_5[3087:3080];
        layer2[62][7:0] = buffer_data_4[3039:3032];
        layer2[62][15:8] = buffer_data_4[3047:3040];
        layer2[62][23:16] = buffer_data_4[3055:3048];
        layer2[62][31:24] = buffer_data_4[3063:3056];
        layer2[62][39:32] = buffer_data_4[3071:3064];
        layer2[62][47:40] = buffer_data_4[3079:3072];
        layer2[62][55:48] = buffer_data_4[3087:3080];
        layer3[62][7:0] = buffer_data_3[3039:3032];
        layer3[62][15:8] = buffer_data_3[3047:3040];
        layer3[62][23:16] = buffer_data_3[3055:3048];
        layer3[62][31:24] = buffer_data_3[3063:3056];
        layer3[62][39:32] = buffer_data_3[3071:3064];
        layer3[62][47:40] = buffer_data_3[3079:3072];
        layer3[62][55:48] = buffer_data_3[3087:3080];
        layer4[62][7:0] = buffer_data_2[3039:3032];
        layer4[62][15:8] = buffer_data_2[3047:3040];
        layer4[62][23:16] = buffer_data_2[3055:3048];
        layer4[62][31:24] = buffer_data_2[3063:3056];
        layer4[62][39:32] = buffer_data_2[3071:3064];
        layer4[62][47:40] = buffer_data_2[3079:3072];
        layer4[62][55:48] = buffer_data_2[3087:3080];
        layer5[62][7:0] = buffer_data_1[3039:3032];
        layer5[62][15:8] = buffer_data_1[3047:3040];
        layer5[62][23:16] = buffer_data_1[3055:3048];
        layer5[62][31:24] = buffer_data_1[3063:3056];
        layer5[62][39:32] = buffer_data_1[3071:3064];
        layer5[62][47:40] = buffer_data_1[3079:3072];
        layer5[62][55:48] = buffer_data_1[3087:3080];
        layer6[62][7:0] = buffer_data_0[3039:3032];
        layer6[62][15:8] = buffer_data_0[3047:3040];
        layer6[62][23:16] = buffer_data_0[3055:3048];
        layer6[62][31:24] = buffer_data_0[3063:3056];
        layer6[62][39:32] = buffer_data_0[3071:3064];
        layer6[62][47:40] = buffer_data_0[3079:3072];
        layer6[62][55:48] = buffer_data_0[3087:3080];
        layer0[63][7:0] = buffer_data_6[3047:3040];
        layer0[63][15:8] = buffer_data_6[3055:3048];
        layer0[63][23:16] = buffer_data_6[3063:3056];
        layer0[63][31:24] = buffer_data_6[3071:3064];
        layer0[63][39:32] = buffer_data_6[3079:3072];
        layer0[63][47:40] = buffer_data_6[3087:3080];
        layer0[63][55:48] = buffer_data_6[3095:3088];
        layer1[63][7:0] = buffer_data_5[3047:3040];
        layer1[63][15:8] = buffer_data_5[3055:3048];
        layer1[63][23:16] = buffer_data_5[3063:3056];
        layer1[63][31:24] = buffer_data_5[3071:3064];
        layer1[63][39:32] = buffer_data_5[3079:3072];
        layer1[63][47:40] = buffer_data_5[3087:3080];
        layer1[63][55:48] = buffer_data_5[3095:3088];
        layer2[63][7:0] = buffer_data_4[3047:3040];
        layer2[63][15:8] = buffer_data_4[3055:3048];
        layer2[63][23:16] = buffer_data_4[3063:3056];
        layer2[63][31:24] = buffer_data_4[3071:3064];
        layer2[63][39:32] = buffer_data_4[3079:3072];
        layer2[63][47:40] = buffer_data_4[3087:3080];
        layer2[63][55:48] = buffer_data_4[3095:3088];
        layer3[63][7:0] = buffer_data_3[3047:3040];
        layer3[63][15:8] = buffer_data_3[3055:3048];
        layer3[63][23:16] = buffer_data_3[3063:3056];
        layer3[63][31:24] = buffer_data_3[3071:3064];
        layer3[63][39:32] = buffer_data_3[3079:3072];
        layer3[63][47:40] = buffer_data_3[3087:3080];
        layer3[63][55:48] = buffer_data_3[3095:3088];
        layer4[63][7:0] = buffer_data_2[3047:3040];
        layer4[63][15:8] = buffer_data_2[3055:3048];
        layer4[63][23:16] = buffer_data_2[3063:3056];
        layer4[63][31:24] = buffer_data_2[3071:3064];
        layer4[63][39:32] = buffer_data_2[3079:3072];
        layer4[63][47:40] = buffer_data_2[3087:3080];
        layer4[63][55:48] = buffer_data_2[3095:3088];
        layer5[63][7:0] = buffer_data_1[3047:3040];
        layer5[63][15:8] = buffer_data_1[3055:3048];
        layer5[63][23:16] = buffer_data_1[3063:3056];
        layer5[63][31:24] = buffer_data_1[3071:3064];
        layer5[63][39:32] = buffer_data_1[3079:3072];
        layer5[63][47:40] = buffer_data_1[3087:3080];
        layer5[63][55:48] = buffer_data_1[3095:3088];
        layer6[63][7:0] = buffer_data_0[3047:3040];
        layer6[63][15:8] = buffer_data_0[3055:3048];
        layer6[63][23:16] = buffer_data_0[3063:3056];
        layer6[63][31:24] = buffer_data_0[3071:3064];
        layer6[63][39:32] = buffer_data_0[3079:3072];
        layer6[63][47:40] = buffer_data_0[3087:3080];
        layer6[63][55:48] = buffer_data_0[3095:3088];
    end
    ST_GAUSSIAN_6: begin
        layer0[0][7:0] = buffer_data_6[3055:3048];
        layer0[0][15:8] = buffer_data_6[3063:3056];
        layer0[0][23:16] = buffer_data_6[3071:3064];
        layer0[0][31:24] = buffer_data_6[3079:3072];
        layer0[0][39:32] = buffer_data_6[3087:3080];
        layer0[0][47:40] = buffer_data_6[3095:3088];
        layer0[0][55:48] = buffer_data_6[3103:3096];
        layer1[0][7:0] = buffer_data_5[3055:3048];
        layer1[0][15:8] = buffer_data_5[3063:3056];
        layer1[0][23:16] = buffer_data_5[3071:3064];
        layer1[0][31:24] = buffer_data_5[3079:3072];
        layer1[0][39:32] = buffer_data_5[3087:3080];
        layer1[0][47:40] = buffer_data_5[3095:3088];
        layer1[0][55:48] = buffer_data_5[3103:3096];
        layer2[0][7:0] = buffer_data_4[3055:3048];
        layer2[0][15:8] = buffer_data_4[3063:3056];
        layer2[0][23:16] = buffer_data_4[3071:3064];
        layer2[0][31:24] = buffer_data_4[3079:3072];
        layer2[0][39:32] = buffer_data_4[3087:3080];
        layer2[0][47:40] = buffer_data_4[3095:3088];
        layer2[0][55:48] = buffer_data_4[3103:3096];
        layer3[0][7:0] = buffer_data_3[3055:3048];
        layer3[0][15:8] = buffer_data_3[3063:3056];
        layer3[0][23:16] = buffer_data_3[3071:3064];
        layer3[0][31:24] = buffer_data_3[3079:3072];
        layer3[0][39:32] = buffer_data_3[3087:3080];
        layer3[0][47:40] = buffer_data_3[3095:3088];
        layer3[0][55:48] = buffer_data_3[3103:3096];
        layer4[0][7:0] = buffer_data_2[3055:3048];
        layer4[0][15:8] = buffer_data_2[3063:3056];
        layer4[0][23:16] = buffer_data_2[3071:3064];
        layer4[0][31:24] = buffer_data_2[3079:3072];
        layer4[0][39:32] = buffer_data_2[3087:3080];
        layer4[0][47:40] = buffer_data_2[3095:3088];
        layer4[0][55:48] = buffer_data_2[3103:3096];
        layer5[0][7:0] = buffer_data_1[3055:3048];
        layer5[0][15:8] = buffer_data_1[3063:3056];
        layer5[0][23:16] = buffer_data_1[3071:3064];
        layer5[0][31:24] = buffer_data_1[3079:3072];
        layer5[0][39:32] = buffer_data_1[3087:3080];
        layer5[0][47:40] = buffer_data_1[3095:3088];
        layer5[0][55:48] = buffer_data_1[3103:3096];
        layer6[0][7:0] = buffer_data_0[3055:3048];
        layer6[0][15:8] = buffer_data_0[3063:3056];
        layer6[0][23:16] = buffer_data_0[3071:3064];
        layer6[0][31:24] = buffer_data_0[3079:3072];
        layer6[0][39:32] = buffer_data_0[3087:3080];
        layer6[0][47:40] = buffer_data_0[3095:3088];
        layer6[0][55:48] = buffer_data_0[3103:3096];
        layer0[1][7:0] = buffer_data_6[3063:3056];
        layer0[1][15:8] = buffer_data_6[3071:3064];
        layer0[1][23:16] = buffer_data_6[3079:3072];
        layer0[1][31:24] = buffer_data_6[3087:3080];
        layer0[1][39:32] = buffer_data_6[3095:3088];
        layer0[1][47:40] = buffer_data_6[3103:3096];
        layer0[1][55:48] = buffer_data_6[3111:3104];
        layer1[1][7:0] = buffer_data_5[3063:3056];
        layer1[1][15:8] = buffer_data_5[3071:3064];
        layer1[1][23:16] = buffer_data_5[3079:3072];
        layer1[1][31:24] = buffer_data_5[3087:3080];
        layer1[1][39:32] = buffer_data_5[3095:3088];
        layer1[1][47:40] = buffer_data_5[3103:3096];
        layer1[1][55:48] = buffer_data_5[3111:3104];
        layer2[1][7:0] = buffer_data_4[3063:3056];
        layer2[1][15:8] = buffer_data_4[3071:3064];
        layer2[1][23:16] = buffer_data_4[3079:3072];
        layer2[1][31:24] = buffer_data_4[3087:3080];
        layer2[1][39:32] = buffer_data_4[3095:3088];
        layer2[1][47:40] = buffer_data_4[3103:3096];
        layer2[1][55:48] = buffer_data_4[3111:3104];
        layer3[1][7:0] = buffer_data_3[3063:3056];
        layer3[1][15:8] = buffer_data_3[3071:3064];
        layer3[1][23:16] = buffer_data_3[3079:3072];
        layer3[1][31:24] = buffer_data_3[3087:3080];
        layer3[1][39:32] = buffer_data_3[3095:3088];
        layer3[1][47:40] = buffer_data_3[3103:3096];
        layer3[1][55:48] = buffer_data_3[3111:3104];
        layer4[1][7:0] = buffer_data_2[3063:3056];
        layer4[1][15:8] = buffer_data_2[3071:3064];
        layer4[1][23:16] = buffer_data_2[3079:3072];
        layer4[1][31:24] = buffer_data_2[3087:3080];
        layer4[1][39:32] = buffer_data_2[3095:3088];
        layer4[1][47:40] = buffer_data_2[3103:3096];
        layer4[1][55:48] = buffer_data_2[3111:3104];
        layer5[1][7:0] = buffer_data_1[3063:3056];
        layer5[1][15:8] = buffer_data_1[3071:3064];
        layer5[1][23:16] = buffer_data_1[3079:3072];
        layer5[1][31:24] = buffer_data_1[3087:3080];
        layer5[1][39:32] = buffer_data_1[3095:3088];
        layer5[1][47:40] = buffer_data_1[3103:3096];
        layer5[1][55:48] = buffer_data_1[3111:3104];
        layer6[1][7:0] = buffer_data_0[3063:3056];
        layer6[1][15:8] = buffer_data_0[3071:3064];
        layer6[1][23:16] = buffer_data_0[3079:3072];
        layer6[1][31:24] = buffer_data_0[3087:3080];
        layer6[1][39:32] = buffer_data_0[3095:3088];
        layer6[1][47:40] = buffer_data_0[3103:3096];
        layer6[1][55:48] = buffer_data_0[3111:3104];
        layer0[2][7:0] = buffer_data_6[3071:3064];
        layer0[2][15:8] = buffer_data_6[3079:3072];
        layer0[2][23:16] = buffer_data_6[3087:3080];
        layer0[2][31:24] = buffer_data_6[3095:3088];
        layer0[2][39:32] = buffer_data_6[3103:3096];
        layer0[2][47:40] = buffer_data_6[3111:3104];
        layer0[2][55:48] = buffer_data_6[3119:3112];
        layer1[2][7:0] = buffer_data_5[3071:3064];
        layer1[2][15:8] = buffer_data_5[3079:3072];
        layer1[2][23:16] = buffer_data_5[3087:3080];
        layer1[2][31:24] = buffer_data_5[3095:3088];
        layer1[2][39:32] = buffer_data_5[3103:3096];
        layer1[2][47:40] = buffer_data_5[3111:3104];
        layer1[2][55:48] = buffer_data_5[3119:3112];
        layer2[2][7:0] = buffer_data_4[3071:3064];
        layer2[2][15:8] = buffer_data_4[3079:3072];
        layer2[2][23:16] = buffer_data_4[3087:3080];
        layer2[2][31:24] = buffer_data_4[3095:3088];
        layer2[2][39:32] = buffer_data_4[3103:3096];
        layer2[2][47:40] = buffer_data_4[3111:3104];
        layer2[2][55:48] = buffer_data_4[3119:3112];
        layer3[2][7:0] = buffer_data_3[3071:3064];
        layer3[2][15:8] = buffer_data_3[3079:3072];
        layer3[2][23:16] = buffer_data_3[3087:3080];
        layer3[2][31:24] = buffer_data_3[3095:3088];
        layer3[2][39:32] = buffer_data_3[3103:3096];
        layer3[2][47:40] = buffer_data_3[3111:3104];
        layer3[2][55:48] = buffer_data_3[3119:3112];
        layer4[2][7:0] = buffer_data_2[3071:3064];
        layer4[2][15:8] = buffer_data_2[3079:3072];
        layer4[2][23:16] = buffer_data_2[3087:3080];
        layer4[2][31:24] = buffer_data_2[3095:3088];
        layer4[2][39:32] = buffer_data_2[3103:3096];
        layer4[2][47:40] = buffer_data_2[3111:3104];
        layer4[2][55:48] = buffer_data_2[3119:3112];
        layer5[2][7:0] = buffer_data_1[3071:3064];
        layer5[2][15:8] = buffer_data_1[3079:3072];
        layer5[2][23:16] = buffer_data_1[3087:3080];
        layer5[2][31:24] = buffer_data_1[3095:3088];
        layer5[2][39:32] = buffer_data_1[3103:3096];
        layer5[2][47:40] = buffer_data_1[3111:3104];
        layer5[2][55:48] = buffer_data_1[3119:3112];
        layer6[2][7:0] = buffer_data_0[3071:3064];
        layer6[2][15:8] = buffer_data_0[3079:3072];
        layer6[2][23:16] = buffer_data_0[3087:3080];
        layer6[2][31:24] = buffer_data_0[3095:3088];
        layer6[2][39:32] = buffer_data_0[3103:3096];
        layer6[2][47:40] = buffer_data_0[3111:3104];
        layer6[2][55:48] = buffer_data_0[3119:3112];
        layer0[3][7:0] = buffer_data_6[3079:3072];
        layer0[3][15:8] = buffer_data_6[3087:3080];
        layer0[3][23:16] = buffer_data_6[3095:3088];
        layer0[3][31:24] = buffer_data_6[3103:3096];
        layer0[3][39:32] = buffer_data_6[3111:3104];
        layer0[3][47:40] = buffer_data_6[3119:3112];
        layer0[3][55:48] = buffer_data_6[3127:3120];
        layer1[3][7:0] = buffer_data_5[3079:3072];
        layer1[3][15:8] = buffer_data_5[3087:3080];
        layer1[3][23:16] = buffer_data_5[3095:3088];
        layer1[3][31:24] = buffer_data_5[3103:3096];
        layer1[3][39:32] = buffer_data_5[3111:3104];
        layer1[3][47:40] = buffer_data_5[3119:3112];
        layer1[3][55:48] = buffer_data_5[3127:3120];
        layer2[3][7:0] = buffer_data_4[3079:3072];
        layer2[3][15:8] = buffer_data_4[3087:3080];
        layer2[3][23:16] = buffer_data_4[3095:3088];
        layer2[3][31:24] = buffer_data_4[3103:3096];
        layer2[3][39:32] = buffer_data_4[3111:3104];
        layer2[3][47:40] = buffer_data_4[3119:3112];
        layer2[3][55:48] = buffer_data_4[3127:3120];
        layer3[3][7:0] = buffer_data_3[3079:3072];
        layer3[3][15:8] = buffer_data_3[3087:3080];
        layer3[3][23:16] = buffer_data_3[3095:3088];
        layer3[3][31:24] = buffer_data_3[3103:3096];
        layer3[3][39:32] = buffer_data_3[3111:3104];
        layer3[3][47:40] = buffer_data_3[3119:3112];
        layer3[3][55:48] = buffer_data_3[3127:3120];
        layer4[3][7:0] = buffer_data_2[3079:3072];
        layer4[3][15:8] = buffer_data_2[3087:3080];
        layer4[3][23:16] = buffer_data_2[3095:3088];
        layer4[3][31:24] = buffer_data_2[3103:3096];
        layer4[3][39:32] = buffer_data_2[3111:3104];
        layer4[3][47:40] = buffer_data_2[3119:3112];
        layer4[3][55:48] = buffer_data_2[3127:3120];
        layer5[3][7:0] = buffer_data_1[3079:3072];
        layer5[3][15:8] = buffer_data_1[3087:3080];
        layer5[3][23:16] = buffer_data_1[3095:3088];
        layer5[3][31:24] = buffer_data_1[3103:3096];
        layer5[3][39:32] = buffer_data_1[3111:3104];
        layer5[3][47:40] = buffer_data_1[3119:3112];
        layer5[3][55:48] = buffer_data_1[3127:3120];
        layer6[3][7:0] = buffer_data_0[3079:3072];
        layer6[3][15:8] = buffer_data_0[3087:3080];
        layer6[3][23:16] = buffer_data_0[3095:3088];
        layer6[3][31:24] = buffer_data_0[3103:3096];
        layer6[3][39:32] = buffer_data_0[3111:3104];
        layer6[3][47:40] = buffer_data_0[3119:3112];
        layer6[3][55:48] = buffer_data_0[3127:3120];
        layer0[4][7:0] = buffer_data_6[3087:3080];
        layer0[4][15:8] = buffer_data_6[3095:3088];
        layer0[4][23:16] = buffer_data_6[3103:3096];
        layer0[4][31:24] = buffer_data_6[3111:3104];
        layer0[4][39:32] = buffer_data_6[3119:3112];
        layer0[4][47:40] = buffer_data_6[3127:3120];
        layer0[4][55:48] = buffer_data_6[3135:3128];
        layer1[4][7:0] = buffer_data_5[3087:3080];
        layer1[4][15:8] = buffer_data_5[3095:3088];
        layer1[4][23:16] = buffer_data_5[3103:3096];
        layer1[4][31:24] = buffer_data_5[3111:3104];
        layer1[4][39:32] = buffer_data_5[3119:3112];
        layer1[4][47:40] = buffer_data_5[3127:3120];
        layer1[4][55:48] = buffer_data_5[3135:3128];
        layer2[4][7:0] = buffer_data_4[3087:3080];
        layer2[4][15:8] = buffer_data_4[3095:3088];
        layer2[4][23:16] = buffer_data_4[3103:3096];
        layer2[4][31:24] = buffer_data_4[3111:3104];
        layer2[4][39:32] = buffer_data_4[3119:3112];
        layer2[4][47:40] = buffer_data_4[3127:3120];
        layer2[4][55:48] = buffer_data_4[3135:3128];
        layer3[4][7:0] = buffer_data_3[3087:3080];
        layer3[4][15:8] = buffer_data_3[3095:3088];
        layer3[4][23:16] = buffer_data_3[3103:3096];
        layer3[4][31:24] = buffer_data_3[3111:3104];
        layer3[4][39:32] = buffer_data_3[3119:3112];
        layer3[4][47:40] = buffer_data_3[3127:3120];
        layer3[4][55:48] = buffer_data_3[3135:3128];
        layer4[4][7:0] = buffer_data_2[3087:3080];
        layer4[4][15:8] = buffer_data_2[3095:3088];
        layer4[4][23:16] = buffer_data_2[3103:3096];
        layer4[4][31:24] = buffer_data_2[3111:3104];
        layer4[4][39:32] = buffer_data_2[3119:3112];
        layer4[4][47:40] = buffer_data_2[3127:3120];
        layer4[4][55:48] = buffer_data_2[3135:3128];
        layer5[4][7:0] = buffer_data_1[3087:3080];
        layer5[4][15:8] = buffer_data_1[3095:3088];
        layer5[4][23:16] = buffer_data_1[3103:3096];
        layer5[4][31:24] = buffer_data_1[3111:3104];
        layer5[4][39:32] = buffer_data_1[3119:3112];
        layer5[4][47:40] = buffer_data_1[3127:3120];
        layer5[4][55:48] = buffer_data_1[3135:3128];
        layer6[4][7:0] = buffer_data_0[3087:3080];
        layer6[4][15:8] = buffer_data_0[3095:3088];
        layer6[4][23:16] = buffer_data_0[3103:3096];
        layer6[4][31:24] = buffer_data_0[3111:3104];
        layer6[4][39:32] = buffer_data_0[3119:3112];
        layer6[4][47:40] = buffer_data_0[3127:3120];
        layer6[4][55:48] = buffer_data_0[3135:3128];
        layer0[5][7:0] = buffer_data_6[3095:3088];
        layer0[5][15:8] = buffer_data_6[3103:3096];
        layer0[5][23:16] = buffer_data_6[3111:3104];
        layer0[5][31:24] = buffer_data_6[3119:3112];
        layer0[5][39:32] = buffer_data_6[3127:3120];
        layer0[5][47:40] = buffer_data_6[3135:3128];
        layer0[5][55:48] = buffer_data_6[3143:3136];
        layer1[5][7:0] = buffer_data_5[3095:3088];
        layer1[5][15:8] = buffer_data_5[3103:3096];
        layer1[5][23:16] = buffer_data_5[3111:3104];
        layer1[5][31:24] = buffer_data_5[3119:3112];
        layer1[5][39:32] = buffer_data_5[3127:3120];
        layer1[5][47:40] = buffer_data_5[3135:3128];
        layer1[5][55:48] = buffer_data_5[3143:3136];
        layer2[5][7:0] = buffer_data_4[3095:3088];
        layer2[5][15:8] = buffer_data_4[3103:3096];
        layer2[5][23:16] = buffer_data_4[3111:3104];
        layer2[5][31:24] = buffer_data_4[3119:3112];
        layer2[5][39:32] = buffer_data_4[3127:3120];
        layer2[5][47:40] = buffer_data_4[3135:3128];
        layer2[5][55:48] = buffer_data_4[3143:3136];
        layer3[5][7:0] = buffer_data_3[3095:3088];
        layer3[5][15:8] = buffer_data_3[3103:3096];
        layer3[5][23:16] = buffer_data_3[3111:3104];
        layer3[5][31:24] = buffer_data_3[3119:3112];
        layer3[5][39:32] = buffer_data_3[3127:3120];
        layer3[5][47:40] = buffer_data_3[3135:3128];
        layer3[5][55:48] = buffer_data_3[3143:3136];
        layer4[5][7:0] = buffer_data_2[3095:3088];
        layer4[5][15:8] = buffer_data_2[3103:3096];
        layer4[5][23:16] = buffer_data_2[3111:3104];
        layer4[5][31:24] = buffer_data_2[3119:3112];
        layer4[5][39:32] = buffer_data_2[3127:3120];
        layer4[5][47:40] = buffer_data_2[3135:3128];
        layer4[5][55:48] = buffer_data_2[3143:3136];
        layer5[5][7:0] = buffer_data_1[3095:3088];
        layer5[5][15:8] = buffer_data_1[3103:3096];
        layer5[5][23:16] = buffer_data_1[3111:3104];
        layer5[5][31:24] = buffer_data_1[3119:3112];
        layer5[5][39:32] = buffer_data_1[3127:3120];
        layer5[5][47:40] = buffer_data_1[3135:3128];
        layer5[5][55:48] = buffer_data_1[3143:3136];
        layer6[5][7:0] = buffer_data_0[3095:3088];
        layer6[5][15:8] = buffer_data_0[3103:3096];
        layer6[5][23:16] = buffer_data_0[3111:3104];
        layer6[5][31:24] = buffer_data_0[3119:3112];
        layer6[5][39:32] = buffer_data_0[3127:3120];
        layer6[5][47:40] = buffer_data_0[3135:3128];
        layer6[5][55:48] = buffer_data_0[3143:3136];
        layer0[6][7:0] = buffer_data_6[3103:3096];
        layer0[6][15:8] = buffer_data_6[3111:3104];
        layer0[6][23:16] = buffer_data_6[3119:3112];
        layer0[6][31:24] = buffer_data_6[3127:3120];
        layer0[6][39:32] = buffer_data_6[3135:3128];
        layer0[6][47:40] = buffer_data_6[3143:3136];
        layer0[6][55:48] = buffer_data_6[3151:3144];
        layer1[6][7:0] = buffer_data_5[3103:3096];
        layer1[6][15:8] = buffer_data_5[3111:3104];
        layer1[6][23:16] = buffer_data_5[3119:3112];
        layer1[6][31:24] = buffer_data_5[3127:3120];
        layer1[6][39:32] = buffer_data_5[3135:3128];
        layer1[6][47:40] = buffer_data_5[3143:3136];
        layer1[6][55:48] = buffer_data_5[3151:3144];
        layer2[6][7:0] = buffer_data_4[3103:3096];
        layer2[6][15:8] = buffer_data_4[3111:3104];
        layer2[6][23:16] = buffer_data_4[3119:3112];
        layer2[6][31:24] = buffer_data_4[3127:3120];
        layer2[6][39:32] = buffer_data_4[3135:3128];
        layer2[6][47:40] = buffer_data_4[3143:3136];
        layer2[6][55:48] = buffer_data_4[3151:3144];
        layer3[6][7:0] = buffer_data_3[3103:3096];
        layer3[6][15:8] = buffer_data_3[3111:3104];
        layer3[6][23:16] = buffer_data_3[3119:3112];
        layer3[6][31:24] = buffer_data_3[3127:3120];
        layer3[6][39:32] = buffer_data_3[3135:3128];
        layer3[6][47:40] = buffer_data_3[3143:3136];
        layer3[6][55:48] = buffer_data_3[3151:3144];
        layer4[6][7:0] = buffer_data_2[3103:3096];
        layer4[6][15:8] = buffer_data_2[3111:3104];
        layer4[6][23:16] = buffer_data_2[3119:3112];
        layer4[6][31:24] = buffer_data_2[3127:3120];
        layer4[6][39:32] = buffer_data_2[3135:3128];
        layer4[6][47:40] = buffer_data_2[3143:3136];
        layer4[6][55:48] = buffer_data_2[3151:3144];
        layer5[6][7:0] = buffer_data_1[3103:3096];
        layer5[6][15:8] = buffer_data_1[3111:3104];
        layer5[6][23:16] = buffer_data_1[3119:3112];
        layer5[6][31:24] = buffer_data_1[3127:3120];
        layer5[6][39:32] = buffer_data_1[3135:3128];
        layer5[6][47:40] = buffer_data_1[3143:3136];
        layer5[6][55:48] = buffer_data_1[3151:3144];
        layer6[6][7:0] = buffer_data_0[3103:3096];
        layer6[6][15:8] = buffer_data_0[3111:3104];
        layer6[6][23:16] = buffer_data_0[3119:3112];
        layer6[6][31:24] = buffer_data_0[3127:3120];
        layer6[6][39:32] = buffer_data_0[3135:3128];
        layer6[6][47:40] = buffer_data_0[3143:3136];
        layer6[6][55:48] = buffer_data_0[3151:3144];
        layer0[7][7:0] = buffer_data_6[3111:3104];
        layer0[7][15:8] = buffer_data_6[3119:3112];
        layer0[7][23:16] = buffer_data_6[3127:3120];
        layer0[7][31:24] = buffer_data_6[3135:3128];
        layer0[7][39:32] = buffer_data_6[3143:3136];
        layer0[7][47:40] = buffer_data_6[3151:3144];
        layer0[7][55:48] = buffer_data_6[3159:3152];
        layer1[7][7:0] = buffer_data_5[3111:3104];
        layer1[7][15:8] = buffer_data_5[3119:3112];
        layer1[7][23:16] = buffer_data_5[3127:3120];
        layer1[7][31:24] = buffer_data_5[3135:3128];
        layer1[7][39:32] = buffer_data_5[3143:3136];
        layer1[7][47:40] = buffer_data_5[3151:3144];
        layer1[7][55:48] = buffer_data_5[3159:3152];
        layer2[7][7:0] = buffer_data_4[3111:3104];
        layer2[7][15:8] = buffer_data_4[3119:3112];
        layer2[7][23:16] = buffer_data_4[3127:3120];
        layer2[7][31:24] = buffer_data_4[3135:3128];
        layer2[7][39:32] = buffer_data_4[3143:3136];
        layer2[7][47:40] = buffer_data_4[3151:3144];
        layer2[7][55:48] = buffer_data_4[3159:3152];
        layer3[7][7:0] = buffer_data_3[3111:3104];
        layer3[7][15:8] = buffer_data_3[3119:3112];
        layer3[7][23:16] = buffer_data_3[3127:3120];
        layer3[7][31:24] = buffer_data_3[3135:3128];
        layer3[7][39:32] = buffer_data_3[3143:3136];
        layer3[7][47:40] = buffer_data_3[3151:3144];
        layer3[7][55:48] = buffer_data_3[3159:3152];
        layer4[7][7:0] = buffer_data_2[3111:3104];
        layer4[7][15:8] = buffer_data_2[3119:3112];
        layer4[7][23:16] = buffer_data_2[3127:3120];
        layer4[7][31:24] = buffer_data_2[3135:3128];
        layer4[7][39:32] = buffer_data_2[3143:3136];
        layer4[7][47:40] = buffer_data_2[3151:3144];
        layer4[7][55:48] = buffer_data_2[3159:3152];
        layer5[7][7:0] = buffer_data_1[3111:3104];
        layer5[7][15:8] = buffer_data_1[3119:3112];
        layer5[7][23:16] = buffer_data_1[3127:3120];
        layer5[7][31:24] = buffer_data_1[3135:3128];
        layer5[7][39:32] = buffer_data_1[3143:3136];
        layer5[7][47:40] = buffer_data_1[3151:3144];
        layer5[7][55:48] = buffer_data_1[3159:3152];
        layer6[7][7:0] = buffer_data_0[3111:3104];
        layer6[7][15:8] = buffer_data_0[3119:3112];
        layer6[7][23:16] = buffer_data_0[3127:3120];
        layer6[7][31:24] = buffer_data_0[3135:3128];
        layer6[7][39:32] = buffer_data_0[3143:3136];
        layer6[7][47:40] = buffer_data_0[3151:3144];
        layer6[7][55:48] = buffer_data_0[3159:3152];
        layer0[8][7:0] = buffer_data_6[3119:3112];
        layer0[8][15:8] = buffer_data_6[3127:3120];
        layer0[8][23:16] = buffer_data_6[3135:3128];
        layer0[8][31:24] = buffer_data_6[3143:3136];
        layer0[8][39:32] = buffer_data_6[3151:3144];
        layer0[8][47:40] = buffer_data_6[3159:3152];
        layer0[8][55:48] = buffer_data_6[3167:3160];
        layer1[8][7:0] = buffer_data_5[3119:3112];
        layer1[8][15:8] = buffer_data_5[3127:3120];
        layer1[8][23:16] = buffer_data_5[3135:3128];
        layer1[8][31:24] = buffer_data_5[3143:3136];
        layer1[8][39:32] = buffer_data_5[3151:3144];
        layer1[8][47:40] = buffer_data_5[3159:3152];
        layer1[8][55:48] = buffer_data_5[3167:3160];
        layer2[8][7:0] = buffer_data_4[3119:3112];
        layer2[8][15:8] = buffer_data_4[3127:3120];
        layer2[8][23:16] = buffer_data_4[3135:3128];
        layer2[8][31:24] = buffer_data_4[3143:3136];
        layer2[8][39:32] = buffer_data_4[3151:3144];
        layer2[8][47:40] = buffer_data_4[3159:3152];
        layer2[8][55:48] = buffer_data_4[3167:3160];
        layer3[8][7:0] = buffer_data_3[3119:3112];
        layer3[8][15:8] = buffer_data_3[3127:3120];
        layer3[8][23:16] = buffer_data_3[3135:3128];
        layer3[8][31:24] = buffer_data_3[3143:3136];
        layer3[8][39:32] = buffer_data_3[3151:3144];
        layer3[8][47:40] = buffer_data_3[3159:3152];
        layer3[8][55:48] = buffer_data_3[3167:3160];
        layer4[8][7:0] = buffer_data_2[3119:3112];
        layer4[8][15:8] = buffer_data_2[3127:3120];
        layer4[8][23:16] = buffer_data_2[3135:3128];
        layer4[8][31:24] = buffer_data_2[3143:3136];
        layer4[8][39:32] = buffer_data_2[3151:3144];
        layer4[8][47:40] = buffer_data_2[3159:3152];
        layer4[8][55:48] = buffer_data_2[3167:3160];
        layer5[8][7:0] = buffer_data_1[3119:3112];
        layer5[8][15:8] = buffer_data_1[3127:3120];
        layer5[8][23:16] = buffer_data_1[3135:3128];
        layer5[8][31:24] = buffer_data_1[3143:3136];
        layer5[8][39:32] = buffer_data_1[3151:3144];
        layer5[8][47:40] = buffer_data_1[3159:3152];
        layer5[8][55:48] = buffer_data_1[3167:3160];
        layer6[8][7:0] = buffer_data_0[3119:3112];
        layer6[8][15:8] = buffer_data_0[3127:3120];
        layer6[8][23:16] = buffer_data_0[3135:3128];
        layer6[8][31:24] = buffer_data_0[3143:3136];
        layer6[8][39:32] = buffer_data_0[3151:3144];
        layer6[8][47:40] = buffer_data_0[3159:3152];
        layer6[8][55:48] = buffer_data_0[3167:3160];
        layer0[9][7:0] = buffer_data_6[3127:3120];
        layer0[9][15:8] = buffer_data_6[3135:3128];
        layer0[9][23:16] = buffer_data_6[3143:3136];
        layer0[9][31:24] = buffer_data_6[3151:3144];
        layer0[9][39:32] = buffer_data_6[3159:3152];
        layer0[9][47:40] = buffer_data_6[3167:3160];
        layer0[9][55:48] = buffer_data_6[3175:3168];
        layer1[9][7:0] = buffer_data_5[3127:3120];
        layer1[9][15:8] = buffer_data_5[3135:3128];
        layer1[9][23:16] = buffer_data_5[3143:3136];
        layer1[9][31:24] = buffer_data_5[3151:3144];
        layer1[9][39:32] = buffer_data_5[3159:3152];
        layer1[9][47:40] = buffer_data_5[3167:3160];
        layer1[9][55:48] = buffer_data_5[3175:3168];
        layer2[9][7:0] = buffer_data_4[3127:3120];
        layer2[9][15:8] = buffer_data_4[3135:3128];
        layer2[9][23:16] = buffer_data_4[3143:3136];
        layer2[9][31:24] = buffer_data_4[3151:3144];
        layer2[9][39:32] = buffer_data_4[3159:3152];
        layer2[9][47:40] = buffer_data_4[3167:3160];
        layer2[9][55:48] = buffer_data_4[3175:3168];
        layer3[9][7:0] = buffer_data_3[3127:3120];
        layer3[9][15:8] = buffer_data_3[3135:3128];
        layer3[9][23:16] = buffer_data_3[3143:3136];
        layer3[9][31:24] = buffer_data_3[3151:3144];
        layer3[9][39:32] = buffer_data_3[3159:3152];
        layer3[9][47:40] = buffer_data_3[3167:3160];
        layer3[9][55:48] = buffer_data_3[3175:3168];
        layer4[9][7:0] = buffer_data_2[3127:3120];
        layer4[9][15:8] = buffer_data_2[3135:3128];
        layer4[9][23:16] = buffer_data_2[3143:3136];
        layer4[9][31:24] = buffer_data_2[3151:3144];
        layer4[9][39:32] = buffer_data_2[3159:3152];
        layer4[9][47:40] = buffer_data_2[3167:3160];
        layer4[9][55:48] = buffer_data_2[3175:3168];
        layer5[9][7:0] = buffer_data_1[3127:3120];
        layer5[9][15:8] = buffer_data_1[3135:3128];
        layer5[9][23:16] = buffer_data_1[3143:3136];
        layer5[9][31:24] = buffer_data_1[3151:3144];
        layer5[9][39:32] = buffer_data_1[3159:3152];
        layer5[9][47:40] = buffer_data_1[3167:3160];
        layer5[9][55:48] = buffer_data_1[3175:3168];
        layer6[9][7:0] = buffer_data_0[3127:3120];
        layer6[9][15:8] = buffer_data_0[3135:3128];
        layer6[9][23:16] = buffer_data_0[3143:3136];
        layer6[9][31:24] = buffer_data_0[3151:3144];
        layer6[9][39:32] = buffer_data_0[3159:3152];
        layer6[9][47:40] = buffer_data_0[3167:3160];
        layer6[9][55:48] = buffer_data_0[3175:3168];
        layer0[10][7:0] = buffer_data_6[3135:3128];
        layer0[10][15:8] = buffer_data_6[3143:3136];
        layer0[10][23:16] = buffer_data_6[3151:3144];
        layer0[10][31:24] = buffer_data_6[3159:3152];
        layer0[10][39:32] = buffer_data_6[3167:3160];
        layer0[10][47:40] = buffer_data_6[3175:3168];
        layer0[10][55:48] = buffer_data_6[3183:3176];
        layer1[10][7:0] = buffer_data_5[3135:3128];
        layer1[10][15:8] = buffer_data_5[3143:3136];
        layer1[10][23:16] = buffer_data_5[3151:3144];
        layer1[10][31:24] = buffer_data_5[3159:3152];
        layer1[10][39:32] = buffer_data_5[3167:3160];
        layer1[10][47:40] = buffer_data_5[3175:3168];
        layer1[10][55:48] = buffer_data_5[3183:3176];
        layer2[10][7:0] = buffer_data_4[3135:3128];
        layer2[10][15:8] = buffer_data_4[3143:3136];
        layer2[10][23:16] = buffer_data_4[3151:3144];
        layer2[10][31:24] = buffer_data_4[3159:3152];
        layer2[10][39:32] = buffer_data_4[3167:3160];
        layer2[10][47:40] = buffer_data_4[3175:3168];
        layer2[10][55:48] = buffer_data_4[3183:3176];
        layer3[10][7:0] = buffer_data_3[3135:3128];
        layer3[10][15:8] = buffer_data_3[3143:3136];
        layer3[10][23:16] = buffer_data_3[3151:3144];
        layer3[10][31:24] = buffer_data_3[3159:3152];
        layer3[10][39:32] = buffer_data_3[3167:3160];
        layer3[10][47:40] = buffer_data_3[3175:3168];
        layer3[10][55:48] = buffer_data_3[3183:3176];
        layer4[10][7:0] = buffer_data_2[3135:3128];
        layer4[10][15:8] = buffer_data_2[3143:3136];
        layer4[10][23:16] = buffer_data_2[3151:3144];
        layer4[10][31:24] = buffer_data_2[3159:3152];
        layer4[10][39:32] = buffer_data_2[3167:3160];
        layer4[10][47:40] = buffer_data_2[3175:3168];
        layer4[10][55:48] = buffer_data_2[3183:3176];
        layer5[10][7:0] = buffer_data_1[3135:3128];
        layer5[10][15:8] = buffer_data_1[3143:3136];
        layer5[10][23:16] = buffer_data_1[3151:3144];
        layer5[10][31:24] = buffer_data_1[3159:3152];
        layer5[10][39:32] = buffer_data_1[3167:3160];
        layer5[10][47:40] = buffer_data_1[3175:3168];
        layer5[10][55:48] = buffer_data_1[3183:3176];
        layer6[10][7:0] = buffer_data_0[3135:3128];
        layer6[10][15:8] = buffer_data_0[3143:3136];
        layer6[10][23:16] = buffer_data_0[3151:3144];
        layer6[10][31:24] = buffer_data_0[3159:3152];
        layer6[10][39:32] = buffer_data_0[3167:3160];
        layer6[10][47:40] = buffer_data_0[3175:3168];
        layer6[10][55:48] = buffer_data_0[3183:3176];
        layer0[11][7:0] = buffer_data_6[3143:3136];
        layer0[11][15:8] = buffer_data_6[3151:3144];
        layer0[11][23:16] = buffer_data_6[3159:3152];
        layer0[11][31:24] = buffer_data_6[3167:3160];
        layer0[11][39:32] = buffer_data_6[3175:3168];
        layer0[11][47:40] = buffer_data_6[3183:3176];
        layer0[11][55:48] = buffer_data_6[3191:3184];
        layer1[11][7:0] = buffer_data_5[3143:3136];
        layer1[11][15:8] = buffer_data_5[3151:3144];
        layer1[11][23:16] = buffer_data_5[3159:3152];
        layer1[11][31:24] = buffer_data_5[3167:3160];
        layer1[11][39:32] = buffer_data_5[3175:3168];
        layer1[11][47:40] = buffer_data_5[3183:3176];
        layer1[11][55:48] = buffer_data_5[3191:3184];
        layer2[11][7:0] = buffer_data_4[3143:3136];
        layer2[11][15:8] = buffer_data_4[3151:3144];
        layer2[11][23:16] = buffer_data_4[3159:3152];
        layer2[11][31:24] = buffer_data_4[3167:3160];
        layer2[11][39:32] = buffer_data_4[3175:3168];
        layer2[11][47:40] = buffer_data_4[3183:3176];
        layer2[11][55:48] = buffer_data_4[3191:3184];
        layer3[11][7:0] = buffer_data_3[3143:3136];
        layer3[11][15:8] = buffer_data_3[3151:3144];
        layer3[11][23:16] = buffer_data_3[3159:3152];
        layer3[11][31:24] = buffer_data_3[3167:3160];
        layer3[11][39:32] = buffer_data_3[3175:3168];
        layer3[11][47:40] = buffer_data_3[3183:3176];
        layer3[11][55:48] = buffer_data_3[3191:3184];
        layer4[11][7:0] = buffer_data_2[3143:3136];
        layer4[11][15:8] = buffer_data_2[3151:3144];
        layer4[11][23:16] = buffer_data_2[3159:3152];
        layer4[11][31:24] = buffer_data_2[3167:3160];
        layer4[11][39:32] = buffer_data_2[3175:3168];
        layer4[11][47:40] = buffer_data_2[3183:3176];
        layer4[11][55:48] = buffer_data_2[3191:3184];
        layer5[11][7:0] = buffer_data_1[3143:3136];
        layer5[11][15:8] = buffer_data_1[3151:3144];
        layer5[11][23:16] = buffer_data_1[3159:3152];
        layer5[11][31:24] = buffer_data_1[3167:3160];
        layer5[11][39:32] = buffer_data_1[3175:3168];
        layer5[11][47:40] = buffer_data_1[3183:3176];
        layer5[11][55:48] = buffer_data_1[3191:3184];
        layer6[11][7:0] = buffer_data_0[3143:3136];
        layer6[11][15:8] = buffer_data_0[3151:3144];
        layer6[11][23:16] = buffer_data_0[3159:3152];
        layer6[11][31:24] = buffer_data_0[3167:3160];
        layer6[11][39:32] = buffer_data_0[3175:3168];
        layer6[11][47:40] = buffer_data_0[3183:3176];
        layer6[11][55:48] = buffer_data_0[3191:3184];
        layer0[12][7:0] = buffer_data_6[3151:3144];
        layer0[12][15:8] = buffer_data_6[3159:3152];
        layer0[12][23:16] = buffer_data_6[3167:3160];
        layer0[12][31:24] = buffer_data_6[3175:3168];
        layer0[12][39:32] = buffer_data_6[3183:3176];
        layer0[12][47:40] = buffer_data_6[3191:3184];
        layer0[12][55:48] = buffer_data_6[3199:3192];
        layer1[12][7:0] = buffer_data_5[3151:3144];
        layer1[12][15:8] = buffer_data_5[3159:3152];
        layer1[12][23:16] = buffer_data_5[3167:3160];
        layer1[12][31:24] = buffer_data_5[3175:3168];
        layer1[12][39:32] = buffer_data_5[3183:3176];
        layer1[12][47:40] = buffer_data_5[3191:3184];
        layer1[12][55:48] = buffer_data_5[3199:3192];
        layer2[12][7:0] = buffer_data_4[3151:3144];
        layer2[12][15:8] = buffer_data_4[3159:3152];
        layer2[12][23:16] = buffer_data_4[3167:3160];
        layer2[12][31:24] = buffer_data_4[3175:3168];
        layer2[12][39:32] = buffer_data_4[3183:3176];
        layer2[12][47:40] = buffer_data_4[3191:3184];
        layer2[12][55:48] = buffer_data_4[3199:3192];
        layer3[12][7:0] = buffer_data_3[3151:3144];
        layer3[12][15:8] = buffer_data_3[3159:3152];
        layer3[12][23:16] = buffer_data_3[3167:3160];
        layer3[12][31:24] = buffer_data_3[3175:3168];
        layer3[12][39:32] = buffer_data_3[3183:3176];
        layer3[12][47:40] = buffer_data_3[3191:3184];
        layer3[12][55:48] = buffer_data_3[3199:3192];
        layer4[12][7:0] = buffer_data_2[3151:3144];
        layer4[12][15:8] = buffer_data_2[3159:3152];
        layer4[12][23:16] = buffer_data_2[3167:3160];
        layer4[12][31:24] = buffer_data_2[3175:3168];
        layer4[12][39:32] = buffer_data_2[3183:3176];
        layer4[12][47:40] = buffer_data_2[3191:3184];
        layer4[12][55:48] = buffer_data_2[3199:3192];
        layer5[12][7:0] = buffer_data_1[3151:3144];
        layer5[12][15:8] = buffer_data_1[3159:3152];
        layer5[12][23:16] = buffer_data_1[3167:3160];
        layer5[12][31:24] = buffer_data_1[3175:3168];
        layer5[12][39:32] = buffer_data_1[3183:3176];
        layer5[12][47:40] = buffer_data_1[3191:3184];
        layer5[12][55:48] = buffer_data_1[3199:3192];
        layer6[12][7:0] = buffer_data_0[3151:3144];
        layer6[12][15:8] = buffer_data_0[3159:3152];
        layer6[12][23:16] = buffer_data_0[3167:3160];
        layer6[12][31:24] = buffer_data_0[3175:3168];
        layer6[12][39:32] = buffer_data_0[3183:3176];
        layer6[12][47:40] = buffer_data_0[3191:3184];
        layer6[12][55:48] = buffer_data_0[3199:3192];
        layer0[13][7:0] = buffer_data_6[3159:3152];
        layer0[13][15:8] = buffer_data_6[3167:3160];
        layer0[13][23:16] = buffer_data_6[3175:3168];
        layer0[13][31:24] = buffer_data_6[3183:3176];
        layer0[13][39:32] = buffer_data_6[3191:3184];
        layer0[13][47:40] = buffer_data_6[3199:3192];
        layer0[13][55:48] = buffer_data_6[3207:3200];
        layer1[13][7:0] = buffer_data_5[3159:3152];
        layer1[13][15:8] = buffer_data_5[3167:3160];
        layer1[13][23:16] = buffer_data_5[3175:3168];
        layer1[13][31:24] = buffer_data_5[3183:3176];
        layer1[13][39:32] = buffer_data_5[3191:3184];
        layer1[13][47:40] = buffer_data_5[3199:3192];
        layer1[13][55:48] = buffer_data_5[3207:3200];
        layer2[13][7:0] = buffer_data_4[3159:3152];
        layer2[13][15:8] = buffer_data_4[3167:3160];
        layer2[13][23:16] = buffer_data_4[3175:3168];
        layer2[13][31:24] = buffer_data_4[3183:3176];
        layer2[13][39:32] = buffer_data_4[3191:3184];
        layer2[13][47:40] = buffer_data_4[3199:3192];
        layer2[13][55:48] = buffer_data_4[3207:3200];
        layer3[13][7:0] = buffer_data_3[3159:3152];
        layer3[13][15:8] = buffer_data_3[3167:3160];
        layer3[13][23:16] = buffer_data_3[3175:3168];
        layer3[13][31:24] = buffer_data_3[3183:3176];
        layer3[13][39:32] = buffer_data_3[3191:3184];
        layer3[13][47:40] = buffer_data_3[3199:3192];
        layer3[13][55:48] = buffer_data_3[3207:3200];
        layer4[13][7:0] = buffer_data_2[3159:3152];
        layer4[13][15:8] = buffer_data_2[3167:3160];
        layer4[13][23:16] = buffer_data_2[3175:3168];
        layer4[13][31:24] = buffer_data_2[3183:3176];
        layer4[13][39:32] = buffer_data_2[3191:3184];
        layer4[13][47:40] = buffer_data_2[3199:3192];
        layer4[13][55:48] = buffer_data_2[3207:3200];
        layer5[13][7:0] = buffer_data_1[3159:3152];
        layer5[13][15:8] = buffer_data_1[3167:3160];
        layer5[13][23:16] = buffer_data_1[3175:3168];
        layer5[13][31:24] = buffer_data_1[3183:3176];
        layer5[13][39:32] = buffer_data_1[3191:3184];
        layer5[13][47:40] = buffer_data_1[3199:3192];
        layer5[13][55:48] = buffer_data_1[3207:3200];
        layer6[13][7:0] = buffer_data_0[3159:3152];
        layer6[13][15:8] = buffer_data_0[3167:3160];
        layer6[13][23:16] = buffer_data_0[3175:3168];
        layer6[13][31:24] = buffer_data_0[3183:3176];
        layer6[13][39:32] = buffer_data_0[3191:3184];
        layer6[13][47:40] = buffer_data_0[3199:3192];
        layer6[13][55:48] = buffer_data_0[3207:3200];
        layer0[14][7:0] = buffer_data_6[3167:3160];
        layer0[14][15:8] = buffer_data_6[3175:3168];
        layer0[14][23:16] = buffer_data_6[3183:3176];
        layer0[14][31:24] = buffer_data_6[3191:3184];
        layer0[14][39:32] = buffer_data_6[3199:3192];
        layer0[14][47:40] = buffer_data_6[3207:3200];
        layer0[14][55:48] = buffer_data_6[3215:3208];
        layer1[14][7:0] = buffer_data_5[3167:3160];
        layer1[14][15:8] = buffer_data_5[3175:3168];
        layer1[14][23:16] = buffer_data_5[3183:3176];
        layer1[14][31:24] = buffer_data_5[3191:3184];
        layer1[14][39:32] = buffer_data_5[3199:3192];
        layer1[14][47:40] = buffer_data_5[3207:3200];
        layer1[14][55:48] = buffer_data_5[3215:3208];
        layer2[14][7:0] = buffer_data_4[3167:3160];
        layer2[14][15:8] = buffer_data_4[3175:3168];
        layer2[14][23:16] = buffer_data_4[3183:3176];
        layer2[14][31:24] = buffer_data_4[3191:3184];
        layer2[14][39:32] = buffer_data_4[3199:3192];
        layer2[14][47:40] = buffer_data_4[3207:3200];
        layer2[14][55:48] = buffer_data_4[3215:3208];
        layer3[14][7:0] = buffer_data_3[3167:3160];
        layer3[14][15:8] = buffer_data_3[3175:3168];
        layer3[14][23:16] = buffer_data_3[3183:3176];
        layer3[14][31:24] = buffer_data_3[3191:3184];
        layer3[14][39:32] = buffer_data_3[3199:3192];
        layer3[14][47:40] = buffer_data_3[3207:3200];
        layer3[14][55:48] = buffer_data_3[3215:3208];
        layer4[14][7:0] = buffer_data_2[3167:3160];
        layer4[14][15:8] = buffer_data_2[3175:3168];
        layer4[14][23:16] = buffer_data_2[3183:3176];
        layer4[14][31:24] = buffer_data_2[3191:3184];
        layer4[14][39:32] = buffer_data_2[3199:3192];
        layer4[14][47:40] = buffer_data_2[3207:3200];
        layer4[14][55:48] = buffer_data_2[3215:3208];
        layer5[14][7:0] = buffer_data_1[3167:3160];
        layer5[14][15:8] = buffer_data_1[3175:3168];
        layer5[14][23:16] = buffer_data_1[3183:3176];
        layer5[14][31:24] = buffer_data_1[3191:3184];
        layer5[14][39:32] = buffer_data_1[3199:3192];
        layer5[14][47:40] = buffer_data_1[3207:3200];
        layer5[14][55:48] = buffer_data_1[3215:3208];
        layer6[14][7:0] = buffer_data_0[3167:3160];
        layer6[14][15:8] = buffer_data_0[3175:3168];
        layer6[14][23:16] = buffer_data_0[3183:3176];
        layer6[14][31:24] = buffer_data_0[3191:3184];
        layer6[14][39:32] = buffer_data_0[3199:3192];
        layer6[14][47:40] = buffer_data_0[3207:3200];
        layer6[14][55:48] = buffer_data_0[3215:3208];
        layer0[15][7:0] = buffer_data_6[3175:3168];
        layer0[15][15:8] = buffer_data_6[3183:3176];
        layer0[15][23:16] = buffer_data_6[3191:3184];
        layer0[15][31:24] = buffer_data_6[3199:3192];
        layer0[15][39:32] = buffer_data_6[3207:3200];
        layer0[15][47:40] = buffer_data_6[3215:3208];
        layer0[15][55:48] = buffer_data_6[3223:3216];
        layer1[15][7:0] = buffer_data_5[3175:3168];
        layer1[15][15:8] = buffer_data_5[3183:3176];
        layer1[15][23:16] = buffer_data_5[3191:3184];
        layer1[15][31:24] = buffer_data_5[3199:3192];
        layer1[15][39:32] = buffer_data_5[3207:3200];
        layer1[15][47:40] = buffer_data_5[3215:3208];
        layer1[15][55:48] = buffer_data_5[3223:3216];
        layer2[15][7:0] = buffer_data_4[3175:3168];
        layer2[15][15:8] = buffer_data_4[3183:3176];
        layer2[15][23:16] = buffer_data_4[3191:3184];
        layer2[15][31:24] = buffer_data_4[3199:3192];
        layer2[15][39:32] = buffer_data_4[3207:3200];
        layer2[15][47:40] = buffer_data_4[3215:3208];
        layer2[15][55:48] = buffer_data_4[3223:3216];
        layer3[15][7:0] = buffer_data_3[3175:3168];
        layer3[15][15:8] = buffer_data_3[3183:3176];
        layer3[15][23:16] = buffer_data_3[3191:3184];
        layer3[15][31:24] = buffer_data_3[3199:3192];
        layer3[15][39:32] = buffer_data_3[3207:3200];
        layer3[15][47:40] = buffer_data_3[3215:3208];
        layer3[15][55:48] = buffer_data_3[3223:3216];
        layer4[15][7:0] = buffer_data_2[3175:3168];
        layer4[15][15:8] = buffer_data_2[3183:3176];
        layer4[15][23:16] = buffer_data_2[3191:3184];
        layer4[15][31:24] = buffer_data_2[3199:3192];
        layer4[15][39:32] = buffer_data_2[3207:3200];
        layer4[15][47:40] = buffer_data_2[3215:3208];
        layer4[15][55:48] = buffer_data_2[3223:3216];
        layer5[15][7:0] = buffer_data_1[3175:3168];
        layer5[15][15:8] = buffer_data_1[3183:3176];
        layer5[15][23:16] = buffer_data_1[3191:3184];
        layer5[15][31:24] = buffer_data_1[3199:3192];
        layer5[15][39:32] = buffer_data_1[3207:3200];
        layer5[15][47:40] = buffer_data_1[3215:3208];
        layer5[15][55:48] = buffer_data_1[3223:3216];
        layer6[15][7:0] = buffer_data_0[3175:3168];
        layer6[15][15:8] = buffer_data_0[3183:3176];
        layer6[15][23:16] = buffer_data_0[3191:3184];
        layer6[15][31:24] = buffer_data_0[3199:3192];
        layer6[15][39:32] = buffer_data_0[3207:3200];
        layer6[15][47:40] = buffer_data_0[3215:3208];
        layer6[15][55:48] = buffer_data_0[3223:3216];
        layer0[16][7:0] = buffer_data_6[3183:3176];
        layer0[16][15:8] = buffer_data_6[3191:3184];
        layer0[16][23:16] = buffer_data_6[3199:3192];
        layer0[16][31:24] = buffer_data_6[3207:3200];
        layer0[16][39:32] = buffer_data_6[3215:3208];
        layer0[16][47:40] = buffer_data_6[3223:3216];
        layer0[16][55:48] = buffer_data_6[3231:3224];
        layer1[16][7:0] = buffer_data_5[3183:3176];
        layer1[16][15:8] = buffer_data_5[3191:3184];
        layer1[16][23:16] = buffer_data_5[3199:3192];
        layer1[16][31:24] = buffer_data_5[3207:3200];
        layer1[16][39:32] = buffer_data_5[3215:3208];
        layer1[16][47:40] = buffer_data_5[3223:3216];
        layer1[16][55:48] = buffer_data_5[3231:3224];
        layer2[16][7:0] = buffer_data_4[3183:3176];
        layer2[16][15:8] = buffer_data_4[3191:3184];
        layer2[16][23:16] = buffer_data_4[3199:3192];
        layer2[16][31:24] = buffer_data_4[3207:3200];
        layer2[16][39:32] = buffer_data_4[3215:3208];
        layer2[16][47:40] = buffer_data_4[3223:3216];
        layer2[16][55:48] = buffer_data_4[3231:3224];
        layer3[16][7:0] = buffer_data_3[3183:3176];
        layer3[16][15:8] = buffer_data_3[3191:3184];
        layer3[16][23:16] = buffer_data_3[3199:3192];
        layer3[16][31:24] = buffer_data_3[3207:3200];
        layer3[16][39:32] = buffer_data_3[3215:3208];
        layer3[16][47:40] = buffer_data_3[3223:3216];
        layer3[16][55:48] = buffer_data_3[3231:3224];
        layer4[16][7:0] = buffer_data_2[3183:3176];
        layer4[16][15:8] = buffer_data_2[3191:3184];
        layer4[16][23:16] = buffer_data_2[3199:3192];
        layer4[16][31:24] = buffer_data_2[3207:3200];
        layer4[16][39:32] = buffer_data_2[3215:3208];
        layer4[16][47:40] = buffer_data_2[3223:3216];
        layer4[16][55:48] = buffer_data_2[3231:3224];
        layer5[16][7:0] = buffer_data_1[3183:3176];
        layer5[16][15:8] = buffer_data_1[3191:3184];
        layer5[16][23:16] = buffer_data_1[3199:3192];
        layer5[16][31:24] = buffer_data_1[3207:3200];
        layer5[16][39:32] = buffer_data_1[3215:3208];
        layer5[16][47:40] = buffer_data_1[3223:3216];
        layer5[16][55:48] = buffer_data_1[3231:3224];
        layer6[16][7:0] = buffer_data_0[3183:3176];
        layer6[16][15:8] = buffer_data_0[3191:3184];
        layer6[16][23:16] = buffer_data_0[3199:3192];
        layer6[16][31:24] = buffer_data_0[3207:3200];
        layer6[16][39:32] = buffer_data_0[3215:3208];
        layer6[16][47:40] = buffer_data_0[3223:3216];
        layer6[16][55:48] = buffer_data_0[3231:3224];
        layer0[17][7:0] = buffer_data_6[3191:3184];
        layer0[17][15:8] = buffer_data_6[3199:3192];
        layer0[17][23:16] = buffer_data_6[3207:3200];
        layer0[17][31:24] = buffer_data_6[3215:3208];
        layer0[17][39:32] = buffer_data_6[3223:3216];
        layer0[17][47:40] = buffer_data_6[3231:3224];
        layer0[17][55:48] = buffer_data_6[3239:3232];
        layer1[17][7:0] = buffer_data_5[3191:3184];
        layer1[17][15:8] = buffer_data_5[3199:3192];
        layer1[17][23:16] = buffer_data_5[3207:3200];
        layer1[17][31:24] = buffer_data_5[3215:3208];
        layer1[17][39:32] = buffer_data_5[3223:3216];
        layer1[17][47:40] = buffer_data_5[3231:3224];
        layer1[17][55:48] = buffer_data_5[3239:3232];
        layer2[17][7:0] = buffer_data_4[3191:3184];
        layer2[17][15:8] = buffer_data_4[3199:3192];
        layer2[17][23:16] = buffer_data_4[3207:3200];
        layer2[17][31:24] = buffer_data_4[3215:3208];
        layer2[17][39:32] = buffer_data_4[3223:3216];
        layer2[17][47:40] = buffer_data_4[3231:3224];
        layer2[17][55:48] = buffer_data_4[3239:3232];
        layer3[17][7:0] = buffer_data_3[3191:3184];
        layer3[17][15:8] = buffer_data_3[3199:3192];
        layer3[17][23:16] = buffer_data_3[3207:3200];
        layer3[17][31:24] = buffer_data_3[3215:3208];
        layer3[17][39:32] = buffer_data_3[3223:3216];
        layer3[17][47:40] = buffer_data_3[3231:3224];
        layer3[17][55:48] = buffer_data_3[3239:3232];
        layer4[17][7:0] = buffer_data_2[3191:3184];
        layer4[17][15:8] = buffer_data_2[3199:3192];
        layer4[17][23:16] = buffer_data_2[3207:3200];
        layer4[17][31:24] = buffer_data_2[3215:3208];
        layer4[17][39:32] = buffer_data_2[3223:3216];
        layer4[17][47:40] = buffer_data_2[3231:3224];
        layer4[17][55:48] = buffer_data_2[3239:3232];
        layer5[17][7:0] = buffer_data_1[3191:3184];
        layer5[17][15:8] = buffer_data_1[3199:3192];
        layer5[17][23:16] = buffer_data_1[3207:3200];
        layer5[17][31:24] = buffer_data_1[3215:3208];
        layer5[17][39:32] = buffer_data_1[3223:3216];
        layer5[17][47:40] = buffer_data_1[3231:3224];
        layer5[17][55:48] = buffer_data_1[3239:3232];
        layer6[17][7:0] = buffer_data_0[3191:3184];
        layer6[17][15:8] = buffer_data_0[3199:3192];
        layer6[17][23:16] = buffer_data_0[3207:3200];
        layer6[17][31:24] = buffer_data_0[3215:3208];
        layer6[17][39:32] = buffer_data_0[3223:3216];
        layer6[17][47:40] = buffer_data_0[3231:3224];
        layer6[17][55:48] = buffer_data_0[3239:3232];
        layer0[18][7:0] = buffer_data_6[3199:3192];
        layer0[18][15:8] = buffer_data_6[3207:3200];
        layer0[18][23:16] = buffer_data_6[3215:3208];
        layer0[18][31:24] = buffer_data_6[3223:3216];
        layer0[18][39:32] = buffer_data_6[3231:3224];
        layer0[18][47:40] = buffer_data_6[3239:3232];
        layer0[18][55:48] = buffer_data_6[3247:3240];
        layer1[18][7:0] = buffer_data_5[3199:3192];
        layer1[18][15:8] = buffer_data_5[3207:3200];
        layer1[18][23:16] = buffer_data_5[3215:3208];
        layer1[18][31:24] = buffer_data_5[3223:3216];
        layer1[18][39:32] = buffer_data_5[3231:3224];
        layer1[18][47:40] = buffer_data_5[3239:3232];
        layer1[18][55:48] = buffer_data_5[3247:3240];
        layer2[18][7:0] = buffer_data_4[3199:3192];
        layer2[18][15:8] = buffer_data_4[3207:3200];
        layer2[18][23:16] = buffer_data_4[3215:3208];
        layer2[18][31:24] = buffer_data_4[3223:3216];
        layer2[18][39:32] = buffer_data_4[3231:3224];
        layer2[18][47:40] = buffer_data_4[3239:3232];
        layer2[18][55:48] = buffer_data_4[3247:3240];
        layer3[18][7:0] = buffer_data_3[3199:3192];
        layer3[18][15:8] = buffer_data_3[3207:3200];
        layer3[18][23:16] = buffer_data_3[3215:3208];
        layer3[18][31:24] = buffer_data_3[3223:3216];
        layer3[18][39:32] = buffer_data_3[3231:3224];
        layer3[18][47:40] = buffer_data_3[3239:3232];
        layer3[18][55:48] = buffer_data_3[3247:3240];
        layer4[18][7:0] = buffer_data_2[3199:3192];
        layer4[18][15:8] = buffer_data_2[3207:3200];
        layer4[18][23:16] = buffer_data_2[3215:3208];
        layer4[18][31:24] = buffer_data_2[3223:3216];
        layer4[18][39:32] = buffer_data_2[3231:3224];
        layer4[18][47:40] = buffer_data_2[3239:3232];
        layer4[18][55:48] = buffer_data_2[3247:3240];
        layer5[18][7:0] = buffer_data_1[3199:3192];
        layer5[18][15:8] = buffer_data_1[3207:3200];
        layer5[18][23:16] = buffer_data_1[3215:3208];
        layer5[18][31:24] = buffer_data_1[3223:3216];
        layer5[18][39:32] = buffer_data_1[3231:3224];
        layer5[18][47:40] = buffer_data_1[3239:3232];
        layer5[18][55:48] = buffer_data_1[3247:3240];
        layer6[18][7:0] = buffer_data_0[3199:3192];
        layer6[18][15:8] = buffer_data_0[3207:3200];
        layer6[18][23:16] = buffer_data_0[3215:3208];
        layer6[18][31:24] = buffer_data_0[3223:3216];
        layer6[18][39:32] = buffer_data_0[3231:3224];
        layer6[18][47:40] = buffer_data_0[3239:3232];
        layer6[18][55:48] = buffer_data_0[3247:3240];
        layer0[19][7:0] = buffer_data_6[3207:3200];
        layer0[19][15:8] = buffer_data_6[3215:3208];
        layer0[19][23:16] = buffer_data_6[3223:3216];
        layer0[19][31:24] = buffer_data_6[3231:3224];
        layer0[19][39:32] = buffer_data_6[3239:3232];
        layer0[19][47:40] = buffer_data_6[3247:3240];
        layer0[19][55:48] = buffer_data_6[3255:3248];
        layer1[19][7:0] = buffer_data_5[3207:3200];
        layer1[19][15:8] = buffer_data_5[3215:3208];
        layer1[19][23:16] = buffer_data_5[3223:3216];
        layer1[19][31:24] = buffer_data_5[3231:3224];
        layer1[19][39:32] = buffer_data_5[3239:3232];
        layer1[19][47:40] = buffer_data_5[3247:3240];
        layer1[19][55:48] = buffer_data_5[3255:3248];
        layer2[19][7:0] = buffer_data_4[3207:3200];
        layer2[19][15:8] = buffer_data_4[3215:3208];
        layer2[19][23:16] = buffer_data_4[3223:3216];
        layer2[19][31:24] = buffer_data_4[3231:3224];
        layer2[19][39:32] = buffer_data_4[3239:3232];
        layer2[19][47:40] = buffer_data_4[3247:3240];
        layer2[19][55:48] = buffer_data_4[3255:3248];
        layer3[19][7:0] = buffer_data_3[3207:3200];
        layer3[19][15:8] = buffer_data_3[3215:3208];
        layer3[19][23:16] = buffer_data_3[3223:3216];
        layer3[19][31:24] = buffer_data_3[3231:3224];
        layer3[19][39:32] = buffer_data_3[3239:3232];
        layer3[19][47:40] = buffer_data_3[3247:3240];
        layer3[19][55:48] = buffer_data_3[3255:3248];
        layer4[19][7:0] = buffer_data_2[3207:3200];
        layer4[19][15:8] = buffer_data_2[3215:3208];
        layer4[19][23:16] = buffer_data_2[3223:3216];
        layer4[19][31:24] = buffer_data_2[3231:3224];
        layer4[19][39:32] = buffer_data_2[3239:3232];
        layer4[19][47:40] = buffer_data_2[3247:3240];
        layer4[19][55:48] = buffer_data_2[3255:3248];
        layer5[19][7:0] = buffer_data_1[3207:3200];
        layer5[19][15:8] = buffer_data_1[3215:3208];
        layer5[19][23:16] = buffer_data_1[3223:3216];
        layer5[19][31:24] = buffer_data_1[3231:3224];
        layer5[19][39:32] = buffer_data_1[3239:3232];
        layer5[19][47:40] = buffer_data_1[3247:3240];
        layer5[19][55:48] = buffer_data_1[3255:3248];
        layer6[19][7:0] = buffer_data_0[3207:3200];
        layer6[19][15:8] = buffer_data_0[3215:3208];
        layer6[19][23:16] = buffer_data_0[3223:3216];
        layer6[19][31:24] = buffer_data_0[3231:3224];
        layer6[19][39:32] = buffer_data_0[3239:3232];
        layer6[19][47:40] = buffer_data_0[3247:3240];
        layer6[19][55:48] = buffer_data_0[3255:3248];
        layer0[20][7:0] = buffer_data_6[3215:3208];
        layer0[20][15:8] = buffer_data_6[3223:3216];
        layer0[20][23:16] = buffer_data_6[3231:3224];
        layer0[20][31:24] = buffer_data_6[3239:3232];
        layer0[20][39:32] = buffer_data_6[3247:3240];
        layer0[20][47:40] = buffer_data_6[3255:3248];
        layer0[20][55:48] = buffer_data_6[3263:3256];
        layer1[20][7:0] = buffer_data_5[3215:3208];
        layer1[20][15:8] = buffer_data_5[3223:3216];
        layer1[20][23:16] = buffer_data_5[3231:3224];
        layer1[20][31:24] = buffer_data_5[3239:3232];
        layer1[20][39:32] = buffer_data_5[3247:3240];
        layer1[20][47:40] = buffer_data_5[3255:3248];
        layer1[20][55:48] = buffer_data_5[3263:3256];
        layer2[20][7:0] = buffer_data_4[3215:3208];
        layer2[20][15:8] = buffer_data_4[3223:3216];
        layer2[20][23:16] = buffer_data_4[3231:3224];
        layer2[20][31:24] = buffer_data_4[3239:3232];
        layer2[20][39:32] = buffer_data_4[3247:3240];
        layer2[20][47:40] = buffer_data_4[3255:3248];
        layer2[20][55:48] = buffer_data_4[3263:3256];
        layer3[20][7:0] = buffer_data_3[3215:3208];
        layer3[20][15:8] = buffer_data_3[3223:3216];
        layer3[20][23:16] = buffer_data_3[3231:3224];
        layer3[20][31:24] = buffer_data_3[3239:3232];
        layer3[20][39:32] = buffer_data_3[3247:3240];
        layer3[20][47:40] = buffer_data_3[3255:3248];
        layer3[20][55:48] = buffer_data_3[3263:3256];
        layer4[20][7:0] = buffer_data_2[3215:3208];
        layer4[20][15:8] = buffer_data_2[3223:3216];
        layer4[20][23:16] = buffer_data_2[3231:3224];
        layer4[20][31:24] = buffer_data_2[3239:3232];
        layer4[20][39:32] = buffer_data_2[3247:3240];
        layer4[20][47:40] = buffer_data_2[3255:3248];
        layer4[20][55:48] = buffer_data_2[3263:3256];
        layer5[20][7:0] = buffer_data_1[3215:3208];
        layer5[20][15:8] = buffer_data_1[3223:3216];
        layer5[20][23:16] = buffer_data_1[3231:3224];
        layer5[20][31:24] = buffer_data_1[3239:3232];
        layer5[20][39:32] = buffer_data_1[3247:3240];
        layer5[20][47:40] = buffer_data_1[3255:3248];
        layer5[20][55:48] = buffer_data_1[3263:3256];
        layer6[20][7:0] = buffer_data_0[3215:3208];
        layer6[20][15:8] = buffer_data_0[3223:3216];
        layer6[20][23:16] = buffer_data_0[3231:3224];
        layer6[20][31:24] = buffer_data_0[3239:3232];
        layer6[20][39:32] = buffer_data_0[3247:3240];
        layer6[20][47:40] = buffer_data_0[3255:3248];
        layer6[20][55:48] = buffer_data_0[3263:3256];
        layer0[21][7:0] = buffer_data_6[3223:3216];
        layer0[21][15:8] = buffer_data_6[3231:3224];
        layer0[21][23:16] = buffer_data_6[3239:3232];
        layer0[21][31:24] = buffer_data_6[3247:3240];
        layer0[21][39:32] = buffer_data_6[3255:3248];
        layer0[21][47:40] = buffer_data_6[3263:3256];
        layer0[21][55:48] = buffer_data_6[3271:3264];
        layer1[21][7:0] = buffer_data_5[3223:3216];
        layer1[21][15:8] = buffer_data_5[3231:3224];
        layer1[21][23:16] = buffer_data_5[3239:3232];
        layer1[21][31:24] = buffer_data_5[3247:3240];
        layer1[21][39:32] = buffer_data_5[3255:3248];
        layer1[21][47:40] = buffer_data_5[3263:3256];
        layer1[21][55:48] = buffer_data_5[3271:3264];
        layer2[21][7:0] = buffer_data_4[3223:3216];
        layer2[21][15:8] = buffer_data_4[3231:3224];
        layer2[21][23:16] = buffer_data_4[3239:3232];
        layer2[21][31:24] = buffer_data_4[3247:3240];
        layer2[21][39:32] = buffer_data_4[3255:3248];
        layer2[21][47:40] = buffer_data_4[3263:3256];
        layer2[21][55:48] = buffer_data_4[3271:3264];
        layer3[21][7:0] = buffer_data_3[3223:3216];
        layer3[21][15:8] = buffer_data_3[3231:3224];
        layer3[21][23:16] = buffer_data_3[3239:3232];
        layer3[21][31:24] = buffer_data_3[3247:3240];
        layer3[21][39:32] = buffer_data_3[3255:3248];
        layer3[21][47:40] = buffer_data_3[3263:3256];
        layer3[21][55:48] = buffer_data_3[3271:3264];
        layer4[21][7:0] = buffer_data_2[3223:3216];
        layer4[21][15:8] = buffer_data_2[3231:3224];
        layer4[21][23:16] = buffer_data_2[3239:3232];
        layer4[21][31:24] = buffer_data_2[3247:3240];
        layer4[21][39:32] = buffer_data_2[3255:3248];
        layer4[21][47:40] = buffer_data_2[3263:3256];
        layer4[21][55:48] = buffer_data_2[3271:3264];
        layer5[21][7:0] = buffer_data_1[3223:3216];
        layer5[21][15:8] = buffer_data_1[3231:3224];
        layer5[21][23:16] = buffer_data_1[3239:3232];
        layer5[21][31:24] = buffer_data_1[3247:3240];
        layer5[21][39:32] = buffer_data_1[3255:3248];
        layer5[21][47:40] = buffer_data_1[3263:3256];
        layer5[21][55:48] = buffer_data_1[3271:3264];
        layer6[21][7:0] = buffer_data_0[3223:3216];
        layer6[21][15:8] = buffer_data_0[3231:3224];
        layer6[21][23:16] = buffer_data_0[3239:3232];
        layer6[21][31:24] = buffer_data_0[3247:3240];
        layer6[21][39:32] = buffer_data_0[3255:3248];
        layer6[21][47:40] = buffer_data_0[3263:3256];
        layer6[21][55:48] = buffer_data_0[3271:3264];
        layer0[22][7:0] = buffer_data_6[3231:3224];
        layer0[22][15:8] = buffer_data_6[3239:3232];
        layer0[22][23:16] = buffer_data_6[3247:3240];
        layer0[22][31:24] = buffer_data_6[3255:3248];
        layer0[22][39:32] = buffer_data_6[3263:3256];
        layer0[22][47:40] = buffer_data_6[3271:3264];
        layer0[22][55:48] = buffer_data_6[3279:3272];
        layer1[22][7:0] = buffer_data_5[3231:3224];
        layer1[22][15:8] = buffer_data_5[3239:3232];
        layer1[22][23:16] = buffer_data_5[3247:3240];
        layer1[22][31:24] = buffer_data_5[3255:3248];
        layer1[22][39:32] = buffer_data_5[3263:3256];
        layer1[22][47:40] = buffer_data_5[3271:3264];
        layer1[22][55:48] = buffer_data_5[3279:3272];
        layer2[22][7:0] = buffer_data_4[3231:3224];
        layer2[22][15:8] = buffer_data_4[3239:3232];
        layer2[22][23:16] = buffer_data_4[3247:3240];
        layer2[22][31:24] = buffer_data_4[3255:3248];
        layer2[22][39:32] = buffer_data_4[3263:3256];
        layer2[22][47:40] = buffer_data_4[3271:3264];
        layer2[22][55:48] = buffer_data_4[3279:3272];
        layer3[22][7:0] = buffer_data_3[3231:3224];
        layer3[22][15:8] = buffer_data_3[3239:3232];
        layer3[22][23:16] = buffer_data_3[3247:3240];
        layer3[22][31:24] = buffer_data_3[3255:3248];
        layer3[22][39:32] = buffer_data_3[3263:3256];
        layer3[22][47:40] = buffer_data_3[3271:3264];
        layer3[22][55:48] = buffer_data_3[3279:3272];
        layer4[22][7:0] = buffer_data_2[3231:3224];
        layer4[22][15:8] = buffer_data_2[3239:3232];
        layer4[22][23:16] = buffer_data_2[3247:3240];
        layer4[22][31:24] = buffer_data_2[3255:3248];
        layer4[22][39:32] = buffer_data_2[3263:3256];
        layer4[22][47:40] = buffer_data_2[3271:3264];
        layer4[22][55:48] = buffer_data_2[3279:3272];
        layer5[22][7:0] = buffer_data_1[3231:3224];
        layer5[22][15:8] = buffer_data_1[3239:3232];
        layer5[22][23:16] = buffer_data_1[3247:3240];
        layer5[22][31:24] = buffer_data_1[3255:3248];
        layer5[22][39:32] = buffer_data_1[3263:3256];
        layer5[22][47:40] = buffer_data_1[3271:3264];
        layer5[22][55:48] = buffer_data_1[3279:3272];
        layer6[22][7:0] = buffer_data_0[3231:3224];
        layer6[22][15:8] = buffer_data_0[3239:3232];
        layer6[22][23:16] = buffer_data_0[3247:3240];
        layer6[22][31:24] = buffer_data_0[3255:3248];
        layer6[22][39:32] = buffer_data_0[3263:3256];
        layer6[22][47:40] = buffer_data_0[3271:3264];
        layer6[22][55:48] = buffer_data_0[3279:3272];
        layer0[23][7:0] = buffer_data_6[3239:3232];
        layer0[23][15:8] = buffer_data_6[3247:3240];
        layer0[23][23:16] = buffer_data_6[3255:3248];
        layer0[23][31:24] = buffer_data_6[3263:3256];
        layer0[23][39:32] = buffer_data_6[3271:3264];
        layer0[23][47:40] = buffer_data_6[3279:3272];
        layer0[23][55:48] = buffer_data_6[3287:3280];
        layer1[23][7:0] = buffer_data_5[3239:3232];
        layer1[23][15:8] = buffer_data_5[3247:3240];
        layer1[23][23:16] = buffer_data_5[3255:3248];
        layer1[23][31:24] = buffer_data_5[3263:3256];
        layer1[23][39:32] = buffer_data_5[3271:3264];
        layer1[23][47:40] = buffer_data_5[3279:3272];
        layer1[23][55:48] = buffer_data_5[3287:3280];
        layer2[23][7:0] = buffer_data_4[3239:3232];
        layer2[23][15:8] = buffer_data_4[3247:3240];
        layer2[23][23:16] = buffer_data_4[3255:3248];
        layer2[23][31:24] = buffer_data_4[3263:3256];
        layer2[23][39:32] = buffer_data_4[3271:3264];
        layer2[23][47:40] = buffer_data_4[3279:3272];
        layer2[23][55:48] = buffer_data_4[3287:3280];
        layer3[23][7:0] = buffer_data_3[3239:3232];
        layer3[23][15:8] = buffer_data_3[3247:3240];
        layer3[23][23:16] = buffer_data_3[3255:3248];
        layer3[23][31:24] = buffer_data_3[3263:3256];
        layer3[23][39:32] = buffer_data_3[3271:3264];
        layer3[23][47:40] = buffer_data_3[3279:3272];
        layer3[23][55:48] = buffer_data_3[3287:3280];
        layer4[23][7:0] = buffer_data_2[3239:3232];
        layer4[23][15:8] = buffer_data_2[3247:3240];
        layer4[23][23:16] = buffer_data_2[3255:3248];
        layer4[23][31:24] = buffer_data_2[3263:3256];
        layer4[23][39:32] = buffer_data_2[3271:3264];
        layer4[23][47:40] = buffer_data_2[3279:3272];
        layer4[23][55:48] = buffer_data_2[3287:3280];
        layer5[23][7:0] = buffer_data_1[3239:3232];
        layer5[23][15:8] = buffer_data_1[3247:3240];
        layer5[23][23:16] = buffer_data_1[3255:3248];
        layer5[23][31:24] = buffer_data_1[3263:3256];
        layer5[23][39:32] = buffer_data_1[3271:3264];
        layer5[23][47:40] = buffer_data_1[3279:3272];
        layer5[23][55:48] = buffer_data_1[3287:3280];
        layer6[23][7:0] = buffer_data_0[3239:3232];
        layer6[23][15:8] = buffer_data_0[3247:3240];
        layer6[23][23:16] = buffer_data_0[3255:3248];
        layer6[23][31:24] = buffer_data_0[3263:3256];
        layer6[23][39:32] = buffer_data_0[3271:3264];
        layer6[23][47:40] = buffer_data_0[3279:3272];
        layer6[23][55:48] = buffer_data_0[3287:3280];
        layer0[24][7:0] = buffer_data_6[3247:3240];
        layer0[24][15:8] = buffer_data_6[3255:3248];
        layer0[24][23:16] = buffer_data_6[3263:3256];
        layer0[24][31:24] = buffer_data_6[3271:3264];
        layer0[24][39:32] = buffer_data_6[3279:3272];
        layer0[24][47:40] = buffer_data_6[3287:3280];
        layer0[24][55:48] = buffer_data_6[3295:3288];
        layer1[24][7:0] = buffer_data_5[3247:3240];
        layer1[24][15:8] = buffer_data_5[3255:3248];
        layer1[24][23:16] = buffer_data_5[3263:3256];
        layer1[24][31:24] = buffer_data_5[3271:3264];
        layer1[24][39:32] = buffer_data_5[3279:3272];
        layer1[24][47:40] = buffer_data_5[3287:3280];
        layer1[24][55:48] = buffer_data_5[3295:3288];
        layer2[24][7:0] = buffer_data_4[3247:3240];
        layer2[24][15:8] = buffer_data_4[3255:3248];
        layer2[24][23:16] = buffer_data_4[3263:3256];
        layer2[24][31:24] = buffer_data_4[3271:3264];
        layer2[24][39:32] = buffer_data_4[3279:3272];
        layer2[24][47:40] = buffer_data_4[3287:3280];
        layer2[24][55:48] = buffer_data_4[3295:3288];
        layer3[24][7:0] = buffer_data_3[3247:3240];
        layer3[24][15:8] = buffer_data_3[3255:3248];
        layer3[24][23:16] = buffer_data_3[3263:3256];
        layer3[24][31:24] = buffer_data_3[3271:3264];
        layer3[24][39:32] = buffer_data_3[3279:3272];
        layer3[24][47:40] = buffer_data_3[3287:3280];
        layer3[24][55:48] = buffer_data_3[3295:3288];
        layer4[24][7:0] = buffer_data_2[3247:3240];
        layer4[24][15:8] = buffer_data_2[3255:3248];
        layer4[24][23:16] = buffer_data_2[3263:3256];
        layer4[24][31:24] = buffer_data_2[3271:3264];
        layer4[24][39:32] = buffer_data_2[3279:3272];
        layer4[24][47:40] = buffer_data_2[3287:3280];
        layer4[24][55:48] = buffer_data_2[3295:3288];
        layer5[24][7:0] = buffer_data_1[3247:3240];
        layer5[24][15:8] = buffer_data_1[3255:3248];
        layer5[24][23:16] = buffer_data_1[3263:3256];
        layer5[24][31:24] = buffer_data_1[3271:3264];
        layer5[24][39:32] = buffer_data_1[3279:3272];
        layer5[24][47:40] = buffer_data_1[3287:3280];
        layer5[24][55:48] = buffer_data_1[3295:3288];
        layer6[24][7:0] = buffer_data_0[3247:3240];
        layer6[24][15:8] = buffer_data_0[3255:3248];
        layer6[24][23:16] = buffer_data_0[3263:3256];
        layer6[24][31:24] = buffer_data_0[3271:3264];
        layer6[24][39:32] = buffer_data_0[3279:3272];
        layer6[24][47:40] = buffer_data_0[3287:3280];
        layer6[24][55:48] = buffer_data_0[3295:3288];
        layer0[25][7:0] = buffer_data_6[3255:3248];
        layer0[25][15:8] = buffer_data_6[3263:3256];
        layer0[25][23:16] = buffer_data_6[3271:3264];
        layer0[25][31:24] = buffer_data_6[3279:3272];
        layer0[25][39:32] = buffer_data_6[3287:3280];
        layer0[25][47:40] = buffer_data_6[3295:3288];
        layer0[25][55:48] = buffer_data_6[3303:3296];
        layer1[25][7:0] = buffer_data_5[3255:3248];
        layer1[25][15:8] = buffer_data_5[3263:3256];
        layer1[25][23:16] = buffer_data_5[3271:3264];
        layer1[25][31:24] = buffer_data_5[3279:3272];
        layer1[25][39:32] = buffer_data_5[3287:3280];
        layer1[25][47:40] = buffer_data_5[3295:3288];
        layer1[25][55:48] = buffer_data_5[3303:3296];
        layer2[25][7:0] = buffer_data_4[3255:3248];
        layer2[25][15:8] = buffer_data_4[3263:3256];
        layer2[25][23:16] = buffer_data_4[3271:3264];
        layer2[25][31:24] = buffer_data_4[3279:3272];
        layer2[25][39:32] = buffer_data_4[3287:3280];
        layer2[25][47:40] = buffer_data_4[3295:3288];
        layer2[25][55:48] = buffer_data_4[3303:3296];
        layer3[25][7:0] = buffer_data_3[3255:3248];
        layer3[25][15:8] = buffer_data_3[3263:3256];
        layer3[25][23:16] = buffer_data_3[3271:3264];
        layer3[25][31:24] = buffer_data_3[3279:3272];
        layer3[25][39:32] = buffer_data_3[3287:3280];
        layer3[25][47:40] = buffer_data_3[3295:3288];
        layer3[25][55:48] = buffer_data_3[3303:3296];
        layer4[25][7:0] = buffer_data_2[3255:3248];
        layer4[25][15:8] = buffer_data_2[3263:3256];
        layer4[25][23:16] = buffer_data_2[3271:3264];
        layer4[25][31:24] = buffer_data_2[3279:3272];
        layer4[25][39:32] = buffer_data_2[3287:3280];
        layer4[25][47:40] = buffer_data_2[3295:3288];
        layer4[25][55:48] = buffer_data_2[3303:3296];
        layer5[25][7:0] = buffer_data_1[3255:3248];
        layer5[25][15:8] = buffer_data_1[3263:3256];
        layer5[25][23:16] = buffer_data_1[3271:3264];
        layer5[25][31:24] = buffer_data_1[3279:3272];
        layer5[25][39:32] = buffer_data_1[3287:3280];
        layer5[25][47:40] = buffer_data_1[3295:3288];
        layer5[25][55:48] = buffer_data_1[3303:3296];
        layer6[25][7:0] = buffer_data_0[3255:3248];
        layer6[25][15:8] = buffer_data_0[3263:3256];
        layer6[25][23:16] = buffer_data_0[3271:3264];
        layer6[25][31:24] = buffer_data_0[3279:3272];
        layer6[25][39:32] = buffer_data_0[3287:3280];
        layer6[25][47:40] = buffer_data_0[3295:3288];
        layer6[25][55:48] = buffer_data_0[3303:3296];
        layer0[26][7:0] = buffer_data_6[3263:3256];
        layer0[26][15:8] = buffer_data_6[3271:3264];
        layer0[26][23:16] = buffer_data_6[3279:3272];
        layer0[26][31:24] = buffer_data_6[3287:3280];
        layer0[26][39:32] = buffer_data_6[3295:3288];
        layer0[26][47:40] = buffer_data_6[3303:3296];
        layer0[26][55:48] = buffer_data_6[3311:3304];
        layer1[26][7:0] = buffer_data_5[3263:3256];
        layer1[26][15:8] = buffer_data_5[3271:3264];
        layer1[26][23:16] = buffer_data_5[3279:3272];
        layer1[26][31:24] = buffer_data_5[3287:3280];
        layer1[26][39:32] = buffer_data_5[3295:3288];
        layer1[26][47:40] = buffer_data_5[3303:3296];
        layer1[26][55:48] = buffer_data_5[3311:3304];
        layer2[26][7:0] = buffer_data_4[3263:3256];
        layer2[26][15:8] = buffer_data_4[3271:3264];
        layer2[26][23:16] = buffer_data_4[3279:3272];
        layer2[26][31:24] = buffer_data_4[3287:3280];
        layer2[26][39:32] = buffer_data_4[3295:3288];
        layer2[26][47:40] = buffer_data_4[3303:3296];
        layer2[26][55:48] = buffer_data_4[3311:3304];
        layer3[26][7:0] = buffer_data_3[3263:3256];
        layer3[26][15:8] = buffer_data_3[3271:3264];
        layer3[26][23:16] = buffer_data_3[3279:3272];
        layer3[26][31:24] = buffer_data_3[3287:3280];
        layer3[26][39:32] = buffer_data_3[3295:3288];
        layer3[26][47:40] = buffer_data_3[3303:3296];
        layer3[26][55:48] = buffer_data_3[3311:3304];
        layer4[26][7:0] = buffer_data_2[3263:3256];
        layer4[26][15:8] = buffer_data_2[3271:3264];
        layer4[26][23:16] = buffer_data_2[3279:3272];
        layer4[26][31:24] = buffer_data_2[3287:3280];
        layer4[26][39:32] = buffer_data_2[3295:3288];
        layer4[26][47:40] = buffer_data_2[3303:3296];
        layer4[26][55:48] = buffer_data_2[3311:3304];
        layer5[26][7:0] = buffer_data_1[3263:3256];
        layer5[26][15:8] = buffer_data_1[3271:3264];
        layer5[26][23:16] = buffer_data_1[3279:3272];
        layer5[26][31:24] = buffer_data_1[3287:3280];
        layer5[26][39:32] = buffer_data_1[3295:3288];
        layer5[26][47:40] = buffer_data_1[3303:3296];
        layer5[26][55:48] = buffer_data_1[3311:3304];
        layer6[26][7:0] = buffer_data_0[3263:3256];
        layer6[26][15:8] = buffer_data_0[3271:3264];
        layer6[26][23:16] = buffer_data_0[3279:3272];
        layer6[26][31:24] = buffer_data_0[3287:3280];
        layer6[26][39:32] = buffer_data_0[3295:3288];
        layer6[26][47:40] = buffer_data_0[3303:3296];
        layer6[26][55:48] = buffer_data_0[3311:3304];
        layer0[27][7:0] = buffer_data_6[3271:3264];
        layer0[27][15:8] = buffer_data_6[3279:3272];
        layer0[27][23:16] = buffer_data_6[3287:3280];
        layer0[27][31:24] = buffer_data_6[3295:3288];
        layer0[27][39:32] = buffer_data_6[3303:3296];
        layer0[27][47:40] = buffer_data_6[3311:3304];
        layer0[27][55:48] = buffer_data_6[3319:3312];
        layer1[27][7:0] = buffer_data_5[3271:3264];
        layer1[27][15:8] = buffer_data_5[3279:3272];
        layer1[27][23:16] = buffer_data_5[3287:3280];
        layer1[27][31:24] = buffer_data_5[3295:3288];
        layer1[27][39:32] = buffer_data_5[3303:3296];
        layer1[27][47:40] = buffer_data_5[3311:3304];
        layer1[27][55:48] = buffer_data_5[3319:3312];
        layer2[27][7:0] = buffer_data_4[3271:3264];
        layer2[27][15:8] = buffer_data_4[3279:3272];
        layer2[27][23:16] = buffer_data_4[3287:3280];
        layer2[27][31:24] = buffer_data_4[3295:3288];
        layer2[27][39:32] = buffer_data_4[3303:3296];
        layer2[27][47:40] = buffer_data_4[3311:3304];
        layer2[27][55:48] = buffer_data_4[3319:3312];
        layer3[27][7:0] = buffer_data_3[3271:3264];
        layer3[27][15:8] = buffer_data_3[3279:3272];
        layer3[27][23:16] = buffer_data_3[3287:3280];
        layer3[27][31:24] = buffer_data_3[3295:3288];
        layer3[27][39:32] = buffer_data_3[3303:3296];
        layer3[27][47:40] = buffer_data_3[3311:3304];
        layer3[27][55:48] = buffer_data_3[3319:3312];
        layer4[27][7:0] = buffer_data_2[3271:3264];
        layer4[27][15:8] = buffer_data_2[3279:3272];
        layer4[27][23:16] = buffer_data_2[3287:3280];
        layer4[27][31:24] = buffer_data_2[3295:3288];
        layer4[27][39:32] = buffer_data_2[3303:3296];
        layer4[27][47:40] = buffer_data_2[3311:3304];
        layer4[27][55:48] = buffer_data_2[3319:3312];
        layer5[27][7:0] = buffer_data_1[3271:3264];
        layer5[27][15:8] = buffer_data_1[3279:3272];
        layer5[27][23:16] = buffer_data_1[3287:3280];
        layer5[27][31:24] = buffer_data_1[3295:3288];
        layer5[27][39:32] = buffer_data_1[3303:3296];
        layer5[27][47:40] = buffer_data_1[3311:3304];
        layer5[27][55:48] = buffer_data_1[3319:3312];
        layer6[27][7:0] = buffer_data_0[3271:3264];
        layer6[27][15:8] = buffer_data_0[3279:3272];
        layer6[27][23:16] = buffer_data_0[3287:3280];
        layer6[27][31:24] = buffer_data_0[3295:3288];
        layer6[27][39:32] = buffer_data_0[3303:3296];
        layer6[27][47:40] = buffer_data_0[3311:3304];
        layer6[27][55:48] = buffer_data_0[3319:3312];
        layer0[28][7:0] = buffer_data_6[3279:3272];
        layer0[28][15:8] = buffer_data_6[3287:3280];
        layer0[28][23:16] = buffer_data_6[3295:3288];
        layer0[28][31:24] = buffer_data_6[3303:3296];
        layer0[28][39:32] = buffer_data_6[3311:3304];
        layer0[28][47:40] = buffer_data_6[3319:3312];
        layer0[28][55:48] = buffer_data_6[3327:3320];
        layer1[28][7:0] = buffer_data_5[3279:3272];
        layer1[28][15:8] = buffer_data_5[3287:3280];
        layer1[28][23:16] = buffer_data_5[3295:3288];
        layer1[28][31:24] = buffer_data_5[3303:3296];
        layer1[28][39:32] = buffer_data_5[3311:3304];
        layer1[28][47:40] = buffer_data_5[3319:3312];
        layer1[28][55:48] = buffer_data_5[3327:3320];
        layer2[28][7:0] = buffer_data_4[3279:3272];
        layer2[28][15:8] = buffer_data_4[3287:3280];
        layer2[28][23:16] = buffer_data_4[3295:3288];
        layer2[28][31:24] = buffer_data_4[3303:3296];
        layer2[28][39:32] = buffer_data_4[3311:3304];
        layer2[28][47:40] = buffer_data_4[3319:3312];
        layer2[28][55:48] = buffer_data_4[3327:3320];
        layer3[28][7:0] = buffer_data_3[3279:3272];
        layer3[28][15:8] = buffer_data_3[3287:3280];
        layer3[28][23:16] = buffer_data_3[3295:3288];
        layer3[28][31:24] = buffer_data_3[3303:3296];
        layer3[28][39:32] = buffer_data_3[3311:3304];
        layer3[28][47:40] = buffer_data_3[3319:3312];
        layer3[28][55:48] = buffer_data_3[3327:3320];
        layer4[28][7:0] = buffer_data_2[3279:3272];
        layer4[28][15:8] = buffer_data_2[3287:3280];
        layer4[28][23:16] = buffer_data_2[3295:3288];
        layer4[28][31:24] = buffer_data_2[3303:3296];
        layer4[28][39:32] = buffer_data_2[3311:3304];
        layer4[28][47:40] = buffer_data_2[3319:3312];
        layer4[28][55:48] = buffer_data_2[3327:3320];
        layer5[28][7:0] = buffer_data_1[3279:3272];
        layer5[28][15:8] = buffer_data_1[3287:3280];
        layer5[28][23:16] = buffer_data_1[3295:3288];
        layer5[28][31:24] = buffer_data_1[3303:3296];
        layer5[28][39:32] = buffer_data_1[3311:3304];
        layer5[28][47:40] = buffer_data_1[3319:3312];
        layer5[28][55:48] = buffer_data_1[3327:3320];
        layer6[28][7:0] = buffer_data_0[3279:3272];
        layer6[28][15:8] = buffer_data_0[3287:3280];
        layer6[28][23:16] = buffer_data_0[3295:3288];
        layer6[28][31:24] = buffer_data_0[3303:3296];
        layer6[28][39:32] = buffer_data_0[3311:3304];
        layer6[28][47:40] = buffer_data_0[3319:3312];
        layer6[28][55:48] = buffer_data_0[3327:3320];
        layer0[29][7:0] = buffer_data_6[3287:3280];
        layer0[29][15:8] = buffer_data_6[3295:3288];
        layer0[29][23:16] = buffer_data_6[3303:3296];
        layer0[29][31:24] = buffer_data_6[3311:3304];
        layer0[29][39:32] = buffer_data_6[3319:3312];
        layer0[29][47:40] = buffer_data_6[3327:3320];
        layer0[29][55:48] = buffer_data_6[3335:3328];
        layer1[29][7:0] = buffer_data_5[3287:3280];
        layer1[29][15:8] = buffer_data_5[3295:3288];
        layer1[29][23:16] = buffer_data_5[3303:3296];
        layer1[29][31:24] = buffer_data_5[3311:3304];
        layer1[29][39:32] = buffer_data_5[3319:3312];
        layer1[29][47:40] = buffer_data_5[3327:3320];
        layer1[29][55:48] = buffer_data_5[3335:3328];
        layer2[29][7:0] = buffer_data_4[3287:3280];
        layer2[29][15:8] = buffer_data_4[3295:3288];
        layer2[29][23:16] = buffer_data_4[3303:3296];
        layer2[29][31:24] = buffer_data_4[3311:3304];
        layer2[29][39:32] = buffer_data_4[3319:3312];
        layer2[29][47:40] = buffer_data_4[3327:3320];
        layer2[29][55:48] = buffer_data_4[3335:3328];
        layer3[29][7:0] = buffer_data_3[3287:3280];
        layer3[29][15:8] = buffer_data_3[3295:3288];
        layer3[29][23:16] = buffer_data_3[3303:3296];
        layer3[29][31:24] = buffer_data_3[3311:3304];
        layer3[29][39:32] = buffer_data_3[3319:3312];
        layer3[29][47:40] = buffer_data_3[3327:3320];
        layer3[29][55:48] = buffer_data_3[3335:3328];
        layer4[29][7:0] = buffer_data_2[3287:3280];
        layer4[29][15:8] = buffer_data_2[3295:3288];
        layer4[29][23:16] = buffer_data_2[3303:3296];
        layer4[29][31:24] = buffer_data_2[3311:3304];
        layer4[29][39:32] = buffer_data_2[3319:3312];
        layer4[29][47:40] = buffer_data_2[3327:3320];
        layer4[29][55:48] = buffer_data_2[3335:3328];
        layer5[29][7:0] = buffer_data_1[3287:3280];
        layer5[29][15:8] = buffer_data_1[3295:3288];
        layer5[29][23:16] = buffer_data_1[3303:3296];
        layer5[29][31:24] = buffer_data_1[3311:3304];
        layer5[29][39:32] = buffer_data_1[3319:3312];
        layer5[29][47:40] = buffer_data_1[3327:3320];
        layer5[29][55:48] = buffer_data_1[3335:3328];
        layer6[29][7:0] = buffer_data_0[3287:3280];
        layer6[29][15:8] = buffer_data_0[3295:3288];
        layer6[29][23:16] = buffer_data_0[3303:3296];
        layer6[29][31:24] = buffer_data_0[3311:3304];
        layer6[29][39:32] = buffer_data_0[3319:3312];
        layer6[29][47:40] = buffer_data_0[3327:3320];
        layer6[29][55:48] = buffer_data_0[3335:3328];
        layer0[30][7:0] = buffer_data_6[3295:3288];
        layer0[30][15:8] = buffer_data_6[3303:3296];
        layer0[30][23:16] = buffer_data_6[3311:3304];
        layer0[30][31:24] = buffer_data_6[3319:3312];
        layer0[30][39:32] = buffer_data_6[3327:3320];
        layer0[30][47:40] = buffer_data_6[3335:3328];
        layer0[30][55:48] = buffer_data_6[3343:3336];
        layer1[30][7:0] = buffer_data_5[3295:3288];
        layer1[30][15:8] = buffer_data_5[3303:3296];
        layer1[30][23:16] = buffer_data_5[3311:3304];
        layer1[30][31:24] = buffer_data_5[3319:3312];
        layer1[30][39:32] = buffer_data_5[3327:3320];
        layer1[30][47:40] = buffer_data_5[3335:3328];
        layer1[30][55:48] = buffer_data_5[3343:3336];
        layer2[30][7:0] = buffer_data_4[3295:3288];
        layer2[30][15:8] = buffer_data_4[3303:3296];
        layer2[30][23:16] = buffer_data_4[3311:3304];
        layer2[30][31:24] = buffer_data_4[3319:3312];
        layer2[30][39:32] = buffer_data_4[3327:3320];
        layer2[30][47:40] = buffer_data_4[3335:3328];
        layer2[30][55:48] = buffer_data_4[3343:3336];
        layer3[30][7:0] = buffer_data_3[3295:3288];
        layer3[30][15:8] = buffer_data_3[3303:3296];
        layer3[30][23:16] = buffer_data_3[3311:3304];
        layer3[30][31:24] = buffer_data_3[3319:3312];
        layer3[30][39:32] = buffer_data_3[3327:3320];
        layer3[30][47:40] = buffer_data_3[3335:3328];
        layer3[30][55:48] = buffer_data_3[3343:3336];
        layer4[30][7:0] = buffer_data_2[3295:3288];
        layer4[30][15:8] = buffer_data_2[3303:3296];
        layer4[30][23:16] = buffer_data_2[3311:3304];
        layer4[30][31:24] = buffer_data_2[3319:3312];
        layer4[30][39:32] = buffer_data_2[3327:3320];
        layer4[30][47:40] = buffer_data_2[3335:3328];
        layer4[30][55:48] = buffer_data_2[3343:3336];
        layer5[30][7:0] = buffer_data_1[3295:3288];
        layer5[30][15:8] = buffer_data_1[3303:3296];
        layer5[30][23:16] = buffer_data_1[3311:3304];
        layer5[30][31:24] = buffer_data_1[3319:3312];
        layer5[30][39:32] = buffer_data_1[3327:3320];
        layer5[30][47:40] = buffer_data_1[3335:3328];
        layer5[30][55:48] = buffer_data_1[3343:3336];
        layer6[30][7:0] = buffer_data_0[3295:3288];
        layer6[30][15:8] = buffer_data_0[3303:3296];
        layer6[30][23:16] = buffer_data_0[3311:3304];
        layer6[30][31:24] = buffer_data_0[3319:3312];
        layer6[30][39:32] = buffer_data_0[3327:3320];
        layer6[30][47:40] = buffer_data_0[3335:3328];
        layer6[30][55:48] = buffer_data_0[3343:3336];
        layer0[31][7:0] = buffer_data_6[3303:3296];
        layer0[31][15:8] = buffer_data_6[3311:3304];
        layer0[31][23:16] = buffer_data_6[3319:3312];
        layer0[31][31:24] = buffer_data_6[3327:3320];
        layer0[31][39:32] = buffer_data_6[3335:3328];
        layer0[31][47:40] = buffer_data_6[3343:3336];
        layer0[31][55:48] = buffer_data_6[3351:3344];
        layer1[31][7:0] = buffer_data_5[3303:3296];
        layer1[31][15:8] = buffer_data_5[3311:3304];
        layer1[31][23:16] = buffer_data_5[3319:3312];
        layer1[31][31:24] = buffer_data_5[3327:3320];
        layer1[31][39:32] = buffer_data_5[3335:3328];
        layer1[31][47:40] = buffer_data_5[3343:3336];
        layer1[31][55:48] = buffer_data_5[3351:3344];
        layer2[31][7:0] = buffer_data_4[3303:3296];
        layer2[31][15:8] = buffer_data_4[3311:3304];
        layer2[31][23:16] = buffer_data_4[3319:3312];
        layer2[31][31:24] = buffer_data_4[3327:3320];
        layer2[31][39:32] = buffer_data_4[3335:3328];
        layer2[31][47:40] = buffer_data_4[3343:3336];
        layer2[31][55:48] = buffer_data_4[3351:3344];
        layer3[31][7:0] = buffer_data_3[3303:3296];
        layer3[31][15:8] = buffer_data_3[3311:3304];
        layer3[31][23:16] = buffer_data_3[3319:3312];
        layer3[31][31:24] = buffer_data_3[3327:3320];
        layer3[31][39:32] = buffer_data_3[3335:3328];
        layer3[31][47:40] = buffer_data_3[3343:3336];
        layer3[31][55:48] = buffer_data_3[3351:3344];
        layer4[31][7:0] = buffer_data_2[3303:3296];
        layer4[31][15:8] = buffer_data_2[3311:3304];
        layer4[31][23:16] = buffer_data_2[3319:3312];
        layer4[31][31:24] = buffer_data_2[3327:3320];
        layer4[31][39:32] = buffer_data_2[3335:3328];
        layer4[31][47:40] = buffer_data_2[3343:3336];
        layer4[31][55:48] = buffer_data_2[3351:3344];
        layer5[31][7:0] = buffer_data_1[3303:3296];
        layer5[31][15:8] = buffer_data_1[3311:3304];
        layer5[31][23:16] = buffer_data_1[3319:3312];
        layer5[31][31:24] = buffer_data_1[3327:3320];
        layer5[31][39:32] = buffer_data_1[3335:3328];
        layer5[31][47:40] = buffer_data_1[3343:3336];
        layer5[31][55:48] = buffer_data_1[3351:3344];
        layer6[31][7:0] = buffer_data_0[3303:3296];
        layer6[31][15:8] = buffer_data_0[3311:3304];
        layer6[31][23:16] = buffer_data_0[3319:3312];
        layer6[31][31:24] = buffer_data_0[3327:3320];
        layer6[31][39:32] = buffer_data_0[3335:3328];
        layer6[31][47:40] = buffer_data_0[3343:3336];
        layer6[31][55:48] = buffer_data_0[3351:3344];
        layer0[32][7:0] = buffer_data_6[3311:3304];
        layer0[32][15:8] = buffer_data_6[3319:3312];
        layer0[32][23:16] = buffer_data_6[3327:3320];
        layer0[32][31:24] = buffer_data_6[3335:3328];
        layer0[32][39:32] = buffer_data_6[3343:3336];
        layer0[32][47:40] = buffer_data_6[3351:3344];
        layer0[32][55:48] = buffer_data_6[3359:3352];
        layer1[32][7:0] = buffer_data_5[3311:3304];
        layer1[32][15:8] = buffer_data_5[3319:3312];
        layer1[32][23:16] = buffer_data_5[3327:3320];
        layer1[32][31:24] = buffer_data_5[3335:3328];
        layer1[32][39:32] = buffer_data_5[3343:3336];
        layer1[32][47:40] = buffer_data_5[3351:3344];
        layer1[32][55:48] = buffer_data_5[3359:3352];
        layer2[32][7:0] = buffer_data_4[3311:3304];
        layer2[32][15:8] = buffer_data_4[3319:3312];
        layer2[32][23:16] = buffer_data_4[3327:3320];
        layer2[32][31:24] = buffer_data_4[3335:3328];
        layer2[32][39:32] = buffer_data_4[3343:3336];
        layer2[32][47:40] = buffer_data_4[3351:3344];
        layer2[32][55:48] = buffer_data_4[3359:3352];
        layer3[32][7:0] = buffer_data_3[3311:3304];
        layer3[32][15:8] = buffer_data_3[3319:3312];
        layer3[32][23:16] = buffer_data_3[3327:3320];
        layer3[32][31:24] = buffer_data_3[3335:3328];
        layer3[32][39:32] = buffer_data_3[3343:3336];
        layer3[32][47:40] = buffer_data_3[3351:3344];
        layer3[32][55:48] = buffer_data_3[3359:3352];
        layer4[32][7:0] = buffer_data_2[3311:3304];
        layer4[32][15:8] = buffer_data_2[3319:3312];
        layer4[32][23:16] = buffer_data_2[3327:3320];
        layer4[32][31:24] = buffer_data_2[3335:3328];
        layer4[32][39:32] = buffer_data_2[3343:3336];
        layer4[32][47:40] = buffer_data_2[3351:3344];
        layer4[32][55:48] = buffer_data_2[3359:3352];
        layer5[32][7:0] = buffer_data_1[3311:3304];
        layer5[32][15:8] = buffer_data_1[3319:3312];
        layer5[32][23:16] = buffer_data_1[3327:3320];
        layer5[32][31:24] = buffer_data_1[3335:3328];
        layer5[32][39:32] = buffer_data_1[3343:3336];
        layer5[32][47:40] = buffer_data_1[3351:3344];
        layer5[32][55:48] = buffer_data_1[3359:3352];
        layer6[32][7:0] = buffer_data_0[3311:3304];
        layer6[32][15:8] = buffer_data_0[3319:3312];
        layer6[32][23:16] = buffer_data_0[3327:3320];
        layer6[32][31:24] = buffer_data_0[3335:3328];
        layer6[32][39:32] = buffer_data_0[3343:3336];
        layer6[32][47:40] = buffer_data_0[3351:3344];
        layer6[32][55:48] = buffer_data_0[3359:3352];
        layer0[33][7:0] = buffer_data_6[3319:3312];
        layer0[33][15:8] = buffer_data_6[3327:3320];
        layer0[33][23:16] = buffer_data_6[3335:3328];
        layer0[33][31:24] = buffer_data_6[3343:3336];
        layer0[33][39:32] = buffer_data_6[3351:3344];
        layer0[33][47:40] = buffer_data_6[3359:3352];
        layer0[33][55:48] = buffer_data_6[3367:3360];
        layer1[33][7:0] = buffer_data_5[3319:3312];
        layer1[33][15:8] = buffer_data_5[3327:3320];
        layer1[33][23:16] = buffer_data_5[3335:3328];
        layer1[33][31:24] = buffer_data_5[3343:3336];
        layer1[33][39:32] = buffer_data_5[3351:3344];
        layer1[33][47:40] = buffer_data_5[3359:3352];
        layer1[33][55:48] = buffer_data_5[3367:3360];
        layer2[33][7:0] = buffer_data_4[3319:3312];
        layer2[33][15:8] = buffer_data_4[3327:3320];
        layer2[33][23:16] = buffer_data_4[3335:3328];
        layer2[33][31:24] = buffer_data_4[3343:3336];
        layer2[33][39:32] = buffer_data_4[3351:3344];
        layer2[33][47:40] = buffer_data_4[3359:3352];
        layer2[33][55:48] = buffer_data_4[3367:3360];
        layer3[33][7:0] = buffer_data_3[3319:3312];
        layer3[33][15:8] = buffer_data_3[3327:3320];
        layer3[33][23:16] = buffer_data_3[3335:3328];
        layer3[33][31:24] = buffer_data_3[3343:3336];
        layer3[33][39:32] = buffer_data_3[3351:3344];
        layer3[33][47:40] = buffer_data_3[3359:3352];
        layer3[33][55:48] = buffer_data_3[3367:3360];
        layer4[33][7:0] = buffer_data_2[3319:3312];
        layer4[33][15:8] = buffer_data_2[3327:3320];
        layer4[33][23:16] = buffer_data_2[3335:3328];
        layer4[33][31:24] = buffer_data_2[3343:3336];
        layer4[33][39:32] = buffer_data_2[3351:3344];
        layer4[33][47:40] = buffer_data_2[3359:3352];
        layer4[33][55:48] = buffer_data_2[3367:3360];
        layer5[33][7:0] = buffer_data_1[3319:3312];
        layer5[33][15:8] = buffer_data_1[3327:3320];
        layer5[33][23:16] = buffer_data_1[3335:3328];
        layer5[33][31:24] = buffer_data_1[3343:3336];
        layer5[33][39:32] = buffer_data_1[3351:3344];
        layer5[33][47:40] = buffer_data_1[3359:3352];
        layer5[33][55:48] = buffer_data_1[3367:3360];
        layer6[33][7:0] = buffer_data_0[3319:3312];
        layer6[33][15:8] = buffer_data_0[3327:3320];
        layer6[33][23:16] = buffer_data_0[3335:3328];
        layer6[33][31:24] = buffer_data_0[3343:3336];
        layer6[33][39:32] = buffer_data_0[3351:3344];
        layer6[33][47:40] = buffer_data_0[3359:3352];
        layer6[33][55:48] = buffer_data_0[3367:3360];
        layer0[34][7:0] = buffer_data_6[3327:3320];
        layer0[34][15:8] = buffer_data_6[3335:3328];
        layer0[34][23:16] = buffer_data_6[3343:3336];
        layer0[34][31:24] = buffer_data_6[3351:3344];
        layer0[34][39:32] = buffer_data_6[3359:3352];
        layer0[34][47:40] = buffer_data_6[3367:3360];
        layer0[34][55:48] = buffer_data_6[3375:3368];
        layer1[34][7:0] = buffer_data_5[3327:3320];
        layer1[34][15:8] = buffer_data_5[3335:3328];
        layer1[34][23:16] = buffer_data_5[3343:3336];
        layer1[34][31:24] = buffer_data_5[3351:3344];
        layer1[34][39:32] = buffer_data_5[3359:3352];
        layer1[34][47:40] = buffer_data_5[3367:3360];
        layer1[34][55:48] = buffer_data_5[3375:3368];
        layer2[34][7:0] = buffer_data_4[3327:3320];
        layer2[34][15:8] = buffer_data_4[3335:3328];
        layer2[34][23:16] = buffer_data_4[3343:3336];
        layer2[34][31:24] = buffer_data_4[3351:3344];
        layer2[34][39:32] = buffer_data_4[3359:3352];
        layer2[34][47:40] = buffer_data_4[3367:3360];
        layer2[34][55:48] = buffer_data_4[3375:3368];
        layer3[34][7:0] = buffer_data_3[3327:3320];
        layer3[34][15:8] = buffer_data_3[3335:3328];
        layer3[34][23:16] = buffer_data_3[3343:3336];
        layer3[34][31:24] = buffer_data_3[3351:3344];
        layer3[34][39:32] = buffer_data_3[3359:3352];
        layer3[34][47:40] = buffer_data_3[3367:3360];
        layer3[34][55:48] = buffer_data_3[3375:3368];
        layer4[34][7:0] = buffer_data_2[3327:3320];
        layer4[34][15:8] = buffer_data_2[3335:3328];
        layer4[34][23:16] = buffer_data_2[3343:3336];
        layer4[34][31:24] = buffer_data_2[3351:3344];
        layer4[34][39:32] = buffer_data_2[3359:3352];
        layer4[34][47:40] = buffer_data_2[3367:3360];
        layer4[34][55:48] = buffer_data_2[3375:3368];
        layer5[34][7:0] = buffer_data_1[3327:3320];
        layer5[34][15:8] = buffer_data_1[3335:3328];
        layer5[34][23:16] = buffer_data_1[3343:3336];
        layer5[34][31:24] = buffer_data_1[3351:3344];
        layer5[34][39:32] = buffer_data_1[3359:3352];
        layer5[34][47:40] = buffer_data_1[3367:3360];
        layer5[34][55:48] = buffer_data_1[3375:3368];
        layer6[34][7:0] = buffer_data_0[3327:3320];
        layer6[34][15:8] = buffer_data_0[3335:3328];
        layer6[34][23:16] = buffer_data_0[3343:3336];
        layer6[34][31:24] = buffer_data_0[3351:3344];
        layer6[34][39:32] = buffer_data_0[3359:3352];
        layer6[34][47:40] = buffer_data_0[3367:3360];
        layer6[34][55:48] = buffer_data_0[3375:3368];
        layer0[35][7:0] = buffer_data_6[3335:3328];
        layer0[35][15:8] = buffer_data_6[3343:3336];
        layer0[35][23:16] = buffer_data_6[3351:3344];
        layer0[35][31:24] = buffer_data_6[3359:3352];
        layer0[35][39:32] = buffer_data_6[3367:3360];
        layer0[35][47:40] = buffer_data_6[3375:3368];
        layer0[35][55:48] = buffer_data_6[3383:3376];
        layer1[35][7:0] = buffer_data_5[3335:3328];
        layer1[35][15:8] = buffer_data_5[3343:3336];
        layer1[35][23:16] = buffer_data_5[3351:3344];
        layer1[35][31:24] = buffer_data_5[3359:3352];
        layer1[35][39:32] = buffer_data_5[3367:3360];
        layer1[35][47:40] = buffer_data_5[3375:3368];
        layer1[35][55:48] = buffer_data_5[3383:3376];
        layer2[35][7:0] = buffer_data_4[3335:3328];
        layer2[35][15:8] = buffer_data_4[3343:3336];
        layer2[35][23:16] = buffer_data_4[3351:3344];
        layer2[35][31:24] = buffer_data_4[3359:3352];
        layer2[35][39:32] = buffer_data_4[3367:3360];
        layer2[35][47:40] = buffer_data_4[3375:3368];
        layer2[35][55:48] = buffer_data_4[3383:3376];
        layer3[35][7:0] = buffer_data_3[3335:3328];
        layer3[35][15:8] = buffer_data_3[3343:3336];
        layer3[35][23:16] = buffer_data_3[3351:3344];
        layer3[35][31:24] = buffer_data_3[3359:3352];
        layer3[35][39:32] = buffer_data_3[3367:3360];
        layer3[35][47:40] = buffer_data_3[3375:3368];
        layer3[35][55:48] = buffer_data_3[3383:3376];
        layer4[35][7:0] = buffer_data_2[3335:3328];
        layer4[35][15:8] = buffer_data_2[3343:3336];
        layer4[35][23:16] = buffer_data_2[3351:3344];
        layer4[35][31:24] = buffer_data_2[3359:3352];
        layer4[35][39:32] = buffer_data_2[3367:3360];
        layer4[35][47:40] = buffer_data_2[3375:3368];
        layer4[35][55:48] = buffer_data_2[3383:3376];
        layer5[35][7:0] = buffer_data_1[3335:3328];
        layer5[35][15:8] = buffer_data_1[3343:3336];
        layer5[35][23:16] = buffer_data_1[3351:3344];
        layer5[35][31:24] = buffer_data_1[3359:3352];
        layer5[35][39:32] = buffer_data_1[3367:3360];
        layer5[35][47:40] = buffer_data_1[3375:3368];
        layer5[35][55:48] = buffer_data_1[3383:3376];
        layer6[35][7:0] = buffer_data_0[3335:3328];
        layer6[35][15:8] = buffer_data_0[3343:3336];
        layer6[35][23:16] = buffer_data_0[3351:3344];
        layer6[35][31:24] = buffer_data_0[3359:3352];
        layer6[35][39:32] = buffer_data_0[3367:3360];
        layer6[35][47:40] = buffer_data_0[3375:3368];
        layer6[35][55:48] = buffer_data_0[3383:3376];
        layer0[36][7:0] = buffer_data_6[3343:3336];
        layer0[36][15:8] = buffer_data_6[3351:3344];
        layer0[36][23:16] = buffer_data_6[3359:3352];
        layer0[36][31:24] = buffer_data_6[3367:3360];
        layer0[36][39:32] = buffer_data_6[3375:3368];
        layer0[36][47:40] = buffer_data_6[3383:3376];
        layer0[36][55:48] = buffer_data_6[3391:3384];
        layer1[36][7:0] = buffer_data_5[3343:3336];
        layer1[36][15:8] = buffer_data_5[3351:3344];
        layer1[36][23:16] = buffer_data_5[3359:3352];
        layer1[36][31:24] = buffer_data_5[3367:3360];
        layer1[36][39:32] = buffer_data_5[3375:3368];
        layer1[36][47:40] = buffer_data_5[3383:3376];
        layer1[36][55:48] = buffer_data_5[3391:3384];
        layer2[36][7:0] = buffer_data_4[3343:3336];
        layer2[36][15:8] = buffer_data_4[3351:3344];
        layer2[36][23:16] = buffer_data_4[3359:3352];
        layer2[36][31:24] = buffer_data_4[3367:3360];
        layer2[36][39:32] = buffer_data_4[3375:3368];
        layer2[36][47:40] = buffer_data_4[3383:3376];
        layer2[36][55:48] = buffer_data_4[3391:3384];
        layer3[36][7:0] = buffer_data_3[3343:3336];
        layer3[36][15:8] = buffer_data_3[3351:3344];
        layer3[36][23:16] = buffer_data_3[3359:3352];
        layer3[36][31:24] = buffer_data_3[3367:3360];
        layer3[36][39:32] = buffer_data_3[3375:3368];
        layer3[36][47:40] = buffer_data_3[3383:3376];
        layer3[36][55:48] = buffer_data_3[3391:3384];
        layer4[36][7:0] = buffer_data_2[3343:3336];
        layer4[36][15:8] = buffer_data_2[3351:3344];
        layer4[36][23:16] = buffer_data_2[3359:3352];
        layer4[36][31:24] = buffer_data_2[3367:3360];
        layer4[36][39:32] = buffer_data_2[3375:3368];
        layer4[36][47:40] = buffer_data_2[3383:3376];
        layer4[36][55:48] = buffer_data_2[3391:3384];
        layer5[36][7:0] = buffer_data_1[3343:3336];
        layer5[36][15:8] = buffer_data_1[3351:3344];
        layer5[36][23:16] = buffer_data_1[3359:3352];
        layer5[36][31:24] = buffer_data_1[3367:3360];
        layer5[36][39:32] = buffer_data_1[3375:3368];
        layer5[36][47:40] = buffer_data_1[3383:3376];
        layer5[36][55:48] = buffer_data_1[3391:3384];
        layer6[36][7:0] = buffer_data_0[3343:3336];
        layer6[36][15:8] = buffer_data_0[3351:3344];
        layer6[36][23:16] = buffer_data_0[3359:3352];
        layer6[36][31:24] = buffer_data_0[3367:3360];
        layer6[36][39:32] = buffer_data_0[3375:3368];
        layer6[36][47:40] = buffer_data_0[3383:3376];
        layer6[36][55:48] = buffer_data_0[3391:3384];
        layer0[37][7:0] = buffer_data_6[3351:3344];
        layer0[37][15:8] = buffer_data_6[3359:3352];
        layer0[37][23:16] = buffer_data_6[3367:3360];
        layer0[37][31:24] = buffer_data_6[3375:3368];
        layer0[37][39:32] = buffer_data_6[3383:3376];
        layer0[37][47:40] = buffer_data_6[3391:3384];
        layer0[37][55:48] = buffer_data_6[3399:3392];
        layer1[37][7:0] = buffer_data_5[3351:3344];
        layer1[37][15:8] = buffer_data_5[3359:3352];
        layer1[37][23:16] = buffer_data_5[3367:3360];
        layer1[37][31:24] = buffer_data_5[3375:3368];
        layer1[37][39:32] = buffer_data_5[3383:3376];
        layer1[37][47:40] = buffer_data_5[3391:3384];
        layer1[37][55:48] = buffer_data_5[3399:3392];
        layer2[37][7:0] = buffer_data_4[3351:3344];
        layer2[37][15:8] = buffer_data_4[3359:3352];
        layer2[37][23:16] = buffer_data_4[3367:3360];
        layer2[37][31:24] = buffer_data_4[3375:3368];
        layer2[37][39:32] = buffer_data_4[3383:3376];
        layer2[37][47:40] = buffer_data_4[3391:3384];
        layer2[37][55:48] = buffer_data_4[3399:3392];
        layer3[37][7:0] = buffer_data_3[3351:3344];
        layer3[37][15:8] = buffer_data_3[3359:3352];
        layer3[37][23:16] = buffer_data_3[3367:3360];
        layer3[37][31:24] = buffer_data_3[3375:3368];
        layer3[37][39:32] = buffer_data_3[3383:3376];
        layer3[37][47:40] = buffer_data_3[3391:3384];
        layer3[37][55:48] = buffer_data_3[3399:3392];
        layer4[37][7:0] = buffer_data_2[3351:3344];
        layer4[37][15:8] = buffer_data_2[3359:3352];
        layer4[37][23:16] = buffer_data_2[3367:3360];
        layer4[37][31:24] = buffer_data_2[3375:3368];
        layer4[37][39:32] = buffer_data_2[3383:3376];
        layer4[37][47:40] = buffer_data_2[3391:3384];
        layer4[37][55:48] = buffer_data_2[3399:3392];
        layer5[37][7:0] = buffer_data_1[3351:3344];
        layer5[37][15:8] = buffer_data_1[3359:3352];
        layer5[37][23:16] = buffer_data_1[3367:3360];
        layer5[37][31:24] = buffer_data_1[3375:3368];
        layer5[37][39:32] = buffer_data_1[3383:3376];
        layer5[37][47:40] = buffer_data_1[3391:3384];
        layer5[37][55:48] = buffer_data_1[3399:3392];
        layer6[37][7:0] = buffer_data_0[3351:3344];
        layer6[37][15:8] = buffer_data_0[3359:3352];
        layer6[37][23:16] = buffer_data_0[3367:3360];
        layer6[37][31:24] = buffer_data_0[3375:3368];
        layer6[37][39:32] = buffer_data_0[3383:3376];
        layer6[37][47:40] = buffer_data_0[3391:3384];
        layer6[37][55:48] = buffer_data_0[3399:3392];
        layer0[38][7:0] = buffer_data_6[3359:3352];
        layer0[38][15:8] = buffer_data_6[3367:3360];
        layer0[38][23:16] = buffer_data_6[3375:3368];
        layer0[38][31:24] = buffer_data_6[3383:3376];
        layer0[38][39:32] = buffer_data_6[3391:3384];
        layer0[38][47:40] = buffer_data_6[3399:3392];
        layer0[38][55:48] = buffer_data_6[3407:3400];
        layer1[38][7:0] = buffer_data_5[3359:3352];
        layer1[38][15:8] = buffer_data_5[3367:3360];
        layer1[38][23:16] = buffer_data_5[3375:3368];
        layer1[38][31:24] = buffer_data_5[3383:3376];
        layer1[38][39:32] = buffer_data_5[3391:3384];
        layer1[38][47:40] = buffer_data_5[3399:3392];
        layer1[38][55:48] = buffer_data_5[3407:3400];
        layer2[38][7:0] = buffer_data_4[3359:3352];
        layer2[38][15:8] = buffer_data_4[3367:3360];
        layer2[38][23:16] = buffer_data_4[3375:3368];
        layer2[38][31:24] = buffer_data_4[3383:3376];
        layer2[38][39:32] = buffer_data_4[3391:3384];
        layer2[38][47:40] = buffer_data_4[3399:3392];
        layer2[38][55:48] = buffer_data_4[3407:3400];
        layer3[38][7:0] = buffer_data_3[3359:3352];
        layer3[38][15:8] = buffer_data_3[3367:3360];
        layer3[38][23:16] = buffer_data_3[3375:3368];
        layer3[38][31:24] = buffer_data_3[3383:3376];
        layer3[38][39:32] = buffer_data_3[3391:3384];
        layer3[38][47:40] = buffer_data_3[3399:3392];
        layer3[38][55:48] = buffer_data_3[3407:3400];
        layer4[38][7:0] = buffer_data_2[3359:3352];
        layer4[38][15:8] = buffer_data_2[3367:3360];
        layer4[38][23:16] = buffer_data_2[3375:3368];
        layer4[38][31:24] = buffer_data_2[3383:3376];
        layer4[38][39:32] = buffer_data_2[3391:3384];
        layer4[38][47:40] = buffer_data_2[3399:3392];
        layer4[38][55:48] = buffer_data_2[3407:3400];
        layer5[38][7:0] = buffer_data_1[3359:3352];
        layer5[38][15:8] = buffer_data_1[3367:3360];
        layer5[38][23:16] = buffer_data_1[3375:3368];
        layer5[38][31:24] = buffer_data_1[3383:3376];
        layer5[38][39:32] = buffer_data_1[3391:3384];
        layer5[38][47:40] = buffer_data_1[3399:3392];
        layer5[38][55:48] = buffer_data_1[3407:3400];
        layer6[38][7:0] = buffer_data_0[3359:3352];
        layer6[38][15:8] = buffer_data_0[3367:3360];
        layer6[38][23:16] = buffer_data_0[3375:3368];
        layer6[38][31:24] = buffer_data_0[3383:3376];
        layer6[38][39:32] = buffer_data_0[3391:3384];
        layer6[38][47:40] = buffer_data_0[3399:3392];
        layer6[38][55:48] = buffer_data_0[3407:3400];
        layer0[39][7:0] = buffer_data_6[3367:3360];
        layer0[39][15:8] = buffer_data_6[3375:3368];
        layer0[39][23:16] = buffer_data_6[3383:3376];
        layer0[39][31:24] = buffer_data_6[3391:3384];
        layer0[39][39:32] = buffer_data_6[3399:3392];
        layer0[39][47:40] = buffer_data_6[3407:3400];
        layer0[39][55:48] = buffer_data_6[3415:3408];
        layer1[39][7:0] = buffer_data_5[3367:3360];
        layer1[39][15:8] = buffer_data_5[3375:3368];
        layer1[39][23:16] = buffer_data_5[3383:3376];
        layer1[39][31:24] = buffer_data_5[3391:3384];
        layer1[39][39:32] = buffer_data_5[3399:3392];
        layer1[39][47:40] = buffer_data_5[3407:3400];
        layer1[39][55:48] = buffer_data_5[3415:3408];
        layer2[39][7:0] = buffer_data_4[3367:3360];
        layer2[39][15:8] = buffer_data_4[3375:3368];
        layer2[39][23:16] = buffer_data_4[3383:3376];
        layer2[39][31:24] = buffer_data_4[3391:3384];
        layer2[39][39:32] = buffer_data_4[3399:3392];
        layer2[39][47:40] = buffer_data_4[3407:3400];
        layer2[39][55:48] = buffer_data_4[3415:3408];
        layer3[39][7:0] = buffer_data_3[3367:3360];
        layer3[39][15:8] = buffer_data_3[3375:3368];
        layer3[39][23:16] = buffer_data_3[3383:3376];
        layer3[39][31:24] = buffer_data_3[3391:3384];
        layer3[39][39:32] = buffer_data_3[3399:3392];
        layer3[39][47:40] = buffer_data_3[3407:3400];
        layer3[39][55:48] = buffer_data_3[3415:3408];
        layer4[39][7:0] = buffer_data_2[3367:3360];
        layer4[39][15:8] = buffer_data_2[3375:3368];
        layer4[39][23:16] = buffer_data_2[3383:3376];
        layer4[39][31:24] = buffer_data_2[3391:3384];
        layer4[39][39:32] = buffer_data_2[3399:3392];
        layer4[39][47:40] = buffer_data_2[3407:3400];
        layer4[39][55:48] = buffer_data_2[3415:3408];
        layer5[39][7:0] = buffer_data_1[3367:3360];
        layer5[39][15:8] = buffer_data_1[3375:3368];
        layer5[39][23:16] = buffer_data_1[3383:3376];
        layer5[39][31:24] = buffer_data_1[3391:3384];
        layer5[39][39:32] = buffer_data_1[3399:3392];
        layer5[39][47:40] = buffer_data_1[3407:3400];
        layer5[39][55:48] = buffer_data_1[3415:3408];
        layer6[39][7:0] = buffer_data_0[3367:3360];
        layer6[39][15:8] = buffer_data_0[3375:3368];
        layer6[39][23:16] = buffer_data_0[3383:3376];
        layer6[39][31:24] = buffer_data_0[3391:3384];
        layer6[39][39:32] = buffer_data_0[3399:3392];
        layer6[39][47:40] = buffer_data_0[3407:3400];
        layer6[39][55:48] = buffer_data_0[3415:3408];
        layer0[40][7:0] = buffer_data_6[3375:3368];
        layer0[40][15:8] = buffer_data_6[3383:3376];
        layer0[40][23:16] = buffer_data_6[3391:3384];
        layer0[40][31:24] = buffer_data_6[3399:3392];
        layer0[40][39:32] = buffer_data_6[3407:3400];
        layer0[40][47:40] = buffer_data_6[3415:3408];
        layer0[40][55:48] = buffer_data_6[3423:3416];
        layer1[40][7:0] = buffer_data_5[3375:3368];
        layer1[40][15:8] = buffer_data_5[3383:3376];
        layer1[40][23:16] = buffer_data_5[3391:3384];
        layer1[40][31:24] = buffer_data_5[3399:3392];
        layer1[40][39:32] = buffer_data_5[3407:3400];
        layer1[40][47:40] = buffer_data_5[3415:3408];
        layer1[40][55:48] = buffer_data_5[3423:3416];
        layer2[40][7:0] = buffer_data_4[3375:3368];
        layer2[40][15:8] = buffer_data_4[3383:3376];
        layer2[40][23:16] = buffer_data_4[3391:3384];
        layer2[40][31:24] = buffer_data_4[3399:3392];
        layer2[40][39:32] = buffer_data_4[3407:3400];
        layer2[40][47:40] = buffer_data_4[3415:3408];
        layer2[40][55:48] = buffer_data_4[3423:3416];
        layer3[40][7:0] = buffer_data_3[3375:3368];
        layer3[40][15:8] = buffer_data_3[3383:3376];
        layer3[40][23:16] = buffer_data_3[3391:3384];
        layer3[40][31:24] = buffer_data_3[3399:3392];
        layer3[40][39:32] = buffer_data_3[3407:3400];
        layer3[40][47:40] = buffer_data_3[3415:3408];
        layer3[40][55:48] = buffer_data_3[3423:3416];
        layer4[40][7:0] = buffer_data_2[3375:3368];
        layer4[40][15:8] = buffer_data_2[3383:3376];
        layer4[40][23:16] = buffer_data_2[3391:3384];
        layer4[40][31:24] = buffer_data_2[3399:3392];
        layer4[40][39:32] = buffer_data_2[3407:3400];
        layer4[40][47:40] = buffer_data_2[3415:3408];
        layer4[40][55:48] = buffer_data_2[3423:3416];
        layer5[40][7:0] = buffer_data_1[3375:3368];
        layer5[40][15:8] = buffer_data_1[3383:3376];
        layer5[40][23:16] = buffer_data_1[3391:3384];
        layer5[40][31:24] = buffer_data_1[3399:3392];
        layer5[40][39:32] = buffer_data_1[3407:3400];
        layer5[40][47:40] = buffer_data_1[3415:3408];
        layer5[40][55:48] = buffer_data_1[3423:3416];
        layer6[40][7:0] = buffer_data_0[3375:3368];
        layer6[40][15:8] = buffer_data_0[3383:3376];
        layer6[40][23:16] = buffer_data_0[3391:3384];
        layer6[40][31:24] = buffer_data_0[3399:3392];
        layer6[40][39:32] = buffer_data_0[3407:3400];
        layer6[40][47:40] = buffer_data_0[3415:3408];
        layer6[40][55:48] = buffer_data_0[3423:3416];
        layer0[41][7:0] = buffer_data_6[3383:3376];
        layer0[41][15:8] = buffer_data_6[3391:3384];
        layer0[41][23:16] = buffer_data_6[3399:3392];
        layer0[41][31:24] = buffer_data_6[3407:3400];
        layer0[41][39:32] = buffer_data_6[3415:3408];
        layer0[41][47:40] = buffer_data_6[3423:3416];
        layer0[41][55:48] = buffer_data_6[3431:3424];
        layer1[41][7:0] = buffer_data_5[3383:3376];
        layer1[41][15:8] = buffer_data_5[3391:3384];
        layer1[41][23:16] = buffer_data_5[3399:3392];
        layer1[41][31:24] = buffer_data_5[3407:3400];
        layer1[41][39:32] = buffer_data_5[3415:3408];
        layer1[41][47:40] = buffer_data_5[3423:3416];
        layer1[41][55:48] = buffer_data_5[3431:3424];
        layer2[41][7:0] = buffer_data_4[3383:3376];
        layer2[41][15:8] = buffer_data_4[3391:3384];
        layer2[41][23:16] = buffer_data_4[3399:3392];
        layer2[41][31:24] = buffer_data_4[3407:3400];
        layer2[41][39:32] = buffer_data_4[3415:3408];
        layer2[41][47:40] = buffer_data_4[3423:3416];
        layer2[41][55:48] = buffer_data_4[3431:3424];
        layer3[41][7:0] = buffer_data_3[3383:3376];
        layer3[41][15:8] = buffer_data_3[3391:3384];
        layer3[41][23:16] = buffer_data_3[3399:3392];
        layer3[41][31:24] = buffer_data_3[3407:3400];
        layer3[41][39:32] = buffer_data_3[3415:3408];
        layer3[41][47:40] = buffer_data_3[3423:3416];
        layer3[41][55:48] = buffer_data_3[3431:3424];
        layer4[41][7:0] = buffer_data_2[3383:3376];
        layer4[41][15:8] = buffer_data_2[3391:3384];
        layer4[41][23:16] = buffer_data_2[3399:3392];
        layer4[41][31:24] = buffer_data_2[3407:3400];
        layer4[41][39:32] = buffer_data_2[3415:3408];
        layer4[41][47:40] = buffer_data_2[3423:3416];
        layer4[41][55:48] = buffer_data_2[3431:3424];
        layer5[41][7:0] = buffer_data_1[3383:3376];
        layer5[41][15:8] = buffer_data_1[3391:3384];
        layer5[41][23:16] = buffer_data_1[3399:3392];
        layer5[41][31:24] = buffer_data_1[3407:3400];
        layer5[41][39:32] = buffer_data_1[3415:3408];
        layer5[41][47:40] = buffer_data_1[3423:3416];
        layer5[41][55:48] = buffer_data_1[3431:3424];
        layer6[41][7:0] = buffer_data_0[3383:3376];
        layer6[41][15:8] = buffer_data_0[3391:3384];
        layer6[41][23:16] = buffer_data_0[3399:3392];
        layer6[41][31:24] = buffer_data_0[3407:3400];
        layer6[41][39:32] = buffer_data_0[3415:3408];
        layer6[41][47:40] = buffer_data_0[3423:3416];
        layer6[41][55:48] = buffer_data_0[3431:3424];
        layer0[42][7:0] = buffer_data_6[3391:3384];
        layer0[42][15:8] = buffer_data_6[3399:3392];
        layer0[42][23:16] = buffer_data_6[3407:3400];
        layer0[42][31:24] = buffer_data_6[3415:3408];
        layer0[42][39:32] = buffer_data_6[3423:3416];
        layer0[42][47:40] = buffer_data_6[3431:3424];
        layer0[42][55:48] = buffer_data_6[3439:3432];
        layer1[42][7:0] = buffer_data_5[3391:3384];
        layer1[42][15:8] = buffer_data_5[3399:3392];
        layer1[42][23:16] = buffer_data_5[3407:3400];
        layer1[42][31:24] = buffer_data_5[3415:3408];
        layer1[42][39:32] = buffer_data_5[3423:3416];
        layer1[42][47:40] = buffer_data_5[3431:3424];
        layer1[42][55:48] = buffer_data_5[3439:3432];
        layer2[42][7:0] = buffer_data_4[3391:3384];
        layer2[42][15:8] = buffer_data_4[3399:3392];
        layer2[42][23:16] = buffer_data_4[3407:3400];
        layer2[42][31:24] = buffer_data_4[3415:3408];
        layer2[42][39:32] = buffer_data_4[3423:3416];
        layer2[42][47:40] = buffer_data_4[3431:3424];
        layer2[42][55:48] = buffer_data_4[3439:3432];
        layer3[42][7:0] = buffer_data_3[3391:3384];
        layer3[42][15:8] = buffer_data_3[3399:3392];
        layer3[42][23:16] = buffer_data_3[3407:3400];
        layer3[42][31:24] = buffer_data_3[3415:3408];
        layer3[42][39:32] = buffer_data_3[3423:3416];
        layer3[42][47:40] = buffer_data_3[3431:3424];
        layer3[42][55:48] = buffer_data_3[3439:3432];
        layer4[42][7:0] = buffer_data_2[3391:3384];
        layer4[42][15:8] = buffer_data_2[3399:3392];
        layer4[42][23:16] = buffer_data_2[3407:3400];
        layer4[42][31:24] = buffer_data_2[3415:3408];
        layer4[42][39:32] = buffer_data_2[3423:3416];
        layer4[42][47:40] = buffer_data_2[3431:3424];
        layer4[42][55:48] = buffer_data_2[3439:3432];
        layer5[42][7:0] = buffer_data_1[3391:3384];
        layer5[42][15:8] = buffer_data_1[3399:3392];
        layer5[42][23:16] = buffer_data_1[3407:3400];
        layer5[42][31:24] = buffer_data_1[3415:3408];
        layer5[42][39:32] = buffer_data_1[3423:3416];
        layer5[42][47:40] = buffer_data_1[3431:3424];
        layer5[42][55:48] = buffer_data_1[3439:3432];
        layer6[42][7:0] = buffer_data_0[3391:3384];
        layer6[42][15:8] = buffer_data_0[3399:3392];
        layer6[42][23:16] = buffer_data_0[3407:3400];
        layer6[42][31:24] = buffer_data_0[3415:3408];
        layer6[42][39:32] = buffer_data_0[3423:3416];
        layer6[42][47:40] = buffer_data_0[3431:3424];
        layer6[42][55:48] = buffer_data_0[3439:3432];
        layer0[43][7:0] = buffer_data_6[3399:3392];
        layer0[43][15:8] = buffer_data_6[3407:3400];
        layer0[43][23:16] = buffer_data_6[3415:3408];
        layer0[43][31:24] = buffer_data_6[3423:3416];
        layer0[43][39:32] = buffer_data_6[3431:3424];
        layer0[43][47:40] = buffer_data_6[3439:3432];
        layer0[43][55:48] = buffer_data_6[3447:3440];
        layer1[43][7:0] = buffer_data_5[3399:3392];
        layer1[43][15:8] = buffer_data_5[3407:3400];
        layer1[43][23:16] = buffer_data_5[3415:3408];
        layer1[43][31:24] = buffer_data_5[3423:3416];
        layer1[43][39:32] = buffer_data_5[3431:3424];
        layer1[43][47:40] = buffer_data_5[3439:3432];
        layer1[43][55:48] = buffer_data_5[3447:3440];
        layer2[43][7:0] = buffer_data_4[3399:3392];
        layer2[43][15:8] = buffer_data_4[3407:3400];
        layer2[43][23:16] = buffer_data_4[3415:3408];
        layer2[43][31:24] = buffer_data_4[3423:3416];
        layer2[43][39:32] = buffer_data_4[3431:3424];
        layer2[43][47:40] = buffer_data_4[3439:3432];
        layer2[43][55:48] = buffer_data_4[3447:3440];
        layer3[43][7:0] = buffer_data_3[3399:3392];
        layer3[43][15:8] = buffer_data_3[3407:3400];
        layer3[43][23:16] = buffer_data_3[3415:3408];
        layer3[43][31:24] = buffer_data_3[3423:3416];
        layer3[43][39:32] = buffer_data_3[3431:3424];
        layer3[43][47:40] = buffer_data_3[3439:3432];
        layer3[43][55:48] = buffer_data_3[3447:3440];
        layer4[43][7:0] = buffer_data_2[3399:3392];
        layer4[43][15:8] = buffer_data_2[3407:3400];
        layer4[43][23:16] = buffer_data_2[3415:3408];
        layer4[43][31:24] = buffer_data_2[3423:3416];
        layer4[43][39:32] = buffer_data_2[3431:3424];
        layer4[43][47:40] = buffer_data_2[3439:3432];
        layer4[43][55:48] = buffer_data_2[3447:3440];
        layer5[43][7:0] = buffer_data_1[3399:3392];
        layer5[43][15:8] = buffer_data_1[3407:3400];
        layer5[43][23:16] = buffer_data_1[3415:3408];
        layer5[43][31:24] = buffer_data_1[3423:3416];
        layer5[43][39:32] = buffer_data_1[3431:3424];
        layer5[43][47:40] = buffer_data_1[3439:3432];
        layer5[43][55:48] = buffer_data_1[3447:3440];
        layer6[43][7:0] = buffer_data_0[3399:3392];
        layer6[43][15:8] = buffer_data_0[3407:3400];
        layer6[43][23:16] = buffer_data_0[3415:3408];
        layer6[43][31:24] = buffer_data_0[3423:3416];
        layer6[43][39:32] = buffer_data_0[3431:3424];
        layer6[43][47:40] = buffer_data_0[3439:3432];
        layer6[43][55:48] = buffer_data_0[3447:3440];
        layer0[44][7:0] = buffer_data_6[3407:3400];
        layer0[44][15:8] = buffer_data_6[3415:3408];
        layer0[44][23:16] = buffer_data_6[3423:3416];
        layer0[44][31:24] = buffer_data_6[3431:3424];
        layer0[44][39:32] = buffer_data_6[3439:3432];
        layer0[44][47:40] = buffer_data_6[3447:3440];
        layer0[44][55:48] = buffer_data_6[3455:3448];
        layer1[44][7:0] = buffer_data_5[3407:3400];
        layer1[44][15:8] = buffer_data_5[3415:3408];
        layer1[44][23:16] = buffer_data_5[3423:3416];
        layer1[44][31:24] = buffer_data_5[3431:3424];
        layer1[44][39:32] = buffer_data_5[3439:3432];
        layer1[44][47:40] = buffer_data_5[3447:3440];
        layer1[44][55:48] = buffer_data_5[3455:3448];
        layer2[44][7:0] = buffer_data_4[3407:3400];
        layer2[44][15:8] = buffer_data_4[3415:3408];
        layer2[44][23:16] = buffer_data_4[3423:3416];
        layer2[44][31:24] = buffer_data_4[3431:3424];
        layer2[44][39:32] = buffer_data_4[3439:3432];
        layer2[44][47:40] = buffer_data_4[3447:3440];
        layer2[44][55:48] = buffer_data_4[3455:3448];
        layer3[44][7:0] = buffer_data_3[3407:3400];
        layer3[44][15:8] = buffer_data_3[3415:3408];
        layer3[44][23:16] = buffer_data_3[3423:3416];
        layer3[44][31:24] = buffer_data_3[3431:3424];
        layer3[44][39:32] = buffer_data_3[3439:3432];
        layer3[44][47:40] = buffer_data_3[3447:3440];
        layer3[44][55:48] = buffer_data_3[3455:3448];
        layer4[44][7:0] = buffer_data_2[3407:3400];
        layer4[44][15:8] = buffer_data_2[3415:3408];
        layer4[44][23:16] = buffer_data_2[3423:3416];
        layer4[44][31:24] = buffer_data_2[3431:3424];
        layer4[44][39:32] = buffer_data_2[3439:3432];
        layer4[44][47:40] = buffer_data_2[3447:3440];
        layer4[44][55:48] = buffer_data_2[3455:3448];
        layer5[44][7:0] = buffer_data_1[3407:3400];
        layer5[44][15:8] = buffer_data_1[3415:3408];
        layer5[44][23:16] = buffer_data_1[3423:3416];
        layer5[44][31:24] = buffer_data_1[3431:3424];
        layer5[44][39:32] = buffer_data_1[3439:3432];
        layer5[44][47:40] = buffer_data_1[3447:3440];
        layer5[44][55:48] = buffer_data_1[3455:3448];
        layer6[44][7:0] = buffer_data_0[3407:3400];
        layer6[44][15:8] = buffer_data_0[3415:3408];
        layer6[44][23:16] = buffer_data_0[3423:3416];
        layer6[44][31:24] = buffer_data_0[3431:3424];
        layer6[44][39:32] = buffer_data_0[3439:3432];
        layer6[44][47:40] = buffer_data_0[3447:3440];
        layer6[44][55:48] = buffer_data_0[3455:3448];
        layer0[45][7:0] = buffer_data_6[3415:3408];
        layer0[45][15:8] = buffer_data_6[3423:3416];
        layer0[45][23:16] = buffer_data_6[3431:3424];
        layer0[45][31:24] = buffer_data_6[3439:3432];
        layer0[45][39:32] = buffer_data_6[3447:3440];
        layer0[45][47:40] = buffer_data_6[3455:3448];
        layer0[45][55:48] = buffer_data_6[3463:3456];
        layer1[45][7:0] = buffer_data_5[3415:3408];
        layer1[45][15:8] = buffer_data_5[3423:3416];
        layer1[45][23:16] = buffer_data_5[3431:3424];
        layer1[45][31:24] = buffer_data_5[3439:3432];
        layer1[45][39:32] = buffer_data_5[3447:3440];
        layer1[45][47:40] = buffer_data_5[3455:3448];
        layer1[45][55:48] = buffer_data_5[3463:3456];
        layer2[45][7:0] = buffer_data_4[3415:3408];
        layer2[45][15:8] = buffer_data_4[3423:3416];
        layer2[45][23:16] = buffer_data_4[3431:3424];
        layer2[45][31:24] = buffer_data_4[3439:3432];
        layer2[45][39:32] = buffer_data_4[3447:3440];
        layer2[45][47:40] = buffer_data_4[3455:3448];
        layer2[45][55:48] = buffer_data_4[3463:3456];
        layer3[45][7:0] = buffer_data_3[3415:3408];
        layer3[45][15:8] = buffer_data_3[3423:3416];
        layer3[45][23:16] = buffer_data_3[3431:3424];
        layer3[45][31:24] = buffer_data_3[3439:3432];
        layer3[45][39:32] = buffer_data_3[3447:3440];
        layer3[45][47:40] = buffer_data_3[3455:3448];
        layer3[45][55:48] = buffer_data_3[3463:3456];
        layer4[45][7:0] = buffer_data_2[3415:3408];
        layer4[45][15:8] = buffer_data_2[3423:3416];
        layer4[45][23:16] = buffer_data_2[3431:3424];
        layer4[45][31:24] = buffer_data_2[3439:3432];
        layer4[45][39:32] = buffer_data_2[3447:3440];
        layer4[45][47:40] = buffer_data_2[3455:3448];
        layer4[45][55:48] = buffer_data_2[3463:3456];
        layer5[45][7:0] = buffer_data_1[3415:3408];
        layer5[45][15:8] = buffer_data_1[3423:3416];
        layer5[45][23:16] = buffer_data_1[3431:3424];
        layer5[45][31:24] = buffer_data_1[3439:3432];
        layer5[45][39:32] = buffer_data_1[3447:3440];
        layer5[45][47:40] = buffer_data_1[3455:3448];
        layer5[45][55:48] = buffer_data_1[3463:3456];
        layer6[45][7:0] = buffer_data_0[3415:3408];
        layer6[45][15:8] = buffer_data_0[3423:3416];
        layer6[45][23:16] = buffer_data_0[3431:3424];
        layer6[45][31:24] = buffer_data_0[3439:3432];
        layer6[45][39:32] = buffer_data_0[3447:3440];
        layer6[45][47:40] = buffer_data_0[3455:3448];
        layer6[45][55:48] = buffer_data_0[3463:3456];
        layer0[46][7:0] = buffer_data_6[3423:3416];
        layer0[46][15:8] = buffer_data_6[3431:3424];
        layer0[46][23:16] = buffer_data_6[3439:3432];
        layer0[46][31:24] = buffer_data_6[3447:3440];
        layer0[46][39:32] = buffer_data_6[3455:3448];
        layer0[46][47:40] = buffer_data_6[3463:3456];
        layer0[46][55:48] = buffer_data_6[3471:3464];
        layer1[46][7:0] = buffer_data_5[3423:3416];
        layer1[46][15:8] = buffer_data_5[3431:3424];
        layer1[46][23:16] = buffer_data_5[3439:3432];
        layer1[46][31:24] = buffer_data_5[3447:3440];
        layer1[46][39:32] = buffer_data_5[3455:3448];
        layer1[46][47:40] = buffer_data_5[3463:3456];
        layer1[46][55:48] = buffer_data_5[3471:3464];
        layer2[46][7:0] = buffer_data_4[3423:3416];
        layer2[46][15:8] = buffer_data_4[3431:3424];
        layer2[46][23:16] = buffer_data_4[3439:3432];
        layer2[46][31:24] = buffer_data_4[3447:3440];
        layer2[46][39:32] = buffer_data_4[3455:3448];
        layer2[46][47:40] = buffer_data_4[3463:3456];
        layer2[46][55:48] = buffer_data_4[3471:3464];
        layer3[46][7:0] = buffer_data_3[3423:3416];
        layer3[46][15:8] = buffer_data_3[3431:3424];
        layer3[46][23:16] = buffer_data_3[3439:3432];
        layer3[46][31:24] = buffer_data_3[3447:3440];
        layer3[46][39:32] = buffer_data_3[3455:3448];
        layer3[46][47:40] = buffer_data_3[3463:3456];
        layer3[46][55:48] = buffer_data_3[3471:3464];
        layer4[46][7:0] = buffer_data_2[3423:3416];
        layer4[46][15:8] = buffer_data_2[3431:3424];
        layer4[46][23:16] = buffer_data_2[3439:3432];
        layer4[46][31:24] = buffer_data_2[3447:3440];
        layer4[46][39:32] = buffer_data_2[3455:3448];
        layer4[46][47:40] = buffer_data_2[3463:3456];
        layer4[46][55:48] = buffer_data_2[3471:3464];
        layer5[46][7:0] = buffer_data_1[3423:3416];
        layer5[46][15:8] = buffer_data_1[3431:3424];
        layer5[46][23:16] = buffer_data_1[3439:3432];
        layer5[46][31:24] = buffer_data_1[3447:3440];
        layer5[46][39:32] = buffer_data_1[3455:3448];
        layer5[46][47:40] = buffer_data_1[3463:3456];
        layer5[46][55:48] = buffer_data_1[3471:3464];
        layer6[46][7:0] = buffer_data_0[3423:3416];
        layer6[46][15:8] = buffer_data_0[3431:3424];
        layer6[46][23:16] = buffer_data_0[3439:3432];
        layer6[46][31:24] = buffer_data_0[3447:3440];
        layer6[46][39:32] = buffer_data_0[3455:3448];
        layer6[46][47:40] = buffer_data_0[3463:3456];
        layer6[46][55:48] = buffer_data_0[3471:3464];
        layer0[47][7:0] = buffer_data_6[3431:3424];
        layer0[47][15:8] = buffer_data_6[3439:3432];
        layer0[47][23:16] = buffer_data_6[3447:3440];
        layer0[47][31:24] = buffer_data_6[3455:3448];
        layer0[47][39:32] = buffer_data_6[3463:3456];
        layer0[47][47:40] = buffer_data_6[3471:3464];
        layer0[47][55:48] = buffer_data_6[3479:3472];
        layer1[47][7:0] = buffer_data_5[3431:3424];
        layer1[47][15:8] = buffer_data_5[3439:3432];
        layer1[47][23:16] = buffer_data_5[3447:3440];
        layer1[47][31:24] = buffer_data_5[3455:3448];
        layer1[47][39:32] = buffer_data_5[3463:3456];
        layer1[47][47:40] = buffer_data_5[3471:3464];
        layer1[47][55:48] = buffer_data_5[3479:3472];
        layer2[47][7:0] = buffer_data_4[3431:3424];
        layer2[47][15:8] = buffer_data_4[3439:3432];
        layer2[47][23:16] = buffer_data_4[3447:3440];
        layer2[47][31:24] = buffer_data_4[3455:3448];
        layer2[47][39:32] = buffer_data_4[3463:3456];
        layer2[47][47:40] = buffer_data_4[3471:3464];
        layer2[47][55:48] = buffer_data_4[3479:3472];
        layer3[47][7:0] = buffer_data_3[3431:3424];
        layer3[47][15:8] = buffer_data_3[3439:3432];
        layer3[47][23:16] = buffer_data_3[3447:3440];
        layer3[47][31:24] = buffer_data_3[3455:3448];
        layer3[47][39:32] = buffer_data_3[3463:3456];
        layer3[47][47:40] = buffer_data_3[3471:3464];
        layer3[47][55:48] = buffer_data_3[3479:3472];
        layer4[47][7:0] = buffer_data_2[3431:3424];
        layer4[47][15:8] = buffer_data_2[3439:3432];
        layer4[47][23:16] = buffer_data_2[3447:3440];
        layer4[47][31:24] = buffer_data_2[3455:3448];
        layer4[47][39:32] = buffer_data_2[3463:3456];
        layer4[47][47:40] = buffer_data_2[3471:3464];
        layer4[47][55:48] = buffer_data_2[3479:3472];
        layer5[47][7:0] = buffer_data_1[3431:3424];
        layer5[47][15:8] = buffer_data_1[3439:3432];
        layer5[47][23:16] = buffer_data_1[3447:3440];
        layer5[47][31:24] = buffer_data_1[3455:3448];
        layer5[47][39:32] = buffer_data_1[3463:3456];
        layer5[47][47:40] = buffer_data_1[3471:3464];
        layer5[47][55:48] = buffer_data_1[3479:3472];
        layer6[47][7:0] = buffer_data_0[3431:3424];
        layer6[47][15:8] = buffer_data_0[3439:3432];
        layer6[47][23:16] = buffer_data_0[3447:3440];
        layer6[47][31:24] = buffer_data_0[3455:3448];
        layer6[47][39:32] = buffer_data_0[3463:3456];
        layer6[47][47:40] = buffer_data_0[3471:3464];
        layer6[47][55:48] = buffer_data_0[3479:3472];
        layer0[48][7:0] = buffer_data_6[3439:3432];
        layer0[48][15:8] = buffer_data_6[3447:3440];
        layer0[48][23:16] = buffer_data_6[3455:3448];
        layer0[48][31:24] = buffer_data_6[3463:3456];
        layer0[48][39:32] = buffer_data_6[3471:3464];
        layer0[48][47:40] = buffer_data_6[3479:3472];
        layer0[48][55:48] = buffer_data_6[3487:3480];
        layer1[48][7:0] = buffer_data_5[3439:3432];
        layer1[48][15:8] = buffer_data_5[3447:3440];
        layer1[48][23:16] = buffer_data_5[3455:3448];
        layer1[48][31:24] = buffer_data_5[3463:3456];
        layer1[48][39:32] = buffer_data_5[3471:3464];
        layer1[48][47:40] = buffer_data_5[3479:3472];
        layer1[48][55:48] = buffer_data_5[3487:3480];
        layer2[48][7:0] = buffer_data_4[3439:3432];
        layer2[48][15:8] = buffer_data_4[3447:3440];
        layer2[48][23:16] = buffer_data_4[3455:3448];
        layer2[48][31:24] = buffer_data_4[3463:3456];
        layer2[48][39:32] = buffer_data_4[3471:3464];
        layer2[48][47:40] = buffer_data_4[3479:3472];
        layer2[48][55:48] = buffer_data_4[3487:3480];
        layer3[48][7:0] = buffer_data_3[3439:3432];
        layer3[48][15:8] = buffer_data_3[3447:3440];
        layer3[48][23:16] = buffer_data_3[3455:3448];
        layer3[48][31:24] = buffer_data_3[3463:3456];
        layer3[48][39:32] = buffer_data_3[3471:3464];
        layer3[48][47:40] = buffer_data_3[3479:3472];
        layer3[48][55:48] = buffer_data_3[3487:3480];
        layer4[48][7:0] = buffer_data_2[3439:3432];
        layer4[48][15:8] = buffer_data_2[3447:3440];
        layer4[48][23:16] = buffer_data_2[3455:3448];
        layer4[48][31:24] = buffer_data_2[3463:3456];
        layer4[48][39:32] = buffer_data_2[3471:3464];
        layer4[48][47:40] = buffer_data_2[3479:3472];
        layer4[48][55:48] = buffer_data_2[3487:3480];
        layer5[48][7:0] = buffer_data_1[3439:3432];
        layer5[48][15:8] = buffer_data_1[3447:3440];
        layer5[48][23:16] = buffer_data_1[3455:3448];
        layer5[48][31:24] = buffer_data_1[3463:3456];
        layer5[48][39:32] = buffer_data_1[3471:3464];
        layer5[48][47:40] = buffer_data_1[3479:3472];
        layer5[48][55:48] = buffer_data_1[3487:3480];
        layer6[48][7:0] = buffer_data_0[3439:3432];
        layer6[48][15:8] = buffer_data_0[3447:3440];
        layer6[48][23:16] = buffer_data_0[3455:3448];
        layer6[48][31:24] = buffer_data_0[3463:3456];
        layer6[48][39:32] = buffer_data_0[3471:3464];
        layer6[48][47:40] = buffer_data_0[3479:3472];
        layer6[48][55:48] = buffer_data_0[3487:3480];
        layer0[49][7:0] = buffer_data_6[3447:3440];
        layer0[49][15:8] = buffer_data_6[3455:3448];
        layer0[49][23:16] = buffer_data_6[3463:3456];
        layer0[49][31:24] = buffer_data_6[3471:3464];
        layer0[49][39:32] = buffer_data_6[3479:3472];
        layer0[49][47:40] = buffer_data_6[3487:3480];
        layer0[49][55:48] = buffer_data_6[3495:3488];
        layer1[49][7:0] = buffer_data_5[3447:3440];
        layer1[49][15:8] = buffer_data_5[3455:3448];
        layer1[49][23:16] = buffer_data_5[3463:3456];
        layer1[49][31:24] = buffer_data_5[3471:3464];
        layer1[49][39:32] = buffer_data_5[3479:3472];
        layer1[49][47:40] = buffer_data_5[3487:3480];
        layer1[49][55:48] = buffer_data_5[3495:3488];
        layer2[49][7:0] = buffer_data_4[3447:3440];
        layer2[49][15:8] = buffer_data_4[3455:3448];
        layer2[49][23:16] = buffer_data_4[3463:3456];
        layer2[49][31:24] = buffer_data_4[3471:3464];
        layer2[49][39:32] = buffer_data_4[3479:3472];
        layer2[49][47:40] = buffer_data_4[3487:3480];
        layer2[49][55:48] = buffer_data_4[3495:3488];
        layer3[49][7:0] = buffer_data_3[3447:3440];
        layer3[49][15:8] = buffer_data_3[3455:3448];
        layer3[49][23:16] = buffer_data_3[3463:3456];
        layer3[49][31:24] = buffer_data_3[3471:3464];
        layer3[49][39:32] = buffer_data_3[3479:3472];
        layer3[49][47:40] = buffer_data_3[3487:3480];
        layer3[49][55:48] = buffer_data_3[3495:3488];
        layer4[49][7:0] = buffer_data_2[3447:3440];
        layer4[49][15:8] = buffer_data_2[3455:3448];
        layer4[49][23:16] = buffer_data_2[3463:3456];
        layer4[49][31:24] = buffer_data_2[3471:3464];
        layer4[49][39:32] = buffer_data_2[3479:3472];
        layer4[49][47:40] = buffer_data_2[3487:3480];
        layer4[49][55:48] = buffer_data_2[3495:3488];
        layer5[49][7:0] = buffer_data_1[3447:3440];
        layer5[49][15:8] = buffer_data_1[3455:3448];
        layer5[49][23:16] = buffer_data_1[3463:3456];
        layer5[49][31:24] = buffer_data_1[3471:3464];
        layer5[49][39:32] = buffer_data_1[3479:3472];
        layer5[49][47:40] = buffer_data_1[3487:3480];
        layer5[49][55:48] = buffer_data_1[3495:3488];
        layer6[49][7:0] = buffer_data_0[3447:3440];
        layer6[49][15:8] = buffer_data_0[3455:3448];
        layer6[49][23:16] = buffer_data_0[3463:3456];
        layer6[49][31:24] = buffer_data_0[3471:3464];
        layer6[49][39:32] = buffer_data_0[3479:3472];
        layer6[49][47:40] = buffer_data_0[3487:3480];
        layer6[49][55:48] = buffer_data_0[3495:3488];
        layer0[50][7:0] = buffer_data_6[3455:3448];
        layer0[50][15:8] = buffer_data_6[3463:3456];
        layer0[50][23:16] = buffer_data_6[3471:3464];
        layer0[50][31:24] = buffer_data_6[3479:3472];
        layer0[50][39:32] = buffer_data_6[3487:3480];
        layer0[50][47:40] = buffer_data_6[3495:3488];
        layer0[50][55:48] = buffer_data_6[3503:3496];
        layer1[50][7:0] = buffer_data_5[3455:3448];
        layer1[50][15:8] = buffer_data_5[3463:3456];
        layer1[50][23:16] = buffer_data_5[3471:3464];
        layer1[50][31:24] = buffer_data_5[3479:3472];
        layer1[50][39:32] = buffer_data_5[3487:3480];
        layer1[50][47:40] = buffer_data_5[3495:3488];
        layer1[50][55:48] = buffer_data_5[3503:3496];
        layer2[50][7:0] = buffer_data_4[3455:3448];
        layer2[50][15:8] = buffer_data_4[3463:3456];
        layer2[50][23:16] = buffer_data_4[3471:3464];
        layer2[50][31:24] = buffer_data_4[3479:3472];
        layer2[50][39:32] = buffer_data_4[3487:3480];
        layer2[50][47:40] = buffer_data_4[3495:3488];
        layer2[50][55:48] = buffer_data_4[3503:3496];
        layer3[50][7:0] = buffer_data_3[3455:3448];
        layer3[50][15:8] = buffer_data_3[3463:3456];
        layer3[50][23:16] = buffer_data_3[3471:3464];
        layer3[50][31:24] = buffer_data_3[3479:3472];
        layer3[50][39:32] = buffer_data_3[3487:3480];
        layer3[50][47:40] = buffer_data_3[3495:3488];
        layer3[50][55:48] = buffer_data_3[3503:3496];
        layer4[50][7:0] = buffer_data_2[3455:3448];
        layer4[50][15:8] = buffer_data_2[3463:3456];
        layer4[50][23:16] = buffer_data_2[3471:3464];
        layer4[50][31:24] = buffer_data_2[3479:3472];
        layer4[50][39:32] = buffer_data_2[3487:3480];
        layer4[50][47:40] = buffer_data_2[3495:3488];
        layer4[50][55:48] = buffer_data_2[3503:3496];
        layer5[50][7:0] = buffer_data_1[3455:3448];
        layer5[50][15:8] = buffer_data_1[3463:3456];
        layer5[50][23:16] = buffer_data_1[3471:3464];
        layer5[50][31:24] = buffer_data_1[3479:3472];
        layer5[50][39:32] = buffer_data_1[3487:3480];
        layer5[50][47:40] = buffer_data_1[3495:3488];
        layer5[50][55:48] = buffer_data_1[3503:3496];
        layer6[50][7:0] = buffer_data_0[3455:3448];
        layer6[50][15:8] = buffer_data_0[3463:3456];
        layer6[50][23:16] = buffer_data_0[3471:3464];
        layer6[50][31:24] = buffer_data_0[3479:3472];
        layer6[50][39:32] = buffer_data_0[3487:3480];
        layer6[50][47:40] = buffer_data_0[3495:3488];
        layer6[50][55:48] = buffer_data_0[3503:3496];
        layer0[51][7:0] = buffer_data_6[3463:3456];
        layer0[51][15:8] = buffer_data_6[3471:3464];
        layer0[51][23:16] = buffer_data_6[3479:3472];
        layer0[51][31:24] = buffer_data_6[3487:3480];
        layer0[51][39:32] = buffer_data_6[3495:3488];
        layer0[51][47:40] = buffer_data_6[3503:3496];
        layer0[51][55:48] = buffer_data_6[3511:3504];
        layer1[51][7:0] = buffer_data_5[3463:3456];
        layer1[51][15:8] = buffer_data_5[3471:3464];
        layer1[51][23:16] = buffer_data_5[3479:3472];
        layer1[51][31:24] = buffer_data_5[3487:3480];
        layer1[51][39:32] = buffer_data_5[3495:3488];
        layer1[51][47:40] = buffer_data_5[3503:3496];
        layer1[51][55:48] = buffer_data_5[3511:3504];
        layer2[51][7:0] = buffer_data_4[3463:3456];
        layer2[51][15:8] = buffer_data_4[3471:3464];
        layer2[51][23:16] = buffer_data_4[3479:3472];
        layer2[51][31:24] = buffer_data_4[3487:3480];
        layer2[51][39:32] = buffer_data_4[3495:3488];
        layer2[51][47:40] = buffer_data_4[3503:3496];
        layer2[51][55:48] = buffer_data_4[3511:3504];
        layer3[51][7:0] = buffer_data_3[3463:3456];
        layer3[51][15:8] = buffer_data_3[3471:3464];
        layer3[51][23:16] = buffer_data_3[3479:3472];
        layer3[51][31:24] = buffer_data_3[3487:3480];
        layer3[51][39:32] = buffer_data_3[3495:3488];
        layer3[51][47:40] = buffer_data_3[3503:3496];
        layer3[51][55:48] = buffer_data_3[3511:3504];
        layer4[51][7:0] = buffer_data_2[3463:3456];
        layer4[51][15:8] = buffer_data_2[3471:3464];
        layer4[51][23:16] = buffer_data_2[3479:3472];
        layer4[51][31:24] = buffer_data_2[3487:3480];
        layer4[51][39:32] = buffer_data_2[3495:3488];
        layer4[51][47:40] = buffer_data_2[3503:3496];
        layer4[51][55:48] = buffer_data_2[3511:3504];
        layer5[51][7:0] = buffer_data_1[3463:3456];
        layer5[51][15:8] = buffer_data_1[3471:3464];
        layer5[51][23:16] = buffer_data_1[3479:3472];
        layer5[51][31:24] = buffer_data_1[3487:3480];
        layer5[51][39:32] = buffer_data_1[3495:3488];
        layer5[51][47:40] = buffer_data_1[3503:3496];
        layer5[51][55:48] = buffer_data_1[3511:3504];
        layer6[51][7:0] = buffer_data_0[3463:3456];
        layer6[51][15:8] = buffer_data_0[3471:3464];
        layer6[51][23:16] = buffer_data_0[3479:3472];
        layer6[51][31:24] = buffer_data_0[3487:3480];
        layer6[51][39:32] = buffer_data_0[3495:3488];
        layer6[51][47:40] = buffer_data_0[3503:3496];
        layer6[51][55:48] = buffer_data_0[3511:3504];
        layer0[52][7:0] = buffer_data_6[3471:3464];
        layer0[52][15:8] = buffer_data_6[3479:3472];
        layer0[52][23:16] = buffer_data_6[3487:3480];
        layer0[52][31:24] = buffer_data_6[3495:3488];
        layer0[52][39:32] = buffer_data_6[3503:3496];
        layer0[52][47:40] = buffer_data_6[3511:3504];
        layer0[52][55:48] = buffer_data_6[3519:3512];
        layer1[52][7:0] = buffer_data_5[3471:3464];
        layer1[52][15:8] = buffer_data_5[3479:3472];
        layer1[52][23:16] = buffer_data_5[3487:3480];
        layer1[52][31:24] = buffer_data_5[3495:3488];
        layer1[52][39:32] = buffer_data_5[3503:3496];
        layer1[52][47:40] = buffer_data_5[3511:3504];
        layer1[52][55:48] = buffer_data_5[3519:3512];
        layer2[52][7:0] = buffer_data_4[3471:3464];
        layer2[52][15:8] = buffer_data_4[3479:3472];
        layer2[52][23:16] = buffer_data_4[3487:3480];
        layer2[52][31:24] = buffer_data_4[3495:3488];
        layer2[52][39:32] = buffer_data_4[3503:3496];
        layer2[52][47:40] = buffer_data_4[3511:3504];
        layer2[52][55:48] = buffer_data_4[3519:3512];
        layer3[52][7:0] = buffer_data_3[3471:3464];
        layer3[52][15:8] = buffer_data_3[3479:3472];
        layer3[52][23:16] = buffer_data_3[3487:3480];
        layer3[52][31:24] = buffer_data_3[3495:3488];
        layer3[52][39:32] = buffer_data_3[3503:3496];
        layer3[52][47:40] = buffer_data_3[3511:3504];
        layer3[52][55:48] = buffer_data_3[3519:3512];
        layer4[52][7:0] = buffer_data_2[3471:3464];
        layer4[52][15:8] = buffer_data_2[3479:3472];
        layer4[52][23:16] = buffer_data_2[3487:3480];
        layer4[52][31:24] = buffer_data_2[3495:3488];
        layer4[52][39:32] = buffer_data_2[3503:3496];
        layer4[52][47:40] = buffer_data_2[3511:3504];
        layer4[52][55:48] = buffer_data_2[3519:3512];
        layer5[52][7:0] = buffer_data_1[3471:3464];
        layer5[52][15:8] = buffer_data_1[3479:3472];
        layer5[52][23:16] = buffer_data_1[3487:3480];
        layer5[52][31:24] = buffer_data_1[3495:3488];
        layer5[52][39:32] = buffer_data_1[3503:3496];
        layer5[52][47:40] = buffer_data_1[3511:3504];
        layer5[52][55:48] = buffer_data_1[3519:3512];
        layer6[52][7:0] = buffer_data_0[3471:3464];
        layer6[52][15:8] = buffer_data_0[3479:3472];
        layer6[52][23:16] = buffer_data_0[3487:3480];
        layer6[52][31:24] = buffer_data_0[3495:3488];
        layer6[52][39:32] = buffer_data_0[3503:3496];
        layer6[52][47:40] = buffer_data_0[3511:3504];
        layer6[52][55:48] = buffer_data_0[3519:3512];
        layer0[53][7:0] = buffer_data_6[3479:3472];
        layer0[53][15:8] = buffer_data_6[3487:3480];
        layer0[53][23:16] = buffer_data_6[3495:3488];
        layer0[53][31:24] = buffer_data_6[3503:3496];
        layer0[53][39:32] = buffer_data_6[3511:3504];
        layer0[53][47:40] = buffer_data_6[3519:3512];
        layer0[53][55:48] = buffer_data_6[3527:3520];
        layer1[53][7:0] = buffer_data_5[3479:3472];
        layer1[53][15:8] = buffer_data_5[3487:3480];
        layer1[53][23:16] = buffer_data_5[3495:3488];
        layer1[53][31:24] = buffer_data_5[3503:3496];
        layer1[53][39:32] = buffer_data_5[3511:3504];
        layer1[53][47:40] = buffer_data_5[3519:3512];
        layer1[53][55:48] = buffer_data_5[3527:3520];
        layer2[53][7:0] = buffer_data_4[3479:3472];
        layer2[53][15:8] = buffer_data_4[3487:3480];
        layer2[53][23:16] = buffer_data_4[3495:3488];
        layer2[53][31:24] = buffer_data_4[3503:3496];
        layer2[53][39:32] = buffer_data_4[3511:3504];
        layer2[53][47:40] = buffer_data_4[3519:3512];
        layer2[53][55:48] = buffer_data_4[3527:3520];
        layer3[53][7:0] = buffer_data_3[3479:3472];
        layer3[53][15:8] = buffer_data_3[3487:3480];
        layer3[53][23:16] = buffer_data_3[3495:3488];
        layer3[53][31:24] = buffer_data_3[3503:3496];
        layer3[53][39:32] = buffer_data_3[3511:3504];
        layer3[53][47:40] = buffer_data_3[3519:3512];
        layer3[53][55:48] = buffer_data_3[3527:3520];
        layer4[53][7:0] = buffer_data_2[3479:3472];
        layer4[53][15:8] = buffer_data_2[3487:3480];
        layer4[53][23:16] = buffer_data_2[3495:3488];
        layer4[53][31:24] = buffer_data_2[3503:3496];
        layer4[53][39:32] = buffer_data_2[3511:3504];
        layer4[53][47:40] = buffer_data_2[3519:3512];
        layer4[53][55:48] = buffer_data_2[3527:3520];
        layer5[53][7:0] = buffer_data_1[3479:3472];
        layer5[53][15:8] = buffer_data_1[3487:3480];
        layer5[53][23:16] = buffer_data_1[3495:3488];
        layer5[53][31:24] = buffer_data_1[3503:3496];
        layer5[53][39:32] = buffer_data_1[3511:3504];
        layer5[53][47:40] = buffer_data_1[3519:3512];
        layer5[53][55:48] = buffer_data_1[3527:3520];
        layer6[53][7:0] = buffer_data_0[3479:3472];
        layer6[53][15:8] = buffer_data_0[3487:3480];
        layer6[53][23:16] = buffer_data_0[3495:3488];
        layer6[53][31:24] = buffer_data_0[3503:3496];
        layer6[53][39:32] = buffer_data_0[3511:3504];
        layer6[53][47:40] = buffer_data_0[3519:3512];
        layer6[53][55:48] = buffer_data_0[3527:3520];
        layer0[54][7:0] = buffer_data_6[3487:3480];
        layer0[54][15:8] = buffer_data_6[3495:3488];
        layer0[54][23:16] = buffer_data_6[3503:3496];
        layer0[54][31:24] = buffer_data_6[3511:3504];
        layer0[54][39:32] = buffer_data_6[3519:3512];
        layer0[54][47:40] = buffer_data_6[3527:3520];
        layer0[54][55:48] = buffer_data_6[3535:3528];
        layer1[54][7:0] = buffer_data_5[3487:3480];
        layer1[54][15:8] = buffer_data_5[3495:3488];
        layer1[54][23:16] = buffer_data_5[3503:3496];
        layer1[54][31:24] = buffer_data_5[3511:3504];
        layer1[54][39:32] = buffer_data_5[3519:3512];
        layer1[54][47:40] = buffer_data_5[3527:3520];
        layer1[54][55:48] = buffer_data_5[3535:3528];
        layer2[54][7:0] = buffer_data_4[3487:3480];
        layer2[54][15:8] = buffer_data_4[3495:3488];
        layer2[54][23:16] = buffer_data_4[3503:3496];
        layer2[54][31:24] = buffer_data_4[3511:3504];
        layer2[54][39:32] = buffer_data_4[3519:3512];
        layer2[54][47:40] = buffer_data_4[3527:3520];
        layer2[54][55:48] = buffer_data_4[3535:3528];
        layer3[54][7:0] = buffer_data_3[3487:3480];
        layer3[54][15:8] = buffer_data_3[3495:3488];
        layer3[54][23:16] = buffer_data_3[3503:3496];
        layer3[54][31:24] = buffer_data_3[3511:3504];
        layer3[54][39:32] = buffer_data_3[3519:3512];
        layer3[54][47:40] = buffer_data_3[3527:3520];
        layer3[54][55:48] = buffer_data_3[3535:3528];
        layer4[54][7:0] = buffer_data_2[3487:3480];
        layer4[54][15:8] = buffer_data_2[3495:3488];
        layer4[54][23:16] = buffer_data_2[3503:3496];
        layer4[54][31:24] = buffer_data_2[3511:3504];
        layer4[54][39:32] = buffer_data_2[3519:3512];
        layer4[54][47:40] = buffer_data_2[3527:3520];
        layer4[54][55:48] = buffer_data_2[3535:3528];
        layer5[54][7:0] = buffer_data_1[3487:3480];
        layer5[54][15:8] = buffer_data_1[3495:3488];
        layer5[54][23:16] = buffer_data_1[3503:3496];
        layer5[54][31:24] = buffer_data_1[3511:3504];
        layer5[54][39:32] = buffer_data_1[3519:3512];
        layer5[54][47:40] = buffer_data_1[3527:3520];
        layer5[54][55:48] = buffer_data_1[3535:3528];
        layer6[54][7:0] = buffer_data_0[3487:3480];
        layer6[54][15:8] = buffer_data_0[3495:3488];
        layer6[54][23:16] = buffer_data_0[3503:3496];
        layer6[54][31:24] = buffer_data_0[3511:3504];
        layer6[54][39:32] = buffer_data_0[3519:3512];
        layer6[54][47:40] = buffer_data_0[3527:3520];
        layer6[54][55:48] = buffer_data_0[3535:3528];
        layer0[55][7:0] = buffer_data_6[3495:3488];
        layer0[55][15:8] = buffer_data_6[3503:3496];
        layer0[55][23:16] = buffer_data_6[3511:3504];
        layer0[55][31:24] = buffer_data_6[3519:3512];
        layer0[55][39:32] = buffer_data_6[3527:3520];
        layer0[55][47:40] = buffer_data_6[3535:3528];
        layer0[55][55:48] = buffer_data_6[3543:3536];
        layer1[55][7:0] = buffer_data_5[3495:3488];
        layer1[55][15:8] = buffer_data_5[3503:3496];
        layer1[55][23:16] = buffer_data_5[3511:3504];
        layer1[55][31:24] = buffer_data_5[3519:3512];
        layer1[55][39:32] = buffer_data_5[3527:3520];
        layer1[55][47:40] = buffer_data_5[3535:3528];
        layer1[55][55:48] = buffer_data_5[3543:3536];
        layer2[55][7:0] = buffer_data_4[3495:3488];
        layer2[55][15:8] = buffer_data_4[3503:3496];
        layer2[55][23:16] = buffer_data_4[3511:3504];
        layer2[55][31:24] = buffer_data_4[3519:3512];
        layer2[55][39:32] = buffer_data_4[3527:3520];
        layer2[55][47:40] = buffer_data_4[3535:3528];
        layer2[55][55:48] = buffer_data_4[3543:3536];
        layer3[55][7:0] = buffer_data_3[3495:3488];
        layer3[55][15:8] = buffer_data_3[3503:3496];
        layer3[55][23:16] = buffer_data_3[3511:3504];
        layer3[55][31:24] = buffer_data_3[3519:3512];
        layer3[55][39:32] = buffer_data_3[3527:3520];
        layer3[55][47:40] = buffer_data_3[3535:3528];
        layer3[55][55:48] = buffer_data_3[3543:3536];
        layer4[55][7:0] = buffer_data_2[3495:3488];
        layer4[55][15:8] = buffer_data_2[3503:3496];
        layer4[55][23:16] = buffer_data_2[3511:3504];
        layer4[55][31:24] = buffer_data_2[3519:3512];
        layer4[55][39:32] = buffer_data_2[3527:3520];
        layer4[55][47:40] = buffer_data_2[3535:3528];
        layer4[55][55:48] = buffer_data_2[3543:3536];
        layer5[55][7:0] = buffer_data_1[3495:3488];
        layer5[55][15:8] = buffer_data_1[3503:3496];
        layer5[55][23:16] = buffer_data_1[3511:3504];
        layer5[55][31:24] = buffer_data_1[3519:3512];
        layer5[55][39:32] = buffer_data_1[3527:3520];
        layer5[55][47:40] = buffer_data_1[3535:3528];
        layer5[55][55:48] = buffer_data_1[3543:3536];
        layer6[55][7:0] = buffer_data_0[3495:3488];
        layer6[55][15:8] = buffer_data_0[3503:3496];
        layer6[55][23:16] = buffer_data_0[3511:3504];
        layer6[55][31:24] = buffer_data_0[3519:3512];
        layer6[55][39:32] = buffer_data_0[3527:3520];
        layer6[55][47:40] = buffer_data_0[3535:3528];
        layer6[55][55:48] = buffer_data_0[3543:3536];
        layer0[56][7:0] = buffer_data_6[3503:3496];
        layer0[56][15:8] = buffer_data_6[3511:3504];
        layer0[56][23:16] = buffer_data_6[3519:3512];
        layer0[56][31:24] = buffer_data_6[3527:3520];
        layer0[56][39:32] = buffer_data_6[3535:3528];
        layer0[56][47:40] = buffer_data_6[3543:3536];
        layer0[56][55:48] = buffer_data_6[3551:3544];
        layer1[56][7:0] = buffer_data_5[3503:3496];
        layer1[56][15:8] = buffer_data_5[3511:3504];
        layer1[56][23:16] = buffer_data_5[3519:3512];
        layer1[56][31:24] = buffer_data_5[3527:3520];
        layer1[56][39:32] = buffer_data_5[3535:3528];
        layer1[56][47:40] = buffer_data_5[3543:3536];
        layer1[56][55:48] = buffer_data_5[3551:3544];
        layer2[56][7:0] = buffer_data_4[3503:3496];
        layer2[56][15:8] = buffer_data_4[3511:3504];
        layer2[56][23:16] = buffer_data_4[3519:3512];
        layer2[56][31:24] = buffer_data_4[3527:3520];
        layer2[56][39:32] = buffer_data_4[3535:3528];
        layer2[56][47:40] = buffer_data_4[3543:3536];
        layer2[56][55:48] = buffer_data_4[3551:3544];
        layer3[56][7:0] = buffer_data_3[3503:3496];
        layer3[56][15:8] = buffer_data_3[3511:3504];
        layer3[56][23:16] = buffer_data_3[3519:3512];
        layer3[56][31:24] = buffer_data_3[3527:3520];
        layer3[56][39:32] = buffer_data_3[3535:3528];
        layer3[56][47:40] = buffer_data_3[3543:3536];
        layer3[56][55:48] = buffer_data_3[3551:3544];
        layer4[56][7:0] = buffer_data_2[3503:3496];
        layer4[56][15:8] = buffer_data_2[3511:3504];
        layer4[56][23:16] = buffer_data_2[3519:3512];
        layer4[56][31:24] = buffer_data_2[3527:3520];
        layer4[56][39:32] = buffer_data_2[3535:3528];
        layer4[56][47:40] = buffer_data_2[3543:3536];
        layer4[56][55:48] = buffer_data_2[3551:3544];
        layer5[56][7:0] = buffer_data_1[3503:3496];
        layer5[56][15:8] = buffer_data_1[3511:3504];
        layer5[56][23:16] = buffer_data_1[3519:3512];
        layer5[56][31:24] = buffer_data_1[3527:3520];
        layer5[56][39:32] = buffer_data_1[3535:3528];
        layer5[56][47:40] = buffer_data_1[3543:3536];
        layer5[56][55:48] = buffer_data_1[3551:3544];
        layer6[56][7:0] = buffer_data_0[3503:3496];
        layer6[56][15:8] = buffer_data_0[3511:3504];
        layer6[56][23:16] = buffer_data_0[3519:3512];
        layer6[56][31:24] = buffer_data_0[3527:3520];
        layer6[56][39:32] = buffer_data_0[3535:3528];
        layer6[56][47:40] = buffer_data_0[3543:3536];
        layer6[56][55:48] = buffer_data_0[3551:3544];
        layer0[57][7:0] = buffer_data_6[3511:3504];
        layer0[57][15:8] = buffer_data_6[3519:3512];
        layer0[57][23:16] = buffer_data_6[3527:3520];
        layer0[57][31:24] = buffer_data_6[3535:3528];
        layer0[57][39:32] = buffer_data_6[3543:3536];
        layer0[57][47:40] = buffer_data_6[3551:3544];
        layer0[57][55:48] = buffer_data_6[3559:3552];
        layer1[57][7:0] = buffer_data_5[3511:3504];
        layer1[57][15:8] = buffer_data_5[3519:3512];
        layer1[57][23:16] = buffer_data_5[3527:3520];
        layer1[57][31:24] = buffer_data_5[3535:3528];
        layer1[57][39:32] = buffer_data_5[3543:3536];
        layer1[57][47:40] = buffer_data_5[3551:3544];
        layer1[57][55:48] = buffer_data_5[3559:3552];
        layer2[57][7:0] = buffer_data_4[3511:3504];
        layer2[57][15:8] = buffer_data_4[3519:3512];
        layer2[57][23:16] = buffer_data_4[3527:3520];
        layer2[57][31:24] = buffer_data_4[3535:3528];
        layer2[57][39:32] = buffer_data_4[3543:3536];
        layer2[57][47:40] = buffer_data_4[3551:3544];
        layer2[57][55:48] = buffer_data_4[3559:3552];
        layer3[57][7:0] = buffer_data_3[3511:3504];
        layer3[57][15:8] = buffer_data_3[3519:3512];
        layer3[57][23:16] = buffer_data_3[3527:3520];
        layer3[57][31:24] = buffer_data_3[3535:3528];
        layer3[57][39:32] = buffer_data_3[3543:3536];
        layer3[57][47:40] = buffer_data_3[3551:3544];
        layer3[57][55:48] = buffer_data_3[3559:3552];
        layer4[57][7:0] = buffer_data_2[3511:3504];
        layer4[57][15:8] = buffer_data_2[3519:3512];
        layer4[57][23:16] = buffer_data_2[3527:3520];
        layer4[57][31:24] = buffer_data_2[3535:3528];
        layer4[57][39:32] = buffer_data_2[3543:3536];
        layer4[57][47:40] = buffer_data_2[3551:3544];
        layer4[57][55:48] = buffer_data_2[3559:3552];
        layer5[57][7:0] = buffer_data_1[3511:3504];
        layer5[57][15:8] = buffer_data_1[3519:3512];
        layer5[57][23:16] = buffer_data_1[3527:3520];
        layer5[57][31:24] = buffer_data_1[3535:3528];
        layer5[57][39:32] = buffer_data_1[3543:3536];
        layer5[57][47:40] = buffer_data_1[3551:3544];
        layer5[57][55:48] = buffer_data_1[3559:3552];
        layer6[57][7:0] = buffer_data_0[3511:3504];
        layer6[57][15:8] = buffer_data_0[3519:3512];
        layer6[57][23:16] = buffer_data_0[3527:3520];
        layer6[57][31:24] = buffer_data_0[3535:3528];
        layer6[57][39:32] = buffer_data_0[3543:3536];
        layer6[57][47:40] = buffer_data_0[3551:3544];
        layer6[57][55:48] = buffer_data_0[3559:3552];
        layer0[58][7:0] = buffer_data_6[3519:3512];
        layer0[58][15:8] = buffer_data_6[3527:3520];
        layer0[58][23:16] = buffer_data_6[3535:3528];
        layer0[58][31:24] = buffer_data_6[3543:3536];
        layer0[58][39:32] = buffer_data_6[3551:3544];
        layer0[58][47:40] = buffer_data_6[3559:3552];
        layer0[58][55:48] = buffer_data_6[3567:3560];
        layer1[58][7:0] = buffer_data_5[3519:3512];
        layer1[58][15:8] = buffer_data_5[3527:3520];
        layer1[58][23:16] = buffer_data_5[3535:3528];
        layer1[58][31:24] = buffer_data_5[3543:3536];
        layer1[58][39:32] = buffer_data_5[3551:3544];
        layer1[58][47:40] = buffer_data_5[3559:3552];
        layer1[58][55:48] = buffer_data_5[3567:3560];
        layer2[58][7:0] = buffer_data_4[3519:3512];
        layer2[58][15:8] = buffer_data_4[3527:3520];
        layer2[58][23:16] = buffer_data_4[3535:3528];
        layer2[58][31:24] = buffer_data_4[3543:3536];
        layer2[58][39:32] = buffer_data_4[3551:3544];
        layer2[58][47:40] = buffer_data_4[3559:3552];
        layer2[58][55:48] = buffer_data_4[3567:3560];
        layer3[58][7:0] = buffer_data_3[3519:3512];
        layer3[58][15:8] = buffer_data_3[3527:3520];
        layer3[58][23:16] = buffer_data_3[3535:3528];
        layer3[58][31:24] = buffer_data_3[3543:3536];
        layer3[58][39:32] = buffer_data_3[3551:3544];
        layer3[58][47:40] = buffer_data_3[3559:3552];
        layer3[58][55:48] = buffer_data_3[3567:3560];
        layer4[58][7:0] = buffer_data_2[3519:3512];
        layer4[58][15:8] = buffer_data_2[3527:3520];
        layer4[58][23:16] = buffer_data_2[3535:3528];
        layer4[58][31:24] = buffer_data_2[3543:3536];
        layer4[58][39:32] = buffer_data_2[3551:3544];
        layer4[58][47:40] = buffer_data_2[3559:3552];
        layer4[58][55:48] = buffer_data_2[3567:3560];
        layer5[58][7:0] = buffer_data_1[3519:3512];
        layer5[58][15:8] = buffer_data_1[3527:3520];
        layer5[58][23:16] = buffer_data_1[3535:3528];
        layer5[58][31:24] = buffer_data_1[3543:3536];
        layer5[58][39:32] = buffer_data_1[3551:3544];
        layer5[58][47:40] = buffer_data_1[3559:3552];
        layer5[58][55:48] = buffer_data_1[3567:3560];
        layer6[58][7:0] = buffer_data_0[3519:3512];
        layer6[58][15:8] = buffer_data_0[3527:3520];
        layer6[58][23:16] = buffer_data_0[3535:3528];
        layer6[58][31:24] = buffer_data_0[3543:3536];
        layer6[58][39:32] = buffer_data_0[3551:3544];
        layer6[58][47:40] = buffer_data_0[3559:3552];
        layer6[58][55:48] = buffer_data_0[3567:3560];
        layer0[59][7:0] = buffer_data_6[3527:3520];
        layer0[59][15:8] = buffer_data_6[3535:3528];
        layer0[59][23:16] = buffer_data_6[3543:3536];
        layer0[59][31:24] = buffer_data_6[3551:3544];
        layer0[59][39:32] = buffer_data_6[3559:3552];
        layer0[59][47:40] = buffer_data_6[3567:3560];
        layer0[59][55:48] = buffer_data_6[3575:3568];
        layer1[59][7:0] = buffer_data_5[3527:3520];
        layer1[59][15:8] = buffer_data_5[3535:3528];
        layer1[59][23:16] = buffer_data_5[3543:3536];
        layer1[59][31:24] = buffer_data_5[3551:3544];
        layer1[59][39:32] = buffer_data_5[3559:3552];
        layer1[59][47:40] = buffer_data_5[3567:3560];
        layer1[59][55:48] = buffer_data_5[3575:3568];
        layer2[59][7:0] = buffer_data_4[3527:3520];
        layer2[59][15:8] = buffer_data_4[3535:3528];
        layer2[59][23:16] = buffer_data_4[3543:3536];
        layer2[59][31:24] = buffer_data_4[3551:3544];
        layer2[59][39:32] = buffer_data_4[3559:3552];
        layer2[59][47:40] = buffer_data_4[3567:3560];
        layer2[59][55:48] = buffer_data_4[3575:3568];
        layer3[59][7:0] = buffer_data_3[3527:3520];
        layer3[59][15:8] = buffer_data_3[3535:3528];
        layer3[59][23:16] = buffer_data_3[3543:3536];
        layer3[59][31:24] = buffer_data_3[3551:3544];
        layer3[59][39:32] = buffer_data_3[3559:3552];
        layer3[59][47:40] = buffer_data_3[3567:3560];
        layer3[59][55:48] = buffer_data_3[3575:3568];
        layer4[59][7:0] = buffer_data_2[3527:3520];
        layer4[59][15:8] = buffer_data_2[3535:3528];
        layer4[59][23:16] = buffer_data_2[3543:3536];
        layer4[59][31:24] = buffer_data_2[3551:3544];
        layer4[59][39:32] = buffer_data_2[3559:3552];
        layer4[59][47:40] = buffer_data_2[3567:3560];
        layer4[59][55:48] = buffer_data_2[3575:3568];
        layer5[59][7:0] = buffer_data_1[3527:3520];
        layer5[59][15:8] = buffer_data_1[3535:3528];
        layer5[59][23:16] = buffer_data_1[3543:3536];
        layer5[59][31:24] = buffer_data_1[3551:3544];
        layer5[59][39:32] = buffer_data_1[3559:3552];
        layer5[59][47:40] = buffer_data_1[3567:3560];
        layer5[59][55:48] = buffer_data_1[3575:3568];
        layer6[59][7:0] = buffer_data_0[3527:3520];
        layer6[59][15:8] = buffer_data_0[3535:3528];
        layer6[59][23:16] = buffer_data_0[3543:3536];
        layer6[59][31:24] = buffer_data_0[3551:3544];
        layer6[59][39:32] = buffer_data_0[3559:3552];
        layer6[59][47:40] = buffer_data_0[3567:3560];
        layer6[59][55:48] = buffer_data_0[3575:3568];
        layer0[60][7:0] = buffer_data_6[3535:3528];
        layer0[60][15:8] = buffer_data_6[3543:3536];
        layer0[60][23:16] = buffer_data_6[3551:3544];
        layer0[60][31:24] = buffer_data_6[3559:3552];
        layer0[60][39:32] = buffer_data_6[3567:3560];
        layer0[60][47:40] = buffer_data_6[3575:3568];
        layer0[60][55:48] = buffer_data_6[3583:3576];
        layer1[60][7:0] = buffer_data_5[3535:3528];
        layer1[60][15:8] = buffer_data_5[3543:3536];
        layer1[60][23:16] = buffer_data_5[3551:3544];
        layer1[60][31:24] = buffer_data_5[3559:3552];
        layer1[60][39:32] = buffer_data_5[3567:3560];
        layer1[60][47:40] = buffer_data_5[3575:3568];
        layer1[60][55:48] = buffer_data_5[3583:3576];
        layer2[60][7:0] = buffer_data_4[3535:3528];
        layer2[60][15:8] = buffer_data_4[3543:3536];
        layer2[60][23:16] = buffer_data_4[3551:3544];
        layer2[60][31:24] = buffer_data_4[3559:3552];
        layer2[60][39:32] = buffer_data_4[3567:3560];
        layer2[60][47:40] = buffer_data_4[3575:3568];
        layer2[60][55:48] = buffer_data_4[3583:3576];
        layer3[60][7:0] = buffer_data_3[3535:3528];
        layer3[60][15:8] = buffer_data_3[3543:3536];
        layer3[60][23:16] = buffer_data_3[3551:3544];
        layer3[60][31:24] = buffer_data_3[3559:3552];
        layer3[60][39:32] = buffer_data_3[3567:3560];
        layer3[60][47:40] = buffer_data_3[3575:3568];
        layer3[60][55:48] = buffer_data_3[3583:3576];
        layer4[60][7:0] = buffer_data_2[3535:3528];
        layer4[60][15:8] = buffer_data_2[3543:3536];
        layer4[60][23:16] = buffer_data_2[3551:3544];
        layer4[60][31:24] = buffer_data_2[3559:3552];
        layer4[60][39:32] = buffer_data_2[3567:3560];
        layer4[60][47:40] = buffer_data_2[3575:3568];
        layer4[60][55:48] = buffer_data_2[3583:3576];
        layer5[60][7:0] = buffer_data_1[3535:3528];
        layer5[60][15:8] = buffer_data_1[3543:3536];
        layer5[60][23:16] = buffer_data_1[3551:3544];
        layer5[60][31:24] = buffer_data_1[3559:3552];
        layer5[60][39:32] = buffer_data_1[3567:3560];
        layer5[60][47:40] = buffer_data_1[3575:3568];
        layer5[60][55:48] = buffer_data_1[3583:3576];
        layer6[60][7:0] = buffer_data_0[3535:3528];
        layer6[60][15:8] = buffer_data_0[3543:3536];
        layer6[60][23:16] = buffer_data_0[3551:3544];
        layer6[60][31:24] = buffer_data_0[3559:3552];
        layer6[60][39:32] = buffer_data_0[3567:3560];
        layer6[60][47:40] = buffer_data_0[3575:3568];
        layer6[60][55:48] = buffer_data_0[3583:3576];
        layer0[61][7:0] = buffer_data_6[3543:3536];
        layer0[61][15:8] = buffer_data_6[3551:3544];
        layer0[61][23:16] = buffer_data_6[3559:3552];
        layer0[61][31:24] = buffer_data_6[3567:3560];
        layer0[61][39:32] = buffer_data_6[3575:3568];
        layer0[61][47:40] = buffer_data_6[3583:3576];
        layer0[61][55:48] = buffer_data_6[3591:3584];
        layer1[61][7:0] = buffer_data_5[3543:3536];
        layer1[61][15:8] = buffer_data_5[3551:3544];
        layer1[61][23:16] = buffer_data_5[3559:3552];
        layer1[61][31:24] = buffer_data_5[3567:3560];
        layer1[61][39:32] = buffer_data_5[3575:3568];
        layer1[61][47:40] = buffer_data_5[3583:3576];
        layer1[61][55:48] = buffer_data_5[3591:3584];
        layer2[61][7:0] = buffer_data_4[3543:3536];
        layer2[61][15:8] = buffer_data_4[3551:3544];
        layer2[61][23:16] = buffer_data_4[3559:3552];
        layer2[61][31:24] = buffer_data_4[3567:3560];
        layer2[61][39:32] = buffer_data_4[3575:3568];
        layer2[61][47:40] = buffer_data_4[3583:3576];
        layer2[61][55:48] = buffer_data_4[3591:3584];
        layer3[61][7:0] = buffer_data_3[3543:3536];
        layer3[61][15:8] = buffer_data_3[3551:3544];
        layer3[61][23:16] = buffer_data_3[3559:3552];
        layer3[61][31:24] = buffer_data_3[3567:3560];
        layer3[61][39:32] = buffer_data_3[3575:3568];
        layer3[61][47:40] = buffer_data_3[3583:3576];
        layer3[61][55:48] = buffer_data_3[3591:3584];
        layer4[61][7:0] = buffer_data_2[3543:3536];
        layer4[61][15:8] = buffer_data_2[3551:3544];
        layer4[61][23:16] = buffer_data_2[3559:3552];
        layer4[61][31:24] = buffer_data_2[3567:3560];
        layer4[61][39:32] = buffer_data_2[3575:3568];
        layer4[61][47:40] = buffer_data_2[3583:3576];
        layer4[61][55:48] = buffer_data_2[3591:3584];
        layer5[61][7:0] = buffer_data_1[3543:3536];
        layer5[61][15:8] = buffer_data_1[3551:3544];
        layer5[61][23:16] = buffer_data_1[3559:3552];
        layer5[61][31:24] = buffer_data_1[3567:3560];
        layer5[61][39:32] = buffer_data_1[3575:3568];
        layer5[61][47:40] = buffer_data_1[3583:3576];
        layer5[61][55:48] = buffer_data_1[3591:3584];
        layer6[61][7:0] = buffer_data_0[3543:3536];
        layer6[61][15:8] = buffer_data_0[3551:3544];
        layer6[61][23:16] = buffer_data_0[3559:3552];
        layer6[61][31:24] = buffer_data_0[3567:3560];
        layer6[61][39:32] = buffer_data_0[3575:3568];
        layer6[61][47:40] = buffer_data_0[3583:3576];
        layer6[61][55:48] = buffer_data_0[3591:3584];
        layer0[62][7:0] = buffer_data_6[3551:3544];
        layer0[62][15:8] = buffer_data_6[3559:3552];
        layer0[62][23:16] = buffer_data_6[3567:3560];
        layer0[62][31:24] = buffer_data_6[3575:3568];
        layer0[62][39:32] = buffer_data_6[3583:3576];
        layer0[62][47:40] = buffer_data_6[3591:3584];
        layer0[62][55:48] = buffer_data_6[3599:3592];
        layer1[62][7:0] = buffer_data_5[3551:3544];
        layer1[62][15:8] = buffer_data_5[3559:3552];
        layer1[62][23:16] = buffer_data_5[3567:3560];
        layer1[62][31:24] = buffer_data_5[3575:3568];
        layer1[62][39:32] = buffer_data_5[3583:3576];
        layer1[62][47:40] = buffer_data_5[3591:3584];
        layer1[62][55:48] = buffer_data_5[3599:3592];
        layer2[62][7:0] = buffer_data_4[3551:3544];
        layer2[62][15:8] = buffer_data_4[3559:3552];
        layer2[62][23:16] = buffer_data_4[3567:3560];
        layer2[62][31:24] = buffer_data_4[3575:3568];
        layer2[62][39:32] = buffer_data_4[3583:3576];
        layer2[62][47:40] = buffer_data_4[3591:3584];
        layer2[62][55:48] = buffer_data_4[3599:3592];
        layer3[62][7:0] = buffer_data_3[3551:3544];
        layer3[62][15:8] = buffer_data_3[3559:3552];
        layer3[62][23:16] = buffer_data_3[3567:3560];
        layer3[62][31:24] = buffer_data_3[3575:3568];
        layer3[62][39:32] = buffer_data_3[3583:3576];
        layer3[62][47:40] = buffer_data_3[3591:3584];
        layer3[62][55:48] = buffer_data_3[3599:3592];
        layer4[62][7:0] = buffer_data_2[3551:3544];
        layer4[62][15:8] = buffer_data_2[3559:3552];
        layer4[62][23:16] = buffer_data_2[3567:3560];
        layer4[62][31:24] = buffer_data_2[3575:3568];
        layer4[62][39:32] = buffer_data_2[3583:3576];
        layer4[62][47:40] = buffer_data_2[3591:3584];
        layer4[62][55:48] = buffer_data_2[3599:3592];
        layer5[62][7:0] = buffer_data_1[3551:3544];
        layer5[62][15:8] = buffer_data_1[3559:3552];
        layer5[62][23:16] = buffer_data_1[3567:3560];
        layer5[62][31:24] = buffer_data_1[3575:3568];
        layer5[62][39:32] = buffer_data_1[3583:3576];
        layer5[62][47:40] = buffer_data_1[3591:3584];
        layer5[62][55:48] = buffer_data_1[3599:3592];
        layer6[62][7:0] = buffer_data_0[3551:3544];
        layer6[62][15:8] = buffer_data_0[3559:3552];
        layer6[62][23:16] = buffer_data_0[3567:3560];
        layer6[62][31:24] = buffer_data_0[3575:3568];
        layer6[62][39:32] = buffer_data_0[3583:3576];
        layer6[62][47:40] = buffer_data_0[3591:3584];
        layer6[62][55:48] = buffer_data_0[3599:3592];
        layer0[63][7:0] = buffer_data_6[3559:3552];
        layer0[63][15:8] = buffer_data_6[3567:3560];
        layer0[63][23:16] = buffer_data_6[3575:3568];
        layer0[63][31:24] = buffer_data_6[3583:3576];
        layer0[63][39:32] = buffer_data_6[3591:3584];
        layer0[63][47:40] = buffer_data_6[3599:3592];
        layer0[63][55:48] = buffer_data_6[3607:3600];
        layer1[63][7:0] = buffer_data_5[3559:3552];
        layer1[63][15:8] = buffer_data_5[3567:3560];
        layer1[63][23:16] = buffer_data_5[3575:3568];
        layer1[63][31:24] = buffer_data_5[3583:3576];
        layer1[63][39:32] = buffer_data_5[3591:3584];
        layer1[63][47:40] = buffer_data_5[3599:3592];
        layer1[63][55:48] = buffer_data_5[3607:3600];
        layer2[63][7:0] = buffer_data_4[3559:3552];
        layer2[63][15:8] = buffer_data_4[3567:3560];
        layer2[63][23:16] = buffer_data_4[3575:3568];
        layer2[63][31:24] = buffer_data_4[3583:3576];
        layer2[63][39:32] = buffer_data_4[3591:3584];
        layer2[63][47:40] = buffer_data_4[3599:3592];
        layer2[63][55:48] = buffer_data_4[3607:3600];
        layer3[63][7:0] = buffer_data_3[3559:3552];
        layer3[63][15:8] = buffer_data_3[3567:3560];
        layer3[63][23:16] = buffer_data_3[3575:3568];
        layer3[63][31:24] = buffer_data_3[3583:3576];
        layer3[63][39:32] = buffer_data_3[3591:3584];
        layer3[63][47:40] = buffer_data_3[3599:3592];
        layer3[63][55:48] = buffer_data_3[3607:3600];
        layer4[63][7:0] = buffer_data_2[3559:3552];
        layer4[63][15:8] = buffer_data_2[3567:3560];
        layer4[63][23:16] = buffer_data_2[3575:3568];
        layer4[63][31:24] = buffer_data_2[3583:3576];
        layer4[63][39:32] = buffer_data_2[3591:3584];
        layer4[63][47:40] = buffer_data_2[3599:3592];
        layer4[63][55:48] = buffer_data_2[3607:3600];
        layer5[63][7:0] = buffer_data_1[3559:3552];
        layer5[63][15:8] = buffer_data_1[3567:3560];
        layer5[63][23:16] = buffer_data_1[3575:3568];
        layer5[63][31:24] = buffer_data_1[3583:3576];
        layer5[63][39:32] = buffer_data_1[3591:3584];
        layer5[63][47:40] = buffer_data_1[3599:3592];
        layer5[63][55:48] = buffer_data_1[3607:3600];
        layer6[63][7:0] = buffer_data_0[3559:3552];
        layer6[63][15:8] = buffer_data_0[3567:3560];
        layer6[63][23:16] = buffer_data_0[3575:3568];
        layer6[63][31:24] = buffer_data_0[3583:3576];
        layer6[63][39:32] = buffer_data_0[3591:3584];
        layer6[63][47:40] = buffer_data_0[3599:3592];
        layer6[63][55:48] = buffer_data_0[3607:3600];
    end
    ST_GAUSSIAN_7: begin
        layer0[0][7:0] = buffer_data_6[3567:3560];
        layer0[0][15:8] = buffer_data_6[3575:3568];
        layer0[0][23:16] = buffer_data_6[3583:3576];
        layer0[0][31:24] = buffer_data_6[3591:3584];
        layer0[0][39:32] = buffer_data_6[3599:3592];
        layer0[0][47:40] = buffer_data_6[3607:3600];
        layer0[0][55:48] = buffer_data_6[3615:3608];
        layer1[0][7:0] = buffer_data_5[3567:3560];
        layer1[0][15:8] = buffer_data_5[3575:3568];
        layer1[0][23:16] = buffer_data_5[3583:3576];
        layer1[0][31:24] = buffer_data_5[3591:3584];
        layer1[0][39:32] = buffer_data_5[3599:3592];
        layer1[0][47:40] = buffer_data_5[3607:3600];
        layer1[0][55:48] = buffer_data_5[3615:3608];
        layer2[0][7:0] = buffer_data_4[3567:3560];
        layer2[0][15:8] = buffer_data_4[3575:3568];
        layer2[0][23:16] = buffer_data_4[3583:3576];
        layer2[0][31:24] = buffer_data_4[3591:3584];
        layer2[0][39:32] = buffer_data_4[3599:3592];
        layer2[0][47:40] = buffer_data_4[3607:3600];
        layer2[0][55:48] = buffer_data_4[3615:3608];
        layer3[0][7:0] = buffer_data_3[3567:3560];
        layer3[0][15:8] = buffer_data_3[3575:3568];
        layer3[0][23:16] = buffer_data_3[3583:3576];
        layer3[0][31:24] = buffer_data_3[3591:3584];
        layer3[0][39:32] = buffer_data_3[3599:3592];
        layer3[0][47:40] = buffer_data_3[3607:3600];
        layer3[0][55:48] = buffer_data_3[3615:3608];
        layer4[0][7:0] = buffer_data_2[3567:3560];
        layer4[0][15:8] = buffer_data_2[3575:3568];
        layer4[0][23:16] = buffer_data_2[3583:3576];
        layer4[0][31:24] = buffer_data_2[3591:3584];
        layer4[0][39:32] = buffer_data_2[3599:3592];
        layer4[0][47:40] = buffer_data_2[3607:3600];
        layer4[0][55:48] = buffer_data_2[3615:3608];
        layer5[0][7:0] = buffer_data_1[3567:3560];
        layer5[0][15:8] = buffer_data_1[3575:3568];
        layer5[0][23:16] = buffer_data_1[3583:3576];
        layer5[0][31:24] = buffer_data_1[3591:3584];
        layer5[0][39:32] = buffer_data_1[3599:3592];
        layer5[0][47:40] = buffer_data_1[3607:3600];
        layer5[0][55:48] = buffer_data_1[3615:3608];
        layer6[0][7:0] = buffer_data_0[3567:3560];
        layer6[0][15:8] = buffer_data_0[3575:3568];
        layer6[0][23:16] = buffer_data_0[3583:3576];
        layer6[0][31:24] = buffer_data_0[3591:3584];
        layer6[0][39:32] = buffer_data_0[3599:3592];
        layer6[0][47:40] = buffer_data_0[3607:3600];
        layer6[0][55:48] = buffer_data_0[3615:3608];
        layer0[1][7:0] = buffer_data_6[3575:3568];
        layer0[1][15:8] = buffer_data_6[3583:3576];
        layer0[1][23:16] = buffer_data_6[3591:3584];
        layer0[1][31:24] = buffer_data_6[3599:3592];
        layer0[1][39:32] = buffer_data_6[3607:3600];
        layer0[1][47:40] = buffer_data_6[3615:3608];
        layer0[1][55:48] = buffer_data_6[3623:3616];
        layer1[1][7:0] = buffer_data_5[3575:3568];
        layer1[1][15:8] = buffer_data_5[3583:3576];
        layer1[1][23:16] = buffer_data_5[3591:3584];
        layer1[1][31:24] = buffer_data_5[3599:3592];
        layer1[1][39:32] = buffer_data_5[3607:3600];
        layer1[1][47:40] = buffer_data_5[3615:3608];
        layer1[1][55:48] = buffer_data_5[3623:3616];
        layer2[1][7:0] = buffer_data_4[3575:3568];
        layer2[1][15:8] = buffer_data_4[3583:3576];
        layer2[1][23:16] = buffer_data_4[3591:3584];
        layer2[1][31:24] = buffer_data_4[3599:3592];
        layer2[1][39:32] = buffer_data_4[3607:3600];
        layer2[1][47:40] = buffer_data_4[3615:3608];
        layer2[1][55:48] = buffer_data_4[3623:3616];
        layer3[1][7:0] = buffer_data_3[3575:3568];
        layer3[1][15:8] = buffer_data_3[3583:3576];
        layer3[1][23:16] = buffer_data_3[3591:3584];
        layer3[1][31:24] = buffer_data_3[3599:3592];
        layer3[1][39:32] = buffer_data_3[3607:3600];
        layer3[1][47:40] = buffer_data_3[3615:3608];
        layer3[1][55:48] = buffer_data_3[3623:3616];
        layer4[1][7:0] = buffer_data_2[3575:3568];
        layer4[1][15:8] = buffer_data_2[3583:3576];
        layer4[1][23:16] = buffer_data_2[3591:3584];
        layer4[1][31:24] = buffer_data_2[3599:3592];
        layer4[1][39:32] = buffer_data_2[3607:3600];
        layer4[1][47:40] = buffer_data_2[3615:3608];
        layer4[1][55:48] = buffer_data_2[3623:3616];
        layer5[1][7:0] = buffer_data_1[3575:3568];
        layer5[1][15:8] = buffer_data_1[3583:3576];
        layer5[1][23:16] = buffer_data_1[3591:3584];
        layer5[1][31:24] = buffer_data_1[3599:3592];
        layer5[1][39:32] = buffer_data_1[3607:3600];
        layer5[1][47:40] = buffer_data_1[3615:3608];
        layer5[1][55:48] = buffer_data_1[3623:3616];
        layer6[1][7:0] = buffer_data_0[3575:3568];
        layer6[1][15:8] = buffer_data_0[3583:3576];
        layer6[1][23:16] = buffer_data_0[3591:3584];
        layer6[1][31:24] = buffer_data_0[3599:3592];
        layer6[1][39:32] = buffer_data_0[3607:3600];
        layer6[1][47:40] = buffer_data_0[3615:3608];
        layer6[1][55:48] = buffer_data_0[3623:3616];
        layer0[2][7:0] = buffer_data_6[3583:3576];
        layer0[2][15:8] = buffer_data_6[3591:3584];
        layer0[2][23:16] = buffer_data_6[3599:3592];
        layer0[2][31:24] = buffer_data_6[3607:3600];
        layer0[2][39:32] = buffer_data_6[3615:3608];
        layer0[2][47:40] = buffer_data_6[3623:3616];
        layer0[2][55:48] = buffer_data_6[3631:3624];
        layer1[2][7:0] = buffer_data_5[3583:3576];
        layer1[2][15:8] = buffer_data_5[3591:3584];
        layer1[2][23:16] = buffer_data_5[3599:3592];
        layer1[2][31:24] = buffer_data_5[3607:3600];
        layer1[2][39:32] = buffer_data_5[3615:3608];
        layer1[2][47:40] = buffer_data_5[3623:3616];
        layer1[2][55:48] = buffer_data_5[3631:3624];
        layer2[2][7:0] = buffer_data_4[3583:3576];
        layer2[2][15:8] = buffer_data_4[3591:3584];
        layer2[2][23:16] = buffer_data_4[3599:3592];
        layer2[2][31:24] = buffer_data_4[3607:3600];
        layer2[2][39:32] = buffer_data_4[3615:3608];
        layer2[2][47:40] = buffer_data_4[3623:3616];
        layer2[2][55:48] = buffer_data_4[3631:3624];
        layer3[2][7:0] = buffer_data_3[3583:3576];
        layer3[2][15:8] = buffer_data_3[3591:3584];
        layer3[2][23:16] = buffer_data_3[3599:3592];
        layer3[2][31:24] = buffer_data_3[3607:3600];
        layer3[2][39:32] = buffer_data_3[3615:3608];
        layer3[2][47:40] = buffer_data_3[3623:3616];
        layer3[2][55:48] = buffer_data_3[3631:3624];
        layer4[2][7:0] = buffer_data_2[3583:3576];
        layer4[2][15:8] = buffer_data_2[3591:3584];
        layer4[2][23:16] = buffer_data_2[3599:3592];
        layer4[2][31:24] = buffer_data_2[3607:3600];
        layer4[2][39:32] = buffer_data_2[3615:3608];
        layer4[2][47:40] = buffer_data_2[3623:3616];
        layer4[2][55:48] = buffer_data_2[3631:3624];
        layer5[2][7:0] = buffer_data_1[3583:3576];
        layer5[2][15:8] = buffer_data_1[3591:3584];
        layer5[2][23:16] = buffer_data_1[3599:3592];
        layer5[2][31:24] = buffer_data_1[3607:3600];
        layer5[2][39:32] = buffer_data_1[3615:3608];
        layer5[2][47:40] = buffer_data_1[3623:3616];
        layer5[2][55:48] = buffer_data_1[3631:3624];
        layer6[2][7:0] = buffer_data_0[3583:3576];
        layer6[2][15:8] = buffer_data_0[3591:3584];
        layer6[2][23:16] = buffer_data_0[3599:3592];
        layer6[2][31:24] = buffer_data_0[3607:3600];
        layer6[2][39:32] = buffer_data_0[3615:3608];
        layer6[2][47:40] = buffer_data_0[3623:3616];
        layer6[2][55:48] = buffer_data_0[3631:3624];
        layer0[3][7:0] = buffer_data_6[3591:3584];
        layer0[3][15:8] = buffer_data_6[3599:3592];
        layer0[3][23:16] = buffer_data_6[3607:3600];
        layer0[3][31:24] = buffer_data_6[3615:3608];
        layer0[3][39:32] = buffer_data_6[3623:3616];
        layer0[3][47:40] = buffer_data_6[3631:3624];
        layer0[3][55:48] = buffer_data_6[3639:3632];
        layer1[3][7:0] = buffer_data_5[3591:3584];
        layer1[3][15:8] = buffer_data_5[3599:3592];
        layer1[3][23:16] = buffer_data_5[3607:3600];
        layer1[3][31:24] = buffer_data_5[3615:3608];
        layer1[3][39:32] = buffer_data_5[3623:3616];
        layer1[3][47:40] = buffer_data_5[3631:3624];
        layer1[3][55:48] = buffer_data_5[3639:3632];
        layer2[3][7:0] = buffer_data_4[3591:3584];
        layer2[3][15:8] = buffer_data_4[3599:3592];
        layer2[3][23:16] = buffer_data_4[3607:3600];
        layer2[3][31:24] = buffer_data_4[3615:3608];
        layer2[3][39:32] = buffer_data_4[3623:3616];
        layer2[3][47:40] = buffer_data_4[3631:3624];
        layer2[3][55:48] = buffer_data_4[3639:3632];
        layer3[3][7:0] = buffer_data_3[3591:3584];
        layer3[3][15:8] = buffer_data_3[3599:3592];
        layer3[3][23:16] = buffer_data_3[3607:3600];
        layer3[3][31:24] = buffer_data_3[3615:3608];
        layer3[3][39:32] = buffer_data_3[3623:3616];
        layer3[3][47:40] = buffer_data_3[3631:3624];
        layer3[3][55:48] = buffer_data_3[3639:3632];
        layer4[3][7:0] = buffer_data_2[3591:3584];
        layer4[3][15:8] = buffer_data_2[3599:3592];
        layer4[3][23:16] = buffer_data_2[3607:3600];
        layer4[3][31:24] = buffer_data_2[3615:3608];
        layer4[3][39:32] = buffer_data_2[3623:3616];
        layer4[3][47:40] = buffer_data_2[3631:3624];
        layer4[3][55:48] = buffer_data_2[3639:3632];
        layer5[3][7:0] = buffer_data_1[3591:3584];
        layer5[3][15:8] = buffer_data_1[3599:3592];
        layer5[3][23:16] = buffer_data_1[3607:3600];
        layer5[3][31:24] = buffer_data_1[3615:3608];
        layer5[3][39:32] = buffer_data_1[3623:3616];
        layer5[3][47:40] = buffer_data_1[3631:3624];
        layer5[3][55:48] = buffer_data_1[3639:3632];
        layer6[3][7:0] = buffer_data_0[3591:3584];
        layer6[3][15:8] = buffer_data_0[3599:3592];
        layer6[3][23:16] = buffer_data_0[3607:3600];
        layer6[3][31:24] = buffer_data_0[3615:3608];
        layer6[3][39:32] = buffer_data_0[3623:3616];
        layer6[3][47:40] = buffer_data_0[3631:3624];
        layer6[3][55:48] = buffer_data_0[3639:3632];
        layer0[4][7:0] = buffer_data_6[3599:3592];
        layer0[4][15:8] = buffer_data_6[3607:3600];
        layer0[4][23:16] = buffer_data_6[3615:3608];
        layer0[4][31:24] = buffer_data_6[3623:3616];
        layer0[4][39:32] = buffer_data_6[3631:3624];
        layer0[4][47:40] = buffer_data_6[3639:3632];
        layer0[4][55:48] = buffer_data_6[3647:3640];
        layer1[4][7:0] = buffer_data_5[3599:3592];
        layer1[4][15:8] = buffer_data_5[3607:3600];
        layer1[4][23:16] = buffer_data_5[3615:3608];
        layer1[4][31:24] = buffer_data_5[3623:3616];
        layer1[4][39:32] = buffer_data_5[3631:3624];
        layer1[4][47:40] = buffer_data_5[3639:3632];
        layer1[4][55:48] = buffer_data_5[3647:3640];
        layer2[4][7:0] = buffer_data_4[3599:3592];
        layer2[4][15:8] = buffer_data_4[3607:3600];
        layer2[4][23:16] = buffer_data_4[3615:3608];
        layer2[4][31:24] = buffer_data_4[3623:3616];
        layer2[4][39:32] = buffer_data_4[3631:3624];
        layer2[4][47:40] = buffer_data_4[3639:3632];
        layer2[4][55:48] = buffer_data_4[3647:3640];
        layer3[4][7:0] = buffer_data_3[3599:3592];
        layer3[4][15:8] = buffer_data_3[3607:3600];
        layer3[4][23:16] = buffer_data_3[3615:3608];
        layer3[4][31:24] = buffer_data_3[3623:3616];
        layer3[4][39:32] = buffer_data_3[3631:3624];
        layer3[4][47:40] = buffer_data_3[3639:3632];
        layer3[4][55:48] = buffer_data_3[3647:3640];
        layer4[4][7:0] = buffer_data_2[3599:3592];
        layer4[4][15:8] = buffer_data_2[3607:3600];
        layer4[4][23:16] = buffer_data_2[3615:3608];
        layer4[4][31:24] = buffer_data_2[3623:3616];
        layer4[4][39:32] = buffer_data_2[3631:3624];
        layer4[4][47:40] = buffer_data_2[3639:3632];
        layer4[4][55:48] = buffer_data_2[3647:3640];
        layer5[4][7:0] = buffer_data_1[3599:3592];
        layer5[4][15:8] = buffer_data_1[3607:3600];
        layer5[4][23:16] = buffer_data_1[3615:3608];
        layer5[4][31:24] = buffer_data_1[3623:3616];
        layer5[4][39:32] = buffer_data_1[3631:3624];
        layer5[4][47:40] = buffer_data_1[3639:3632];
        layer5[4][55:48] = buffer_data_1[3647:3640];
        layer6[4][7:0] = buffer_data_0[3599:3592];
        layer6[4][15:8] = buffer_data_0[3607:3600];
        layer6[4][23:16] = buffer_data_0[3615:3608];
        layer6[4][31:24] = buffer_data_0[3623:3616];
        layer6[4][39:32] = buffer_data_0[3631:3624];
        layer6[4][47:40] = buffer_data_0[3639:3632];
        layer6[4][55:48] = buffer_data_0[3647:3640];
        layer0[5][7:0] = buffer_data_6[3607:3600];
        layer0[5][15:8] = buffer_data_6[3615:3608];
        layer0[5][23:16] = buffer_data_6[3623:3616];
        layer0[5][31:24] = buffer_data_6[3631:3624];
        layer0[5][39:32] = buffer_data_6[3639:3632];
        layer0[5][47:40] = buffer_data_6[3647:3640];
        layer0[5][55:48] = buffer_data_6[3655:3648];
        layer1[5][7:0] = buffer_data_5[3607:3600];
        layer1[5][15:8] = buffer_data_5[3615:3608];
        layer1[5][23:16] = buffer_data_5[3623:3616];
        layer1[5][31:24] = buffer_data_5[3631:3624];
        layer1[5][39:32] = buffer_data_5[3639:3632];
        layer1[5][47:40] = buffer_data_5[3647:3640];
        layer1[5][55:48] = buffer_data_5[3655:3648];
        layer2[5][7:0] = buffer_data_4[3607:3600];
        layer2[5][15:8] = buffer_data_4[3615:3608];
        layer2[5][23:16] = buffer_data_4[3623:3616];
        layer2[5][31:24] = buffer_data_4[3631:3624];
        layer2[5][39:32] = buffer_data_4[3639:3632];
        layer2[5][47:40] = buffer_data_4[3647:3640];
        layer2[5][55:48] = buffer_data_4[3655:3648];
        layer3[5][7:0] = buffer_data_3[3607:3600];
        layer3[5][15:8] = buffer_data_3[3615:3608];
        layer3[5][23:16] = buffer_data_3[3623:3616];
        layer3[5][31:24] = buffer_data_3[3631:3624];
        layer3[5][39:32] = buffer_data_3[3639:3632];
        layer3[5][47:40] = buffer_data_3[3647:3640];
        layer3[5][55:48] = buffer_data_3[3655:3648];
        layer4[5][7:0] = buffer_data_2[3607:3600];
        layer4[5][15:8] = buffer_data_2[3615:3608];
        layer4[5][23:16] = buffer_data_2[3623:3616];
        layer4[5][31:24] = buffer_data_2[3631:3624];
        layer4[5][39:32] = buffer_data_2[3639:3632];
        layer4[5][47:40] = buffer_data_2[3647:3640];
        layer4[5][55:48] = buffer_data_2[3655:3648];
        layer5[5][7:0] = buffer_data_1[3607:3600];
        layer5[5][15:8] = buffer_data_1[3615:3608];
        layer5[5][23:16] = buffer_data_1[3623:3616];
        layer5[5][31:24] = buffer_data_1[3631:3624];
        layer5[5][39:32] = buffer_data_1[3639:3632];
        layer5[5][47:40] = buffer_data_1[3647:3640];
        layer5[5][55:48] = buffer_data_1[3655:3648];
        layer6[5][7:0] = buffer_data_0[3607:3600];
        layer6[5][15:8] = buffer_data_0[3615:3608];
        layer6[5][23:16] = buffer_data_0[3623:3616];
        layer6[5][31:24] = buffer_data_0[3631:3624];
        layer6[5][39:32] = buffer_data_0[3639:3632];
        layer6[5][47:40] = buffer_data_0[3647:3640];
        layer6[5][55:48] = buffer_data_0[3655:3648];
        layer0[6][7:0] = buffer_data_6[3615:3608];
        layer0[6][15:8] = buffer_data_6[3623:3616];
        layer0[6][23:16] = buffer_data_6[3631:3624];
        layer0[6][31:24] = buffer_data_6[3639:3632];
        layer0[6][39:32] = buffer_data_6[3647:3640];
        layer0[6][47:40] = buffer_data_6[3655:3648];
        layer0[6][55:48] = buffer_data_6[3663:3656];
        layer1[6][7:0] = buffer_data_5[3615:3608];
        layer1[6][15:8] = buffer_data_5[3623:3616];
        layer1[6][23:16] = buffer_data_5[3631:3624];
        layer1[6][31:24] = buffer_data_5[3639:3632];
        layer1[6][39:32] = buffer_data_5[3647:3640];
        layer1[6][47:40] = buffer_data_5[3655:3648];
        layer1[6][55:48] = buffer_data_5[3663:3656];
        layer2[6][7:0] = buffer_data_4[3615:3608];
        layer2[6][15:8] = buffer_data_4[3623:3616];
        layer2[6][23:16] = buffer_data_4[3631:3624];
        layer2[6][31:24] = buffer_data_4[3639:3632];
        layer2[6][39:32] = buffer_data_4[3647:3640];
        layer2[6][47:40] = buffer_data_4[3655:3648];
        layer2[6][55:48] = buffer_data_4[3663:3656];
        layer3[6][7:0] = buffer_data_3[3615:3608];
        layer3[6][15:8] = buffer_data_3[3623:3616];
        layer3[6][23:16] = buffer_data_3[3631:3624];
        layer3[6][31:24] = buffer_data_3[3639:3632];
        layer3[6][39:32] = buffer_data_3[3647:3640];
        layer3[6][47:40] = buffer_data_3[3655:3648];
        layer3[6][55:48] = buffer_data_3[3663:3656];
        layer4[6][7:0] = buffer_data_2[3615:3608];
        layer4[6][15:8] = buffer_data_2[3623:3616];
        layer4[6][23:16] = buffer_data_2[3631:3624];
        layer4[6][31:24] = buffer_data_2[3639:3632];
        layer4[6][39:32] = buffer_data_2[3647:3640];
        layer4[6][47:40] = buffer_data_2[3655:3648];
        layer4[6][55:48] = buffer_data_2[3663:3656];
        layer5[6][7:0] = buffer_data_1[3615:3608];
        layer5[6][15:8] = buffer_data_1[3623:3616];
        layer5[6][23:16] = buffer_data_1[3631:3624];
        layer5[6][31:24] = buffer_data_1[3639:3632];
        layer5[6][39:32] = buffer_data_1[3647:3640];
        layer5[6][47:40] = buffer_data_1[3655:3648];
        layer5[6][55:48] = buffer_data_1[3663:3656];
        layer6[6][7:0] = buffer_data_0[3615:3608];
        layer6[6][15:8] = buffer_data_0[3623:3616];
        layer6[6][23:16] = buffer_data_0[3631:3624];
        layer6[6][31:24] = buffer_data_0[3639:3632];
        layer6[6][39:32] = buffer_data_0[3647:3640];
        layer6[6][47:40] = buffer_data_0[3655:3648];
        layer6[6][55:48] = buffer_data_0[3663:3656];
        layer0[7][7:0] = buffer_data_6[3623:3616];
        layer0[7][15:8] = buffer_data_6[3631:3624];
        layer0[7][23:16] = buffer_data_6[3639:3632];
        layer0[7][31:24] = buffer_data_6[3647:3640];
        layer0[7][39:32] = buffer_data_6[3655:3648];
        layer0[7][47:40] = buffer_data_6[3663:3656];
        layer0[7][55:48] = buffer_data_6[3671:3664];
        layer1[7][7:0] = buffer_data_5[3623:3616];
        layer1[7][15:8] = buffer_data_5[3631:3624];
        layer1[7][23:16] = buffer_data_5[3639:3632];
        layer1[7][31:24] = buffer_data_5[3647:3640];
        layer1[7][39:32] = buffer_data_5[3655:3648];
        layer1[7][47:40] = buffer_data_5[3663:3656];
        layer1[7][55:48] = buffer_data_5[3671:3664];
        layer2[7][7:0] = buffer_data_4[3623:3616];
        layer2[7][15:8] = buffer_data_4[3631:3624];
        layer2[7][23:16] = buffer_data_4[3639:3632];
        layer2[7][31:24] = buffer_data_4[3647:3640];
        layer2[7][39:32] = buffer_data_4[3655:3648];
        layer2[7][47:40] = buffer_data_4[3663:3656];
        layer2[7][55:48] = buffer_data_4[3671:3664];
        layer3[7][7:0] = buffer_data_3[3623:3616];
        layer3[7][15:8] = buffer_data_3[3631:3624];
        layer3[7][23:16] = buffer_data_3[3639:3632];
        layer3[7][31:24] = buffer_data_3[3647:3640];
        layer3[7][39:32] = buffer_data_3[3655:3648];
        layer3[7][47:40] = buffer_data_3[3663:3656];
        layer3[7][55:48] = buffer_data_3[3671:3664];
        layer4[7][7:0] = buffer_data_2[3623:3616];
        layer4[7][15:8] = buffer_data_2[3631:3624];
        layer4[7][23:16] = buffer_data_2[3639:3632];
        layer4[7][31:24] = buffer_data_2[3647:3640];
        layer4[7][39:32] = buffer_data_2[3655:3648];
        layer4[7][47:40] = buffer_data_2[3663:3656];
        layer4[7][55:48] = buffer_data_2[3671:3664];
        layer5[7][7:0] = buffer_data_1[3623:3616];
        layer5[7][15:8] = buffer_data_1[3631:3624];
        layer5[7][23:16] = buffer_data_1[3639:3632];
        layer5[7][31:24] = buffer_data_1[3647:3640];
        layer5[7][39:32] = buffer_data_1[3655:3648];
        layer5[7][47:40] = buffer_data_1[3663:3656];
        layer5[7][55:48] = buffer_data_1[3671:3664];
        layer6[7][7:0] = buffer_data_0[3623:3616];
        layer6[7][15:8] = buffer_data_0[3631:3624];
        layer6[7][23:16] = buffer_data_0[3639:3632];
        layer6[7][31:24] = buffer_data_0[3647:3640];
        layer6[7][39:32] = buffer_data_0[3655:3648];
        layer6[7][47:40] = buffer_data_0[3663:3656];
        layer6[7][55:48] = buffer_data_0[3671:3664];
        layer0[8][7:0] = buffer_data_6[3631:3624];
        layer0[8][15:8] = buffer_data_6[3639:3632];
        layer0[8][23:16] = buffer_data_6[3647:3640];
        layer0[8][31:24] = buffer_data_6[3655:3648];
        layer0[8][39:32] = buffer_data_6[3663:3656];
        layer0[8][47:40] = buffer_data_6[3671:3664];
        layer0[8][55:48] = buffer_data_6[3679:3672];
        layer1[8][7:0] = buffer_data_5[3631:3624];
        layer1[8][15:8] = buffer_data_5[3639:3632];
        layer1[8][23:16] = buffer_data_5[3647:3640];
        layer1[8][31:24] = buffer_data_5[3655:3648];
        layer1[8][39:32] = buffer_data_5[3663:3656];
        layer1[8][47:40] = buffer_data_5[3671:3664];
        layer1[8][55:48] = buffer_data_5[3679:3672];
        layer2[8][7:0] = buffer_data_4[3631:3624];
        layer2[8][15:8] = buffer_data_4[3639:3632];
        layer2[8][23:16] = buffer_data_4[3647:3640];
        layer2[8][31:24] = buffer_data_4[3655:3648];
        layer2[8][39:32] = buffer_data_4[3663:3656];
        layer2[8][47:40] = buffer_data_4[3671:3664];
        layer2[8][55:48] = buffer_data_4[3679:3672];
        layer3[8][7:0] = buffer_data_3[3631:3624];
        layer3[8][15:8] = buffer_data_3[3639:3632];
        layer3[8][23:16] = buffer_data_3[3647:3640];
        layer3[8][31:24] = buffer_data_3[3655:3648];
        layer3[8][39:32] = buffer_data_3[3663:3656];
        layer3[8][47:40] = buffer_data_3[3671:3664];
        layer3[8][55:48] = buffer_data_3[3679:3672];
        layer4[8][7:0] = buffer_data_2[3631:3624];
        layer4[8][15:8] = buffer_data_2[3639:3632];
        layer4[8][23:16] = buffer_data_2[3647:3640];
        layer4[8][31:24] = buffer_data_2[3655:3648];
        layer4[8][39:32] = buffer_data_2[3663:3656];
        layer4[8][47:40] = buffer_data_2[3671:3664];
        layer4[8][55:48] = buffer_data_2[3679:3672];
        layer5[8][7:0] = buffer_data_1[3631:3624];
        layer5[8][15:8] = buffer_data_1[3639:3632];
        layer5[8][23:16] = buffer_data_1[3647:3640];
        layer5[8][31:24] = buffer_data_1[3655:3648];
        layer5[8][39:32] = buffer_data_1[3663:3656];
        layer5[8][47:40] = buffer_data_1[3671:3664];
        layer5[8][55:48] = buffer_data_1[3679:3672];
        layer6[8][7:0] = buffer_data_0[3631:3624];
        layer6[8][15:8] = buffer_data_0[3639:3632];
        layer6[8][23:16] = buffer_data_0[3647:3640];
        layer6[8][31:24] = buffer_data_0[3655:3648];
        layer6[8][39:32] = buffer_data_0[3663:3656];
        layer6[8][47:40] = buffer_data_0[3671:3664];
        layer6[8][55:48] = buffer_data_0[3679:3672];
        layer0[9][7:0] = buffer_data_6[3639:3632];
        layer0[9][15:8] = buffer_data_6[3647:3640];
        layer0[9][23:16] = buffer_data_6[3655:3648];
        layer0[9][31:24] = buffer_data_6[3663:3656];
        layer0[9][39:32] = buffer_data_6[3671:3664];
        layer0[9][47:40] = buffer_data_6[3679:3672];
        layer0[9][55:48] = buffer_data_6[3687:3680];
        layer1[9][7:0] = buffer_data_5[3639:3632];
        layer1[9][15:8] = buffer_data_5[3647:3640];
        layer1[9][23:16] = buffer_data_5[3655:3648];
        layer1[9][31:24] = buffer_data_5[3663:3656];
        layer1[9][39:32] = buffer_data_5[3671:3664];
        layer1[9][47:40] = buffer_data_5[3679:3672];
        layer1[9][55:48] = buffer_data_5[3687:3680];
        layer2[9][7:0] = buffer_data_4[3639:3632];
        layer2[9][15:8] = buffer_data_4[3647:3640];
        layer2[9][23:16] = buffer_data_4[3655:3648];
        layer2[9][31:24] = buffer_data_4[3663:3656];
        layer2[9][39:32] = buffer_data_4[3671:3664];
        layer2[9][47:40] = buffer_data_4[3679:3672];
        layer2[9][55:48] = buffer_data_4[3687:3680];
        layer3[9][7:0] = buffer_data_3[3639:3632];
        layer3[9][15:8] = buffer_data_3[3647:3640];
        layer3[9][23:16] = buffer_data_3[3655:3648];
        layer3[9][31:24] = buffer_data_3[3663:3656];
        layer3[9][39:32] = buffer_data_3[3671:3664];
        layer3[9][47:40] = buffer_data_3[3679:3672];
        layer3[9][55:48] = buffer_data_3[3687:3680];
        layer4[9][7:0] = buffer_data_2[3639:3632];
        layer4[9][15:8] = buffer_data_2[3647:3640];
        layer4[9][23:16] = buffer_data_2[3655:3648];
        layer4[9][31:24] = buffer_data_2[3663:3656];
        layer4[9][39:32] = buffer_data_2[3671:3664];
        layer4[9][47:40] = buffer_data_2[3679:3672];
        layer4[9][55:48] = buffer_data_2[3687:3680];
        layer5[9][7:0] = buffer_data_1[3639:3632];
        layer5[9][15:8] = buffer_data_1[3647:3640];
        layer5[9][23:16] = buffer_data_1[3655:3648];
        layer5[9][31:24] = buffer_data_1[3663:3656];
        layer5[9][39:32] = buffer_data_1[3671:3664];
        layer5[9][47:40] = buffer_data_1[3679:3672];
        layer5[9][55:48] = buffer_data_1[3687:3680];
        layer6[9][7:0] = buffer_data_0[3639:3632];
        layer6[9][15:8] = buffer_data_0[3647:3640];
        layer6[9][23:16] = buffer_data_0[3655:3648];
        layer6[9][31:24] = buffer_data_0[3663:3656];
        layer6[9][39:32] = buffer_data_0[3671:3664];
        layer6[9][47:40] = buffer_data_0[3679:3672];
        layer6[9][55:48] = buffer_data_0[3687:3680];
        layer0[10][7:0] = buffer_data_6[3647:3640];
        layer0[10][15:8] = buffer_data_6[3655:3648];
        layer0[10][23:16] = buffer_data_6[3663:3656];
        layer0[10][31:24] = buffer_data_6[3671:3664];
        layer0[10][39:32] = buffer_data_6[3679:3672];
        layer0[10][47:40] = buffer_data_6[3687:3680];
        layer0[10][55:48] = buffer_data_6[3695:3688];
        layer1[10][7:0] = buffer_data_5[3647:3640];
        layer1[10][15:8] = buffer_data_5[3655:3648];
        layer1[10][23:16] = buffer_data_5[3663:3656];
        layer1[10][31:24] = buffer_data_5[3671:3664];
        layer1[10][39:32] = buffer_data_5[3679:3672];
        layer1[10][47:40] = buffer_data_5[3687:3680];
        layer1[10][55:48] = buffer_data_5[3695:3688];
        layer2[10][7:0] = buffer_data_4[3647:3640];
        layer2[10][15:8] = buffer_data_4[3655:3648];
        layer2[10][23:16] = buffer_data_4[3663:3656];
        layer2[10][31:24] = buffer_data_4[3671:3664];
        layer2[10][39:32] = buffer_data_4[3679:3672];
        layer2[10][47:40] = buffer_data_4[3687:3680];
        layer2[10][55:48] = buffer_data_4[3695:3688];
        layer3[10][7:0] = buffer_data_3[3647:3640];
        layer3[10][15:8] = buffer_data_3[3655:3648];
        layer3[10][23:16] = buffer_data_3[3663:3656];
        layer3[10][31:24] = buffer_data_3[3671:3664];
        layer3[10][39:32] = buffer_data_3[3679:3672];
        layer3[10][47:40] = buffer_data_3[3687:3680];
        layer3[10][55:48] = buffer_data_3[3695:3688];
        layer4[10][7:0] = buffer_data_2[3647:3640];
        layer4[10][15:8] = buffer_data_2[3655:3648];
        layer4[10][23:16] = buffer_data_2[3663:3656];
        layer4[10][31:24] = buffer_data_2[3671:3664];
        layer4[10][39:32] = buffer_data_2[3679:3672];
        layer4[10][47:40] = buffer_data_2[3687:3680];
        layer4[10][55:48] = buffer_data_2[3695:3688];
        layer5[10][7:0] = buffer_data_1[3647:3640];
        layer5[10][15:8] = buffer_data_1[3655:3648];
        layer5[10][23:16] = buffer_data_1[3663:3656];
        layer5[10][31:24] = buffer_data_1[3671:3664];
        layer5[10][39:32] = buffer_data_1[3679:3672];
        layer5[10][47:40] = buffer_data_1[3687:3680];
        layer5[10][55:48] = buffer_data_1[3695:3688];
        layer6[10][7:0] = buffer_data_0[3647:3640];
        layer6[10][15:8] = buffer_data_0[3655:3648];
        layer6[10][23:16] = buffer_data_0[3663:3656];
        layer6[10][31:24] = buffer_data_0[3671:3664];
        layer6[10][39:32] = buffer_data_0[3679:3672];
        layer6[10][47:40] = buffer_data_0[3687:3680];
        layer6[10][55:48] = buffer_data_0[3695:3688];
        layer0[11][7:0] = buffer_data_6[3655:3648];
        layer0[11][15:8] = buffer_data_6[3663:3656];
        layer0[11][23:16] = buffer_data_6[3671:3664];
        layer0[11][31:24] = buffer_data_6[3679:3672];
        layer0[11][39:32] = buffer_data_6[3687:3680];
        layer0[11][47:40] = buffer_data_6[3695:3688];
        layer0[11][55:48] = buffer_data_6[3703:3696];
        layer1[11][7:0] = buffer_data_5[3655:3648];
        layer1[11][15:8] = buffer_data_5[3663:3656];
        layer1[11][23:16] = buffer_data_5[3671:3664];
        layer1[11][31:24] = buffer_data_5[3679:3672];
        layer1[11][39:32] = buffer_data_5[3687:3680];
        layer1[11][47:40] = buffer_data_5[3695:3688];
        layer1[11][55:48] = buffer_data_5[3703:3696];
        layer2[11][7:0] = buffer_data_4[3655:3648];
        layer2[11][15:8] = buffer_data_4[3663:3656];
        layer2[11][23:16] = buffer_data_4[3671:3664];
        layer2[11][31:24] = buffer_data_4[3679:3672];
        layer2[11][39:32] = buffer_data_4[3687:3680];
        layer2[11][47:40] = buffer_data_4[3695:3688];
        layer2[11][55:48] = buffer_data_4[3703:3696];
        layer3[11][7:0] = buffer_data_3[3655:3648];
        layer3[11][15:8] = buffer_data_3[3663:3656];
        layer3[11][23:16] = buffer_data_3[3671:3664];
        layer3[11][31:24] = buffer_data_3[3679:3672];
        layer3[11][39:32] = buffer_data_3[3687:3680];
        layer3[11][47:40] = buffer_data_3[3695:3688];
        layer3[11][55:48] = buffer_data_3[3703:3696];
        layer4[11][7:0] = buffer_data_2[3655:3648];
        layer4[11][15:8] = buffer_data_2[3663:3656];
        layer4[11][23:16] = buffer_data_2[3671:3664];
        layer4[11][31:24] = buffer_data_2[3679:3672];
        layer4[11][39:32] = buffer_data_2[3687:3680];
        layer4[11][47:40] = buffer_data_2[3695:3688];
        layer4[11][55:48] = buffer_data_2[3703:3696];
        layer5[11][7:0] = buffer_data_1[3655:3648];
        layer5[11][15:8] = buffer_data_1[3663:3656];
        layer5[11][23:16] = buffer_data_1[3671:3664];
        layer5[11][31:24] = buffer_data_1[3679:3672];
        layer5[11][39:32] = buffer_data_1[3687:3680];
        layer5[11][47:40] = buffer_data_1[3695:3688];
        layer5[11][55:48] = buffer_data_1[3703:3696];
        layer6[11][7:0] = buffer_data_0[3655:3648];
        layer6[11][15:8] = buffer_data_0[3663:3656];
        layer6[11][23:16] = buffer_data_0[3671:3664];
        layer6[11][31:24] = buffer_data_0[3679:3672];
        layer6[11][39:32] = buffer_data_0[3687:3680];
        layer6[11][47:40] = buffer_data_0[3695:3688];
        layer6[11][55:48] = buffer_data_0[3703:3696];
        layer0[12][7:0] = buffer_data_6[3663:3656];
        layer0[12][15:8] = buffer_data_6[3671:3664];
        layer0[12][23:16] = buffer_data_6[3679:3672];
        layer0[12][31:24] = buffer_data_6[3687:3680];
        layer0[12][39:32] = buffer_data_6[3695:3688];
        layer0[12][47:40] = buffer_data_6[3703:3696];
        layer0[12][55:48] = buffer_data_6[3711:3704];
        layer1[12][7:0] = buffer_data_5[3663:3656];
        layer1[12][15:8] = buffer_data_5[3671:3664];
        layer1[12][23:16] = buffer_data_5[3679:3672];
        layer1[12][31:24] = buffer_data_5[3687:3680];
        layer1[12][39:32] = buffer_data_5[3695:3688];
        layer1[12][47:40] = buffer_data_5[3703:3696];
        layer1[12][55:48] = buffer_data_5[3711:3704];
        layer2[12][7:0] = buffer_data_4[3663:3656];
        layer2[12][15:8] = buffer_data_4[3671:3664];
        layer2[12][23:16] = buffer_data_4[3679:3672];
        layer2[12][31:24] = buffer_data_4[3687:3680];
        layer2[12][39:32] = buffer_data_4[3695:3688];
        layer2[12][47:40] = buffer_data_4[3703:3696];
        layer2[12][55:48] = buffer_data_4[3711:3704];
        layer3[12][7:0] = buffer_data_3[3663:3656];
        layer3[12][15:8] = buffer_data_3[3671:3664];
        layer3[12][23:16] = buffer_data_3[3679:3672];
        layer3[12][31:24] = buffer_data_3[3687:3680];
        layer3[12][39:32] = buffer_data_3[3695:3688];
        layer3[12][47:40] = buffer_data_3[3703:3696];
        layer3[12][55:48] = buffer_data_3[3711:3704];
        layer4[12][7:0] = buffer_data_2[3663:3656];
        layer4[12][15:8] = buffer_data_2[3671:3664];
        layer4[12][23:16] = buffer_data_2[3679:3672];
        layer4[12][31:24] = buffer_data_2[3687:3680];
        layer4[12][39:32] = buffer_data_2[3695:3688];
        layer4[12][47:40] = buffer_data_2[3703:3696];
        layer4[12][55:48] = buffer_data_2[3711:3704];
        layer5[12][7:0] = buffer_data_1[3663:3656];
        layer5[12][15:8] = buffer_data_1[3671:3664];
        layer5[12][23:16] = buffer_data_1[3679:3672];
        layer5[12][31:24] = buffer_data_1[3687:3680];
        layer5[12][39:32] = buffer_data_1[3695:3688];
        layer5[12][47:40] = buffer_data_1[3703:3696];
        layer5[12][55:48] = buffer_data_1[3711:3704];
        layer6[12][7:0] = buffer_data_0[3663:3656];
        layer6[12][15:8] = buffer_data_0[3671:3664];
        layer6[12][23:16] = buffer_data_0[3679:3672];
        layer6[12][31:24] = buffer_data_0[3687:3680];
        layer6[12][39:32] = buffer_data_0[3695:3688];
        layer6[12][47:40] = buffer_data_0[3703:3696];
        layer6[12][55:48] = buffer_data_0[3711:3704];
        layer0[13][7:0] = buffer_data_6[3671:3664];
        layer0[13][15:8] = buffer_data_6[3679:3672];
        layer0[13][23:16] = buffer_data_6[3687:3680];
        layer0[13][31:24] = buffer_data_6[3695:3688];
        layer0[13][39:32] = buffer_data_6[3703:3696];
        layer0[13][47:40] = buffer_data_6[3711:3704];
        layer0[13][55:48] = buffer_data_6[3719:3712];
        layer1[13][7:0] = buffer_data_5[3671:3664];
        layer1[13][15:8] = buffer_data_5[3679:3672];
        layer1[13][23:16] = buffer_data_5[3687:3680];
        layer1[13][31:24] = buffer_data_5[3695:3688];
        layer1[13][39:32] = buffer_data_5[3703:3696];
        layer1[13][47:40] = buffer_data_5[3711:3704];
        layer1[13][55:48] = buffer_data_5[3719:3712];
        layer2[13][7:0] = buffer_data_4[3671:3664];
        layer2[13][15:8] = buffer_data_4[3679:3672];
        layer2[13][23:16] = buffer_data_4[3687:3680];
        layer2[13][31:24] = buffer_data_4[3695:3688];
        layer2[13][39:32] = buffer_data_4[3703:3696];
        layer2[13][47:40] = buffer_data_4[3711:3704];
        layer2[13][55:48] = buffer_data_4[3719:3712];
        layer3[13][7:0] = buffer_data_3[3671:3664];
        layer3[13][15:8] = buffer_data_3[3679:3672];
        layer3[13][23:16] = buffer_data_3[3687:3680];
        layer3[13][31:24] = buffer_data_3[3695:3688];
        layer3[13][39:32] = buffer_data_3[3703:3696];
        layer3[13][47:40] = buffer_data_3[3711:3704];
        layer3[13][55:48] = buffer_data_3[3719:3712];
        layer4[13][7:0] = buffer_data_2[3671:3664];
        layer4[13][15:8] = buffer_data_2[3679:3672];
        layer4[13][23:16] = buffer_data_2[3687:3680];
        layer4[13][31:24] = buffer_data_2[3695:3688];
        layer4[13][39:32] = buffer_data_2[3703:3696];
        layer4[13][47:40] = buffer_data_2[3711:3704];
        layer4[13][55:48] = buffer_data_2[3719:3712];
        layer5[13][7:0] = buffer_data_1[3671:3664];
        layer5[13][15:8] = buffer_data_1[3679:3672];
        layer5[13][23:16] = buffer_data_1[3687:3680];
        layer5[13][31:24] = buffer_data_1[3695:3688];
        layer5[13][39:32] = buffer_data_1[3703:3696];
        layer5[13][47:40] = buffer_data_1[3711:3704];
        layer5[13][55:48] = buffer_data_1[3719:3712];
        layer6[13][7:0] = buffer_data_0[3671:3664];
        layer6[13][15:8] = buffer_data_0[3679:3672];
        layer6[13][23:16] = buffer_data_0[3687:3680];
        layer6[13][31:24] = buffer_data_0[3695:3688];
        layer6[13][39:32] = buffer_data_0[3703:3696];
        layer6[13][47:40] = buffer_data_0[3711:3704];
        layer6[13][55:48] = buffer_data_0[3719:3712];
        layer0[14][7:0] = buffer_data_6[3679:3672];
        layer0[14][15:8] = buffer_data_6[3687:3680];
        layer0[14][23:16] = buffer_data_6[3695:3688];
        layer0[14][31:24] = buffer_data_6[3703:3696];
        layer0[14][39:32] = buffer_data_6[3711:3704];
        layer0[14][47:40] = buffer_data_6[3719:3712];
        layer0[14][55:48] = buffer_data_6[3727:3720];
        layer1[14][7:0] = buffer_data_5[3679:3672];
        layer1[14][15:8] = buffer_data_5[3687:3680];
        layer1[14][23:16] = buffer_data_5[3695:3688];
        layer1[14][31:24] = buffer_data_5[3703:3696];
        layer1[14][39:32] = buffer_data_5[3711:3704];
        layer1[14][47:40] = buffer_data_5[3719:3712];
        layer1[14][55:48] = buffer_data_5[3727:3720];
        layer2[14][7:0] = buffer_data_4[3679:3672];
        layer2[14][15:8] = buffer_data_4[3687:3680];
        layer2[14][23:16] = buffer_data_4[3695:3688];
        layer2[14][31:24] = buffer_data_4[3703:3696];
        layer2[14][39:32] = buffer_data_4[3711:3704];
        layer2[14][47:40] = buffer_data_4[3719:3712];
        layer2[14][55:48] = buffer_data_4[3727:3720];
        layer3[14][7:0] = buffer_data_3[3679:3672];
        layer3[14][15:8] = buffer_data_3[3687:3680];
        layer3[14][23:16] = buffer_data_3[3695:3688];
        layer3[14][31:24] = buffer_data_3[3703:3696];
        layer3[14][39:32] = buffer_data_3[3711:3704];
        layer3[14][47:40] = buffer_data_3[3719:3712];
        layer3[14][55:48] = buffer_data_3[3727:3720];
        layer4[14][7:0] = buffer_data_2[3679:3672];
        layer4[14][15:8] = buffer_data_2[3687:3680];
        layer4[14][23:16] = buffer_data_2[3695:3688];
        layer4[14][31:24] = buffer_data_2[3703:3696];
        layer4[14][39:32] = buffer_data_2[3711:3704];
        layer4[14][47:40] = buffer_data_2[3719:3712];
        layer4[14][55:48] = buffer_data_2[3727:3720];
        layer5[14][7:0] = buffer_data_1[3679:3672];
        layer5[14][15:8] = buffer_data_1[3687:3680];
        layer5[14][23:16] = buffer_data_1[3695:3688];
        layer5[14][31:24] = buffer_data_1[3703:3696];
        layer5[14][39:32] = buffer_data_1[3711:3704];
        layer5[14][47:40] = buffer_data_1[3719:3712];
        layer5[14][55:48] = buffer_data_1[3727:3720];
        layer6[14][7:0] = buffer_data_0[3679:3672];
        layer6[14][15:8] = buffer_data_0[3687:3680];
        layer6[14][23:16] = buffer_data_0[3695:3688];
        layer6[14][31:24] = buffer_data_0[3703:3696];
        layer6[14][39:32] = buffer_data_0[3711:3704];
        layer6[14][47:40] = buffer_data_0[3719:3712];
        layer6[14][55:48] = buffer_data_0[3727:3720];
        layer0[15][7:0] = buffer_data_6[3687:3680];
        layer0[15][15:8] = buffer_data_6[3695:3688];
        layer0[15][23:16] = buffer_data_6[3703:3696];
        layer0[15][31:24] = buffer_data_6[3711:3704];
        layer0[15][39:32] = buffer_data_6[3719:3712];
        layer0[15][47:40] = buffer_data_6[3727:3720];
        layer0[15][55:48] = buffer_data_6[3735:3728];
        layer1[15][7:0] = buffer_data_5[3687:3680];
        layer1[15][15:8] = buffer_data_5[3695:3688];
        layer1[15][23:16] = buffer_data_5[3703:3696];
        layer1[15][31:24] = buffer_data_5[3711:3704];
        layer1[15][39:32] = buffer_data_5[3719:3712];
        layer1[15][47:40] = buffer_data_5[3727:3720];
        layer1[15][55:48] = buffer_data_5[3735:3728];
        layer2[15][7:0] = buffer_data_4[3687:3680];
        layer2[15][15:8] = buffer_data_4[3695:3688];
        layer2[15][23:16] = buffer_data_4[3703:3696];
        layer2[15][31:24] = buffer_data_4[3711:3704];
        layer2[15][39:32] = buffer_data_4[3719:3712];
        layer2[15][47:40] = buffer_data_4[3727:3720];
        layer2[15][55:48] = buffer_data_4[3735:3728];
        layer3[15][7:0] = buffer_data_3[3687:3680];
        layer3[15][15:8] = buffer_data_3[3695:3688];
        layer3[15][23:16] = buffer_data_3[3703:3696];
        layer3[15][31:24] = buffer_data_3[3711:3704];
        layer3[15][39:32] = buffer_data_3[3719:3712];
        layer3[15][47:40] = buffer_data_3[3727:3720];
        layer3[15][55:48] = buffer_data_3[3735:3728];
        layer4[15][7:0] = buffer_data_2[3687:3680];
        layer4[15][15:8] = buffer_data_2[3695:3688];
        layer4[15][23:16] = buffer_data_2[3703:3696];
        layer4[15][31:24] = buffer_data_2[3711:3704];
        layer4[15][39:32] = buffer_data_2[3719:3712];
        layer4[15][47:40] = buffer_data_2[3727:3720];
        layer4[15][55:48] = buffer_data_2[3735:3728];
        layer5[15][7:0] = buffer_data_1[3687:3680];
        layer5[15][15:8] = buffer_data_1[3695:3688];
        layer5[15][23:16] = buffer_data_1[3703:3696];
        layer5[15][31:24] = buffer_data_1[3711:3704];
        layer5[15][39:32] = buffer_data_1[3719:3712];
        layer5[15][47:40] = buffer_data_1[3727:3720];
        layer5[15][55:48] = buffer_data_1[3735:3728];
        layer6[15][7:0] = buffer_data_0[3687:3680];
        layer6[15][15:8] = buffer_data_0[3695:3688];
        layer6[15][23:16] = buffer_data_0[3703:3696];
        layer6[15][31:24] = buffer_data_0[3711:3704];
        layer6[15][39:32] = buffer_data_0[3719:3712];
        layer6[15][47:40] = buffer_data_0[3727:3720];
        layer6[15][55:48] = buffer_data_0[3735:3728];
        layer0[16][7:0] = buffer_data_6[3695:3688];
        layer0[16][15:8] = buffer_data_6[3703:3696];
        layer0[16][23:16] = buffer_data_6[3711:3704];
        layer0[16][31:24] = buffer_data_6[3719:3712];
        layer0[16][39:32] = buffer_data_6[3727:3720];
        layer0[16][47:40] = buffer_data_6[3735:3728];
        layer0[16][55:48] = buffer_data_6[3743:3736];
        layer1[16][7:0] = buffer_data_5[3695:3688];
        layer1[16][15:8] = buffer_data_5[3703:3696];
        layer1[16][23:16] = buffer_data_5[3711:3704];
        layer1[16][31:24] = buffer_data_5[3719:3712];
        layer1[16][39:32] = buffer_data_5[3727:3720];
        layer1[16][47:40] = buffer_data_5[3735:3728];
        layer1[16][55:48] = buffer_data_5[3743:3736];
        layer2[16][7:0] = buffer_data_4[3695:3688];
        layer2[16][15:8] = buffer_data_4[3703:3696];
        layer2[16][23:16] = buffer_data_4[3711:3704];
        layer2[16][31:24] = buffer_data_4[3719:3712];
        layer2[16][39:32] = buffer_data_4[3727:3720];
        layer2[16][47:40] = buffer_data_4[3735:3728];
        layer2[16][55:48] = buffer_data_4[3743:3736];
        layer3[16][7:0] = buffer_data_3[3695:3688];
        layer3[16][15:8] = buffer_data_3[3703:3696];
        layer3[16][23:16] = buffer_data_3[3711:3704];
        layer3[16][31:24] = buffer_data_3[3719:3712];
        layer3[16][39:32] = buffer_data_3[3727:3720];
        layer3[16][47:40] = buffer_data_3[3735:3728];
        layer3[16][55:48] = buffer_data_3[3743:3736];
        layer4[16][7:0] = buffer_data_2[3695:3688];
        layer4[16][15:8] = buffer_data_2[3703:3696];
        layer4[16][23:16] = buffer_data_2[3711:3704];
        layer4[16][31:24] = buffer_data_2[3719:3712];
        layer4[16][39:32] = buffer_data_2[3727:3720];
        layer4[16][47:40] = buffer_data_2[3735:3728];
        layer4[16][55:48] = buffer_data_2[3743:3736];
        layer5[16][7:0] = buffer_data_1[3695:3688];
        layer5[16][15:8] = buffer_data_1[3703:3696];
        layer5[16][23:16] = buffer_data_1[3711:3704];
        layer5[16][31:24] = buffer_data_1[3719:3712];
        layer5[16][39:32] = buffer_data_1[3727:3720];
        layer5[16][47:40] = buffer_data_1[3735:3728];
        layer5[16][55:48] = buffer_data_1[3743:3736];
        layer6[16][7:0] = buffer_data_0[3695:3688];
        layer6[16][15:8] = buffer_data_0[3703:3696];
        layer6[16][23:16] = buffer_data_0[3711:3704];
        layer6[16][31:24] = buffer_data_0[3719:3712];
        layer6[16][39:32] = buffer_data_0[3727:3720];
        layer6[16][47:40] = buffer_data_0[3735:3728];
        layer6[16][55:48] = buffer_data_0[3743:3736];
        layer0[17][7:0] = buffer_data_6[3703:3696];
        layer0[17][15:8] = buffer_data_6[3711:3704];
        layer0[17][23:16] = buffer_data_6[3719:3712];
        layer0[17][31:24] = buffer_data_6[3727:3720];
        layer0[17][39:32] = buffer_data_6[3735:3728];
        layer0[17][47:40] = buffer_data_6[3743:3736];
        layer0[17][55:48] = buffer_data_6[3751:3744];
        layer1[17][7:0] = buffer_data_5[3703:3696];
        layer1[17][15:8] = buffer_data_5[3711:3704];
        layer1[17][23:16] = buffer_data_5[3719:3712];
        layer1[17][31:24] = buffer_data_5[3727:3720];
        layer1[17][39:32] = buffer_data_5[3735:3728];
        layer1[17][47:40] = buffer_data_5[3743:3736];
        layer1[17][55:48] = buffer_data_5[3751:3744];
        layer2[17][7:0] = buffer_data_4[3703:3696];
        layer2[17][15:8] = buffer_data_4[3711:3704];
        layer2[17][23:16] = buffer_data_4[3719:3712];
        layer2[17][31:24] = buffer_data_4[3727:3720];
        layer2[17][39:32] = buffer_data_4[3735:3728];
        layer2[17][47:40] = buffer_data_4[3743:3736];
        layer2[17][55:48] = buffer_data_4[3751:3744];
        layer3[17][7:0] = buffer_data_3[3703:3696];
        layer3[17][15:8] = buffer_data_3[3711:3704];
        layer3[17][23:16] = buffer_data_3[3719:3712];
        layer3[17][31:24] = buffer_data_3[3727:3720];
        layer3[17][39:32] = buffer_data_3[3735:3728];
        layer3[17][47:40] = buffer_data_3[3743:3736];
        layer3[17][55:48] = buffer_data_3[3751:3744];
        layer4[17][7:0] = buffer_data_2[3703:3696];
        layer4[17][15:8] = buffer_data_2[3711:3704];
        layer4[17][23:16] = buffer_data_2[3719:3712];
        layer4[17][31:24] = buffer_data_2[3727:3720];
        layer4[17][39:32] = buffer_data_2[3735:3728];
        layer4[17][47:40] = buffer_data_2[3743:3736];
        layer4[17][55:48] = buffer_data_2[3751:3744];
        layer5[17][7:0] = buffer_data_1[3703:3696];
        layer5[17][15:8] = buffer_data_1[3711:3704];
        layer5[17][23:16] = buffer_data_1[3719:3712];
        layer5[17][31:24] = buffer_data_1[3727:3720];
        layer5[17][39:32] = buffer_data_1[3735:3728];
        layer5[17][47:40] = buffer_data_1[3743:3736];
        layer5[17][55:48] = buffer_data_1[3751:3744];
        layer6[17][7:0] = buffer_data_0[3703:3696];
        layer6[17][15:8] = buffer_data_0[3711:3704];
        layer6[17][23:16] = buffer_data_0[3719:3712];
        layer6[17][31:24] = buffer_data_0[3727:3720];
        layer6[17][39:32] = buffer_data_0[3735:3728];
        layer6[17][47:40] = buffer_data_0[3743:3736];
        layer6[17][55:48] = buffer_data_0[3751:3744];
        layer0[18][7:0] = buffer_data_6[3711:3704];
        layer0[18][15:8] = buffer_data_6[3719:3712];
        layer0[18][23:16] = buffer_data_6[3727:3720];
        layer0[18][31:24] = buffer_data_6[3735:3728];
        layer0[18][39:32] = buffer_data_6[3743:3736];
        layer0[18][47:40] = buffer_data_6[3751:3744];
        layer0[18][55:48] = buffer_data_6[3759:3752];
        layer1[18][7:0] = buffer_data_5[3711:3704];
        layer1[18][15:8] = buffer_data_5[3719:3712];
        layer1[18][23:16] = buffer_data_5[3727:3720];
        layer1[18][31:24] = buffer_data_5[3735:3728];
        layer1[18][39:32] = buffer_data_5[3743:3736];
        layer1[18][47:40] = buffer_data_5[3751:3744];
        layer1[18][55:48] = buffer_data_5[3759:3752];
        layer2[18][7:0] = buffer_data_4[3711:3704];
        layer2[18][15:8] = buffer_data_4[3719:3712];
        layer2[18][23:16] = buffer_data_4[3727:3720];
        layer2[18][31:24] = buffer_data_4[3735:3728];
        layer2[18][39:32] = buffer_data_4[3743:3736];
        layer2[18][47:40] = buffer_data_4[3751:3744];
        layer2[18][55:48] = buffer_data_4[3759:3752];
        layer3[18][7:0] = buffer_data_3[3711:3704];
        layer3[18][15:8] = buffer_data_3[3719:3712];
        layer3[18][23:16] = buffer_data_3[3727:3720];
        layer3[18][31:24] = buffer_data_3[3735:3728];
        layer3[18][39:32] = buffer_data_3[3743:3736];
        layer3[18][47:40] = buffer_data_3[3751:3744];
        layer3[18][55:48] = buffer_data_3[3759:3752];
        layer4[18][7:0] = buffer_data_2[3711:3704];
        layer4[18][15:8] = buffer_data_2[3719:3712];
        layer4[18][23:16] = buffer_data_2[3727:3720];
        layer4[18][31:24] = buffer_data_2[3735:3728];
        layer4[18][39:32] = buffer_data_2[3743:3736];
        layer4[18][47:40] = buffer_data_2[3751:3744];
        layer4[18][55:48] = buffer_data_2[3759:3752];
        layer5[18][7:0] = buffer_data_1[3711:3704];
        layer5[18][15:8] = buffer_data_1[3719:3712];
        layer5[18][23:16] = buffer_data_1[3727:3720];
        layer5[18][31:24] = buffer_data_1[3735:3728];
        layer5[18][39:32] = buffer_data_1[3743:3736];
        layer5[18][47:40] = buffer_data_1[3751:3744];
        layer5[18][55:48] = buffer_data_1[3759:3752];
        layer6[18][7:0] = buffer_data_0[3711:3704];
        layer6[18][15:8] = buffer_data_0[3719:3712];
        layer6[18][23:16] = buffer_data_0[3727:3720];
        layer6[18][31:24] = buffer_data_0[3735:3728];
        layer6[18][39:32] = buffer_data_0[3743:3736];
        layer6[18][47:40] = buffer_data_0[3751:3744];
        layer6[18][55:48] = buffer_data_0[3759:3752];
        layer0[19][7:0] = buffer_data_6[3719:3712];
        layer0[19][15:8] = buffer_data_6[3727:3720];
        layer0[19][23:16] = buffer_data_6[3735:3728];
        layer0[19][31:24] = buffer_data_6[3743:3736];
        layer0[19][39:32] = buffer_data_6[3751:3744];
        layer0[19][47:40] = buffer_data_6[3759:3752];
        layer0[19][55:48] = buffer_data_6[3767:3760];
        layer1[19][7:0] = buffer_data_5[3719:3712];
        layer1[19][15:8] = buffer_data_5[3727:3720];
        layer1[19][23:16] = buffer_data_5[3735:3728];
        layer1[19][31:24] = buffer_data_5[3743:3736];
        layer1[19][39:32] = buffer_data_5[3751:3744];
        layer1[19][47:40] = buffer_data_5[3759:3752];
        layer1[19][55:48] = buffer_data_5[3767:3760];
        layer2[19][7:0] = buffer_data_4[3719:3712];
        layer2[19][15:8] = buffer_data_4[3727:3720];
        layer2[19][23:16] = buffer_data_4[3735:3728];
        layer2[19][31:24] = buffer_data_4[3743:3736];
        layer2[19][39:32] = buffer_data_4[3751:3744];
        layer2[19][47:40] = buffer_data_4[3759:3752];
        layer2[19][55:48] = buffer_data_4[3767:3760];
        layer3[19][7:0] = buffer_data_3[3719:3712];
        layer3[19][15:8] = buffer_data_3[3727:3720];
        layer3[19][23:16] = buffer_data_3[3735:3728];
        layer3[19][31:24] = buffer_data_3[3743:3736];
        layer3[19][39:32] = buffer_data_3[3751:3744];
        layer3[19][47:40] = buffer_data_3[3759:3752];
        layer3[19][55:48] = buffer_data_3[3767:3760];
        layer4[19][7:0] = buffer_data_2[3719:3712];
        layer4[19][15:8] = buffer_data_2[3727:3720];
        layer4[19][23:16] = buffer_data_2[3735:3728];
        layer4[19][31:24] = buffer_data_2[3743:3736];
        layer4[19][39:32] = buffer_data_2[3751:3744];
        layer4[19][47:40] = buffer_data_2[3759:3752];
        layer4[19][55:48] = buffer_data_2[3767:3760];
        layer5[19][7:0] = buffer_data_1[3719:3712];
        layer5[19][15:8] = buffer_data_1[3727:3720];
        layer5[19][23:16] = buffer_data_1[3735:3728];
        layer5[19][31:24] = buffer_data_1[3743:3736];
        layer5[19][39:32] = buffer_data_1[3751:3744];
        layer5[19][47:40] = buffer_data_1[3759:3752];
        layer5[19][55:48] = buffer_data_1[3767:3760];
        layer6[19][7:0] = buffer_data_0[3719:3712];
        layer6[19][15:8] = buffer_data_0[3727:3720];
        layer6[19][23:16] = buffer_data_0[3735:3728];
        layer6[19][31:24] = buffer_data_0[3743:3736];
        layer6[19][39:32] = buffer_data_0[3751:3744];
        layer6[19][47:40] = buffer_data_0[3759:3752];
        layer6[19][55:48] = buffer_data_0[3767:3760];
        layer0[20][7:0] = buffer_data_6[3727:3720];
        layer0[20][15:8] = buffer_data_6[3735:3728];
        layer0[20][23:16] = buffer_data_6[3743:3736];
        layer0[20][31:24] = buffer_data_6[3751:3744];
        layer0[20][39:32] = buffer_data_6[3759:3752];
        layer0[20][47:40] = buffer_data_6[3767:3760];
        layer0[20][55:48] = buffer_data_6[3775:3768];
        layer1[20][7:0] = buffer_data_5[3727:3720];
        layer1[20][15:8] = buffer_data_5[3735:3728];
        layer1[20][23:16] = buffer_data_5[3743:3736];
        layer1[20][31:24] = buffer_data_5[3751:3744];
        layer1[20][39:32] = buffer_data_5[3759:3752];
        layer1[20][47:40] = buffer_data_5[3767:3760];
        layer1[20][55:48] = buffer_data_5[3775:3768];
        layer2[20][7:0] = buffer_data_4[3727:3720];
        layer2[20][15:8] = buffer_data_4[3735:3728];
        layer2[20][23:16] = buffer_data_4[3743:3736];
        layer2[20][31:24] = buffer_data_4[3751:3744];
        layer2[20][39:32] = buffer_data_4[3759:3752];
        layer2[20][47:40] = buffer_data_4[3767:3760];
        layer2[20][55:48] = buffer_data_4[3775:3768];
        layer3[20][7:0] = buffer_data_3[3727:3720];
        layer3[20][15:8] = buffer_data_3[3735:3728];
        layer3[20][23:16] = buffer_data_3[3743:3736];
        layer3[20][31:24] = buffer_data_3[3751:3744];
        layer3[20][39:32] = buffer_data_3[3759:3752];
        layer3[20][47:40] = buffer_data_3[3767:3760];
        layer3[20][55:48] = buffer_data_3[3775:3768];
        layer4[20][7:0] = buffer_data_2[3727:3720];
        layer4[20][15:8] = buffer_data_2[3735:3728];
        layer4[20][23:16] = buffer_data_2[3743:3736];
        layer4[20][31:24] = buffer_data_2[3751:3744];
        layer4[20][39:32] = buffer_data_2[3759:3752];
        layer4[20][47:40] = buffer_data_2[3767:3760];
        layer4[20][55:48] = buffer_data_2[3775:3768];
        layer5[20][7:0] = buffer_data_1[3727:3720];
        layer5[20][15:8] = buffer_data_1[3735:3728];
        layer5[20][23:16] = buffer_data_1[3743:3736];
        layer5[20][31:24] = buffer_data_1[3751:3744];
        layer5[20][39:32] = buffer_data_1[3759:3752];
        layer5[20][47:40] = buffer_data_1[3767:3760];
        layer5[20][55:48] = buffer_data_1[3775:3768];
        layer6[20][7:0] = buffer_data_0[3727:3720];
        layer6[20][15:8] = buffer_data_0[3735:3728];
        layer6[20][23:16] = buffer_data_0[3743:3736];
        layer6[20][31:24] = buffer_data_0[3751:3744];
        layer6[20][39:32] = buffer_data_0[3759:3752];
        layer6[20][47:40] = buffer_data_0[3767:3760];
        layer6[20][55:48] = buffer_data_0[3775:3768];
        layer0[21][7:0] = buffer_data_6[3735:3728];
        layer0[21][15:8] = buffer_data_6[3743:3736];
        layer0[21][23:16] = buffer_data_6[3751:3744];
        layer0[21][31:24] = buffer_data_6[3759:3752];
        layer0[21][39:32] = buffer_data_6[3767:3760];
        layer0[21][47:40] = buffer_data_6[3775:3768];
        layer0[21][55:48] = buffer_data_6[3783:3776];
        layer1[21][7:0] = buffer_data_5[3735:3728];
        layer1[21][15:8] = buffer_data_5[3743:3736];
        layer1[21][23:16] = buffer_data_5[3751:3744];
        layer1[21][31:24] = buffer_data_5[3759:3752];
        layer1[21][39:32] = buffer_data_5[3767:3760];
        layer1[21][47:40] = buffer_data_5[3775:3768];
        layer1[21][55:48] = buffer_data_5[3783:3776];
        layer2[21][7:0] = buffer_data_4[3735:3728];
        layer2[21][15:8] = buffer_data_4[3743:3736];
        layer2[21][23:16] = buffer_data_4[3751:3744];
        layer2[21][31:24] = buffer_data_4[3759:3752];
        layer2[21][39:32] = buffer_data_4[3767:3760];
        layer2[21][47:40] = buffer_data_4[3775:3768];
        layer2[21][55:48] = buffer_data_4[3783:3776];
        layer3[21][7:0] = buffer_data_3[3735:3728];
        layer3[21][15:8] = buffer_data_3[3743:3736];
        layer3[21][23:16] = buffer_data_3[3751:3744];
        layer3[21][31:24] = buffer_data_3[3759:3752];
        layer3[21][39:32] = buffer_data_3[3767:3760];
        layer3[21][47:40] = buffer_data_3[3775:3768];
        layer3[21][55:48] = buffer_data_3[3783:3776];
        layer4[21][7:0] = buffer_data_2[3735:3728];
        layer4[21][15:8] = buffer_data_2[3743:3736];
        layer4[21][23:16] = buffer_data_2[3751:3744];
        layer4[21][31:24] = buffer_data_2[3759:3752];
        layer4[21][39:32] = buffer_data_2[3767:3760];
        layer4[21][47:40] = buffer_data_2[3775:3768];
        layer4[21][55:48] = buffer_data_2[3783:3776];
        layer5[21][7:0] = buffer_data_1[3735:3728];
        layer5[21][15:8] = buffer_data_1[3743:3736];
        layer5[21][23:16] = buffer_data_1[3751:3744];
        layer5[21][31:24] = buffer_data_1[3759:3752];
        layer5[21][39:32] = buffer_data_1[3767:3760];
        layer5[21][47:40] = buffer_data_1[3775:3768];
        layer5[21][55:48] = buffer_data_1[3783:3776];
        layer6[21][7:0] = buffer_data_0[3735:3728];
        layer6[21][15:8] = buffer_data_0[3743:3736];
        layer6[21][23:16] = buffer_data_0[3751:3744];
        layer6[21][31:24] = buffer_data_0[3759:3752];
        layer6[21][39:32] = buffer_data_0[3767:3760];
        layer6[21][47:40] = buffer_data_0[3775:3768];
        layer6[21][55:48] = buffer_data_0[3783:3776];
        layer0[22][7:0] = buffer_data_6[3743:3736];
        layer0[22][15:8] = buffer_data_6[3751:3744];
        layer0[22][23:16] = buffer_data_6[3759:3752];
        layer0[22][31:24] = buffer_data_6[3767:3760];
        layer0[22][39:32] = buffer_data_6[3775:3768];
        layer0[22][47:40] = buffer_data_6[3783:3776];
        layer0[22][55:48] = buffer_data_6[3791:3784];
        layer1[22][7:0] = buffer_data_5[3743:3736];
        layer1[22][15:8] = buffer_data_5[3751:3744];
        layer1[22][23:16] = buffer_data_5[3759:3752];
        layer1[22][31:24] = buffer_data_5[3767:3760];
        layer1[22][39:32] = buffer_data_5[3775:3768];
        layer1[22][47:40] = buffer_data_5[3783:3776];
        layer1[22][55:48] = buffer_data_5[3791:3784];
        layer2[22][7:0] = buffer_data_4[3743:3736];
        layer2[22][15:8] = buffer_data_4[3751:3744];
        layer2[22][23:16] = buffer_data_4[3759:3752];
        layer2[22][31:24] = buffer_data_4[3767:3760];
        layer2[22][39:32] = buffer_data_4[3775:3768];
        layer2[22][47:40] = buffer_data_4[3783:3776];
        layer2[22][55:48] = buffer_data_4[3791:3784];
        layer3[22][7:0] = buffer_data_3[3743:3736];
        layer3[22][15:8] = buffer_data_3[3751:3744];
        layer3[22][23:16] = buffer_data_3[3759:3752];
        layer3[22][31:24] = buffer_data_3[3767:3760];
        layer3[22][39:32] = buffer_data_3[3775:3768];
        layer3[22][47:40] = buffer_data_3[3783:3776];
        layer3[22][55:48] = buffer_data_3[3791:3784];
        layer4[22][7:0] = buffer_data_2[3743:3736];
        layer4[22][15:8] = buffer_data_2[3751:3744];
        layer4[22][23:16] = buffer_data_2[3759:3752];
        layer4[22][31:24] = buffer_data_2[3767:3760];
        layer4[22][39:32] = buffer_data_2[3775:3768];
        layer4[22][47:40] = buffer_data_2[3783:3776];
        layer4[22][55:48] = buffer_data_2[3791:3784];
        layer5[22][7:0] = buffer_data_1[3743:3736];
        layer5[22][15:8] = buffer_data_1[3751:3744];
        layer5[22][23:16] = buffer_data_1[3759:3752];
        layer5[22][31:24] = buffer_data_1[3767:3760];
        layer5[22][39:32] = buffer_data_1[3775:3768];
        layer5[22][47:40] = buffer_data_1[3783:3776];
        layer5[22][55:48] = buffer_data_1[3791:3784];
        layer6[22][7:0] = buffer_data_0[3743:3736];
        layer6[22][15:8] = buffer_data_0[3751:3744];
        layer6[22][23:16] = buffer_data_0[3759:3752];
        layer6[22][31:24] = buffer_data_0[3767:3760];
        layer6[22][39:32] = buffer_data_0[3775:3768];
        layer6[22][47:40] = buffer_data_0[3783:3776];
        layer6[22][55:48] = buffer_data_0[3791:3784];
        layer0[23][7:0] = buffer_data_6[3751:3744];
        layer0[23][15:8] = buffer_data_6[3759:3752];
        layer0[23][23:16] = buffer_data_6[3767:3760];
        layer0[23][31:24] = buffer_data_6[3775:3768];
        layer0[23][39:32] = buffer_data_6[3783:3776];
        layer0[23][47:40] = buffer_data_6[3791:3784];
        layer0[23][55:48] = buffer_data_6[3799:3792];
        layer1[23][7:0] = buffer_data_5[3751:3744];
        layer1[23][15:8] = buffer_data_5[3759:3752];
        layer1[23][23:16] = buffer_data_5[3767:3760];
        layer1[23][31:24] = buffer_data_5[3775:3768];
        layer1[23][39:32] = buffer_data_5[3783:3776];
        layer1[23][47:40] = buffer_data_5[3791:3784];
        layer1[23][55:48] = buffer_data_5[3799:3792];
        layer2[23][7:0] = buffer_data_4[3751:3744];
        layer2[23][15:8] = buffer_data_4[3759:3752];
        layer2[23][23:16] = buffer_data_4[3767:3760];
        layer2[23][31:24] = buffer_data_4[3775:3768];
        layer2[23][39:32] = buffer_data_4[3783:3776];
        layer2[23][47:40] = buffer_data_4[3791:3784];
        layer2[23][55:48] = buffer_data_4[3799:3792];
        layer3[23][7:0] = buffer_data_3[3751:3744];
        layer3[23][15:8] = buffer_data_3[3759:3752];
        layer3[23][23:16] = buffer_data_3[3767:3760];
        layer3[23][31:24] = buffer_data_3[3775:3768];
        layer3[23][39:32] = buffer_data_3[3783:3776];
        layer3[23][47:40] = buffer_data_3[3791:3784];
        layer3[23][55:48] = buffer_data_3[3799:3792];
        layer4[23][7:0] = buffer_data_2[3751:3744];
        layer4[23][15:8] = buffer_data_2[3759:3752];
        layer4[23][23:16] = buffer_data_2[3767:3760];
        layer4[23][31:24] = buffer_data_2[3775:3768];
        layer4[23][39:32] = buffer_data_2[3783:3776];
        layer4[23][47:40] = buffer_data_2[3791:3784];
        layer4[23][55:48] = buffer_data_2[3799:3792];
        layer5[23][7:0] = buffer_data_1[3751:3744];
        layer5[23][15:8] = buffer_data_1[3759:3752];
        layer5[23][23:16] = buffer_data_1[3767:3760];
        layer5[23][31:24] = buffer_data_1[3775:3768];
        layer5[23][39:32] = buffer_data_1[3783:3776];
        layer5[23][47:40] = buffer_data_1[3791:3784];
        layer5[23][55:48] = buffer_data_1[3799:3792];
        layer6[23][7:0] = buffer_data_0[3751:3744];
        layer6[23][15:8] = buffer_data_0[3759:3752];
        layer6[23][23:16] = buffer_data_0[3767:3760];
        layer6[23][31:24] = buffer_data_0[3775:3768];
        layer6[23][39:32] = buffer_data_0[3783:3776];
        layer6[23][47:40] = buffer_data_0[3791:3784];
        layer6[23][55:48] = buffer_data_0[3799:3792];
        layer0[24][7:0] = buffer_data_6[3759:3752];
        layer0[24][15:8] = buffer_data_6[3767:3760];
        layer0[24][23:16] = buffer_data_6[3775:3768];
        layer0[24][31:24] = buffer_data_6[3783:3776];
        layer0[24][39:32] = buffer_data_6[3791:3784];
        layer0[24][47:40] = buffer_data_6[3799:3792];
        layer0[24][55:48] = buffer_data_6[3807:3800];
        layer1[24][7:0] = buffer_data_5[3759:3752];
        layer1[24][15:8] = buffer_data_5[3767:3760];
        layer1[24][23:16] = buffer_data_5[3775:3768];
        layer1[24][31:24] = buffer_data_5[3783:3776];
        layer1[24][39:32] = buffer_data_5[3791:3784];
        layer1[24][47:40] = buffer_data_5[3799:3792];
        layer1[24][55:48] = buffer_data_5[3807:3800];
        layer2[24][7:0] = buffer_data_4[3759:3752];
        layer2[24][15:8] = buffer_data_4[3767:3760];
        layer2[24][23:16] = buffer_data_4[3775:3768];
        layer2[24][31:24] = buffer_data_4[3783:3776];
        layer2[24][39:32] = buffer_data_4[3791:3784];
        layer2[24][47:40] = buffer_data_4[3799:3792];
        layer2[24][55:48] = buffer_data_4[3807:3800];
        layer3[24][7:0] = buffer_data_3[3759:3752];
        layer3[24][15:8] = buffer_data_3[3767:3760];
        layer3[24][23:16] = buffer_data_3[3775:3768];
        layer3[24][31:24] = buffer_data_3[3783:3776];
        layer3[24][39:32] = buffer_data_3[3791:3784];
        layer3[24][47:40] = buffer_data_3[3799:3792];
        layer3[24][55:48] = buffer_data_3[3807:3800];
        layer4[24][7:0] = buffer_data_2[3759:3752];
        layer4[24][15:8] = buffer_data_2[3767:3760];
        layer4[24][23:16] = buffer_data_2[3775:3768];
        layer4[24][31:24] = buffer_data_2[3783:3776];
        layer4[24][39:32] = buffer_data_2[3791:3784];
        layer4[24][47:40] = buffer_data_2[3799:3792];
        layer4[24][55:48] = buffer_data_2[3807:3800];
        layer5[24][7:0] = buffer_data_1[3759:3752];
        layer5[24][15:8] = buffer_data_1[3767:3760];
        layer5[24][23:16] = buffer_data_1[3775:3768];
        layer5[24][31:24] = buffer_data_1[3783:3776];
        layer5[24][39:32] = buffer_data_1[3791:3784];
        layer5[24][47:40] = buffer_data_1[3799:3792];
        layer5[24][55:48] = buffer_data_1[3807:3800];
        layer6[24][7:0] = buffer_data_0[3759:3752];
        layer6[24][15:8] = buffer_data_0[3767:3760];
        layer6[24][23:16] = buffer_data_0[3775:3768];
        layer6[24][31:24] = buffer_data_0[3783:3776];
        layer6[24][39:32] = buffer_data_0[3791:3784];
        layer6[24][47:40] = buffer_data_0[3799:3792];
        layer6[24][55:48] = buffer_data_0[3807:3800];
        layer0[25][7:0] = buffer_data_6[3767:3760];
        layer0[25][15:8] = buffer_data_6[3775:3768];
        layer0[25][23:16] = buffer_data_6[3783:3776];
        layer0[25][31:24] = buffer_data_6[3791:3784];
        layer0[25][39:32] = buffer_data_6[3799:3792];
        layer0[25][47:40] = buffer_data_6[3807:3800];
        layer0[25][55:48] = buffer_data_6[3815:3808];
        layer1[25][7:0] = buffer_data_5[3767:3760];
        layer1[25][15:8] = buffer_data_5[3775:3768];
        layer1[25][23:16] = buffer_data_5[3783:3776];
        layer1[25][31:24] = buffer_data_5[3791:3784];
        layer1[25][39:32] = buffer_data_5[3799:3792];
        layer1[25][47:40] = buffer_data_5[3807:3800];
        layer1[25][55:48] = buffer_data_5[3815:3808];
        layer2[25][7:0] = buffer_data_4[3767:3760];
        layer2[25][15:8] = buffer_data_4[3775:3768];
        layer2[25][23:16] = buffer_data_4[3783:3776];
        layer2[25][31:24] = buffer_data_4[3791:3784];
        layer2[25][39:32] = buffer_data_4[3799:3792];
        layer2[25][47:40] = buffer_data_4[3807:3800];
        layer2[25][55:48] = buffer_data_4[3815:3808];
        layer3[25][7:0] = buffer_data_3[3767:3760];
        layer3[25][15:8] = buffer_data_3[3775:3768];
        layer3[25][23:16] = buffer_data_3[3783:3776];
        layer3[25][31:24] = buffer_data_3[3791:3784];
        layer3[25][39:32] = buffer_data_3[3799:3792];
        layer3[25][47:40] = buffer_data_3[3807:3800];
        layer3[25][55:48] = buffer_data_3[3815:3808];
        layer4[25][7:0] = buffer_data_2[3767:3760];
        layer4[25][15:8] = buffer_data_2[3775:3768];
        layer4[25][23:16] = buffer_data_2[3783:3776];
        layer4[25][31:24] = buffer_data_2[3791:3784];
        layer4[25][39:32] = buffer_data_2[3799:3792];
        layer4[25][47:40] = buffer_data_2[3807:3800];
        layer4[25][55:48] = buffer_data_2[3815:3808];
        layer5[25][7:0] = buffer_data_1[3767:3760];
        layer5[25][15:8] = buffer_data_1[3775:3768];
        layer5[25][23:16] = buffer_data_1[3783:3776];
        layer5[25][31:24] = buffer_data_1[3791:3784];
        layer5[25][39:32] = buffer_data_1[3799:3792];
        layer5[25][47:40] = buffer_data_1[3807:3800];
        layer5[25][55:48] = buffer_data_1[3815:3808];
        layer6[25][7:0] = buffer_data_0[3767:3760];
        layer6[25][15:8] = buffer_data_0[3775:3768];
        layer6[25][23:16] = buffer_data_0[3783:3776];
        layer6[25][31:24] = buffer_data_0[3791:3784];
        layer6[25][39:32] = buffer_data_0[3799:3792];
        layer6[25][47:40] = buffer_data_0[3807:3800];
        layer6[25][55:48] = buffer_data_0[3815:3808];
        layer0[26][7:0] = buffer_data_6[3775:3768];
        layer0[26][15:8] = buffer_data_6[3783:3776];
        layer0[26][23:16] = buffer_data_6[3791:3784];
        layer0[26][31:24] = buffer_data_6[3799:3792];
        layer0[26][39:32] = buffer_data_6[3807:3800];
        layer0[26][47:40] = buffer_data_6[3815:3808];
        layer0[26][55:48] = buffer_data_6[3823:3816];
        layer1[26][7:0] = buffer_data_5[3775:3768];
        layer1[26][15:8] = buffer_data_5[3783:3776];
        layer1[26][23:16] = buffer_data_5[3791:3784];
        layer1[26][31:24] = buffer_data_5[3799:3792];
        layer1[26][39:32] = buffer_data_5[3807:3800];
        layer1[26][47:40] = buffer_data_5[3815:3808];
        layer1[26][55:48] = buffer_data_5[3823:3816];
        layer2[26][7:0] = buffer_data_4[3775:3768];
        layer2[26][15:8] = buffer_data_4[3783:3776];
        layer2[26][23:16] = buffer_data_4[3791:3784];
        layer2[26][31:24] = buffer_data_4[3799:3792];
        layer2[26][39:32] = buffer_data_4[3807:3800];
        layer2[26][47:40] = buffer_data_4[3815:3808];
        layer2[26][55:48] = buffer_data_4[3823:3816];
        layer3[26][7:0] = buffer_data_3[3775:3768];
        layer3[26][15:8] = buffer_data_3[3783:3776];
        layer3[26][23:16] = buffer_data_3[3791:3784];
        layer3[26][31:24] = buffer_data_3[3799:3792];
        layer3[26][39:32] = buffer_data_3[3807:3800];
        layer3[26][47:40] = buffer_data_3[3815:3808];
        layer3[26][55:48] = buffer_data_3[3823:3816];
        layer4[26][7:0] = buffer_data_2[3775:3768];
        layer4[26][15:8] = buffer_data_2[3783:3776];
        layer4[26][23:16] = buffer_data_2[3791:3784];
        layer4[26][31:24] = buffer_data_2[3799:3792];
        layer4[26][39:32] = buffer_data_2[3807:3800];
        layer4[26][47:40] = buffer_data_2[3815:3808];
        layer4[26][55:48] = buffer_data_2[3823:3816];
        layer5[26][7:0] = buffer_data_1[3775:3768];
        layer5[26][15:8] = buffer_data_1[3783:3776];
        layer5[26][23:16] = buffer_data_1[3791:3784];
        layer5[26][31:24] = buffer_data_1[3799:3792];
        layer5[26][39:32] = buffer_data_1[3807:3800];
        layer5[26][47:40] = buffer_data_1[3815:3808];
        layer5[26][55:48] = buffer_data_1[3823:3816];
        layer6[26][7:0] = buffer_data_0[3775:3768];
        layer6[26][15:8] = buffer_data_0[3783:3776];
        layer6[26][23:16] = buffer_data_0[3791:3784];
        layer6[26][31:24] = buffer_data_0[3799:3792];
        layer6[26][39:32] = buffer_data_0[3807:3800];
        layer6[26][47:40] = buffer_data_0[3815:3808];
        layer6[26][55:48] = buffer_data_0[3823:3816];
        layer0[27][7:0] = buffer_data_6[3783:3776];
        layer0[27][15:8] = buffer_data_6[3791:3784];
        layer0[27][23:16] = buffer_data_6[3799:3792];
        layer0[27][31:24] = buffer_data_6[3807:3800];
        layer0[27][39:32] = buffer_data_6[3815:3808];
        layer0[27][47:40] = buffer_data_6[3823:3816];
        layer0[27][55:48] = buffer_data_6[3831:3824];
        layer1[27][7:0] = buffer_data_5[3783:3776];
        layer1[27][15:8] = buffer_data_5[3791:3784];
        layer1[27][23:16] = buffer_data_5[3799:3792];
        layer1[27][31:24] = buffer_data_5[3807:3800];
        layer1[27][39:32] = buffer_data_5[3815:3808];
        layer1[27][47:40] = buffer_data_5[3823:3816];
        layer1[27][55:48] = buffer_data_5[3831:3824];
        layer2[27][7:0] = buffer_data_4[3783:3776];
        layer2[27][15:8] = buffer_data_4[3791:3784];
        layer2[27][23:16] = buffer_data_4[3799:3792];
        layer2[27][31:24] = buffer_data_4[3807:3800];
        layer2[27][39:32] = buffer_data_4[3815:3808];
        layer2[27][47:40] = buffer_data_4[3823:3816];
        layer2[27][55:48] = buffer_data_4[3831:3824];
        layer3[27][7:0] = buffer_data_3[3783:3776];
        layer3[27][15:8] = buffer_data_3[3791:3784];
        layer3[27][23:16] = buffer_data_3[3799:3792];
        layer3[27][31:24] = buffer_data_3[3807:3800];
        layer3[27][39:32] = buffer_data_3[3815:3808];
        layer3[27][47:40] = buffer_data_3[3823:3816];
        layer3[27][55:48] = buffer_data_3[3831:3824];
        layer4[27][7:0] = buffer_data_2[3783:3776];
        layer4[27][15:8] = buffer_data_2[3791:3784];
        layer4[27][23:16] = buffer_data_2[3799:3792];
        layer4[27][31:24] = buffer_data_2[3807:3800];
        layer4[27][39:32] = buffer_data_2[3815:3808];
        layer4[27][47:40] = buffer_data_2[3823:3816];
        layer4[27][55:48] = buffer_data_2[3831:3824];
        layer5[27][7:0] = buffer_data_1[3783:3776];
        layer5[27][15:8] = buffer_data_1[3791:3784];
        layer5[27][23:16] = buffer_data_1[3799:3792];
        layer5[27][31:24] = buffer_data_1[3807:3800];
        layer5[27][39:32] = buffer_data_1[3815:3808];
        layer5[27][47:40] = buffer_data_1[3823:3816];
        layer5[27][55:48] = buffer_data_1[3831:3824];
        layer6[27][7:0] = buffer_data_0[3783:3776];
        layer6[27][15:8] = buffer_data_0[3791:3784];
        layer6[27][23:16] = buffer_data_0[3799:3792];
        layer6[27][31:24] = buffer_data_0[3807:3800];
        layer6[27][39:32] = buffer_data_0[3815:3808];
        layer6[27][47:40] = buffer_data_0[3823:3816];
        layer6[27][55:48] = buffer_data_0[3831:3824];
        layer0[28][7:0] = buffer_data_6[3791:3784];
        layer0[28][15:8] = buffer_data_6[3799:3792];
        layer0[28][23:16] = buffer_data_6[3807:3800];
        layer0[28][31:24] = buffer_data_6[3815:3808];
        layer0[28][39:32] = buffer_data_6[3823:3816];
        layer0[28][47:40] = buffer_data_6[3831:3824];
        layer0[28][55:48] = buffer_data_6[3839:3832];
        layer1[28][7:0] = buffer_data_5[3791:3784];
        layer1[28][15:8] = buffer_data_5[3799:3792];
        layer1[28][23:16] = buffer_data_5[3807:3800];
        layer1[28][31:24] = buffer_data_5[3815:3808];
        layer1[28][39:32] = buffer_data_5[3823:3816];
        layer1[28][47:40] = buffer_data_5[3831:3824];
        layer1[28][55:48] = buffer_data_5[3839:3832];
        layer2[28][7:0] = buffer_data_4[3791:3784];
        layer2[28][15:8] = buffer_data_4[3799:3792];
        layer2[28][23:16] = buffer_data_4[3807:3800];
        layer2[28][31:24] = buffer_data_4[3815:3808];
        layer2[28][39:32] = buffer_data_4[3823:3816];
        layer2[28][47:40] = buffer_data_4[3831:3824];
        layer2[28][55:48] = buffer_data_4[3839:3832];
        layer3[28][7:0] = buffer_data_3[3791:3784];
        layer3[28][15:8] = buffer_data_3[3799:3792];
        layer3[28][23:16] = buffer_data_3[3807:3800];
        layer3[28][31:24] = buffer_data_3[3815:3808];
        layer3[28][39:32] = buffer_data_3[3823:3816];
        layer3[28][47:40] = buffer_data_3[3831:3824];
        layer3[28][55:48] = buffer_data_3[3839:3832];
        layer4[28][7:0] = buffer_data_2[3791:3784];
        layer4[28][15:8] = buffer_data_2[3799:3792];
        layer4[28][23:16] = buffer_data_2[3807:3800];
        layer4[28][31:24] = buffer_data_2[3815:3808];
        layer4[28][39:32] = buffer_data_2[3823:3816];
        layer4[28][47:40] = buffer_data_2[3831:3824];
        layer4[28][55:48] = buffer_data_2[3839:3832];
        layer5[28][7:0] = buffer_data_1[3791:3784];
        layer5[28][15:8] = buffer_data_1[3799:3792];
        layer5[28][23:16] = buffer_data_1[3807:3800];
        layer5[28][31:24] = buffer_data_1[3815:3808];
        layer5[28][39:32] = buffer_data_1[3823:3816];
        layer5[28][47:40] = buffer_data_1[3831:3824];
        layer5[28][55:48] = buffer_data_1[3839:3832];
        layer6[28][7:0] = buffer_data_0[3791:3784];
        layer6[28][15:8] = buffer_data_0[3799:3792];
        layer6[28][23:16] = buffer_data_0[3807:3800];
        layer6[28][31:24] = buffer_data_0[3815:3808];
        layer6[28][39:32] = buffer_data_0[3823:3816];
        layer6[28][47:40] = buffer_data_0[3831:3824];
        layer6[28][55:48] = buffer_data_0[3839:3832];
        layer0[29][7:0] = buffer_data_6[3799:3792];
        layer0[29][15:8] = buffer_data_6[3807:3800];
        layer0[29][23:16] = buffer_data_6[3815:3808];
        layer0[29][31:24] = buffer_data_6[3823:3816];
        layer0[29][39:32] = buffer_data_6[3831:3824];
        layer0[29][47:40] = buffer_data_6[3839:3832];
        layer0[29][55:48] = buffer_data_6[3847:3840];
        layer1[29][7:0] = buffer_data_5[3799:3792];
        layer1[29][15:8] = buffer_data_5[3807:3800];
        layer1[29][23:16] = buffer_data_5[3815:3808];
        layer1[29][31:24] = buffer_data_5[3823:3816];
        layer1[29][39:32] = buffer_data_5[3831:3824];
        layer1[29][47:40] = buffer_data_5[3839:3832];
        layer1[29][55:48] = buffer_data_5[3847:3840];
        layer2[29][7:0] = buffer_data_4[3799:3792];
        layer2[29][15:8] = buffer_data_4[3807:3800];
        layer2[29][23:16] = buffer_data_4[3815:3808];
        layer2[29][31:24] = buffer_data_4[3823:3816];
        layer2[29][39:32] = buffer_data_4[3831:3824];
        layer2[29][47:40] = buffer_data_4[3839:3832];
        layer2[29][55:48] = buffer_data_4[3847:3840];
        layer3[29][7:0] = buffer_data_3[3799:3792];
        layer3[29][15:8] = buffer_data_3[3807:3800];
        layer3[29][23:16] = buffer_data_3[3815:3808];
        layer3[29][31:24] = buffer_data_3[3823:3816];
        layer3[29][39:32] = buffer_data_3[3831:3824];
        layer3[29][47:40] = buffer_data_3[3839:3832];
        layer3[29][55:48] = buffer_data_3[3847:3840];
        layer4[29][7:0] = buffer_data_2[3799:3792];
        layer4[29][15:8] = buffer_data_2[3807:3800];
        layer4[29][23:16] = buffer_data_2[3815:3808];
        layer4[29][31:24] = buffer_data_2[3823:3816];
        layer4[29][39:32] = buffer_data_2[3831:3824];
        layer4[29][47:40] = buffer_data_2[3839:3832];
        layer4[29][55:48] = buffer_data_2[3847:3840];
        layer5[29][7:0] = buffer_data_1[3799:3792];
        layer5[29][15:8] = buffer_data_1[3807:3800];
        layer5[29][23:16] = buffer_data_1[3815:3808];
        layer5[29][31:24] = buffer_data_1[3823:3816];
        layer5[29][39:32] = buffer_data_1[3831:3824];
        layer5[29][47:40] = buffer_data_1[3839:3832];
        layer5[29][55:48] = buffer_data_1[3847:3840];
        layer6[29][7:0] = buffer_data_0[3799:3792];
        layer6[29][15:8] = buffer_data_0[3807:3800];
        layer6[29][23:16] = buffer_data_0[3815:3808];
        layer6[29][31:24] = buffer_data_0[3823:3816];
        layer6[29][39:32] = buffer_data_0[3831:3824];
        layer6[29][47:40] = buffer_data_0[3839:3832];
        layer6[29][55:48] = buffer_data_0[3847:3840];
        layer0[30][7:0] = buffer_data_6[3807:3800];
        layer0[30][15:8] = buffer_data_6[3815:3808];
        layer0[30][23:16] = buffer_data_6[3823:3816];
        layer0[30][31:24] = buffer_data_6[3831:3824];
        layer0[30][39:32] = buffer_data_6[3839:3832];
        layer0[30][47:40] = buffer_data_6[3847:3840];
        layer0[30][55:48] = buffer_data_6[3855:3848];
        layer1[30][7:0] = buffer_data_5[3807:3800];
        layer1[30][15:8] = buffer_data_5[3815:3808];
        layer1[30][23:16] = buffer_data_5[3823:3816];
        layer1[30][31:24] = buffer_data_5[3831:3824];
        layer1[30][39:32] = buffer_data_5[3839:3832];
        layer1[30][47:40] = buffer_data_5[3847:3840];
        layer1[30][55:48] = buffer_data_5[3855:3848];
        layer2[30][7:0] = buffer_data_4[3807:3800];
        layer2[30][15:8] = buffer_data_4[3815:3808];
        layer2[30][23:16] = buffer_data_4[3823:3816];
        layer2[30][31:24] = buffer_data_4[3831:3824];
        layer2[30][39:32] = buffer_data_4[3839:3832];
        layer2[30][47:40] = buffer_data_4[3847:3840];
        layer2[30][55:48] = buffer_data_4[3855:3848];
        layer3[30][7:0] = buffer_data_3[3807:3800];
        layer3[30][15:8] = buffer_data_3[3815:3808];
        layer3[30][23:16] = buffer_data_3[3823:3816];
        layer3[30][31:24] = buffer_data_3[3831:3824];
        layer3[30][39:32] = buffer_data_3[3839:3832];
        layer3[30][47:40] = buffer_data_3[3847:3840];
        layer3[30][55:48] = buffer_data_3[3855:3848];
        layer4[30][7:0] = buffer_data_2[3807:3800];
        layer4[30][15:8] = buffer_data_2[3815:3808];
        layer4[30][23:16] = buffer_data_2[3823:3816];
        layer4[30][31:24] = buffer_data_2[3831:3824];
        layer4[30][39:32] = buffer_data_2[3839:3832];
        layer4[30][47:40] = buffer_data_2[3847:3840];
        layer4[30][55:48] = buffer_data_2[3855:3848];
        layer5[30][7:0] = buffer_data_1[3807:3800];
        layer5[30][15:8] = buffer_data_1[3815:3808];
        layer5[30][23:16] = buffer_data_1[3823:3816];
        layer5[30][31:24] = buffer_data_1[3831:3824];
        layer5[30][39:32] = buffer_data_1[3839:3832];
        layer5[30][47:40] = buffer_data_1[3847:3840];
        layer5[30][55:48] = buffer_data_1[3855:3848];
        layer6[30][7:0] = buffer_data_0[3807:3800];
        layer6[30][15:8] = buffer_data_0[3815:3808];
        layer6[30][23:16] = buffer_data_0[3823:3816];
        layer6[30][31:24] = buffer_data_0[3831:3824];
        layer6[30][39:32] = buffer_data_0[3839:3832];
        layer6[30][47:40] = buffer_data_0[3847:3840];
        layer6[30][55:48] = buffer_data_0[3855:3848];
        layer0[31][7:0] = buffer_data_6[3815:3808];
        layer0[31][15:8] = buffer_data_6[3823:3816];
        layer0[31][23:16] = buffer_data_6[3831:3824];
        layer0[31][31:24] = buffer_data_6[3839:3832];
        layer0[31][39:32] = buffer_data_6[3847:3840];
        layer0[31][47:40] = buffer_data_6[3855:3848];
        layer0[31][55:48] = buffer_data_6[3863:3856];
        layer1[31][7:0] = buffer_data_5[3815:3808];
        layer1[31][15:8] = buffer_data_5[3823:3816];
        layer1[31][23:16] = buffer_data_5[3831:3824];
        layer1[31][31:24] = buffer_data_5[3839:3832];
        layer1[31][39:32] = buffer_data_5[3847:3840];
        layer1[31][47:40] = buffer_data_5[3855:3848];
        layer1[31][55:48] = buffer_data_5[3863:3856];
        layer2[31][7:0] = buffer_data_4[3815:3808];
        layer2[31][15:8] = buffer_data_4[3823:3816];
        layer2[31][23:16] = buffer_data_4[3831:3824];
        layer2[31][31:24] = buffer_data_4[3839:3832];
        layer2[31][39:32] = buffer_data_4[3847:3840];
        layer2[31][47:40] = buffer_data_4[3855:3848];
        layer2[31][55:48] = buffer_data_4[3863:3856];
        layer3[31][7:0] = buffer_data_3[3815:3808];
        layer3[31][15:8] = buffer_data_3[3823:3816];
        layer3[31][23:16] = buffer_data_3[3831:3824];
        layer3[31][31:24] = buffer_data_3[3839:3832];
        layer3[31][39:32] = buffer_data_3[3847:3840];
        layer3[31][47:40] = buffer_data_3[3855:3848];
        layer3[31][55:48] = buffer_data_3[3863:3856];
        layer4[31][7:0] = buffer_data_2[3815:3808];
        layer4[31][15:8] = buffer_data_2[3823:3816];
        layer4[31][23:16] = buffer_data_2[3831:3824];
        layer4[31][31:24] = buffer_data_2[3839:3832];
        layer4[31][39:32] = buffer_data_2[3847:3840];
        layer4[31][47:40] = buffer_data_2[3855:3848];
        layer4[31][55:48] = buffer_data_2[3863:3856];
        layer5[31][7:0] = buffer_data_1[3815:3808];
        layer5[31][15:8] = buffer_data_1[3823:3816];
        layer5[31][23:16] = buffer_data_1[3831:3824];
        layer5[31][31:24] = buffer_data_1[3839:3832];
        layer5[31][39:32] = buffer_data_1[3847:3840];
        layer5[31][47:40] = buffer_data_1[3855:3848];
        layer5[31][55:48] = buffer_data_1[3863:3856];
        layer6[31][7:0] = buffer_data_0[3815:3808];
        layer6[31][15:8] = buffer_data_0[3823:3816];
        layer6[31][23:16] = buffer_data_0[3831:3824];
        layer6[31][31:24] = buffer_data_0[3839:3832];
        layer6[31][39:32] = buffer_data_0[3847:3840];
        layer6[31][47:40] = buffer_data_0[3855:3848];
        layer6[31][55:48] = buffer_data_0[3863:3856];
        layer0[32][7:0] = buffer_data_6[3823:3816];
        layer0[32][15:8] = buffer_data_6[3831:3824];
        layer0[32][23:16] = buffer_data_6[3839:3832];
        layer0[32][31:24] = buffer_data_6[3847:3840];
        layer0[32][39:32] = buffer_data_6[3855:3848];
        layer0[32][47:40] = buffer_data_6[3863:3856];
        layer0[32][55:48] = buffer_data_6[3871:3864];
        layer1[32][7:0] = buffer_data_5[3823:3816];
        layer1[32][15:8] = buffer_data_5[3831:3824];
        layer1[32][23:16] = buffer_data_5[3839:3832];
        layer1[32][31:24] = buffer_data_5[3847:3840];
        layer1[32][39:32] = buffer_data_5[3855:3848];
        layer1[32][47:40] = buffer_data_5[3863:3856];
        layer1[32][55:48] = buffer_data_5[3871:3864];
        layer2[32][7:0] = buffer_data_4[3823:3816];
        layer2[32][15:8] = buffer_data_4[3831:3824];
        layer2[32][23:16] = buffer_data_4[3839:3832];
        layer2[32][31:24] = buffer_data_4[3847:3840];
        layer2[32][39:32] = buffer_data_4[3855:3848];
        layer2[32][47:40] = buffer_data_4[3863:3856];
        layer2[32][55:48] = buffer_data_4[3871:3864];
        layer3[32][7:0] = buffer_data_3[3823:3816];
        layer3[32][15:8] = buffer_data_3[3831:3824];
        layer3[32][23:16] = buffer_data_3[3839:3832];
        layer3[32][31:24] = buffer_data_3[3847:3840];
        layer3[32][39:32] = buffer_data_3[3855:3848];
        layer3[32][47:40] = buffer_data_3[3863:3856];
        layer3[32][55:48] = buffer_data_3[3871:3864];
        layer4[32][7:0] = buffer_data_2[3823:3816];
        layer4[32][15:8] = buffer_data_2[3831:3824];
        layer4[32][23:16] = buffer_data_2[3839:3832];
        layer4[32][31:24] = buffer_data_2[3847:3840];
        layer4[32][39:32] = buffer_data_2[3855:3848];
        layer4[32][47:40] = buffer_data_2[3863:3856];
        layer4[32][55:48] = buffer_data_2[3871:3864];
        layer5[32][7:0] = buffer_data_1[3823:3816];
        layer5[32][15:8] = buffer_data_1[3831:3824];
        layer5[32][23:16] = buffer_data_1[3839:3832];
        layer5[32][31:24] = buffer_data_1[3847:3840];
        layer5[32][39:32] = buffer_data_1[3855:3848];
        layer5[32][47:40] = buffer_data_1[3863:3856];
        layer5[32][55:48] = buffer_data_1[3871:3864];
        layer6[32][7:0] = buffer_data_0[3823:3816];
        layer6[32][15:8] = buffer_data_0[3831:3824];
        layer6[32][23:16] = buffer_data_0[3839:3832];
        layer6[32][31:24] = buffer_data_0[3847:3840];
        layer6[32][39:32] = buffer_data_0[3855:3848];
        layer6[32][47:40] = buffer_data_0[3863:3856];
        layer6[32][55:48] = buffer_data_0[3871:3864];
        layer0[33][7:0] = buffer_data_6[3831:3824];
        layer0[33][15:8] = buffer_data_6[3839:3832];
        layer0[33][23:16] = buffer_data_6[3847:3840];
        layer0[33][31:24] = buffer_data_6[3855:3848];
        layer0[33][39:32] = buffer_data_6[3863:3856];
        layer0[33][47:40] = buffer_data_6[3871:3864];
        layer0[33][55:48] = buffer_data_6[3879:3872];
        layer1[33][7:0] = buffer_data_5[3831:3824];
        layer1[33][15:8] = buffer_data_5[3839:3832];
        layer1[33][23:16] = buffer_data_5[3847:3840];
        layer1[33][31:24] = buffer_data_5[3855:3848];
        layer1[33][39:32] = buffer_data_5[3863:3856];
        layer1[33][47:40] = buffer_data_5[3871:3864];
        layer1[33][55:48] = buffer_data_5[3879:3872];
        layer2[33][7:0] = buffer_data_4[3831:3824];
        layer2[33][15:8] = buffer_data_4[3839:3832];
        layer2[33][23:16] = buffer_data_4[3847:3840];
        layer2[33][31:24] = buffer_data_4[3855:3848];
        layer2[33][39:32] = buffer_data_4[3863:3856];
        layer2[33][47:40] = buffer_data_4[3871:3864];
        layer2[33][55:48] = buffer_data_4[3879:3872];
        layer3[33][7:0] = buffer_data_3[3831:3824];
        layer3[33][15:8] = buffer_data_3[3839:3832];
        layer3[33][23:16] = buffer_data_3[3847:3840];
        layer3[33][31:24] = buffer_data_3[3855:3848];
        layer3[33][39:32] = buffer_data_3[3863:3856];
        layer3[33][47:40] = buffer_data_3[3871:3864];
        layer3[33][55:48] = buffer_data_3[3879:3872];
        layer4[33][7:0] = buffer_data_2[3831:3824];
        layer4[33][15:8] = buffer_data_2[3839:3832];
        layer4[33][23:16] = buffer_data_2[3847:3840];
        layer4[33][31:24] = buffer_data_2[3855:3848];
        layer4[33][39:32] = buffer_data_2[3863:3856];
        layer4[33][47:40] = buffer_data_2[3871:3864];
        layer4[33][55:48] = buffer_data_2[3879:3872];
        layer5[33][7:0] = buffer_data_1[3831:3824];
        layer5[33][15:8] = buffer_data_1[3839:3832];
        layer5[33][23:16] = buffer_data_1[3847:3840];
        layer5[33][31:24] = buffer_data_1[3855:3848];
        layer5[33][39:32] = buffer_data_1[3863:3856];
        layer5[33][47:40] = buffer_data_1[3871:3864];
        layer5[33][55:48] = buffer_data_1[3879:3872];
        layer6[33][7:0] = buffer_data_0[3831:3824];
        layer6[33][15:8] = buffer_data_0[3839:3832];
        layer6[33][23:16] = buffer_data_0[3847:3840];
        layer6[33][31:24] = buffer_data_0[3855:3848];
        layer6[33][39:32] = buffer_data_0[3863:3856];
        layer6[33][47:40] = buffer_data_0[3871:3864];
        layer6[33][55:48] = buffer_data_0[3879:3872];
        layer0[34][7:0] = buffer_data_6[3839:3832];
        layer0[34][15:8] = buffer_data_6[3847:3840];
        layer0[34][23:16] = buffer_data_6[3855:3848];
        layer0[34][31:24] = buffer_data_6[3863:3856];
        layer0[34][39:32] = buffer_data_6[3871:3864];
        layer0[34][47:40] = buffer_data_6[3879:3872];
        layer0[34][55:48] = buffer_data_6[3887:3880];
        layer1[34][7:0] = buffer_data_5[3839:3832];
        layer1[34][15:8] = buffer_data_5[3847:3840];
        layer1[34][23:16] = buffer_data_5[3855:3848];
        layer1[34][31:24] = buffer_data_5[3863:3856];
        layer1[34][39:32] = buffer_data_5[3871:3864];
        layer1[34][47:40] = buffer_data_5[3879:3872];
        layer1[34][55:48] = buffer_data_5[3887:3880];
        layer2[34][7:0] = buffer_data_4[3839:3832];
        layer2[34][15:8] = buffer_data_4[3847:3840];
        layer2[34][23:16] = buffer_data_4[3855:3848];
        layer2[34][31:24] = buffer_data_4[3863:3856];
        layer2[34][39:32] = buffer_data_4[3871:3864];
        layer2[34][47:40] = buffer_data_4[3879:3872];
        layer2[34][55:48] = buffer_data_4[3887:3880];
        layer3[34][7:0] = buffer_data_3[3839:3832];
        layer3[34][15:8] = buffer_data_3[3847:3840];
        layer3[34][23:16] = buffer_data_3[3855:3848];
        layer3[34][31:24] = buffer_data_3[3863:3856];
        layer3[34][39:32] = buffer_data_3[3871:3864];
        layer3[34][47:40] = buffer_data_3[3879:3872];
        layer3[34][55:48] = buffer_data_3[3887:3880];
        layer4[34][7:0] = buffer_data_2[3839:3832];
        layer4[34][15:8] = buffer_data_2[3847:3840];
        layer4[34][23:16] = buffer_data_2[3855:3848];
        layer4[34][31:24] = buffer_data_2[3863:3856];
        layer4[34][39:32] = buffer_data_2[3871:3864];
        layer4[34][47:40] = buffer_data_2[3879:3872];
        layer4[34][55:48] = buffer_data_2[3887:3880];
        layer5[34][7:0] = buffer_data_1[3839:3832];
        layer5[34][15:8] = buffer_data_1[3847:3840];
        layer5[34][23:16] = buffer_data_1[3855:3848];
        layer5[34][31:24] = buffer_data_1[3863:3856];
        layer5[34][39:32] = buffer_data_1[3871:3864];
        layer5[34][47:40] = buffer_data_1[3879:3872];
        layer5[34][55:48] = buffer_data_1[3887:3880];
        layer6[34][7:0] = buffer_data_0[3839:3832];
        layer6[34][15:8] = buffer_data_0[3847:3840];
        layer6[34][23:16] = buffer_data_0[3855:3848];
        layer6[34][31:24] = buffer_data_0[3863:3856];
        layer6[34][39:32] = buffer_data_0[3871:3864];
        layer6[34][47:40] = buffer_data_0[3879:3872];
        layer6[34][55:48] = buffer_data_0[3887:3880];
        layer0[35][7:0] = buffer_data_6[3847:3840];
        layer0[35][15:8] = buffer_data_6[3855:3848];
        layer0[35][23:16] = buffer_data_6[3863:3856];
        layer0[35][31:24] = buffer_data_6[3871:3864];
        layer0[35][39:32] = buffer_data_6[3879:3872];
        layer0[35][47:40] = buffer_data_6[3887:3880];
        layer0[35][55:48] = buffer_data_6[3895:3888];
        layer1[35][7:0] = buffer_data_5[3847:3840];
        layer1[35][15:8] = buffer_data_5[3855:3848];
        layer1[35][23:16] = buffer_data_5[3863:3856];
        layer1[35][31:24] = buffer_data_5[3871:3864];
        layer1[35][39:32] = buffer_data_5[3879:3872];
        layer1[35][47:40] = buffer_data_5[3887:3880];
        layer1[35][55:48] = buffer_data_5[3895:3888];
        layer2[35][7:0] = buffer_data_4[3847:3840];
        layer2[35][15:8] = buffer_data_4[3855:3848];
        layer2[35][23:16] = buffer_data_4[3863:3856];
        layer2[35][31:24] = buffer_data_4[3871:3864];
        layer2[35][39:32] = buffer_data_4[3879:3872];
        layer2[35][47:40] = buffer_data_4[3887:3880];
        layer2[35][55:48] = buffer_data_4[3895:3888];
        layer3[35][7:0] = buffer_data_3[3847:3840];
        layer3[35][15:8] = buffer_data_3[3855:3848];
        layer3[35][23:16] = buffer_data_3[3863:3856];
        layer3[35][31:24] = buffer_data_3[3871:3864];
        layer3[35][39:32] = buffer_data_3[3879:3872];
        layer3[35][47:40] = buffer_data_3[3887:3880];
        layer3[35][55:48] = buffer_data_3[3895:3888];
        layer4[35][7:0] = buffer_data_2[3847:3840];
        layer4[35][15:8] = buffer_data_2[3855:3848];
        layer4[35][23:16] = buffer_data_2[3863:3856];
        layer4[35][31:24] = buffer_data_2[3871:3864];
        layer4[35][39:32] = buffer_data_2[3879:3872];
        layer4[35][47:40] = buffer_data_2[3887:3880];
        layer4[35][55:48] = buffer_data_2[3895:3888];
        layer5[35][7:0] = buffer_data_1[3847:3840];
        layer5[35][15:8] = buffer_data_1[3855:3848];
        layer5[35][23:16] = buffer_data_1[3863:3856];
        layer5[35][31:24] = buffer_data_1[3871:3864];
        layer5[35][39:32] = buffer_data_1[3879:3872];
        layer5[35][47:40] = buffer_data_1[3887:3880];
        layer5[35][55:48] = buffer_data_1[3895:3888];
        layer6[35][7:0] = buffer_data_0[3847:3840];
        layer6[35][15:8] = buffer_data_0[3855:3848];
        layer6[35][23:16] = buffer_data_0[3863:3856];
        layer6[35][31:24] = buffer_data_0[3871:3864];
        layer6[35][39:32] = buffer_data_0[3879:3872];
        layer6[35][47:40] = buffer_data_0[3887:3880];
        layer6[35][55:48] = buffer_data_0[3895:3888];
        layer0[36][7:0] = buffer_data_6[3855:3848];
        layer0[36][15:8] = buffer_data_6[3863:3856];
        layer0[36][23:16] = buffer_data_6[3871:3864];
        layer0[36][31:24] = buffer_data_6[3879:3872];
        layer0[36][39:32] = buffer_data_6[3887:3880];
        layer0[36][47:40] = buffer_data_6[3895:3888];
        layer0[36][55:48] = buffer_data_6[3903:3896];
        layer1[36][7:0] = buffer_data_5[3855:3848];
        layer1[36][15:8] = buffer_data_5[3863:3856];
        layer1[36][23:16] = buffer_data_5[3871:3864];
        layer1[36][31:24] = buffer_data_5[3879:3872];
        layer1[36][39:32] = buffer_data_5[3887:3880];
        layer1[36][47:40] = buffer_data_5[3895:3888];
        layer1[36][55:48] = buffer_data_5[3903:3896];
        layer2[36][7:0] = buffer_data_4[3855:3848];
        layer2[36][15:8] = buffer_data_4[3863:3856];
        layer2[36][23:16] = buffer_data_4[3871:3864];
        layer2[36][31:24] = buffer_data_4[3879:3872];
        layer2[36][39:32] = buffer_data_4[3887:3880];
        layer2[36][47:40] = buffer_data_4[3895:3888];
        layer2[36][55:48] = buffer_data_4[3903:3896];
        layer3[36][7:0] = buffer_data_3[3855:3848];
        layer3[36][15:8] = buffer_data_3[3863:3856];
        layer3[36][23:16] = buffer_data_3[3871:3864];
        layer3[36][31:24] = buffer_data_3[3879:3872];
        layer3[36][39:32] = buffer_data_3[3887:3880];
        layer3[36][47:40] = buffer_data_3[3895:3888];
        layer3[36][55:48] = buffer_data_3[3903:3896];
        layer4[36][7:0] = buffer_data_2[3855:3848];
        layer4[36][15:8] = buffer_data_2[3863:3856];
        layer4[36][23:16] = buffer_data_2[3871:3864];
        layer4[36][31:24] = buffer_data_2[3879:3872];
        layer4[36][39:32] = buffer_data_2[3887:3880];
        layer4[36][47:40] = buffer_data_2[3895:3888];
        layer4[36][55:48] = buffer_data_2[3903:3896];
        layer5[36][7:0] = buffer_data_1[3855:3848];
        layer5[36][15:8] = buffer_data_1[3863:3856];
        layer5[36][23:16] = buffer_data_1[3871:3864];
        layer5[36][31:24] = buffer_data_1[3879:3872];
        layer5[36][39:32] = buffer_data_1[3887:3880];
        layer5[36][47:40] = buffer_data_1[3895:3888];
        layer5[36][55:48] = buffer_data_1[3903:3896];
        layer6[36][7:0] = buffer_data_0[3855:3848];
        layer6[36][15:8] = buffer_data_0[3863:3856];
        layer6[36][23:16] = buffer_data_0[3871:3864];
        layer6[36][31:24] = buffer_data_0[3879:3872];
        layer6[36][39:32] = buffer_data_0[3887:3880];
        layer6[36][47:40] = buffer_data_0[3895:3888];
        layer6[36][55:48] = buffer_data_0[3903:3896];
        layer0[37][7:0] = buffer_data_6[3863:3856];
        layer0[37][15:8] = buffer_data_6[3871:3864];
        layer0[37][23:16] = buffer_data_6[3879:3872];
        layer0[37][31:24] = buffer_data_6[3887:3880];
        layer0[37][39:32] = buffer_data_6[3895:3888];
        layer0[37][47:40] = buffer_data_6[3903:3896];
        layer0[37][55:48] = buffer_data_6[3911:3904];
        layer1[37][7:0] = buffer_data_5[3863:3856];
        layer1[37][15:8] = buffer_data_5[3871:3864];
        layer1[37][23:16] = buffer_data_5[3879:3872];
        layer1[37][31:24] = buffer_data_5[3887:3880];
        layer1[37][39:32] = buffer_data_5[3895:3888];
        layer1[37][47:40] = buffer_data_5[3903:3896];
        layer1[37][55:48] = buffer_data_5[3911:3904];
        layer2[37][7:0] = buffer_data_4[3863:3856];
        layer2[37][15:8] = buffer_data_4[3871:3864];
        layer2[37][23:16] = buffer_data_4[3879:3872];
        layer2[37][31:24] = buffer_data_4[3887:3880];
        layer2[37][39:32] = buffer_data_4[3895:3888];
        layer2[37][47:40] = buffer_data_4[3903:3896];
        layer2[37][55:48] = buffer_data_4[3911:3904];
        layer3[37][7:0] = buffer_data_3[3863:3856];
        layer3[37][15:8] = buffer_data_3[3871:3864];
        layer3[37][23:16] = buffer_data_3[3879:3872];
        layer3[37][31:24] = buffer_data_3[3887:3880];
        layer3[37][39:32] = buffer_data_3[3895:3888];
        layer3[37][47:40] = buffer_data_3[3903:3896];
        layer3[37][55:48] = buffer_data_3[3911:3904];
        layer4[37][7:0] = buffer_data_2[3863:3856];
        layer4[37][15:8] = buffer_data_2[3871:3864];
        layer4[37][23:16] = buffer_data_2[3879:3872];
        layer4[37][31:24] = buffer_data_2[3887:3880];
        layer4[37][39:32] = buffer_data_2[3895:3888];
        layer4[37][47:40] = buffer_data_2[3903:3896];
        layer4[37][55:48] = buffer_data_2[3911:3904];
        layer5[37][7:0] = buffer_data_1[3863:3856];
        layer5[37][15:8] = buffer_data_1[3871:3864];
        layer5[37][23:16] = buffer_data_1[3879:3872];
        layer5[37][31:24] = buffer_data_1[3887:3880];
        layer5[37][39:32] = buffer_data_1[3895:3888];
        layer5[37][47:40] = buffer_data_1[3903:3896];
        layer5[37][55:48] = buffer_data_1[3911:3904];
        layer6[37][7:0] = buffer_data_0[3863:3856];
        layer6[37][15:8] = buffer_data_0[3871:3864];
        layer6[37][23:16] = buffer_data_0[3879:3872];
        layer6[37][31:24] = buffer_data_0[3887:3880];
        layer6[37][39:32] = buffer_data_0[3895:3888];
        layer6[37][47:40] = buffer_data_0[3903:3896];
        layer6[37][55:48] = buffer_data_0[3911:3904];
        layer0[38][7:0] = buffer_data_6[3871:3864];
        layer0[38][15:8] = buffer_data_6[3879:3872];
        layer0[38][23:16] = buffer_data_6[3887:3880];
        layer0[38][31:24] = buffer_data_6[3895:3888];
        layer0[38][39:32] = buffer_data_6[3903:3896];
        layer0[38][47:40] = buffer_data_6[3911:3904];
        layer0[38][55:48] = buffer_data_6[3919:3912];
        layer1[38][7:0] = buffer_data_5[3871:3864];
        layer1[38][15:8] = buffer_data_5[3879:3872];
        layer1[38][23:16] = buffer_data_5[3887:3880];
        layer1[38][31:24] = buffer_data_5[3895:3888];
        layer1[38][39:32] = buffer_data_5[3903:3896];
        layer1[38][47:40] = buffer_data_5[3911:3904];
        layer1[38][55:48] = buffer_data_5[3919:3912];
        layer2[38][7:0] = buffer_data_4[3871:3864];
        layer2[38][15:8] = buffer_data_4[3879:3872];
        layer2[38][23:16] = buffer_data_4[3887:3880];
        layer2[38][31:24] = buffer_data_4[3895:3888];
        layer2[38][39:32] = buffer_data_4[3903:3896];
        layer2[38][47:40] = buffer_data_4[3911:3904];
        layer2[38][55:48] = buffer_data_4[3919:3912];
        layer3[38][7:0] = buffer_data_3[3871:3864];
        layer3[38][15:8] = buffer_data_3[3879:3872];
        layer3[38][23:16] = buffer_data_3[3887:3880];
        layer3[38][31:24] = buffer_data_3[3895:3888];
        layer3[38][39:32] = buffer_data_3[3903:3896];
        layer3[38][47:40] = buffer_data_3[3911:3904];
        layer3[38][55:48] = buffer_data_3[3919:3912];
        layer4[38][7:0] = buffer_data_2[3871:3864];
        layer4[38][15:8] = buffer_data_2[3879:3872];
        layer4[38][23:16] = buffer_data_2[3887:3880];
        layer4[38][31:24] = buffer_data_2[3895:3888];
        layer4[38][39:32] = buffer_data_2[3903:3896];
        layer4[38][47:40] = buffer_data_2[3911:3904];
        layer4[38][55:48] = buffer_data_2[3919:3912];
        layer5[38][7:0] = buffer_data_1[3871:3864];
        layer5[38][15:8] = buffer_data_1[3879:3872];
        layer5[38][23:16] = buffer_data_1[3887:3880];
        layer5[38][31:24] = buffer_data_1[3895:3888];
        layer5[38][39:32] = buffer_data_1[3903:3896];
        layer5[38][47:40] = buffer_data_1[3911:3904];
        layer5[38][55:48] = buffer_data_1[3919:3912];
        layer6[38][7:0] = buffer_data_0[3871:3864];
        layer6[38][15:8] = buffer_data_0[3879:3872];
        layer6[38][23:16] = buffer_data_0[3887:3880];
        layer6[38][31:24] = buffer_data_0[3895:3888];
        layer6[38][39:32] = buffer_data_0[3903:3896];
        layer6[38][47:40] = buffer_data_0[3911:3904];
        layer6[38][55:48] = buffer_data_0[3919:3912];
        layer0[39][7:0] = buffer_data_6[3879:3872];
        layer0[39][15:8] = buffer_data_6[3887:3880];
        layer0[39][23:16] = buffer_data_6[3895:3888];
        layer0[39][31:24] = buffer_data_6[3903:3896];
        layer0[39][39:32] = buffer_data_6[3911:3904];
        layer0[39][47:40] = buffer_data_6[3919:3912];
        layer0[39][55:48] = buffer_data_6[3927:3920];
        layer1[39][7:0] = buffer_data_5[3879:3872];
        layer1[39][15:8] = buffer_data_5[3887:3880];
        layer1[39][23:16] = buffer_data_5[3895:3888];
        layer1[39][31:24] = buffer_data_5[3903:3896];
        layer1[39][39:32] = buffer_data_5[3911:3904];
        layer1[39][47:40] = buffer_data_5[3919:3912];
        layer1[39][55:48] = buffer_data_5[3927:3920];
        layer2[39][7:0] = buffer_data_4[3879:3872];
        layer2[39][15:8] = buffer_data_4[3887:3880];
        layer2[39][23:16] = buffer_data_4[3895:3888];
        layer2[39][31:24] = buffer_data_4[3903:3896];
        layer2[39][39:32] = buffer_data_4[3911:3904];
        layer2[39][47:40] = buffer_data_4[3919:3912];
        layer2[39][55:48] = buffer_data_4[3927:3920];
        layer3[39][7:0] = buffer_data_3[3879:3872];
        layer3[39][15:8] = buffer_data_3[3887:3880];
        layer3[39][23:16] = buffer_data_3[3895:3888];
        layer3[39][31:24] = buffer_data_3[3903:3896];
        layer3[39][39:32] = buffer_data_3[3911:3904];
        layer3[39][47:40] = buffer_data_3[3919:3912];
        layer3[39][55:48] = buffer_data_3[3927:3920];
        layer4[39][7:0] = buffer_data_2[3879:3872];
        layer4[39][15:8] = buffer_data_2[3887:3880];
        layer4[39][23:16] = buffer_data_2[3895:3888];
        layer4[39][31:24] = buffer_data_2[3903:3896];
        layer4[39][39:32] = buffer_data_2[3911:3904];
        layer4[39][47:40] = buffer_data_2[3919:3912];
        layer4[39][55:48] = buffer_data_2[3927:3920];
        layer5[39][7:0] = buffer_data_1[3879:3872];
        layer5[39][15:8] = buffer_data_1[3887:3880];
        layer5[39][23:16] = buffer_data_1[3895:3888];
        layer5[39][31:24] = buffer_data_1[3903:3896];
        layer5[39][39:32] = buffer_data_1[3911:3904];
        layer5[39][47:40] = buffer_data_1[3919:3912];
        layer5[39][55:48] = buffer_data_1[3927:3920];
        layer6[39][7:0] = buffer_data_0[3879:3872];
        layer6[39][15:8] = buffer_data_0[3887:3880];
        layer6[39][23:16] = buffer_data_0[3895:3888];
        layer6[39][31:24] = buffer_data_0[3903:3896];
        layer6[39][39:32] = buffer_data_0[3911:3904];
        layer6[39][47:40] = buffer_data_0[3919:3912];
        layer6[39][55:48] = buffer_data_0[3927:3920];
        layer0[40][7:0] = buffer_data_6[3887:3880];
        layer0[40][15:8] = buffer_data_6[3895:3888];
        layer0[40][23:16] = buffer_data_6[3903:3896];
        layer0[40][31:24] = buffer_data_6[3911:3904];
        layer0[40][39:32] = buffer_data_6[3919:3912];
        layer0[40][47:40] = buffer_data_6[3927:3920];
        layer0[40][55:48] = buffer_data_6[3935:3928];
        layer1[40][7:0] = buffer_data_5[3887:3880];
        layer1[40][15:8] = buffer_data_5[3895:3888];
        layer1[40][23:16] = buffer_data_5[3903:3896];
        layer1[40][31:24] = buffer_data_5[3911:3904];
        layer1[40][39:32] = buffer_data_5[3919:3912];
        layer1[40][47:40] = buffer_data_5[3927:3920];
        layer1[40][55:48] = buffer_data_5[3935:3928];
        layer2[40][7:0] = buffer_data_4[3887:3880];
        layer2[40][15:8] = buffer_data_4[3895:3888];
        layer2[40][23:16] = buffer_data_4[3903:3896];
        layer2[40][31:24] = buffer_data_4[3911:3904];
        layer2[40][39:32] = buffer_data_4[3919:3912];
        layer2[40][47:40] = buffer_data_4[3927:3920];
        layer2[40][55:48] = buffer_data_4[3935:3928];
        layer3[40][7:0] = buffer_data_3[3887:3880];
        layer3[40][15:8] = buffer_data_3[3895:3888];
        layer3[40][23:16] = buffer_data_3[3903:3896];
        layer3[40][31:24] = buffer_data_3[3911:3904];
        layer3[40][39:32] = buffer_data_3[3919:3912];
        layer3[40][47:40] = buffer_data_3[3927:3920];
        layer3[40][55:48] = buffer_data_3[3935:3928];
        layer4[40][7:0] = buffer_data_2[3887:3880];
        layer4[40][15:8] = buffer_data_2[3895:3888];
        layer4[40][23:16] = buffer_data_2[3903:3896];
        layer4[40][31:24] = buffer_data_2[3911:3904];
        layer4[40][39:32] = buffer_data_2[3919:3912];
        layer4[40][47:40] = buffer_data_2[3927:3920];
        layer4[40][55:48] = buffer_data_2[3935:3928];
        layer5[40][7:0] = buffer_data_1[3887:3880];
        layer5[40][15:8] = buffer_data_1[3895:3888];
        layer5[40][23:16] = buffer_data_1[3903:3896];
        layer5[40][31:24] = buffer_data_1[3911:3904];
        layer5[40][39:32] = buffer_data_1[3919:3912];
        layer5[40][47:40] = buffer_data_1[3927:3920];
        layer5[40][55:48] = buffer_data_1[3935:3928];
        layer6[40][7:0] = buffer_data_0[3887:3880];
        layer6[40][15:8] = buffer_data_0[3895:3888];
        layer6[40][23:16] = buffer_data_0[3903:3896];
        layer6[40][31:24] = buffer_data_0[3911:3904];
        layer6[40][39:32] = buffer_data_0[3919:3912];
        layer6[40][47:40] = buffer_data_0[3927:3920];
        layer6[40][55:48] = buffer_data_0[3935:3928];
        layer0[41][7:0] = buffer_data_6[3895:3888];
        layer0[41][15:8] = buffer_data_6[3903:3896];
        layer0[41][23:16] = buffer_data_6[3911:3904];
        layer0[41][31:24] = buffer_data_6[3919:3912];
        layer0[41][39:32] = buffer_data_6[3927:3920];
        layer0[41][47:40] = buffer_data_6[3935:3928];
        layer0[41][55:48] = buffer_data_6[3943:3936];
        layer1[41][7:0] = buffer_data_5[3895:3888];
        layer1[41][15:8] = buffer_data_5[3903:3896];
        layer1[41][23:16] = buffer_data_5[3911:3904];
        layer1[41][31:24] = buffer_data_5[3919:3912];
        layer1[41][39:32] = buffer_data_5[3927:3920];
        layer1[41][47:40] = buffer_data_5[3935:3928];
        layer1[41][55:48] = buffer_data_5[3943:3936];
        layer2[41][7:0] = buffer_data_4[3895:3888];
        layer2[41][15:8] = buffer_data_4[3903:3896];
        layer2[41][23:16] = buffer_data_4[3911:3904];
        layer2[41][31:24] = buffer_data_4[3919:3912];
        layer2[41][39:32] = buffer_data_4[3927:3920];
        layer2[41][47:40] = buffer_data_4[3935:3928];
        layer2[41][55:48] = buffer_data_4[3943:3936];
        layer3[41][7:0] = buffer_data_3[3895:3888];
        layer3[41][15:8] = buffer_data_3[3903:3896];
        layer3[41][23:16] = buffer_data_3[3911:3904];
        layer3[41][31:24] = buffer_data_3[3919:3912];
        layer3[41][39:32] = buffer_data_3[3927:3920];
        layer3[41][47:40] = buffer_data_3[3935:3928];
        layer3[41][55:48] = buffer_data_3[3943:3936];
        layer4[41][7:0] = buffer_data_2[3895:3888];
        layer4[41][15:8] = buffer_data_2[3903:3896];
        layer4[41][23:16] = buffer_data_2[3911:3904];
        layer4[41][31:24] = buffer_data_2[3919:3912];
        layer4[41][39:32] = buffer_data_2[3927:3920];
        layer4[41][47:40] = buffer_data_2[3935:3928];
        layer4[41][55:48] = buffer_data_2[3943:3936];
        layer5[41][7:0] = buffer_data_1[3895:3888];
        layer5[41][15:8] = buffer_data_1[3903:3896];
        layer5[41][23:16] = buffer_data_1[3911:3904];
        layer5[41][31:24] = buffer_data_1[3919:3912];
        layer5[41][39:32] = buffer_data_1[3927:3920];
        layer5[41][47:40] = buffer_data_1[3935:3928];
        layer5[41][55:48] = buffer_data_1[3943:3936];
        layer6[41][7:0] = buffer_data_0[3895:3888];
        layer6[41][15:8] = buffer_data_0[3903:3896];
        layer6[41][23:16] = buffer_data_0[3911:3904];
        layer6[41][31:24] = buffer_data_0[3919:3912];
        layer6[41][39:32] = buffer_data_0[3927:3920];
        layer6[41][47:40] = buffer_data_0[3935:3928];
        layer6[41][55:48] = buffer_data_0[3943:3936];
        layer0[42][7:0] = buffer_data_6[3903:3896];
        layer0[42][15:8] = buffer_data_6[3911:3904];
        layer0[42][23:16] = buffer_data_6[3919:3912];
        layer0[42][31:24] = buffer_data_6[3927:3920];
        layer0[42][39:32] = buffer_data_6[3935:3928];
        layer0[42][47:40] = buffer_data_6[3943:3936];
        layer0[42][55:48] = buffer_data_6[3951:3944];
        layer1[42][7:0] = buffer_data_5[3903:3896];
        layer1[42][15:8] = buffer_data_5[3911:3904];
        layer1[42][23:16] = buffer_data_5[3919:3912];
        layer1[42][31:24] = buffer_data_5[3927:3920];
        layer1[42][39:32] = buffer_data_5[3935:3928];
        layer1[42][47:40] = buffer_data_5[3943:3936];
        layer1[42][55:48] = buffer_data_5[3951:3944];
        layer2[42][7:0] = buffer_data_4[3903:3896];
        layer2[42][15:8] = buffer_data_4[3911:3904];
        layer2[42][23:16] = buffer_data_4[3919:3912];
        layer2[42][31:24] = buffer_data_4[3927:3920];
        layer2[42][39:32] = buffer_data_4[3935:3928];
        layer2[42][47:40] = buffer_data_4[3943:3936];
        layer2[42][55:48] = buffer_data_4[3951:3944];
        layer3[42][7:0] = buffer_data_3[3903:3896];
        layer3[42][15:8] = buffer_data_3[3911:3904];
        layer3[42][23:16] = buffer_data_3[3919:3912];
        layer3[42][31:24] = buffer_data_3[3927:3920];
        layer3[42][39:32] = buffer_data_3[3935:3928];
        layer3[42][47:40] = buffer_data_3[3943:3936];
        layer3[42][55:48] = buffer_data_3[3951:3944];
        layer4[42][7:0] = buffer_data_2[3903:3896];
        layer4[42][15:8] = buffer_data_2[3911:3904];
        layer4[42][23:16] = buffer_data_2[3919:3912];
        layer4[42][31:24] = buffer_data_2[3927:3920];
        layer4[42][39:32] = buffer_data_2[3935:3928];
        layer4[42][47:40] = buffer_data_2[3943:3936];
        layer4[42][55:48] = buffer_data_2[3951:3944];
        layer5[42][7:0] = buffer_data_1[3903:3896];
        layer5[42][15:8] = buffer_data_1[3911:3904];
        layer5[42][23:16] = buffer_data_1[3919:3912];
        layer5[42][31:24] = buffer_data_1[3927:3920];
        layer5[42][39:32] = buffer_data_1[3935:3928];
        layer5[42][47:40] = buffer_data_1[3943:3936];
        layer5[42][55:48] = buffer_data_1[3951:3944];
        layer6[42][7:0] = buffer_data_0[3903:3896];
        layer6[42][15:8] = buffer_data_0[3911:3904];
        layer6[42][23:16] = buffer_data_0[3919:3912];
        layer6[42][31:24] = buffer_data_0[3927:3920];
        layer6[42][39:32] = buffer_data_0[3935:3928];
        layer6[42][47:40] = buffer_data_0[3943:3936];
        layer6[42][55:48] = buffer_data_0[3951:3944];
        layer0[43][7:0] = buffer_data_6[3911:3904];
        layer0[43][15:8] = buffer_data_6[3919:3912];
        layer0[43][23:16] = buffer_data_6[3927:3920];
        layer0[43][31:24] = buffer_data_6[3935:3928];
        layer0[43][39:32] = buffer_data_6[3943:3936];
        layer0[43][47:40] = buffer_data_6[3951:3944];
        layer0[43][55:48] = buffer_data_6[3959:3952];
        layer1[43][7:0] = buffer_data_5[3911:3904];
        layer1[43][15:8] = buffer_data_5[3919:3912];
        layer1[43][23:16] = buffer_data_5[3927:3920];
        layer1[43][31:24] = buffer_data_5[3935:3928];
        layer1[43][39:32] = buffer_data_5[3943:3936];
        layer1[43][47:40] = buffer_data_5[3951:3944];
        layer1[43][55:48] = buffer_data_5[3959:3952];
        layer2[43][7:0] = buffer_data_4[3911:3904];
        layer2[43][15:8] = buffer_data_4[3919:3912];
        layer2[43][23:16] = buffer_data_4[3927:3920];
        layer2[43][31:24] = buffer_data_4[3935:3928];
        layer2[43][39:32] = buffer_data_4[3943:3936];
        layer2[43][47:40] = buffer_data_4[3951:3944];
        layer2[43][55:48] = buffer_data_4[3959:3952];
        layer3[43][7:0] = buffer_data_3[3911:3904];
        layer3[43][15:8] = buffer_data_3[3919:3912];
        layer3[43][23:16] = buffer_data_3[3927:3920];
        layer3[43][31:24] = buffer_data_3[3935:3928];
        layer3[43][39:32] = buffer_data_3[3943:3936];
        layer3[43][47:40] = buffer_data_3[3951:3944];
        layer3[43][55:48] = buffer_data_3[3959:3952];
        layer4[43][7:0] = buffer_data_2[3911:3904];
        layer4[43][15:8] = buffer_data_2[3919:3912];
        layer4[43][23:16] = buffer_data_2[3927:3920];
        layer4[43][31:24] = buffer_data_2[3935:3928];
        layer4[43][39:32] = buffer_data_2[3943:3936];
        layer4[43][47:40] = buffer_data_2[3951:3944];
        layer4[43][55:48] = buffer_data_2[3959:3952];
        layer5[43][7:0] = buffer_data_1[3911:3904];
        layer5[43][15:8] = buffer_data_1[3919:3912];
        layer5[43][23:16] = buffer_data_1[3927:3920];
        layer5[43][31:24] = buffer_data_1[3935:3928];
        layer5[43][39:32] = buffer_data_1[3943:3936];
        layer5[43][47:40] = buffer_data_1[3951:3944];
        layer5[43][55:48] = buffer_data_1[3959:3952];
        layer6[43][7:0] = buffer_data_0[3911:3904];
        layer6[43][15:8] = buffer_data_0[3919:3912];
        layer6[43][23:16] = buffer_data_0[3927:3920];
        layer6[43][31:24] = buffer_data_0[3935:3928];
        layer6[43][39:32] = buffer_data_0[3943:3936];
        layer6[43][47:40] = buffer_data_0[3951:3944];
        layer6[43][55:48] = buffer_data_0[3959:3952];
        layer0[44][7:0] = buffer_data_6[3919:3912];
        layer0[44][15:8] = buffer_data_6[3927:3920];
        layer0[44][23:16] = buffer_data_6[3935:3928];
        layer0[44][31:24] = buffer_data_6[3943:3936];
        layer0[44][39:32] = buffer_data_6[3951:3944];
        layer0[44][47:40] = buffer_data_6[3959:3952];
        layer0[44][55:48] = buffer_data_6[3967:3960];
        layer1[44][7:0] = buffer_data_5[3919:3912];
        layer1[44][15:8] = buffer_data_5[3927:3920];
        layer1[44][23:16] = buffer_data_5[3935:3928];
        layer1[44][31:24] = buffer_data_5[3943:3936];
        layer1[44][39:32] = buffer_data_5[3951:3944];
        layer1[44][47:40] = buffer_data_5[3959:3952];
        layer1[44][55:48] = buffer_data_5[3967:3960];
        layer2[44][7:0] = buffer_data_4[3919:3912];
        layer2[44][15:8] = buffer_data_4[3927:3920];
        layer2[44][23:16] = buffer_data_4[3935:3928];
        layer2[44][31:24] = buffer_data_4[3943:3936];
        layer2[44][39:32] = buffer_data_4[3951:3944];
        layer2[44][47:40] = buffer_data_4[3959:3952];
        layer2[44][55:48] = buffer_data_4[3967:3960];
        layer3[44][7:0] = buffer_data_3[3919:3912];
        layer3[44][15:8] = buffer_data_3[3927:3920];
        layer3[44][23:16] = buffer_data_3[3935:3928];
        layer3[44][31:24] = buffer_data_3[3943:3936];
        layer3[44][39:32] = buffer_data_3[3951:3944];
        layer3[44][47:40] = buffer_data_3[3959:3952];
        layer3[44][55:48] = buffer_data_3[3967:3960];
        layer4[44][7:0] = buffer_data_2[3919:3912];
        layer4[44][15:8] = buffer_data_2[3927:3920];
        layer4[44][23:16] = buffer_data_2[3935:3928];
        layer4[44][31:24] = buffer_data_2[3943:3936];
        layer4[44][39:32] = buffer_data_2[3951:3944];
        layer4[44][47:40] = buffer_data_2[3959:3952];
        layer4[44][55:48] = buffer_data_2[3967:3960];
        layer5[44][7:0] = buffer_data_1[3919:3912];
        layer5[44][15:8] = buffer_data_1[3927:3920];
        layer5[44][23:16] = buffer_data_1[3935:3928];
        layer5[44][31:24] = buffer_data_1[3943:3936];
        layer5[44][39:32] = buffer_data_1[3951:3944];
        layer5[44][47:40] = buffer_data_1[3959:3952];
        layer5[44][55:48] = buffer_data_1[3967:3960];
        layer6[44][7:0] = buffer_data_0[3919:3912];
        layer6[44][15:8] = buffer_data_0[3927:3920];
        layer6[44][23:16] = buffer_data_0[3935:3928];
        layer6[44][31:24] = buffer_data_0[3943:3936];
        layer6[44][39:32] = buffer_data_0[3951:3944];
        layer6[44][47:40] = buffer_data_0[3959:3952];
        layer6[44][55:48] = buffer_data_0[3967:3960];
        layer0[45][7:0] = buffer_data_6[3927:3920];
        layer0[45][15:8] = buffer_data_6[3935:3928];
        layer0[45][23:16] = buffer_data_6[3943:3936];
        layer0[45][31:24] = buffer_data_6[3951:3944];
        layer0[45][39:32] = buffer_data_6[3959:3952];
        layer0[45][47:40] = buffer_data_6[3967:3960];
        layer0[45][55:48] = buffer_data_6[3975:3968];
        layer1[45][7:0] = buffer_data_5[3927:3920];
        layer1[45][15:8] = buffer_data_5[3935:3928];
        layer1[45][23:16] = buffer_data_5[3943:3936];
        layer1[45][31:24] = buffer_data_5[3951:3944];
        layer1[45][39:32] = buffer_data_5[3959:3952];
        layer1[45][47:40] = buffer_data_5[3967:3960];
        layer1[45][55:48] = buffer_data_5[3975:3968];
        layer2[45][7:0] = buffer_data_4[3927:3920];
        layer2[45][15:8] = buffer_data_4[3935:3928];
        layer2[45][23:16] = buffer_data_4[3943:3936];
        layer2[45][31:24] = buffer_data_4[3951:3944];
        layer2[45][39:32] = buffer_data_4[3959:3952];
        layer2[45][47:40] = buffer_data_4[3967:3960];
        layer2[45][55:48] = buffer_data_4[3975:3968];
        layer3[45][7:0] = buffer_data_3[3927:3920];
        layer3[45][15:8] = buffer_data_3[3935:3928];
        layer3[45][23:16] = buffer_data_3[3943:3936];
        layer3[45][31:24] = buffer_data_3[3951:3944];
        layer3[45][39:32] = buffer_data_3[3959:3952];
        layer3[45][47:40] = buffer_data_3[3967:3960];
        layer3[45][55:48] = buffer_data_3[3975:3968];
        layer4[45][7:0] = buffer_data_2[3927:3920];
        layer4[45][15:8] = buffer_data_2[3935:3928];
        layer4[45][23:16] = buffer_data_2[3943:3936];
        layer4[45][31:24] = buffer_data_2[3951:3944];
        layer4[45][39:32] = buffer_data_2[3959:3952];
        layer4[45][47:40] = buffer_data_2[3967:3960];
        layer4[45][55:48] = buffer_data_2[3975:3968];
        layer5[45][7:0] = buffer_data_1[3927:3920];
        layer5[45][15:8] = buffer_data_1[3935:3928];
        layer5[45][23:16] = buffer_data_1[3943:3936];
        layer5[45][31:24] = buffer_data_1[3951:3944];
        layer5[45][39:32] = buffer_data_1[3959:3952];
        layer5[45][47:40] = buffer_data_1[3967:3960];
        layer5[45][55:48] = buffer_data_1[3975:3968];
        layer6[45][7:0] = buffer_data_0[3927:3920];
        layer6[45][15:8] = buffer_data_0[3935:3928];
        layer6[45][23:16] = buffer_data_0[3943:3936];
        layer6[45][31:24] = buffer_data_0[3951:3944];
        layer6[45][39:32] = buffer_data_0[3959:3952];
        layer6[45][47:40] = buffer_data_0[3967:3960];
        layer6[45][55:48] = buffer_data_0[3975:3968];
        layer0[46][7:0] = buffer_data_6[3935:3928];
        layer0[46][15:8] = buffer_data_6[3943:3936];
        layer0[46][23:16] = buffer_data_6[3951:3944];
        layer0[46][31:24] = buffer_data_6[3959:3952];
        layer0[46][39:32] = buffer_data_6[3967:3960];
        layer0[46][47:40] = buffer_data_6[3975:3968];
        layer0[46][55:48] = buffer_data_6[3983:3976];
        layer1[46][7:0] = buffer_data_5[3935:3928];
        layer1[46][15:8] = buffer_data_5[3943:3936];
        layer1[46][23:16] = buffer_data_5[3951:3944];
        layer1[46][31:24] = buffer_data_5[3959:3952];
        layer1[46][39:32] = buffer_data_5[3967:3960];
        layer1[46][47:40] = buffer_data_5[3975:3968];
        layer1[46][55:48] = buffer_data_5[3983:3976];
        layer2[46][7:0] = buffer_data_4[3935:3928];
        layer2[46][15:8] = buffer_data_4[3943:3936];
        layer2[46][23:16] = buffer_data_4[3951:3944];
        layer2[46][31:24] = buffer_data_4[3959:3952];
        layer2[46][39:32] = buffer_data_4[3967:3960];
        layer2[46][47:40] = buffer_data_4[3975:3968];
        layer2[46][55:48] = buffer_data_4[3983:3976];
        layer3[46][7:0] = buffer_data_3[3935:3928];
        layer3[46][15:8] = buffer_data_3[3943:3936];
        layer3[46][23:16] = buffer_data_3[3951:3944];
        layer3[46][31:24] = buffer_data_3[3959:3952];
        layer3[46][39:32] = buffer_data_3[3967:3960];
        layer3[46][47:40] = buffer_data_3[3975:3968];
        layer3[46][55:48] = buffer_data_3[3983:3976];
        layer4[46][7:0] = buffer_data_2[3935:3928];
        layer4[46][15:8] = buffer_data_2[3943:3936];
        layer4[46][23:16] = buffer_data_2[3951:3944];
        layer4[46][31:24] = buffer_data_2[3959:3952];
        layer4[46][39:32] = buffer_data_2[3967:3960];
        layer4[46][47:40] = buffer_data_2[3975:3968];
        layer4[46][55:48] = buffer_data_2[3983:3976];
        layer5[46][7:0] = buffer_data_1[3935:3928];
        layer5[46][15:8] = buffer_data_1[3943:3936];
        layer5[46][23:16] = buffer_data_1[3951:3944];
        layer5[46][31:24] = buffer_data_1[3959:3952];
        layer5[46][39:32] = buffer_data_1[3967:3960];
        layer5[46][47:40] = buffer_data_1[3975:3968];
        layer5[46][55:48] = buffer_data_1[3983:3976];
        layer6[46][7:0] = buffer_data_0[3935:3928];
        layer6[46][15:8] = buffer_data_0[3943:3936];
        layer6[46][23:16] = buffer_data_0[3951:3944];
        layer6[46][31:24] = buffer_data_0[3959:3952];
        layer6[46][39:32] = buffer_data_0[3967:3960];
        layer6[46][47:40] = buffer_data_0[3975:3968];
        layer6[46][55:48] = buffer_data_0[3983:3976];
        layer0[47][7:0] = buffer_data_6[3943:3936];
        layer0[47][15:8] = buffer_data_6[3951:3944];
        layer0[47][23:16] = buffer_data_6[3959:3952];
        layer0[47][31:24] = buffer_data_6[3967:3960];
        layer0[47][39:32] = buffer_data_6[3975:3968];
        layer0[47][47:40] = buffer_data_6[3983:3976];
        layer0[47][55:48] = buffer_data_6[3991:3984];
        layer1[47][7:0] = buffer_data_5[3943:3936];
        layer1[47][15:8] = buffer_data_5[3951:3944];
        layer1[47][23:16] = buffer_data_5[3959:3952];
        layer1[47][31:24] = buffer_data_5[3967:3960];
        layer1[47][39:32] = buffer_data_5[3975:3968];
        layer1[47][47:40] = buffer_data_5[3983:3976];
        layer1[47][55:48] = buffer_data_5[3991:3984];
        layer2[47][7:0] = buffer_data_4[3943:3936];
        layer2[47][15:8] = buffer_data_4[3951:3944];
        layer2[47][23:16] = buffer_data_4[3959:3952];
        layer2[47][31:24] = buffer_data_4[3967:3960];
        layer2[47][39:32] = buffer_data_4[3975:3968];
        layer2[47][47:40] = buffer_data_4[3983:3976];
        layer2[47][55:48] = buffer_data_4[3991:3984];
        layer3[47][7:0] = buffer_data_3[3943:3936];
        layer3[47][15:8] = buffer_data_3[3951:3944];
        layer3[47][23:16] = buffer_data_3[3959:3952];
        layer3[47][31:24] = buffer_data_3[3967:3960];
        layer3[47][39:32] = buffer_data_3[3975:3968];
        layer3[47][47:40] = buffer_data_3[3983:3976];
        layer3[47][55:48] = buffer_data_3[3991:3984];
        layer4[47][7:0] = buffer_data_2[3943:3936];
        layer4[47][15:8] = buffer_data_2[3951:3944];
        layer4[47][23:16] = buffer_data_2[3959:3952];
        layer4[47][31:24] = buffer_data_2[3967:3960];
        layer4[47][39:32] = buffer_data_2[3975:3968];
        layer4[47][47:40] = buffer_data_2[3983:3976];
        layer4[47][55:48] = buffer_data_2[3991:3984];
        layer5[47][7:0] = buffer_data_1[3943:3936];
        layer5[47][15:8] = buffer_data_1[3951:3944];
        layer5[47][23:16] = buffer_data_1[3959:3952];
        layer5[47][31:24] = buffer_data_1[3967:3960];
        layer5[47][39:32] = buffer_data_1[3975:3968];
        layer5[47][47:40] = buffer_data_1[3983:3976];
        layer5[47][55:48] = buffer_data_1[3991:3984];
        layer6[47][7:0] = buffer_data_0[3943:3936];
        layer6[47][15:8] = buffer_data_0[3951:3944];
        layer6[47][23:16] = buffer_data_0[3959:3952];
        layer6[47][31:24] = buffer_data_0[3967:3960];
        layer6[47][39:32] = buffer_data_0[3975:3968];
        layer6[47][47:40] = buffer_data_0[3983:3976];
        layer6[47][55:48] = buffer_data_0[3991:3984];
        layer0[48][7:0] = buffer_data_6[3951:3944];
        layer0[48][15:8] = buffer_data_6[3959:3952];
        layer0[48][23:16] = buffer_data_6[3967:3960];
        layer0[48][31:24] = buffer_data_6[3975:3968];
        layer0[48][39:32] = buffer_data_6[3983:3976];
        layer0[48][47:40] = buffer_data_6[3991:3984];
        layer0[48][55:48] = buffer_data_6[3999:3992];
        layer1[48][7:0] = buffer_data_5[3951:3944];
        layer1[48][15:8] = buffer_data_5[3959:3952];
        layer1[48][23:16] = buffer_data_5[3967:3960];
        layer1[48][31:24] = buffer_data_5[3975:3968];
        layer1[48][39:32] = buffer_data_5[3983:3976];
        layer1[48][47:40] = buffer_data_5[3991:3984];
        layer1[48][55:48] = buffer_data_5[3999:3992];
        layer2[48][7:0] = buffer_data_4[3951:3944];
        layer2[48][15:8] = buffer_data_4[3959:3952];
        layer2[48][23:16] = buffer_data_4[3967:3960];
        layer2[48][31:24] = buffer_data_4[3975:3968];
        layer2[48][39:32] = buffer_data_4[3983:3976];
        layer2[48][47:40] = buffer_data_4[3991:3984];
        layer2[48][55:48] = buffer_data_4[3999:3992];
        layer3[48][7:0] = buffer_data_3[3951:3944];
        layer3[48][15:8] = buffer_data_3[3959:3952];
        layer3[48][23:16] = buffer_data_3[3967:3960];
        layer3[48][31:24] = buffer_data_3[3975:3968];
        layer3[48][39:32] = buffer_data_3[3983:3976];
        layer3[48][47:40] = buffer_data_3[3991:3984];
        layer3[48][55:48] = buffer_data_3[3999:3992];
        layer4[48][7:0] = buffer_data_2[3951:3944];
        layer4[48][15:8] = buffer_data_2[3959:3952];
        layer4[48][23:16] = buffer_data_2[3967:3960];
        layer4[48][31:24] = buffer_data_2[3975:3968];
        layer4[48][39:32] = buffer_data_2[3983:3976];
        layer4[48][47:40] = buffer_data_2[3991:3984];
        layer4[48][55:48] = buffer_data_2[3999:3992];
        layer5[48][7:0] = buffer_data_1[3951:3944];
        layer5[48][15:8] = buffer_data_1[3959:3952];
        layer5[48][23:16] = buffer_data_1[3967:3960];
        layer5[48][31:24] = buffer_data_1[3975:3968];
        layer5[48][39:32] = buffer_data_1[3983:3976];
        layer5[48][47:40] = buffer_data_1[3991:3984];
        layer5[48][55:48] = buffer_data_1[3999:3992];
        layer6[48][7:0] = buffer_data_0[3951:3944];
        layer6[48][15:8] = buffer_data_0[3959:3952];
        layer6[48][23:16] = buffer_data_0[3967:3960];
        layer6[48][31:24] = buffer_data_0[3975:3968];
        layer6[48][39:32] = buffer_data_0[3983:3976];
        layer6[48][47:40] = buffer_data_0[3991:3984];
        layer6[48][55:48] = buffer_data_0[3999:3992];
        layer0[49][7:0] = buffer_data_6[3959:3952];
        layer0[49][15:8] = buffer_data_6[3967:3960];
        layer0[49][23:16] = buffer_data_6[3975:3968];
        layer0[49][31:24] = buffer_data_6[3983:3976];
        layer0[49][39:32] = buffer_data_6[3991:3984];
        layer0[49][47:40] = buffer_data_6[3999:3992];
        layer0[49][55:48] = buffer_data_6[4007:4000];
        layer1[49][7:0] = buffer_data_5[3959:3952];
        layer1[49][15:8] = buffer_data_5[3967:3960];
        layer1[49][23:16] = buffer_data_5[3975:3968];
        layer1[49][31:24] = buffer_data_5[3983:3976];
        layer1[49][39:32] = buffer_data_5[3991:3984];
        layer1[49][47:40] = buffer_data_5[3999:3992];
        layer1[49][55:48] = buffer_data_5[4007:4000];
        layer2[49][7:0] = buffer_data_4[3959:3952];
        layer2[49][15:8] = buffer_data_4[3967:3960];
        layer2[49][23:16] = buffer_data_4[3975:3968];
        layer2[49][31:24] = buffer_data_4[3983:3976];
        layer2[49][39:32] = buffer_data_4[3991:3984];
        layer2[49][47:40] = buffer_data_4[3999:3992];
        layer2[49][55:48] = buffer_data_4[4007:4000];
        layer3[49][7:0] = buffer_data_3[3959:3952];
        layer3[49][15:8] = buffer_data_3[3967:3960];
        layer3[49][23:16] = buffer_data_3[3975:3968];
        layer3[49][31:24] = buffer_data_3[3983:3976];
        layer3[49][39:32] = buffer_data_3[3991:3984];
        layer3[49][47:40] = buffer_data_3[3999:3992];
        layer3[49][55:48] = buffer_data_3[4007:4000];
        layer4[49][7:0] = buffer_data_2[3959:3952];
        layer4[49][15:8] = buffer_data_2[3967:3960];
        layer4[49][23:16] = buffer_data_2[3975:3968];
        layer4[49][31:24] = buffer_data_2[3983:3976];
        layer4[49][39:32] = buffer_data_2[3991:3984];
        layer4[49][47:40] = buffer_data_2[3999:3992];
        layer4[49][55:48] = buffer_data_2[4007:4000];
        layer5[49][7:0] = buffer_data_1[3959:3952];
        layer5[49][15:8] = buffer_data_1[3967:3960];
        layer5[49][23:16] = buffer_data_1[3975:3968];
        layer5[49][31:24] = buffer_data_1[3983:3976];
        layer5[49][39:32] = buffer_data_1[3991:3984];
        layer5[49][47:40] = buffer_data_1[3999:3992];
        layer5[49][55:48] = buffer_data_1[4007:4000];
        layer6[49][7:0] = buffer_data_0[3959:3952];
        layer6[49][15:8] = buffer_data_0[3967:3960];
        layer6[49][23:16] = buffer_data_0[3975:3968];
        layer6[49][31:24] = buffer_data_0[3983:3976];
        layer6[49][39:32] = buffer_data_0[3991:3984];
        layer6[49][47:40] = buffer_data_0[3999:3992];
        layer6[49][55:48] = buffer_data_0[4007:4000];
        layer0[50][7:0] = buffer_data_6[3967:3960];
        layer0[50][15:8] = buffer_data_6[3975:3968];
        layer0[50][23:16] = buffer_data_6[3983:3976];
        layer0[50][31:24] = buffer_data_6[3991:3984];
        layer0[50][39:32] = buffer_data_6[3999:3992];
        layer0[50][47:40] = buffer_data_6[4007:4000];
        layer0[50][55:48] = buffer_data_6[4015:4008];
        layer1[50][7:0] = buffer_data_5[3967:3960];
        layer1[50][15:8] = buffer_data_5[3975:3968];
        layer1[50][23:16] = buffer_data_5[3983:3976];
        layer1[50][31:24] = buffer_data_5[3991:3984];
        layer1[50][39:32] = buffer_data_5[3999:3992];
        layer1[50][47:40] = buffer_data_5[4007:4000];
        layer1[50][55:48] = buffer_data_5[4015:4008];
        layer2[50][7:0] = buffer_data_4[3967:3960];
        layer2[50][15:8] = buffer_data_4[3975:3968];
        layer2[50][23:16] = buffer_data_4[3983:3976];
        layer2[50][31:24] = buffer_data_4[3991:3984];
        layer2[50][39:32] = buffer_data_4[3999:3992];
        layer2[50][47:40] = buffer_data_4[4007:4000];
        layer2[50][55:48] = buffer_data_4[4015:4008];
        layer3[50][7:0] = buffer_data_3[3967:3960];
        layer3[50][15:8] = buffer_data_3[3975:3968];
        layer3[50][23:16] = buffer_data_3[3983:3976];
        layer3[50][31:24] = buffer_data_3[3991:3984];
        layer3[50][39:32] = buffer_data_3[3999:3992];
        layer3[50][47:40] = buffer_data_3[4007:4000];
        layer3[50][55:48] = buffer_data_3[4015:4008];
        layer4[50][7:0] = buffer_data_2[3967:3960];
        layer4[50][15:8] = buffer_data_2[3975:3968];
        layer4[50][23:16] = buffer_data_2[3983:3976];
        layer4[50][31:24] = buffer_data_2[3991:3984];
        layer4[50][39:32] = buffer_data_2[3999:3992];
        layer4[50][47:40] = buffer_data_2[4007:4000];
        layer4[50][55:48] = buffer_data_2[4015:4008];
        layer5[50][7:0] = buffer_data_1[3967:3960];
        layer5[50][15:8] = buffer_data_1[3975:3968];
        layer5[50][23:16] = buffer_data_1[3983:3976];
        layer5[50][31:24] = buffer_data_1[3991:3984];
        layer5[50][39:32] = buffer_data_1[3999:3992];
        layer5[50][47:40] = buffer_data_1[4007:4000];
        layer5[50][55:48] = buffer_data_1[4015:4008];
        layer6[50][7:0] = buffer_data_0[3967:3960];
        layer6[50][15:8] = buffer_data_0[3975:3968];
        layer6[50][23:16] = buffer_data_0[3983:3976];
        layer6[50][31:24] = buffer_data_0[3991:3984];
        layer6[50][39:32] = buffer_data_0[3999:3992];
        layer6[50][47:40] = buffer_data_0[4007:4000];
        layer6[50][55:48] = buffer_data_0[4015:4008];
        layer0[51][7:0] = buffer_data_6[3975:3968];
        layer0[51][15:8] = buffer_data_6[3983:3976];
        layer0[51][23:16] = buffer_data_6[3991:3984];
        layer0[51][31:24] = buffer_data_6[3999:3992];
        layer0[51][39:32] = buffer_data_6[4007:4000];
        layer0[51][47:40] = buffer_data_6[4015:4008];
        layer0[51][55:48] = buffer_data_6[4023:4016];
        layer1[51][7:0] = buffer_data_5[3975:3968];
        layer1[51][15:8] = buffer_data_5[3983:3976];
        layer1[51][23:16] = buffer_data_5[3991:3984];
        layer1[51][31:24] = buffer_data_5[3999:3992];
        layer1[51][39:32] = buffer_data_5[4007:4000];
        layer1[51][47:40] = buffer_data_5[4015:4008];
        layer1[51][55:48] = buffer_data_5[4023:4016];
        layer2[51][7:0] = buffer_data_4[3975:3968];
        layer2[51][15:8] = buffer_data_4[3983:3976];
        layer2[51][23:16] = buffer_data_4[3991:3984];
        layer2[51][31:24] = buffer_data_4[3999:3992];
        layer2[51][39:32] = buffer_data_4[4007:4000];
        layer2[51][47:40] = buffer_data_4[4015:4008];
        layer2[51][55:48] = buffer_data_4[4023:4016];
        layer3[51][7:0] = buffer_data_3[3975:3968];
        layer3[51][15:8] = buffer_data_3[3983:3976];
        layer3[51][23:16] = buffer_data_3[3991:3984];
        layer3[51][31:24] = buffer_data_3[3999:3992];
        layer3[51][39:32] = buffer_data_3[4007:4000];
        layer3[51][47:40] = buffer_data_3[4015:4008];
        layer3[51][55:48] = buffer_data_3[4023:4016];
        layer4[51][7:0] = buffer_data_2[3975:3968];
        layer4[51][15:8] = buffer_data_2[3983:3976];
        layer4[51][23:16] = buffer_data_2[3991:3984];
        layer4[51][31:24] = buffer_data_2[3999:3992];
        layer4[51][39:32] = buffer_data_2[4007:4000];
        layer4[51][47:40] = buffer_data_2[4015:4008];
        layer4[51][55:48] = buffer_data_2[4023:4016];
        layer5[51][7:0] = buffer_data_1[3975:3968];
        layer5[51][15:8] = buffer_data_1[3983:3976];
        layer5[51][23:16] = buffer_data_1[3991:3984];
        layer5[51][31:24] = buffer_data_1[3999:3992];
        layer5[51][39:32] = buffer_data_1[4007:4000];
        layer5[51][47:40] = buffer_data_1[4015:4008];
        layer5[51][55:48] = buffer_data_1[4023:4016];
        layer6[51][7:0] = buffer_data_0[3975:3968];
        layer6[51][15:8] = buffer_data_0[3983:3976];
        layer6[51][23:16] = buffer_data_0[3991:3984];
        layer6[51][31:24] = buffer_data_0[3999:3992];
        layer6[51][39:32] = buffer_data_0[4007:4000];
        layer6[51][47:40] = buffer_data_0[4015:4008];
        layer6[51][55:48] = buffer_data_0[4023:4016];
        layer0[52][7:0] = buffer_data_6[3983:3976];
        layer0[52][15:8] = buffer_data_6[3991:3984];
        layer0[52][23:16] = buffer_data_6[3999:3992];
        layer0[52][31:24] = buffer_data_6[4007:4000];
        layer0[52][39:32] = buffer_data_6[4015:4008];
        layer0[52][47:40] = buffer_data_6[4023:4016];
        layer0[52][55:48] = buffer_data_6[4031:4024];
        layer1[52][7:0] = buffer_data_5[3983:3976];
        layer1[52][15:8] = buffer_data_5[3991:3984];
        layer1[52][23:16] = buffer_data_5[3999:3992];
        layer1[52][31:24] = buffer_data_5[4007:4000];
        layer1[52][39:32] = buffer_data_5[4015:4008];
        layer1[52][47:40] = buffer_data_5[4023:4016];
        layer1[52][55:48] = buffer_data_5[4031:4024];
        layer2[52][7:0] = buffer_data_4[3983:3976];
        layer2[52][15:8] = buffer_data_4[3991:3984];
        layer2[52][23:16] = buffer_data_4[3999:3992];
        layer2[52][31:24] = buffer_data_4[4007:4000];
        layer2[52][39:32] = buffer_data_4[4015:4008];
        layer2[52][47:40] = buffer_data_4[4023:4016];
        layer2[52][55:48] = buffer_data_4[4031:4024];
        layer3[52][7:0] = buffer_data_3[3983:3976];
        layer3[52][15:8] = buffer_data_3[3991:3984];
        layer3[52][23:16] = buffer_data_3[3999:3992];
        layer3[52][31:24] = buffer_data_3[4007:4000];
        layer3[52][39:32] = buffer_data_3[4015:4008];
        layer3[52][47:40] = buffer_data_3[4023:4016];
        layer3[52][55:48] = buffer_data_3[4031:4024];
        layer4[52][7:0] = buffer_data_2[3983:3976];
        layer4[52][15:8] = buffer_data_2[3991:3984];
        layer4[52][23:16] = buffer_data_2[3999:3992];
        layer4[52][31:24] = buffer_data_2[4007:4000];
        layer4[52][39:32] = buffer_data_2[4015:4008];
        layer4[52][47:40] = buffer_data_2[4023:4016];
        layer4[52][55:48] = buffer_data_2[4031:4024];
        layer5[52][7:0] = buffer_data_1[3983:3976];
        layer5[52][15:8] = buffer_data_1[3991:3984];
        layer5[52][23:16] = buffer_data_1[3999:3992];
        layer5[52][31:24] = buffer_data_1[4007:4000];
        layer5[52][39:32] = buffer_data_1[4015:4008];
        layer5[52][47:40] = buffer_data_1[4023:4016];
        layer5[52][55:48] = buffer_data_1[4031:4024];
        layer6[52][7:0] = buffer_data_0[3983:3976];
        layer6[52][15:8] = buffer_data_0[3991:3984];
        layer6[52][23:16] = buffer_data_0[3999:3992];
        layer6[52][31:24] = buffer_data_0[4007:4000];
        layer6[52][39:32] = buffer_data_0[4015:4008];
        layer6[52][47:40] = buffer_data_0[4023:4016];
        layer6[52][55:48] = buffer_data_0[4031:4024];
        layer0[53][7:0] = buffer_data_6[3991:3984];
        layer0[53][15:8] = buffer_data_6[3999:3992];
        layer0[53][23:16] = buffer_data_6[4007:4000];
        layer0[53][31:24] = buffer_data_6[4015:4008];
        layer0[53][39:32] = buffer_data_6[4023:4016];
        layer0[53][47:40] = buffer_data_6[4031:4024];
        layer0[53][55:48] = buffer_data_6[4039:4032];
        layer1[53][7:0] = buffer_data_5[3991:3984];
        layer1[53][15:8] = buffer_data_5[3999:3992];
        layer1[53][23:16] = buffer_data_5[4007:4000];
        layer1[53][31:24] = buffer_data_5[4015:4008];
        layer1[53][39:32] = buffer_data_5[4023:4016];
        layer1[53][47:40] = buffer_data_5[4031:4024];
        layer1[53][55:48] = buffer_data_5[4039:4032];
        layer2[53][7:0] = buffer_data_4[3991:3984];
        layer2[53][15:8] = buffer_data_4[3999:3992];
        layer2[53][23:16] = buffer_data_4[4007:4000];
        layer2[53][31:24] = buffer_data_4[4015:4008];
        layer2[53][39:32] = buffer_data_4[4023:4016];
        layer2[53][47:40] = buffer_data_4[4031:4024];
        layer2[53][55:48] = buffer_data_4[4039:4032];
        layer3[53][7:0] = buffer_data_3[3991:3984];
        layer3[53][15:8] = buffer_data_3[3999:3992];
        layer3[53][23:16] = buffer_data_3[4007:4000];
        layer3[53][31:24] = buffer_data_3[4015:4008];
        layer3[53][39:32] = buffer_data_3[4023:4016];
        layer3[53][47:40] = buffer_data_3[4031:4024];
        layer3[53][55:48] = buffer_data_3[4039:4032];
        layer4[53][7:0] = buffer_data_2[3991:3984];
        layer4[53][15:8] = buffer_data_2[3999:3992];
        layer4[53][23:16] = buffer_data_2[4007:4000];
        layer4[53][31:24] = buffer_data_2[4015:4008];
        layer4[53][39:32] = buffer_data_2[4023:4016];
        layer4[53][47:40] = buffer_data_2[4031:4024];
        layer4[53][55:48] = buffer_data_2[4039:4032];
        layer5[53][7:0] = buffer_data_1[3991:3984];
        layer5[53][15:8] = buffer_data_1[3999:3992];
        layer5[53][23:16] = buffer_data_1[4007:4000];
        layer5[53][31:24] = buffer_data_1[4015:4008];
        layer5[53][39:32] = buffer_data_1[4023:4016];
        layer5[53][47:40] = buffer_data_1[4031:4024];
        layer5[53][55:48] = buffer_data_1[4039:4032];
        layer6[53][7:0] = buffer_data_0[3991:3984];
        layer6[53][15:8] = buffer_data_0[3999:3992];
        layer6[53][23:16] = buffer_data_0[4007:4000];
        layer6[53][31:24] = buffer_data_0[4015:4008];
        layer6[53][39:32] = buffer_data_0[4023:4016];
        layer6[53][47:40] = buffer_data_0[4031:4024];
        layer6[53][55:48] = buffer_data_0[4039:4032];
        layer0[54][7:0] = buffer_data_6[3999:3992];
        layer0[54][15:8] = buffer_data_6[4007:4000];
        layer0[54][23:16] = buffer_data_6[4015:4008];
        layer0[54][31:24] = buffer_data_6[4023:4016];
        layer0[54][39:32] = buffer_data_6[4031:4024];
        layer0[54][47:40] = buffer_data_6[4039:4032];
        layer0[54][55:48] = buffer_data_6[4047:4040];
        layer1[54][7:0] = buffer_data_5[3999:3992];
        layer1[54][15:8] = buffer_data_5[4007:4000];
        layer1[54][23:16] = buffer_data_5[4015:4008];
        layer1[54][31:24] = buffer_data_5[4023:4016];
        layer1[54][39:32] = buffer_data_5[4031:4024];
        layer1[54][47:40] = buffer_data_5[4039:4032];
        layer1[54][55:48] = buffer_data_5[4047:4040];
        layer2[54][7:0] = buffer_data_4[3999:3992];
        layer2[54][15:8] = buffer_data_4[4007:4000];
        layer2[54][23:16] = buffer_data_4[4015:4008];
        layer2[54][31:24] = buffer_data_4[4023:4016];
        layer2[54][39:32] = buffer_data_4[4031:4024];
        layer2[54][47:40] = buffer_data_4[4039:4032];
        layer2[54][55:48] = buffer_data_4[4047:4040];
        layer3[54][7:0] = buffer_data_3[3999:3992];
        layer3[54][15:8] = buffer_data_3[4007:4000];
        layer3[54][23:16] = buffer_data_3[4015:4008];
        layer3[54][31:24] = buffer_data_3[4023:4016];
        layer3[54][39:32] = buffer_data_3[4031:4024];
        layer3[54][47:40] = buffer_data_3[4039:4032];
        layer3[54][55:48] = buffer_data_3[4047:4040];
        layer4[54][7:0] = buffer_data_2[3999:3992];
        layer4[54][15:8] = buffer_data_2[4007:4000];
        layer4[54][23:16] = buffer_data_2[4015:4008];
        layer4[54][31:24] = buffer_data_2[4023:4016];
        layer4[54][39:32] = buffer_data_2[4031:4024];
        layer4[54][47:40] = buffer_data_2[4039:4032];
        layer4[54][55:48] = buffer_data_2[4047:4040];
        layer5[54][7:0] = buffer_data_1[3999:3992];
        layer5[54][15:8] = buffer_data_1[4007:4000];
        layer5[54][23:16] = buffer_data_1[4015:4008];
        layer5[54][31:24] = buffer_data_1[4023:4016];
        layer5[54][39:32] = buffer_data_1[4031:4024];
        layer5[54][47:40] = buffer_data_1[4039:4032];
        layer5[54][55:48] = buffer_data_1[4047:4040];
        layer6[54][7:0] = buffer_data_0[3999:3992];
        layer6[54][15:8] = buffer_data_0[4007:4000];
        layer6[54][23:16] = buffer_data_0[4015:4008];
        layer6[54][31:24] = buffer_data_0[4023:4016];
        layer6[54][39:32] = buffer_data_0[4031:4024];
        layer6[54][47:40] = buffer_data_0[4039:4032];
        layer6[54][55:48] = buffer_data_0[4047:4040];
        layer0[55][7:0] = buffer_data_6[4007:4000];
        layer0[55][15:8] = buffer_data_6[4015:4008];
        layer0[55][23:16] = buffer_data_6[4023:4016];
        layer0[55][31:24] = buffer_data_6[4031:4024];
        layer0[55][39:32] = buffer_data_6[4039:4032];
        layer0[55][47:40] = buffer_data_6[4047:4040];
        layer0[55][55:48] = buffer_data_6[4055:4048];
        layer1[55][7:0] = buffer_data_5[4007:4000];
        layer1[55][15:8] = buffer_data_5[4015:4008];
        layer1[55][23:16] = buffer_data_5[4023:4016];
        layer1[55][31:24] = buffer_data_5[4031:4024];
        layer1[55][39:32] = buffer_data_5[4039:4032];
        layer1[55][47:40] = buffer_data_5[4047:4040];
        layer1[55][55:48] = buffer_data_5[4055:4048];
        layer2[55][7:0] = buffer_data_4[4007:4000];
        layer2[55][15:8] = buffer_data_4[4015:4008];
        layer2[55][23:16] = buffer_data_4[4023:4016];
        layer2[55][31:24] = buffer_data_4[4031:4024];
        layer2[55][39:32] = buffer_data_4[4039:4032];
        layer2[55][47:40] = buffer_data_4[4047:4040];
        layer2[55][55:48] = buffer_data_4[4055:4048];
        layer3[55][7:0] = buffer_data_3[4007:4000];
        layer3[55][15:8] = buffer_data_3[4015:4008];
        layer3[55][23:16] = buffer_data_3[4023:4016];
        layer3[55][31:24] = buffer_data_3[4031:4024];
        layer3[55][39:32] = buffer_data_3[4039:4032];
        layer3[55][47:40] = buffer_data_3[4047:4040];
        layer3[55][55:48] = buffer_data_3[4055:4048];
        layer4[55][7:0] = buffer_data_2[4007:4000];
        layer4[55][15:8] = buffer_data_2[4015:4008];
        layer4[55][23:16] = buffer_data_2[4023:4016];
        layer4[55][31:24] = buffer_data_2[4031:4024];
        layer4[55][39:32] = buffer_data_2[4039:4032];
        layer4[55][47:40] = buffer_data_2[4047:4040];
        layer4[55][55:48] = buffer_data_2[4055:4048];
        layer5[55][7:0] = buffer_data_1[4007:4000];
        layer5[55][15:8] = buffer_data_1[4015:4008];
        layer5[55][23:16] = buffer_data_1[4023:4016];
        layer5[55][31:24] = buffer_data_1[4031:4024];
        layer5[55][39:32] = buffer_data_1[4039:4032];
        layer5[55][47:40] = buffer_data_1[4047:4040];
        layer5[55][55:48] = buffer_data_1[4055:4048];
        layer6[55][7:0] = buffer_data_0[4007:4000];
        layer6[55][15:8] = buffer_data_0[4015:4008];
        layer6[55][23:16] = buffer_data_0[4023:4016];
        layer6[55][31:24] = buffer_data_0[4031:4024];
        layer6[55][39:32] = buffer_data_0[4039:4032];
        layer6[55][47:40] = buffer_data_0[4047:4040];
        layer6[55][55:48] = buffer_data_0[4055:4048];
        layer0[56][7:0] = buffer_data_6[4015:4008];
        layer0[56][15:8] = buffer_data_6[4023:4016];
        layer0[56][23:16] = buffer_data_6[4031:4024];
        layer0[56][31:24] = buffer_data_6[4039:4032];
        layer0[56][39:32] = buffer_data_6[4047:4040];
        layer0[56][47:40] = buffer_data_6[4055:4048];
        layer0[56][55:48] = buffer_data_6[4063:4056];
        layer1[56][7:0] = buffer_data_5[4015:4008];
        layer1[56][15:8] = buffer_data_5[4023:4016];
        layer1[56][23:16] = buffer_data_5[4031:4024];
        layer1[56][31:24] = buffer_data_5[4039:4032];
        layer1[56][39:32] = buffer_data_5[4047:4040];
        layer1[56][47:40] = buffer_data_5[4055:4048];
        layer1[56][55:48] = buffer_data_5[4063:4056];
        layer2[56][7:0] = buffer_data_4[4015:4008];
        layer2[56][15:8] = buffer_data_4[4023:4016];
        layer2[56][23:16] = buffer_data_4[4031:4024];
        layer2[56][31:24] = buffer_data_4[4039:4032];
        layer2[56][39:32] = buffer_data_4[4047:4040];
        layer2[56][47:40] = buffer_data_4[4055:4048];
        layer2[56][55:48] = buffer_data_4[4063:4056];
        layer3[56][7:0] = buffer_data_3[4015:4008];
        layer3[56][15:8] = buffer_data_3[4023:4016];
        layer3[56][23:16] = buffer_data_3[4031:4024];
        layer3[56][31:24] = buffer_data_3[4039:4032];
        layer3[56][39:32] = buffer_data_3[4047:4040];
        layer3[56][47:40] = buffer_data_3[4055:4048];
        layer3[56][55:48] = buffer_data_3[4063:4056];
        layer4[56][7:0] = buffer_data_2[4015:4008];
        layer4[56][15:8] = buffer_data_2[4023:4016];
        layer4[56][23:16] = buffer_data_2[4031:4024];
        layer4[56][31:24] = buffer_data_2[4039:4032];
        layer4[56][39:32] = buffer_data_2[4047:4040];
        layer4[56][47:40] = buffer_data_2[4055:4048];
        layer4[56][55:48] = buffer_data_2[4063:4056];
        layer5[56][7:0] = buffer_data_1[4015:4008];
        layer5[56][15:8] = buffer_data_1[4023:4016];
        layer5[56][23:16] = buffer_data_1[4031:4024];
        layer5[56][31:24] = buffer_data_1[4039:4032];
        layer5[56][39:32] = buffer_data_1[4047:4040];
        layer5[56][47:40] = buffer_data_1[4055:4048];
        layer5[56][55:48] = buffer_data_1[4063:4056];
        layer6[56][7:0] = buffer_data_0[4015:4008];
        layer6[56][15:8] = buffer_data_0[4023:4016];
        layer6[56][23:16] = buffer_data_0[4031:4024];
        layer6[56][31:24] = buffer_data_0[4039:4032];
        layer6[56][39:32] = buffer_data_0[4047:4040];
        layer6[56][47:40] = buffer_data_0[4055:4048];
        layer6[56][55:48] = buffer_data_0[4063:4056];
        layer0[57][7:0] = buffer_data_6[4023:4016];
        layer0[57][15:8] = buffer_data_6[4031:4024];
        layer0[57][23:16] = buffer_data_6[4039:4032];
        layer0[57][31:24] = buffer_data_6[4047:4040];
        layer0[57][39:32] = buffer_data_6[4055:4048];
        layer0[57][47:40] = buffer_data_6[4063:4056];
        layer0[57][55:48] = buffer_data_6[4071:4064];
        layer1[57][7:0] = buffer_data_5[4023:4016];
        layer1[57][15:8] = buffer_data_5[4031:4024];
        layer1[57][23:16] = buffer_data_5[4039:4032];
        layer1[57][31:24] = buffer_data_5[4047:4040];
        layer1[57][39:32] = buffer_data_5[4055:4048];
        layer1[57][47:40] = buffer_data_5[4063:4056];
        layer1[57][55:48] = buffer_data_5[4071:4064];
        layer2[57][7:0] = buffer_data_4[4023:4016];
        layer2[57][15:8] = buffer_data_4[4031:4024];
        layer2[57][23:16] = buffer_data_4[4039:4032];
        layer2[57][31:24] = buffer_data_4[4047:4040];
        layer2[57][39:32] = buffer_data_4[4055:4048];
        layer2[57][47:40] = buffer_data_4[4063:4056];
        layer2[57][55:48] = buffer_data_4[4071:4064];
        layer3[57][7:0] = buffer_data_3[4023:4016];
        layer3[57][15:8] = buffer_data_3[4031:4024];
        layer3[57][23:16] = buffer_data_3[4039:4032];
        layer3[57][31:24] = buffer_data_3[4047:4040];
        layer3[57][39:32] = buffer_data_3[4055:4048];
        layer3[57][47:40] = buffer_data_3[4063:4056];
        layer3[57][55:48] = buffer_data_3[4071:4064];
        layer4[57][7:0] = buffer_data_2[4023:4016];
        layer4[57][15:8] = buffer_data_2[4031:4024];
        layer4[57][23:16] = buffer_data_2[4039:4032];
        layer4[57][31:24] = buffer_data_2[4047:4040];
        layer4[57][39:32] = buffer_data_2[4055:4048];
        layer4[57][47:40] = buffer_data_2[4063:4056];
        layer4[57][55:48] = buffer_data_2[4071:4064];
        layer5[57][7:0] = buffer_data_1[4023:4016];
        layer5[57][15:8] = buffer_data_1[4031:4024];
        layer5[57][23:16] = buffer_data_1[4039:4032];
        layer5[57][31:24] = buffer_data_1[4047:4040];
        layer5[57][39:32] = buffer_data_1[4055:4048];
        layer5[57][47:40] = buffer_data_1[4063:4056];
        layer5[57][55:48] = buffer_data_1[4071:4064];
        layer6[57][7:0] = buffer_data_0[4023:4016];
        layer6[57][15:8] = buffer_data_0[4031:4024];
        layer6[57][23:16] = buffer_data_0[4039:4032];
        layer6[57][31:24] = buffer_data_0[4047:4040];
        layer6[57][39:32] = buffer_data_0[4055:4048];
        layer6[57][47:40] = buffer_data_0[4063:4056];
        layer6[57][55:48] = buffer_data_0[4071:4064];
        layer0[58][7:0] = buffer_data_6[4031:4024];
        layer0[58][15:8] = buffer_data_6[4039:4032];
        layer0[58][23:16] = buffer_data_6[4047:4040];
        layer0[58][31:24] = buffer_data_6[4055:4048];
        layer0[58][39:32] = buffer_data_6[4063:4056];
        layer0[58][47:40] = buffer_data_6[4071:4064];
        layer0[58][55:48] = buffer_data_6[4079:4072];
        layer1[58][7:0] = buffer_data_5[4031:4024];
        layer1[58][15:8] = buffer_data_5[4039:4032];
        layer1[58][23:16] = buffer_data_5[4047:4040];
        layer1[58][31:24] = buffer_data_5[4055:4048];
        layer1[58][39:32] = buffer_data_5[4063:4056];
        layer1[58][47:40] = buffer_data_5[4071:4064];
        layer1[58][55:48] = buffer_data_5[4079:4072];
        layer2[58][7:0] = buffer_data_4[4031:4024];
        layer2[58][15:8] = buffer_data_4[4039:4032];
        layer2[58][23:16] = buffer_data_4[4047:4040];
        layer2[58][31:24] = buffer_data_4[4055:4048];
        layer2[58][39:32] = buffer_data_4[4063:4056];
        layer2[58][47:40] = buffer_data_4[4071:4064];
        layer2[58][55:48] = buffer_data_4[4079:4072];
        layer3[58][7:0] = buffer_data_3[4031:4024];
        layer3[58][15:8] = buffer_data_3[4039:4032];
        layer3[58][23:16] = buffer_data_3[4047:4040];
        layer3[58][31:24] = buffer_data_3[4055:4048];
        layer3[58][39:32] = buffer_data_3[4063:4056];
        layer3[58][47:40] = buffer_data_3[4071:4064];
        layer3[58][55:48] = buffer_data_3[4079:4072];
        layer4[58][7:0] = buffer_data_2[4031:4024];
        layer4[58][15:8] = buffer_data_2[4039:4032];
        layer4[58][23:16] = buffer_data_2[4047:4040];
        layer4[58][31:24] = buffer_data_2[4055:4048];
        layer4[58][39:32] = buffer_data_2[4063:4056];
        layer4[58][47:40] = buffer_data_2[4071:4064];
        layer4[58][55:48] = buffer_data_2[4079:4072];
        layer5[58][7:0] = buffer_data_1[4031:4024];
        layer5[58][15:8] = buffer_data_1[4039:4032];
        layer5[58][23:16] = buffer_data_1[4047:4040];
        layer5[58][31:24] = buffer_data_1[4055:4048];
        layer5[58][39:32] = buffer_data_1[4063:4056];
        layer5[58][47:40] = buffer_data_1[4071:4064];
        layer5[58][55:48] = buffer_data_1[4079:4072];
        layer6[58][7:0] = buffer_data_0[4031:4024];
        layer6[58][15:8] = buffer_data_0[4039:4032];
        layer6[58][23:16] = buffer_data_0[4047:4040];
        layer6[58][31:24] = buffer_data_0[4055:4048];
        layer6[58][39:32] = buffer_data_0[4063:4056];
        layer6[58][47:40] = buffer_data_0[4071:4064];
        layer6[58][55:48] = buffer_data_0[4079:4072];
        layer0[59][7:0] = buffer_data_6[4039:4032];
        layer0[59][15:8] = buffer_data_6[4047:4040];
        layer0[59][23:16] = buffer_data_6[4055:4048];
        layer0[59][31:24] = buffer_data_6[4063:4056];
        layer0[59][39:32] = buffer_data_6[4071:4064];
        layer0[59][47:40] = buffer_data_6[4079:4072];
        layer0[59][55:48] = buffer_data_6[4087:4080];
        layer1[59][7:0] = buffer_data_5[4039:4032];
        layer1[59][15:8] = buffer_data_5[4047:4040];
        layer1[59][23:16] = buffer_data_5[4055:4048];
        layer1[59][31:24] = buffer_data_5[4063:4056];
        layer1[59][39:32] = buffer_data_5[4071:4064];
        layer1[59][47:40] = buffer_data_5[4079:4072];
        layer1[59][55:48] = buffer_data_5[4087:4080];
        layer2[59][7:0] = buffer_data_4[4039:4032];
        layer2[59][15:8] = buffer_data_4[4047:4040];
        layer2[59][23:16] = buffer_data_4[4055:4048];
        layer2[59][31:24] = buffer_data_4[4063:4056];
        layer2[59][39:32] = buffer_data_4[4071:4064];
        layer2[59][47:40] = buffer_data_4[4079:4072];
        layer2[59][55:48] = buffer_data_4[4087:4080];
        layer3[59][7:0] = buffer_data_3[4039:4032];
        layer3[59][15:8] = buffer_data_3[4047:4040];
        layer3[59][23:16] = buffer_data_3[4055:4048];
        layer3[59][31:24] = buffer_data_3[4063:4056];
        layer3[59][39:32] = buffer_data_3[4071:4064];
        layer3[59][47:40] = buffer_data_3[4079:4072];
        layer3[59][55:48] = buffer_data_3[4087:4080];
        layer4[59][7:0] = buffer_data_2[4039:4032];
        layer4[59][15:8] = buffer_data_2[4047:4040];
        layer4[59][23:16] = buffer_data_2[4055:4048];
        layer4[59][31:24] = buffer_data_2[4063:4056];
        layer4[59][39:32] = buffer_data_2[4071:4064];
        layer4[59][47:40] = buffer_data_2[4079:4072];
        layer4[59][55:48] = buffer_data_2[4087:4080];
        layer5[59][7:0] = buffer_data_1[4039:4032];
        layer5[59][15:8] = buffer_data_1[4047:4040];
        layer5[59][23:16] = buffer_data_1[4055:4048];
        layer5[59][31:24] = buffer_data_1[4063:4056];
        layer5[59][39:32] = buffer_data_1[4071:4064];
        layer5[59][47:40] = buffer_data_1[4079:4072];
        layer5[59][55:48] = buffer_data_1[4087:4080];
        layer6[59][7:0] = buffer_data_0[4039:4032];
        layer6[59][15:8] = buffer_data_0[4047:4040];
        layer6[59][23:16] = buffer_data_0[4055:4048];
        layer6[59][31:24] = buffer_data_0[4063:4056];
        layer6[59][39:32] = buffer_data_0[4071:4064];
        layer6[59][47:40] = buffer_data_0[4079:4072];
        layer6[59][55:48] = buffer_data_0[4087:4080];
        layer0[60][7:0] = buffer_data_6[4047:4040];
        layer0[60][15:8] = buffer_data_6[4055:4048];
        layer0[60][23:16] = buffer_data_6[4063:4056];
        layer0[60][31:24] = buffer_data_6[4071:4064];
        layer0[60][39:32] = buffer_data_6[4079:4072];
        layer0[60][47:40] = buffer_data_6[4087:4080];
        layer0[60][55:48] = buffer_data_6[4095:4088];
        layer1[60][7:0] = buffer_data_5[4047:4040];
        layer1[60][15:8] = buffer_data_5[4055:4048];
        layer1[60][23:16] = buffer_data_5[4063:4056];
        layer1[60][31:24] = buffer_data_5[4071:4064];
        layer1[60][39:32] = buffer_data_5[4079:4072];
        layer1[60][47:40] = buffer_data_5[4087:4080];
        layer1[60][55:48] = buffer_data_5[4095:4088];
        layer2[60][7:0] = buffer_data_4[4047:4040];
        layer2[60][15:8] = buffer_data_4[4055:4048];
        layer2[60][23:16] = buffer_data_4[4063:4056];
        layer2[60][31:24] = buffer_data_4[4071:4064];
        layer2[60][39:32] = buffer_data_4[4079:4072];
        layer2[60][47:40] = buffer_data_4[4087:4080];
        layer2[60][55:48] = buffer_data_4[4095:4088];
        layer3[60][7:0] = buffer_data_3[4047:4040];
        layer3[60][15:8] = buffer_data_3[4055:4048];
        layer3[60][23:16] = buffer_data_3[4063:4056];
        layer3[60][31:24] = buffer_data_3[4071:4064];
        layer3[60][39:32] = buffer_data_3[4079:4072];
        layer3[60][47:40] = buffer_data_3[4087:4080];
        layer3[60][55:48] = buffer_data_3[4095:4088];
        layer4[60][7:0] = buffer_data_2[4047:4040];
        layer4[60][15:8] = buffer_data_2[4055:4048];
        layer4[60][23:16] = buffer_data_2[4063:4056];
        layer4[60][31:24] = buffer_data_2[4071:4064];
        layer4[60][39:32] = buffer_data_2[4079:4072];
        layer4[60][47:40] = buffer_data_2[4087:4080];
        layer4[60][55:48] = buffer_data_2[4095:4088];
        layer5[60][7:0] = buffer_data_1[4047:4040];
        layer5[60][15:8] = buffer_data_1[4055:4048];
        layer5[60][23:16] = buffer_data_1[4063:4056];
        layer5[60][31:24] = buffer_data_1[4071:4064];
        layer5[60][39:32] = buffer_data_1[4079:4072];
        layer5[60][47:40] = buffer_data_1[4087:4080];
        layer5[60][55:48] = buffer_data_1[4095:4088];
        layer6[60][7:0] = buffer_data_0[4047:4040];
        layer6[60][15:8] = buffer_data_0[4055:4048];
        layer6[60][23:16] = buffer_data_0[4063:4056];
        layer6[60][31:24] = buffer_data_0[4071:4064];
        layer6[60][39:32] = buffer_data_0[4079:4072];
        layer6[60][47:40] = buffer_data_0[4087:4080];
        layer6[60][55:48] = buffer_data_0[4095:4088];
        layer0[61][7:0] = buffer_data_6[4055:4048];
        layer0[61][15:8] = buffer_data_6[4063:4056];
        layer0[61][23:16] = buffer_data_6[4071:4064];
        layer0[61][31:24] = buffer_data_6[4079:4072];
        layer0[61][39:32] = buffer_data_6[4087:4080];
        layer0[61][47:40] = buffer_data_6[4095:4088];
        layer0[61][55:48] = buffer_data_6[4103:4096];
        layer1[61][7:0] = buffer_data_5[4055:4048];
        layer1[61][15:8] = buffer_data_5[4063:4056];
        layer1[61][23:16] = buffer_data_5[4071:4064];
        layer1[61][31:24] = buffer_data_5[4079:4072];
        layer1[61][39:32] = buffer_data_5[4087:4080];
        layer1[61][47:40] = buffer_data_5[4095:4088];
        layer1[61][55:48] = buffer_data_5[4103:4096];
        layer2[61][7:0] = buffer_data_4[4055:4048];
        layer2[61][15:8] = buffer_data_4[4063:4056];
        layer2[61][23:16] = buffer_data_4[4071:4064];
        layer2[61][31:24] = buffer_data_4[4079:4072];
        layer2[61][39:32] = buffer_data_4[4087:4080];
        layer2[61][47:40] = buffer_data_4[4095:4088];
        layer2[61][55:48] = buffer_data_4[4103:4096];
        layer3[61][7:0] = buffer_data_3[4055:4048];
        layer3[61][15:8] = buffer_data_3[4063:4056];
        layer3[61][23:16] = buffer_data_3[4071:4064];
        layer3[61][31:24] = buffer_data_3[4079:4072];
        layer3[61][39:32] = buffer_data_3[4087:4080];
        layer3[61][47:40] = buffer_data_3[4095:4088];
        layer3[61][55:48] = buffer_data_3[4103:4096];
        layer4[61][7:0] = buffer_data_2[4055:4048];
        layer4[61][15:8] = buffer_data_2[4063:4056];
        layer4[61][23:16] = buffer_data_2[4071:4064];
        layer4[61][31:24] = buffer_data_2[4079:4072];
        layer4[61][39:32] = buffer_data_2[4087:4080];
        layer4[61][47:40] = buffer_data_2[4095:4088];
        layer4[61][55:48] = buffer_data_2[4103:4096];
        layer5[61][7:0] = buffer_data_1[4055:4048];
        layer5[61][15:8] = buffer_data_1[4063:4056];
        layer5[61][23:16] = buffer_data_1[4071:4064];
        layer5[61][31:24] = buffer_data_1[4079:4072];
        layer5[61][39:32] = buffer_data_1[4087:4080];
        layer5[61][47:40] = buffer_data_1[4095:4088];
        layer5[61][55:48] = buffer_data_1[4103:4096];
        layer6[61][7:0] = buffer_data_0[4055:4048];
        layer6[61][15:8] = buffer_data_0[4063:4056];
        layer6[61][23:16] = buffer_data_0[4071:4064];
        layer6[61][31:24] = buffer_data_0[4079:4072];
        layer6[61][39:32] = buffer_data_0[4087:4080];
        layer6[61][47:40] = buffer_data_0[4095:4088];
        layer6[61][55:48] = buffer_data_0[4103:4096];
        layer0[62][7:0] = buffer_data_6[4063:4056];
        layer0[62][15:8] = buffer_data_6[4071:4064];
        layer0[62][23:16] = buffer_data_6[4079:4072];
        layer0[62][31:24] = buffer_data_6[4087:4080];
        layer0[62][39:32] = buffer_data_6[4095:4088];
        layer0[62][47:40] = buffer_data_6[4103:4096];
        layer0[62][55:48] = buffer_data_6[4111:4104];
        layer1[62][7:0] = buffer_data_5[4063:4056];
        layer1[62][15:8] = buffer_data_5[4071:4064];
        layer1[62][23:16] = buffer_data_5[4079:4072];
        layer1[62][31:24] = buffer_data_5[4087:4080];
        layer1[62][39:32] = buffer_data_5[4095:4088];
        layer1[62][47:40] = buffer_data_5[4103:4096];
        layer1[62][55:48] = buffer_data_5[4111:4104];
        layer2[62][7:0] = buffer_data_4[4063:4056];
        layer2[62][15:8] = buffer_data_4[4071:4064];
        layer2[62][23:16] = buffer_data_4[4079:4072];
        layer2[62][31:24] = buffer_data_4[4087:4080];
        layer2[62][39:32] = buffer_data_4[4095:4088];
        layer2[62][47:40] = buffer_data_4[4103:4096];
        layer2[62][55:48] = buffer_data_4[4111:4104];
        layer3[62][7:0] = buffer_data_3[4063:4056];
        layer3[62][15:8] = buffer_data_3[4071:4064];
        layer3[62][23:16] = buffer_data_3[4079:4072];
        layer3[62][31:24] = buffer_data_3[4087:4080];
        layer3[62][39:32] = buffer_data_3[4095:4088];
        layer3[62][47:40] = buffer_data_3[4103:4096];
        layer3[62][55:48] = buffer_data_3[4111:4104];
        layer4[62][7:0] = buffer_data_2[4063:4056];
        layer4[62][15:8] = buffer_data_2[4071:4064];
        layer4[62][23:16] = buffer_data_2[4079:4072];
        layer4[62][31:24] = buffer_data_2[4087:4080];
        layer4[62][39:32] = buffer_data_2[4095:4088];
        layer4[62][47:40] = buffer_data_2[4103:4096];
        layer4[62][55:48] = buffer_data_2[4111:4104];
        layer5[62][7:0] = buffer_data_1[4063:4056];
        layer5[62][15:8] = buffer_data_1[4071:4064];
        layer5[62][23:16] = buffer_data_1[4079:4072];
        layer5[62][31:24] = buffer_data_1[4087:4080];
        layer5[62][39:32] = buffer_data_1[4095:4088];
        layer5[62][47:40] = buffer_data_1[4103:4096];
        layer5[62][55:48] = buffer_data_1[4111:4104];
        layer6[62][7:0] = buffer_data_0[4063:4056];
        layer6[62][15:8] = buffer_data_0[4071:4064];
        layer6[62][23:16] = buffer_data_0[4079:4072];
        layer6[62][31:24] = buffer_data_0[4087:4080];
        layer6[62][39:32] = buffer_data_0[4095:4088];
        layer6[62][47:40] = buffer_data_0[4103:4096];
        layer6[62][55:48] = buffer_data_0[4111:4104];
        layer0[63][7:0] = buffer_data_6[4071:4064];
        layer0[63][15:8] = buffer_data_6[4079:4072];
        layer0[63][23:16] = buffer_data_6[4087:4080];
        layer0[63][31:24] = buffer_data_6[4095:4088];
        layer0[63][39:32] = buffer_data_6[4103:4096];
        layer0[63][47:40] = buffer_data_6[4111:4104];
        layer0[63][55:48] = buffer_data_6[4119:4112];
        layer1[63][7:0] = buffer_data_5[4071:4064];
        layer1[63][15:8] = buffer_data_5[4079:4072];
        layer1[63][23:16] = buffer_data_5[4087:4080];
        layer1[63][31:24] = buffer_data_5[4095:4088];
        layer1[63][39:32] = buffer_data_5[4103:4096];
        layer1[63][47:40] = buffer_data_5[4111:4104];
        layer1[63][55:48] = buffer_data_5[4119:4112];
        layer2[63][7:0] = buffer_data_4[4071:4064];
        layer2[63][15:8] = buffer_data_4[4079:4072];
        layer2[63][23:16] = buffer_data_4[4087:4080];
        layer2[63][31:24] = buffer_data_4[4095:4088];
        layer2[63][39:32] = buffer_data_4[4103:4096];
        layer2[63][47:40] = buffer_data_4[4111:4104];
        layer2[63][55:48] = buffer_data_4[4119:4112];
        layer3[63][7:0] = buffer_data_3[4071:4064];
        layer3[63][15:8] = buffer_data_3[4079:4072];
        layer3[63][23:16] = buffer_data_3[4087:4080];
        layer3[63][31:24] = buffer_data_3[4095:4088];
        layer3[63][39:32] = buffer_data_3[4103:4096];
        layer3[63][47:40] = buffer_data_3[4111:4104];
        layer3[63][55:48] = buffer_data_3[4119:4112];
        layer4[63][7:0] = buffer_data_2[4071:4064];
        layer4[63][15:8] = buffer_data_2[4079:4072];
        layer4[63][23:16] = buffer_data_2[4087:4080];
        layer4[63][31:24] = buffer_data_2[4095:4088];
        layer4[63][39:32] = buffer_data_2[4103:4096];
        layer4[63][47:40] = buffer_data_2[4111:4104];
        layer4[63][55:48] = buffer_data_2[4119:4112];
        layer5[63][7:0] = buffer_data_1[4071:4064];
        layer5[63][15:8] = buffer_data_1[4079:4072];
        layer5[63][23:16] = buffer_data_1[4087:4080];
        layer5[63][31:24] = buffer_data_1[4095:4088];
        layer5[63][39:32] = buffer_data_1[4103:4096];
        layer5[63][47:40] = buffer_data_1[4111:4104];
        layer5[63][55:48] = buffer_data_1[4119:4112];
        layer6[63][7:0] = buffer_data_0[4071:4064];
        layer6[63][15:8] = buffer_data_0[4079:4072];
        layer6[63][23:16] = buffer_data_0[4087:4080];
        layer6[63][31:24] = buffer_data_0[4095:4088];
        layer6[63][39:32] = buffer_data_0[4103:4096];
        layer6[63][47:40] = buffer_data_0[4111:4104];
        layer6[63][55:48] = buffer_data_0[4119:4112];
    end
    ST_GAUSSIAN_8: begin
        layer0[0][7:0] = buffer_data_6[4079:4072];
        layer0[0][15:8] = buffer_data_6[4087:4080];
        layer0[0][23:16] = buffer_data_6[4095:4088];
        layer0[0][31:24] = buffer_data_6[4103:4096];
        layer0[0][39:32] = buffer_data_6[4111:4104];
        layer0[0][47:40] = buffer_data_6[4119:4112];
        layer0[0][55:48] = buffer_data_6[4127:4120];
        layer1[0][7:0] = buffer_data_5[4079:4072];
        layer1[0][15:8] = buffer_data_5[4087:4080];
        layer1[0][23:16] = buffer_data_5[4095:4088];
        layer1[0][31:24] = buffer_data_5[4103:4096];
        layer1[0][39:32] = buffer_data_5[4111:4104];
        layer1[0][47:40] = buffer_data_5[4119:4112];
        layer1[0][55:48] = buffer_data_5[4127:4120];
        layer2[0][7:0] = buffer_data_4[4079:4072];
        layer2[0][15:8] = buffer_data_4[4087:4080];
        layer2[0][23:16] = buffer_data_4[4095:4088];
        layer2[0][31:24] = buffer_data_4[4103:4096];
        layer2[0][39:32] = buffer_data_4[4111:4104];
        layer2[0][47:40] = buffer_data_4[4119:4112];
        layer2[0][55:48] = buffer_data_4[4127:4120];
        layer3[0][7:0] = buffer_data_3[4079:4072];
        layer3[0][15:8] = buffer_data_3[4087:4080];
        layer3[0][23:16] = buffer_data_3[4095:4088];
        layer3[0][31:24] = buffer_data_3[4103:4096];
        layer3[0][39:32] = buffer_data_3[4111:4104];
        layer3[0][47:40] = buffer_data_3[4119:4112];
        layer3[0][55:48] = buffer_data_3[4127:4120];
        layer4[0][7:0] = buffer_data_2[4079:4072];
        layer4[0][15:8] = buffer_data_2[4087:4080];
        layer4[0][23:16] = buffer_data_2[4095:4088];
        layer4[0][31:24] = buffer_data_2[4103:4096];
        layer4[0][39:32] = buffer_data_2[4111:4104];
        layer4[0][47:40] = buffer_data_2[4119:4112];
        layer4[0][55:48] = buffer_data_2[4127:4120];
        layer5[0][7:0] = buffer_data_1[4079:4072];
        layer5[0][15:8] = buffer_data_1[4087:4080];
        layer5[0][23:16] = buffer_data_1[4095:4088];
        layer5[0][31:24] = buffer_data_1[4103:4096];
        layer5[0][39:32] = buffer_data_1[4111:4104];
        layer5[0][47:40] = buffer_data_1[4119:4112];
        layer5[0][55:48] = buffer_data_1[4127:4120];
        layer6[0][7:0] = buffer_data_0[4079:4072];
        layer6[0][15:8] = buffer_data_0[4087:4080];
        layer6[0][23:16] = buffer_data_0[4095:4088];
        layer6[0][31:24] = buffer_data_0[4103:4096];
        layer6[0][39:32] = buffer_data_0[4111:4104];
        layer6[0][47:40] = buffer_data_0[4119:4112];
        layer6[0][55:48] = buffer_data_0[4127:4120];
        layer0[1][7:0] = buffer_data_6[4087:4080];
        layer0[1][15:8] = buffer_data_6[4095:4088];
        layer0[1][23:16] = buffer_data_6[4103:4096];
        layer0[1][31:24] = buffer_data_6[4111:4104];
        layer0[1][39:32] = buffer_data_6[4119:4112];
        layer0[1][47:40] = buffer_data_6[4127:4120];
        layer0[1][55:48] = buffer_data_6[4135:4128];
        layer1[1][7:0] = buffer_data_5[4087:4080];
        layer1[1][15:8] = buffer_data_5[4095:4088];
        layer1[1][23:16] = buffer_data_5[4103:4096];
        layer1[1][31:24] = buffer_data_5[4111:4104];
        layer1[1][39:32] = buffer_data_5[4119:4112];
        layer1[1][47:40] = buffer_data_5[4127:4120];
        layer1[1][55:48] = buffer_data_5[4135:4128];
        layer2[1][7:0] = buffer_data_4[4087:4080];
        layer2[1][15:8] = buffer_data_4[4095:4088];
        layer2[1][23:16] = buffer_data_4[4103:4096];
        layer2[1][31:24] = buffer_data_4[4111:4104];
        layer2[1][39:32] = buffer_data_4[4119:4112];
        layer2[1][47:40] = buffer_data_4[4127:4120];
        layer2[1][55:48] = buffer_data_4[4135:4128];
        layer3[1][7:0] = buffer_data_3[4087:4080];
        layer3[1][15:8] = buffer_data_3[4095:4088];
        layer3[1][23:16] = buffer_data_3[4103:4096];
        layer3[1][31:24] = buffer_data_3[4111:4104];
        layer3[1][39:32] = buffer_data_3[4119:4112];
        layer3[1][47:40] = buffer_data_3[4127:4120];
        layer3[1][55:48] = buffer_data_3[4135:4128];
        layer4[1][7:0] = buffer_data_2[4087:4080];
        layer4[1][15:8] = buffer_data_2[4095:4088];
        layer4[1][23:16] = buffer_data_2[4103:4096];
        layer4[1][31:24] = buffer_data_2[4111:4104];
        layer4[1][39:32] = buffer_data_2[4119:4112];
        layer4[1][47:40] = buffer_data_2[4127:4120];
        layer4[1][55:48] = buffer_data_2[4135:4128];
        layer5[1][7:0] = buffer_data_1[4087:4080];
        layer5[1][15:8] = buffer_data_1[4095:4088];
        layer5[1][23:16] = buffer_data_1[4103:4096];
        layer5[1][31:24] = buffer_data_1[4111:4104];
        layer5[1][39:32] = buffer_data_1[4119:4112];
        layer5[1][47:40] = buffer_data_1[4127:4120];
        layer5[1][55:48] = buffer_data_1[4135:4128];
        layer6[1][7:0] = buffer_data_0[4087:4080];
        layer6[1][15:8] = buffer_data_0[4095:4088];
        layer6[1][23:16] = buffer_data_0[4103:4096];
        layer6[1][31:24] = buffer_data_0[4111:4104];
        layer6[1][39:32] = buffer_data_0[4119:4112];
        layer6[1][47:40] = buffer_data_0[4127:4120];
        layer6[1][55:48] = buffer_data_0[4135:4128];
        layer0[2][7:0] = buffer_data_6[4095:4088];
        layer0[2][15:8] = buffer_data_6[4103:4096];
        layer0[2][23:16] = buffer_data_6[4111:4104];
        layer0[2][31:24] = buffer_data_6[4119:4112];
        layer0[2][39:32] = buffer_data_6[4127:4120];
        layer0[2][47:40] = buffer_data_6[4135:4128];
        layer0[2][55:48] = buffer_data_6[4143:4136];
        layer1[2][7:0] = buffer_data_5[4095:4088];
        layer1[2][15:8] = buffer_data_5[4103:4096];
        layer1[2][23:16] = buffer_data_5[4111:4104];
        layer1[2][31:24] = buffer_data_5[4119:4112];
        layer1[2][39:32] = buffer_data_5[4127:4120];
        layer1[2][47:40] = buffer_data_5[4135:4128];
        layer1[2][55:48] = buffer_data_5[4143:4136];
        layer2[2][7:0] = buffer_data_4[4095:4088];
        layer2[2][15:8] = buffer_data_4[4103:4096];
        layer2[2][23:16] = buffer_data_4[4111:4104];
        layer2[2][31:24] = buffer_data_4[4119:4112];
        layer2[2][39:32] = buffer_data_4[4127:4120];
        layer2[2][47:40] = buffer_data_4[4135:4128];
        layer2[2][55:48] = buffer_data_4[4143:4136];
        layer3[2][7:0] = buffer_data_3[4095:4088];
        layer3[2][15:8] = buffer_data_3[4103:4096];
        layer3[2][23:16] = buffer_data_3[4111:4104];
        layer3[2][31:24] = buffer_data_3[4119:4112];
        layer3[2][39:32] = buffer_data_3[4127:4120];
        layer3[2][47:40] = buffer_data_3[4135:4128];
        layer3[2][55:48] = buffer_data_3[4143:4136];
        layer4[2][7:0] = buffer_data_2[4095:4088];
        layer4[2][15:8] = buffer_data_2[4103:4096];
        layer4[2][23:16] = buffer_data_2[4111:4104];
        layer4[2][31:24] = buffer_data_2[4119:4112];
        layer4[2][39:32] = buffer_data_2[4127:4120];
        layer4[2][47:40] = buffer_data_2[4135:4128];
        layer4[2][55:48] = buffer_data_2[4143:4136];
        layer5[2][7:0] = buffer_data_1[4095:4088];
        layer5[2][15:8] = buffer_data_1[4103:4096];
        layer5[2][23:16] = buffer_data_1[4111:4104];
        layer5[2][31:24] = buffer_data_1[4119:4112];
        layer5[2][39:32] = buffer_data_1[4127:4120];
        layer5[2][47:40] = buffer_data_1[4135:4128];
        layer5[2][55:48] = buffer_data_1[4143:4136];
        layer6[2][7:0] = buffer_data_0[4095:4088];
        layer6[2][15:8] = buffer_data_0[4103:4096];
        layer6[2][23:16] = buffer_data_0[4111:4104];
        layer6[2][31:24] = buffer_data_0[4119:4112];
        layer6[2][39:32] = buffer_data_0[4127:4120];
        layer6[2][47:40] = buffer_data_0[4135:4128];
        layer6[2][55:48] = buffer_data_0[4143:4136];
        layer0[3][7:0] = buffer_data_6[4103:4096];
        layer0[3][15:8] = buffer_data_6[4111:4104];
        layer0[3][23:16] = buffer_data_6[4119:4112];
        layer0[3][31:24] = buffer_data_6[4127:4120];
        layer0[3][39:32] = buffer_data_6[4135:4128];
        layer0[3][47:40] = buffer_data_6[4143:4136];
        layer0[3][55:48] = buffer_data_6[4151:4144];
        layer1[3][7:0] = buffer_data_5[4103:4096];
        layer1[3][15:8] = buffer_data_5[4111:4104];
        layer1[3][23:16] = buffer_data_5[4119:4112];
        layer1[3][31:24] = buffer_data_5[4127:4120];
        layer1[3][39:32] = buffer_data_5[4135:4128];
        layer1[3][47:40] = buffer_data_5[4143:4136];
        layer1[3][55:48] = buffer_data_5[4151:4144];
        layer2[3][7:0] = buffer_data_4[4103:4096];
        layer2[3][15:8] = buffer_data_4[4111:4104];
        layer2[3][23:16] = buffer_data_4[4119:4112];
        layer2[3][31:24] = buffer_data_4[4127:4120];
        layer2[3][39:32] = buffer_data_4[4135:4128];
        layer2[3][47:40] = buffer_data_4[4143:4136];
        layer2[3][55:48] = buffer_data_4[4151:4144];
        layer3[3][7:0] = buffer_data_3[4103:4096];
        layer3[3][15:8] = buffer_data_3[4111:4104];
        layer3[3][23:16] = buffer_data_3[4119:4112];
        layer3[3][31:24] = buffer_data_3[4127:4120];
        layer3[3][39:32] = buffer_data_3[4135:4128];
        layer3[3][47:40] = buffer_data_3[4143:4136];
        layer3[3][55:48] = buffer_data_3[4151:4144];
        layer4[3][7:0] = buffer_data_2[4103:4096];
        layer4[3][15:8] = buffer_data_2[4111:4104];
        layer4[3][23:16] = buffer_data_2[4119:4112];
        layer4[3][31:24] = buffer_data_2[4127:4120];
        layer4[3][39:32] = buffer_data_2[4135:4128];
        layer4[3][47:40] = buffer_data_2[4143:4136];
        layer4[3][55:48] = buffer_data_2[4151:4144];
        layer5[3][7:0] = buffer_data_1[4103:4096];
        layer5[3][15:8] = buffer_data_1[4111:4104];
        layer5[3][23:16] = buffer_data_1[4119:4112];
        layer5[3][31:24] = buffer_data_1[4127:4120];
        layer5[3][39:32] = buffer_data_1[4135:4128];
        layer5[3][47:40] = buffer_data_1[4143:4136];
        layer5[3][55:48] = buffer_data_1[4151:4144];
        layer6[3][7:0] = buffer_data_0[4103:4096];
        layer6[3][15:8] = buffer_data_0[4111:4104];
        layer6[3][23:16] = buffer_data_0[4119:4112];
        layer6[3][31:24] = buffer_data_0[4127:4120];
        layer6[3][39:32] = buffer_data_0[4135:4128];
        layer6[3][47:40] = buffer_data_0[4143:4136];
        layer6[3][55:48] = buffer_data_0[4151:4144];
        layer0[4][7:0] = buffer_data_6[4111:4104];
        layer0[4][15:8] = buffer_data_6[4119:4112];
        layer0[4][23:16] = buffer_data_6[4127:4120];
        layer0[4][31:24] = buffer_data_6[4135:4128];
        layer0[4][39:32] = buffer_data_6[4143:4136];
        layer0[4][47:40] = buffer_data_6[4151:4144];
        layer0[4][55:48] = buffer_data_6[4159:4152];
        layer1[4][7:0] = buffer_data_5[4111:4104];
        layer1[4][15:8] = buffer_data_5[4119:4112];
        layer1[4][23:16] = buffer_data_5[4127:4120];
        layer1[4][31:24] = buffer_data_5[4135:4128];
        layer1[4][39:32] = buffer_data_5[4143:4136];
        layer1[4][47:40] = buffer_data_5[4151:4144];
        layer1[4][55:48] = buffer_data_5[4159:4152];
        layer2[4][7:0] = buffer_data_4[4111:4104];
        layer2[4][15:8] = buffer_data_4[4119:4112];
        layer2[4][23:16] = buffer_data_4[4127:4120];
        layer2[4][31:24] = buffer_data_4[4135:4128];
        layer2[4][39:32] = buffer_data_4[4143:4136];
        layer2[4][47:40] = buffer_data_4[4151:4144];
        layer2[4][55:48] = buffer_data_4[4159:4152];
        layer3[4][7:0] = buffer_data_3[4111:4104];
        layer3[4][15:8] = buffer_data_3[4119:4112];
        layer3[4][23:16] = buffer_data_3[4127:4120];
        layer3[4][31:24] = buffer_data_3[4135:4128];
        layer3[4][39:32] = buffer_data_3[4143:4136];
        layer3[4][47:40] = buffer_data_3[4151:4144];
        layer3[4][55:48] = buffer_data_3[4159:4152];
        layer4[4][7:0] = buffer_data_2[4111:4104];
        layer4[4][15:8] = buffer_data_2[4119:4112];
        layer4[4][23:16] = buffer_data_2[4127:4120];
        layer4[4][31:24] = buffer_data_2[4135:4128];
        layer4[4][39:32] = buffer_data_2[4143:4136];
        layer4[4][47:40] = buffer_data_2[4151:4144];
        layer4[4][55:48] = buffer_data_2[4159:4152];
        layer5[4][7:0] = buffer_data_1[4111:4104];
        layer5[4][15:8] = buffer_data_1[4119:4112];
        layer5[4][23:16] = buffer_data_1[4127:4120];
        layer5[4][31:24] = buffer_data_1[4135:4128];
        layer5[4][39:32] = buffer_data_1[4143:4136];
        layer5[4][47:40] = buffer_data_1[4151:4144];
        layer5[4][55:48] = buffer_data_1[4159:4152];
        layer6[4][7:0] = buffer_data_0[4111:4104];
        layer6[4][15:8] = buffer_data_0[4119:4112];
        layer6[4][23:16] = buffer_data_0[4127:4120];
        layer6[4][31:24] = buffer_data_0[4135:4128];
        layer6[4][39:32] = buffer_data_0[4143:4136];
        layer6[4][47:40] = buffer_data_0[4151:4144];
        layer6[4][55:48] = buffer_data_0[4159:4152];
        layer0[5][7:0] = buffer_data_6[4119:4112];
        layer0[5][15:8] = buffer_data_6[4127:4120];
        layer0[5][23:16] = buffer_data_6[4135:4128];
        layer0[5][31:24] = buffer_data_6[4143:4136];
        layer0[5][39:32] = buffer_data_6[4151:4144];
        layer0[5][47:40] = buffer_data_6[4159:4152];
        layer0[5][55:48] = buffer_data_6[4167:4160];
        layer1[5][7:0] = buffer_data_5[4119:4112];
        layer1[5][15:8] = buffer_data_5[4127:4120];
        layer1[5][23:16] = buffer_data_5[4135:4128];
        layer1[5][31:24] = buffer_data_5[4143:4136];
        layer1[5][39:32] = buffer_data_5[4151:4144];
        layer1[5][47:40] = buffer_data_5[4159:4152];
        layer1[5][55:48] = buffer_data_5[4167:4160];
        layer2[5][7:0] = buffer_data_4[4119:4112];
        layer2[5][15:8] = buffer_data_4[4127:4120];
        layer2[5][23:16] = buffer_data_4[4135:4128];
        layer2[5][31:24] = buffer_data_4[4143:4136];
        layer2[5][39:32] = buffer_data_4[4151:4144];
        layer2[5][47:40] = buffer_data_4[4159:4152];
        layer2[5][55:48] = buffer_data_4[4167:4160];
        layer3[5][7:0] = buffer_data_3[4119:4112];
        layer3[5][15:8] = buffer_data_3[4127:4120];
        layer3[5][23:16] = buffer_data_3[4135:4128];
        layer3[5][31:24] = buffer_data_3[4143:4136];
        layer3[5][39:32] = buffer_data_3[4151:4144];
        layer3[5][47:40] = buffer_data_3[4159:4152];
        layer3[5][55:48] = buffer_data_3[4167:4160];
        layer4[5][7:0] = buffer_data_2[4119:4112];
        layer4[5][15:8] = buffer_data_2[4127:4120];
        layer4[5][23:16] = buffer_data_2[4135:4128];
        layer4[5][31:24] = buffer_data_2[4143:4136];
        layer4[5][39:32] = buffer_data_2[4151:4144];
        layer4[5][47:40] = buffer_data_2[4159:4152];
        layer4[5][55:48] = buffer_data_2[4167:4160];
        layer5[5][7:0] = buffer_data_1[4119:4112];
        layer5[5][15:8] = buffer_data_1[4127:4120];
        layer5[5][23:16] = buffer_data_1[4135:4128];
        layer5[5][31:24] = buffer_data_1[4143:4136];
        layer5[5][39:32] = buffer_data_1[4151:4144];
        layer5[5][47:40] = buffer_data_1[4159:4152];
        layer5[5][55:48] = buffer_data_1[4167:4160];
        layer6[5][7:0] = buffer_data_0[4119:4112];
        layer6[5][15:8] = buffer_data_0[4127:4120];
        layer6[5][23:16] = buffer_data_0[4135:4128];
        layer6[5][31:24] = buffer_data_0[4143:4136];
        layer6[5][39:32] = buffer_data_0[4151:4144];
        layer6[5][47:40] = buffer_data_0[4159:4152];
        layer6[5][55:48] = buffer_data_0[4167:4160];
        layer0[6][7:0] = buffer_data_6[4127:4120];
        layer0[6][15:8] = buffer_data_6[4135:4128];
        layer0[6][23:16] = buffer_data_6[4143:4136];
        layer0[6][31:24] = buffer_data_6[4151:4144];
        layer0[6][39:32] = buffer_data_6[4159:4152];
        layer0[6][47:40] = buffer_data_6[4167:4160];
        layer0[6][55:48] = buffer_data_6[4175:4168];
        layer1[6][7:0] = buffer_data_5[4127:4120];
        layer1[6][15:8] = buffer_data_5[4135:4128];
        layer1[6][23:16] = buffer_data_5[4143:4136];
        layer1[6][31:24] = buffer_data_5[4151:4144];
        layer1[6][39:32] = buffer_data_5[4159:4152];
        layer1[6][47:40] = buffer_data_5[4167:4160];
        layer1[6][55:48] = buffer_data_5[4175:4168];
        layer2[6][7:0] = buffer_data_4[4127:4120];
        layer2[6][15:8] = buffer_data_4[4135:4128];
        layer2[6][23:16] = buffer_data_4[4143:4136];
        layer2[6][31:24] = buffer_data_4[4151:4144];
        layer2[6][39:32] = buffer_data_4[4159:4152];
        layer2[6][47:40] = buffer_data_4[4167:4160];
        layer2[6][55:48] = buffer_data_4[4175:4168];
        layer3[6][7:0] = buffer_data_3[4127:4120];
        layer3[6][15:8] = buffer_data_3[4135:4128];
        layer3[6][23:16] = buffer_data_3[4143:4136];
        layer3[6][31:24] = buffer_data_3[4151:4144];
        layer3[6][39:32] = buffer_data_3[4159:4152];
        layer3[6][47:40] = buffer_data_3[4167:4160];
        layer3[6][55:48] = buffer_data_3[4175:4168];
        layer4[6][7:0] = buffer_data_2[4127:4120];
        layer4[6][15:8] = buffer_data_2[4135:4128];
        layer4[6][23:16] = buffer_data_2[4143:4136];
        layer4[6][31:24] = buffer_data_2[4151:4144];
        layer4[6][39:32] = buffer_data_2[4159:4152];
        layer4[6][47:40] = buffer_data_2[4167:4160];
        layer4[6][55:48] = buffer_data_2[4175:4168];
        layer5[6][7:0] = buffer_data_1[4127:4120];
        layer5[6][15:8] = buffer_data_1[4135:4128];
        layer5[6][23:16] = buffer_data_1[4143:4136];
        layer5[6][31:24] = buffer_data_1[4151:4144];
        layer5[6][39:32] = buffer_data_1[4159:4152];
        layer5[6][47:40] = buffer_data_1[4167:4160];
        layer5[6][55:48] = buffer_data_1[4175:4168];
        layer6[6][7:0] = buffer_data_0[4127:4120];
        layer6[6][15:8] = buffer_data_0[4135:4128];
        layer6[6][23:16] = buffer_data_0[4143:4136];
        layer6[6][31:24] = buffer_data_0[4151:4144];
        layer6[6][39:32] = buffer_data_0[4159:4152];
        layer6[6][47:40] = buffer_data_0[4167:4160];
        layer6[6][55:48] = buffer_data_0[4175:4168];
        layer0[7][7:0] = buffer_data_6[4135:4128];
        layer0[7][15:8] = buffer_data_6[4143:4136];
        layer0[7][23:16] = buffer_data_6[4151:4144];
        layer0[7][31:24] = buffer_data_6[4159:4152];
        layer0[7][39:32] = buffer_data_6[4167:4160];
        layer0[7][47:40] = buffer_data_6[4175:4168];
        layer0[7][55:48] = buffer_data_6[4183:4176];
        layer1[7][7:0] = buffer_data_5[4135:4128];
        layer1[7][15:8] = buffer_data_5[4143:4136];
        layer1[7][23:16] = buffer_data_5[4151:4144];
        layer1[7][31:24] = buffer_data_5[4159:4152];
        layer1[7][39:32] = buffer_data_5[4167:4160];
        layer1[7][47:40] = buffer_data_5[4175:4168];
        layer1[7][55:48] = buffer_data_5[4183:4176];
        layer2[7][7:0] = buffer_data_4[4135:4128];
        layer2[7][15:8] = buffer_data_4[4143:4136];
        layer2[7][23:16] = buffer_data_4[4151:4144];
        layer2[7][31:24] = buffer_data_4[4159:4152];
        layer2[7][39:32] = buffer_data_4[4167:4160];
        layer2[7][47:40] = buffer_data_4[4175:4168];
        layer2[7][55:48] = buffer_data_4[4183:4176];
        layer3[7][7:0] = buffer_data_3[4135:4128];
        layer3[7][15:8] = buffer_data_3[4143:4136];
        layer3[7][23:16] = buffer_data_3[4151:4144];
        layer3[7][31:24] = buffer_data_3[4159:4152];
        layer3[7][39:32] = buffer_data_3[4167:4160];
        layer3[7][47:40] = buffer_data_3[4175:4168];
        layer3[7][55:48] = buffer_data_3[4183:4176];
        layer4[7][7:0] = buffer_data_2[4135:4128];
        layer4[7][15:8] = buffer_data_2[4143:4136];
        layer4[7][23:16] = buffer_data_2[4151:4144];
        layer4[7][31:24] = buffer_data_2[4159:4152];
        layer4[7][39:32] = buffer_data_2[4167:4160];
        layer4[7][47:40] = buffer_data_2[4175:4168];
        layer4[7][55:48] = buffer_data_2[4183:4176];
        layer5[7][7:0] = buffer_data_1[4135:4128];
        layer5[7][15:8] = buffer_data_1[4143:4136];
        layer5[7][23:16] = buffer_data_1[4151:4144];
        layer5[7][31:24] = buffer_data_1[4159:4152];
        layer5[7][39:32] = buffer_data_1[4167:4160];
        layer5[7][47:40] = buffer_data_1[4175:4168];
        layer5[7][55:48] = buffer_data_1[4183:4176];
        layer6[7][7:0] = buffer_data_0[4135:4128];
        layer6[7][15:8] = buffer_data_0[4143:4136];
        layer6[7][23:16] = buffer_data_0[4151:4144];
        layer6[7][31:24] = buffer_data_0[4159:4152];
        layer6[7][39:32] = buffer_data_0[4167:4160];
        layer6[7][47:40] = buffer_data_0[4175:4168];
        layer6[7][55:48] = buffer_data_0[4183:4176];
        layer0[8][7:0] = buffer_data_6[4143:4136];
        layer0[8][15:8] = buffer_data_6[4151:4144];
        layer0[8][23:16] = buffer_data_6[4159:4152];
        layer0[8][31:24] = buffer_data_6[4167:4160];
        layer0[8][39:32] = buffer_data_6[4175:4168];
        layer0[8][47:40] = buffer_data_6[4183:4176];
        layer0[8][55:48] = buffer_data_6[4191:4184];
        layer1[8][7:0] = buffer_data_5[4143:4136];
        layer1[8][15:8] = buffer_data_5[4151:4144];
        layer1[8][23:16] = buffer_data_5[4159:4152];
        layer1[8][31:24] = buffer_data_5[4167:4160];
        layer1[8][39:32] = buffer_data_5[4175:4168];
        layer1[8][47:40] = buffer_data_5[4183:4176];
        layer1[8][55:48] = buffer_data_5[4191:4184];
        layer2[8][7:0] = buffer_data_4[4143:4136];
        layer2[8][15:8] = buffer_data_4[4151:4144];
        layer2[8][23:16] = buffer_data_4[4159:4152];
        layer2[8][31:24] = buffer_data_4[4167:4160];
        layer2[8][39:32] = buffer_data_4[4175:4168];
        layer2[8][47:40] = buffer_data_4[4183:4176];
        layer2[8][55:48] = buffer_data_4[4191:4184];
        layer3[8][7:0] = buffer_data_3[4143:4136];
        layer3[8][15:8] = buffer_data_3[4151:4144];
        layer3[8][23:16] = buffer_data_3[4159:4152];
        layer3[8][31:24] = buffer_data_3[4167:4160];
        layer3[8][39:32] = buffer_data_3[4175:4168];
        layer3[8][47:40] = buffer_data_3[4183:4176];
        layer3[8][55:48] = buffer_data_3[4191:4184];
        layer4[8][7:0] = buffer_data_2[4143:4136];
        layer4[8][15:8] = buffer_data_2[4151:4144];
        layer4[8][23:16] = buffer_data_2[4159:4152];
        layer4[8][31:24] = buffer_data_2[4167:4160];
        layer4[8][39:32] = buffer_data_2[4175:4168];
        layer4[8][47:40] = buffer_data_2[4183:4176];
        layer4[8][55:48] = buffer_data_2[4191:4184];
        layer5[8][7:0] = buffer_data_1[4143:4136];
        layer5[8][15:8] = buffer_data_1[4151:4144];
        layer5[8][23:16] = buffer_data_1[4159:4152];
        layer5[8][31:24] = buffer_data_1[4167:4160];
        layer5[8][39:32] = buffer_data_1[4175:4168];
        layer5[8][47:40] = buffer_data_1[4183:4176];
        layer5[8][55:48] = buffer_data_1[4191:4184];
        layer6[8][7:0] = buffer_data_0[4143:4136];
        layer6[8][15:8] = buffer_data_0[4151:4144];
        layer6[8][23:16] = buffer_data_0[4159:4152];
        layer6[8][31:24] = buffer_data_0[4167:4160];
        layer6[8][39:32] = buffer_data_0[4175:4168];
        layer6[8][47:40] = buffer_data_0[4183:4176];
        layer6[8][55:48] = buffer_data_0[4191:4184];
        layer0[9][7:0] = buffer_data_6[4151:4144];
        layer0[9][15:8] = buffer_data_6[4159:4152];
        layer0[9][23:16] = buffer_data_6[4167:4160];
        layer0[9][31:24] = buffer_data_6[4175:4168];
        layer0[9][39:32] = buffer_data_6[4183:4176];
        layer0[9][47:40] = buffer_data_6[4191:4184];
        layer0[9][55:48] = buffer_data_6[4199:4192];
        layer1[9][7:0] = buffer_data_5[4151:4144];
        layer1[9][15:8] = buffer_data_5[4159:4152];
        layer1[9][23:16] = buffer_data_5[4167:4160];
        layer1[9][31:24] = buffer_data_5[4175:4168];
        layer1[9][39:32] = buffer_data_5[4183:4176];
        layer1[9][47:40] = buffer_data_5[4191:4184];
        layer1[9][55:48] = buffer_data_5[4199:4192];
        layer2[9][7:0] = buffer_data_4[4151:4144];
        layer2[9][15:8] = buffer_data_4[4159:4152];
        layer2[9][23:16] = buffer_data_4[4167:4160];
        layer2[9][31:24] = buffer_data_4[4175:4168];
        layer2[9][39:32] = buffer_data_4[4183:4176];
        layer2[9][47:40] = buffer_data_4[4191:4184];
        layer2[9][55:48] = buffer_data_4[4199:4192];
        layer3[9][7:0] = buffer_data_3[4151:4144];
        layer3[9][15:8] = buffer_data_3[4159:4152];
        layer3[9][23:16] = buffer_data_3[4167:4160];
        layer3[9][31:24] = buffer_data_3[4175:4168];
        layer3[9][39:32] = buffer_data_3[4183:4176];
        layer3[9][47:40] = buffer_data_3[4191:4184];
        layer3[9][55:48] = buffer_data_3[4199:4192];
        layer4[9][7:0] = buffer_data_2[4151:4144];
        layer4[9][15:8] = buffer_data_2[4159:4152];
        layer4[9][23:16] = buffer_data_2[4167:4160];
        layer4[9][31:24] = buffer_data_2[4175:4168];
        layer4[9][39:32] = buffer_data_2[4183:4176];
        layer4[9][47:40] = buffer_data_2[4191:4184];
        layer4[9][55:48] = buffer_data_2[4199:4192];
        layer5[9][7:0] = buffer_data_1[4151:4144];
        layer5[9][15:8] = buffer_data_1[4159:4152];
        layer5[9][23:16] = buffer_data_1[4167:4160];
        layer5[9][31:24] = buffer_data_1[4175:4168];
        layer5[9][39:32] = buffer_data_1[4183:4176];
        layer5[9][47:40] = buffer_data_1[4191:4184];
        layer5[9][55:48] = buffer_data_1[4199:4192];
        layer6[9][7:0] = buffer_data_0[4151:4144];
        layer6[9][15:8] = buffer_data_0[4159:4152];
        layer6[9][23:16] = buffer_data_0[4167:4160];
        layer6[9][31:24] = buffer_data_0[4175:4168];
        layer6[9][39:32] = buffer_data_0[4183:4176];
        layer6[9][47:40] = buffer_data_0[4191:4184];
        layer6[9][55:48] = buffer_data_0[4199:4192];
        layer0[10][7:0] = buffer_data_6[4159:4152];
        layer0[10][15:8] = buffer_data_6[4167:4160];
        layer0[10][23:16] = buffer_data_6[4175:4168];
        layer0[10][31:24] = buffer_data_6[4183:4176];
        layer0[10][39:32] = buffer_data_6[4191:4184];
        layer0[10][47:40] = buffer_data_6[4199:4192];
        layer0[10][55:48] = buffer_data_6[4207:4200];
        layer1[10][7:0] = buffer_data_5[4159:4152];
        layer1[10][15:8] = buffer_data_5[4167:4160];
        layer1[10][23:16] = buffer_data_5[4175:4168];
        layer1[10][31:24] = buffer_data_5[4183:4176];
        layer1[10][39:32] = buffer_data_5[4191:4184];
        layer1[10][47:40] = buffer_data_5[4199:4192];
        layer1[10][55:48] = buffer_data_5[4207:4200];
        layer2[10][7:0] = buffer_data_4[4159:4152];
        layer2[10][15:8] = buffer_data_4[4167:4160];
        layer2[10][23:16] = buffer_data_4[4175:4168];
        layer2[10][31:24] = buffer_data_4[4183:4176];
        layer2[10][39:32] = buffer_data_4[4191:4184];
        layer2[10][47:40] = buffer_data_4[4199:4192];
        layer2[10][55:48] = buffer_data_4[4207:4200];
        layer3[10][7:0] = buffer_data_3[4159:4152];
        layer3[10][15:8] = buffer_data_3[4167:4160];
        layer3[10][23:16] = buffer_data_3[4175:4168];
        layer3[10][31:24] = buffer_data_3[4183:4176];
        layer3[10][39:32] = buffer_data_3[4191:4184];
        layer3[10][47:40] = buffer_data_3[4199:4192];
        layer3[10][55:48] = buffer_data_3[4207:4200];
        layer4[10][7:0] = buffer_data_2[4159:4152];
        layer4[10][15:8] = buffer_data_2[4167:4160];
        layer4[10][23:16] = buffer_data_2[4175:4168];
        layer4[10][31:24] = buffer_data_2[4183:4176];
        layer4[10][39:32] = buffer_data_2[4191:4184];
        layer4[10][47:40] = buffer_data_2[4199:4192];
        layer4[10][55:48] = buffer_data_2[4207:4200];
        layer5[10][7:0] = buffer_data_1[4159:4152];
        layer5[10][15:8] = buffer_data_1[4167:4160];
        layer5[10][23:16] = buffer_data_1[4175:4168];
        layer5[10][31:24] = buffer_data_1[4183:4176];
        layer5[10][39:32] = buffer_data_1[4191:4184];
        layer5[10][47:40] = buffer_data_1[4199:4192];
        layer5[10][55:48] = buffer_data_1[4207:4200];
        layer6[10][7:0] = buffer_data_0[4159:4152];
        layer6[10][15:8] = buffer_data_0[4167:4160];
        layer6[10][23:16] = buffer_data_0[4175:4168];
        layer6[10][31:24] = buffer_data_0[4183:4176];
        layer6[10][39:32] = buffer_data_0[4191:4184];
        layer6[10][47:40] = buffer_data_0[4199:4192];
        layer6[10][55:48] = buffer_data_0[4207:4200];
        layer0[11][7:0] = buffer_data_6[4167:4160];
        layer0[11][15:8] = buffer_data_6[4175:4168];
        layer0[11][23:16] = buffer_data_6[4183:4176];
        layer0[11][31:24] = buffer_data_6[4191:4184];
        layer0[11][39:32] = buffer_data_6[4199:4192];
        layer0[11][47:40] = buffer_data_6[4207:4200];
        layer0[11][55:48] = buffer_data_6[4215:4208];
        layer1[11][7:0] = buffer_data_5[4167:4160];
        layer1[11][15:8] = buffer_data_5[4175:4168];
        layer1[11][23:16] = buffer_data_5[4183:4176];
        layer1[11][31:24] = buffer_data_5[4191:4184];
        layer1[11][39:32] = buffer_data_5[4199:4192];
        layer1[11][47:40] = buffer_data_5[4207:4200];
        layer1[11][55:48] = buffer_data_5[4215:4208];
        layer2[11][7:0] = buffer_data_4[4167:4160];
        layer2[11][15:8] = buffer_data_4[4175:4168];
        layer2[11][23:16] = buffer_data_4[4183:4176];
        layer2[11][31:24] = buffer_data_4[4191:4184];
        layer2[11][39:32] = buffer_data_4[4199:4192];
        layer2[11][47:40] = buffer_data_4[4207:4200];
        layer2[11][55:48] = buffer_data_4[4215:4208];
        layer3[11][7:0] = buffer_data_3[4167:4160];
        layer3[11][15:8] = buffer_data_3[4175:4168];
        layer3[11][23:16] = buffer_data_3[4183:4176];
        layer3[11][31:24] = buffer_data_3[4191:4184];
        layer3[11][39:32] = buffer_data_3[4199:4192];
        layer3[11][47:40] = buffer_data_3[4207:4200];
        layer3[11][55:48] = buffer_data_3[4215:4208];
        layer4[11][7:0] = buffer_data_2[4167:4160];
        layer4[11][15:8] = buffer_data_2[4175:4168];
        layer4[11][23:16] = buffer_data_2[4183:4176];
        layer4[11][31:24] = buffer_data_2[4191:4184];
        layer4[11][39:32] = buffer_data_2[4199:4192];
        layer4[11][47:40] = buffer_data_2[4207:4200];
        layer4[11][55:48] = buffer_data_2[4215:4208];
        layer5[11][7:0] = buffer_data_1[4167:4160];
        layer5[11][15:8] = buffer_data_1[4175:4168];
        layer5[11][23:16] = buffer_data_1[4183:4176];
        layer5[11][31:24] = buffer_data_1[4191:4184];
        layer5[11][39:32] = buffer_data_1[4199:4192];
        layer5[11][47:40] = buffer_data_1[4207:4200];
        layer5[11][55:48] = buffer_data_1[4215:4208];
        layer6[11][7:0] = buffer_data_0[4167:4160];
        layer6[11][15:8] = buffer_data_0[4175:4168];
        layer6[11][23:16] = buffer_data_0[4183:4176];
        layer6[11][31:24] = buffer_data_0[4191:4184];
        layer6[11][39:32] = buffer_data_0[4199:4192];
        layer6[11][47:40] = buffer_data_0[4207:4200];
        layer6[11][55:48] = buffer_data_0[4215:4208];
        layer0[12][7:0] = buffer_data_6[4175:4168];
        layer0[12][15:8] = buffer_data_6[4183:4176];
        layer0[12][23:16] = buffer_data_6[4191:4184];
        layer0[12][31:24] = buffer_data_6[4199:4192];
        layer0[12][39:32] = buffer_data_6[4207:4200];
        layer0[12][47:40] = buffer_data_6[4215:4208];
        layer0[12][55:48] = buffer_data_6[4223:4216];
        layer1[12][7:0] = buffer_data_5[4175:4168];
        layer1[12][15:8] = buffer_data_5[4183:4176];
        layer1[12][23:16] = buffer_data_5[4191:4184];
        layer1[12][31:24] = buffer_data_5[4199:4192];
        layer1[12][39:32] = buffer_data_5[4207:4200];
        layer1[12][47:40] = buffer_data_5[4215:4208];
        layer1[12][55:48] = buffer_data_5[4223:4216];
        layer2[12][7:0] = buffer_data_4[4175:4168];
        layer2[12][15:8] = buffer_data_4[4183:4176];
        layer2[12][23:16] = buffer_data_4[4191:4184];
        layer2[12][31:24] = buffer_data_4[4199:4192];
        layer2[12][39:32] = buffer_data_4[4207:4200];
        layer2[12][47:40] = buffer_data_4[4215:4208];
        layer2[12][55:48] = buffer_data_4[4223:4216];
        layer3[12][7:0] = buffer_data_3[4175:4168];
        layer3[12][15:8] = buffer_data_3[4183:4176];
        layer3[12][23:16] = buffer_data_3[4191:4184];
        layer3[12][31:24] = buffer_data_3[4199:4192];
        layer3[12][39:32] = buffer_data_3[4207:4200];
        layer3[12][47:40] = buffer_data_3[4215:4208];
        layer3[12][55:48] = buffer_data_3[4223:4216];
        layer4[12][7:0] = buffer_data_2[4175:4168];
        layer4[12][15:8] = buffer_data_2[4183:4176];
        layer4[12][23:16] = buffer_data_2[4191:4184];
        layer4[12][31:24] = buffer_data_2[4199:4192];
        layer4[12][39:32] = buffer_data_2[4207:4200];
        layer4[12][47:40] = buffer_data_2[4215:4208];
        layer4[12][55:48] = buffer_data_2[4223:4216];
        layer5[12][7:0] = buffer_data_1[4175:4168];
        layer5[12][15:8] = buffer_data_1[4183:4176];
        layer5[12][23:16] = buffer_data_1[4191:4184];
        layer5[12][31:24] = buffer_data_1[4199:4192];
        layer5[12][39:32] = buffer_data_1[4207:4200];
        layer5[12][47:40] = buffer_data_1[4215:4208];
        layer5[12][55:48] = buffer_data_1[4223:4216];
        layer6[12][7:0] = buffer_data_0[4175:4168];
        layer6[12][15:8] = buffer_data_0[4183:4176];
        layer6[12][23:16] = buffer_data_0[4191:4184];
        layer6[12][31:24] = buffer_data_0[4199:4192];
        layer6[12][39:32] = buffer_data_0[4207:4200];
        layer6[12][47:40] = buffer_data_0[4215:4208];
        layer6[12][55:48] = buffer_data_0[4223:4216];
        layer0[13][7:0] = buffer_data_6[4183:4176];
        layer0[13][15:8] = buffer_data_6[4191:4184];
        layer0[13][23:16] = buffer_data_6[4199:4192];
        layer0[13][31:24] = buffer_data_6[4207:4200];
        layer0[13][39:32] = buffer_data_6[4215:4208];
        layer0[13][47:40] = buffer_data_6[4223:4216];
        layer0[13][55:48] = buffer_data_6[4231:4224];
        layer1[13][7:0] = buffer_data_5[4183:4176];
        layer1[13][15:8] = buffer_data_5[4191:4184];
        layer1[13][23:16] = buffer_data_5[4199:4192];
        layer1[13][31:24] = buffer_data_5[4207:4200];
        layer1[13][39:32] = buffer_data_5[4215:4208];
        layer1[13][47:40] = buffer_data_5[4223:4216];
        layer1[13][55:48] = buffer_data_5[4231:4224];
        layer2[13][7:0] = buffer_data_4[4183:4176];
        layer2[13][15:8] = buffer_data_4[4191:4184];
        layer2[13][23:16] = buffer_data_4[4199:4192];
        layer2[13][31:24] = buffer_data_4[4207:4200];
        layer2[13][39:32] = buffer_data_4[4215:4208];
        layer2[13][47:40] = buffer_data_4[4223:4216];
        layer2[13][55:48] = buffer_data_4[4231:4224];
        layer3[13][7:0] = buffer_data_3[4183:4176];
        layer3[13][15:8] = buffer_data_3[4191:4184];
        layer3[13][23:16] = buffer_data_3[4199:4192];
        layer3[13][31:24] = buffer_data_3[4207:4200];
        layer3[13][39:32] = buffer_data_3[4215:4208];
        layer3[13][47:40] = buffer_data_3[4223:4216];
        layer3[13][55:48] = buffer_data_3[4231:4224];
        layer4[13][7:0] = buffer_data_2[4183:4176];
        layer4[13][15:8] = buffer_data_2[4191:4184];
        layer4[13][23:16] = buffer_data_2[4199:4192];
        layer4[13][31:24] = buffer_data_2[4207:4200];
        layer4[13][39:32] = buffer_data_2[4215:4208];
        layer4[13][47:40] = buffer_data_2[4223:4216];
        layer4[13][55:48] = buffer_data_2[4231:4224];
        layer5[13][7:0] = buffer_data_1[4183:4176];
        layer5[13][15:8] = buffer_data_1[4191:4184];
        layer5[13][23:16] = buffer_data_1[4199:4192];
        layer5[13][31:24] = buffer_data_1[4207:4200];
        layer5[13][39:32] = buffer_data_1[4215:4208];
        layer5[13][47:40] = buffer_data_1[4223:4216];
        layer5[13][55:48] = buffer_data_1[4231:4224];
        layer6[13][7:0] = buffer_data_0[4183:4176];
        layer6[13][15:8] = buffer_data_0[4191:4184];
        layer6[13][23:16] = buffer_data_0[4199:4192];
        layer6[13][31:24] = buffer_data_0[4207:4200];
        layer6[13][39:32] = buffer_data_0[4215:4208];
        layer6[13][47:40] = buffer_data_0[4223:4216];
        layer6[13][55:48] = buffer_data_0[4231:4224];
        layer0[14][7:0] = buffer_data_6[4191:4184];
        layer0[14][15:8] = buffer_data_6[4199:4192];
        layer0[14][23:16] = buffer_data_6[4207:4200];
        layer0[14][31:24] = buffer_data_6[4215:4208];
        layer0[14][39:32] = buffer_data_6[4223:4216];
        layer0[14][47:40] = buffer_data_6[4231:4224];
        layer0[14][55:48] = buffer_data_6[4239:4232];
        layer1[14][7:0] = buffer_data_5[4191:4184];
        layer1[14][15:8] = buffer_data_5[4199:4192];
        layer1[14][23:16] = buffer_data_5[4207:4200];
        layer1[14][31:24] = buffer_data_5[4215:4208];
        layer1[14][39:32] = buffer_data_5[4223:4216];
        layer1[14][47:40] = buffer_data_5[4231:4224];
        layer1[14][55:48] = buffer_data_5[4239:4232];
        layer2[14][7:0] = buffer_data_4[4191:4184];
        layer2[14][15:8] = buffer_data_4[4199:4192];
        layer2[14][23:16] = buffer_data_4[4207:4200];
        layer2[14][31:24] = buffer_data_4[4215:4208];
        layer2[14][39:32] = buffer_data_4[4223:4216];
        layer2[14][47:40] = buffer_data_4[4231:4224];
        layer2[14][55:48] = buffer_data_4[4239:4232];
        layer3[14][7:0] = buffer_data_3[4191:4184];
        layer3[14][15:8] = buffer_data_3[4199:4192];
        layer3[14][23:16] = buffer_data_3[4207:4200];
        layer3[14][31:24] = buffer_data_3[4215:4208];
        layer3[14][39:32] = buffer_data_3[4223:4216];
        layer3[14][47:40] = buffer_data_3[4231:4224];
        layer3[14][55:48] = buffer_data_3[4239:4232];
        layer4[14][7:0] = buffer_data_2[4191:4184];
        layer4[14][15:8] = buffer_data_2[4199:4192];
        layer4[14][23:16] = buffer_data_2[4207:4200];
        layer4[14][31:24] = buffer_data_2[4215:4208];
        layer4[14][39:32] = buffer_data_2[4223:4216];
        layer4[14][47:40] = buffer_data_2[4231:4224];
        layer4[14][55:48] = buffer_data_2[4239:4232];
        layer5[14][7:0] = buffer_data_1[4191:4184];
        layer5[14][15:8] = buffer_data_1[4199:4192];
        layer5[14][23:16] = buffer_data_1[4207:4200];
        layer5[14][31:24] = buffer_data_1[4215:4208];
        layer5[14][39:32] = buffer_data_1[4223:4216];
        layer5[14][47:40] = buffer_data_1[4231:4224];
        layer5[14][55:48] = buffer_data_1[4239:4232];
        layer6[14][7:0] = buffer_data_0[4191:4184];
        layer6[14][15:8] = buffer_data_0[4199:4192];
        layer6[14][23:16] = buffer_data_0[4207:4200];
        layer6[14][31:24] = buffer_data_0[4215:4208];
        layer6[14][39:32] = buffer_data_0[4223:4216];
        layer6[14][47:40] = buffer_data_0[4231:4224];
        layer6[14][55:48] = buffer_data_0[4239:4232];
        layer0[15][7:0] = buffer_data_6[4199:4192];
        layer0[15][15:8] = buffer_data_6[4207:4200];
        layer0[15][23:16] = buffer_data_6[4215:4208];
        layer0[15][31:24] = buffer_data_6[4223:4216];
        layer0[15][39:32] = buffer_data_6[4231:4224];
        layer0[15][47:40] = buffer_data_6[4239:4232];
        layer0[15][55:48] = buffer_data_6[4247:4240];
        layer1[15][7:0] = buffer_data_5[4199:4192];
        layer1[15][15:8] = buffer_data_5[4207:4200];
        layer1[15][23:16] = buffer_data_5[4215:4208];
        layer1[15][31:24] = buffer_data_5[4223:4216];
        layer1[15][39:32] = buffer_data_5[4231:4224];
        layer1[15][47:40] = buffer_data_5[4239:4232];
        layer1[15][55:48] = buffer_data_5[4247:4240];
        layer2[15][7:0] = buffer_data_4[4199:4192];
        layer2[15][15:8] = buffer_data_4[4207:4200];
        layer2[15][23:16] = buffer_data_4[4215:4208];
        layer2[15][31:24] = buffer_data_4[4223:4216];
        layer2[15][39:32] = buffer_data_4[4231:4224];
        layer2[15][47:40] = buffer_data_4[4239:4232];
        layer2[15][55:48] = buffer_data_4[4247:4240];
        layer3[15][7:0] = buffer_data_3[4199:4192];
        layer3[15][15:8] = buffer_data_3[4207:4200];
        layer3[15][23:16] = buffer_data_3[4215:4208];
        layer3[15][31:24] = buffer_data_3[4223:4216];
        layer3[15][39:32] = buffer_data_3[4231:4224];
        layer3[15][47:40] = buffer_data_3[4239:4232];
        layer3[15][55:48] = buffer_data_3[4247:4240];
        layer4[15][7:0] = buffer_data_2[4199:4192];
        layer4[15][15:8] = buffer_data_2[4207:4200];
        layer4[15][23:16] = buffer_data_2[4215:4208];
        layer4[15][31:24] = buffer_data_2[4223:4216];
        layer4[15][39:32] = buffer_data_2[4231:4224];
        layer4[15][47:40] = buffer_data_2[4239:4232];
        layer4[15][55:48] = buffer_data_2[4247:4240];
        layer5[15][7:0] = buffer_data_1[4199:4192];
        layer5[15][15:8] = buffer_data_1[4207:4200];
        layer5[15][23:16] = buffer_data_1[4215:4208];
        layer5[15][31:24] = buffer_data_1[4223:4216];
        layer5[15][39:32] = buffer_data_1[4231:4224];
        layer5[15][47:40] = buffer_data_1[4239:4232];
        layer5[15][55:48] = buffer_data_1[4247:4240];
        layer6[15][7:0] = buffer_data_0[4199:4192];
        layer6[15][15:8] = buffer_data_0[4207:4200];
        layer6[15][23:16] = buffer_data_0[4215:4208];
        layer6[15][31:24] = buffer_data_0[4223:4216];
        layer6[15][39:32] = buffer_data_0[4231:4224];
        layer6[15][47:40] = buffer_data_0[4239:4232];
        layer6[15][55:48] = buffer_data_0[4247:4240];
        layer0[16][7:0] = buffer_data_6[4207:4200];
        layer0[16][15:8] = buffer_data_6[4215:4208];
        layer0[16][23:16] = buffer_data_6[4223:4216];
        layer0[16][31:24] = buffer_data_6[4231:4224];
        layer0[16][39:32] = buffer_data_6[4239:4232];
        layer0[16][47:40] = buffer_data_6[4247:4240];
        layer0[16][55:48] = buffer_data_6[4255:4248];
        layer1[16][7:0] = buffer_data_5[4207:4200];
        layer1[16][15:8] = buffer_data_5[4215:4208];
        layer1[16][23:16] = buffer_data_5[4223:4216];
        layer1[16][31:24] = buffer_data_5[4231:4224];
        layer1[16][39:32] = buffer_data_5[4239:4232];
        layer1[16][47:40] = buffer_data_5[4247:4240];
        layer1[16][55:48] = buffer_data_5[4255:4248];
        layer2[16][7:0] = buffer_data_4[4207:4200];
        layer2[16][15:8] = buffer_data_4[4215:4208];
        layer2[16][23:16] = buffer_data_4[4223:4216];
        layer2[16][31:24] = buffer_data_4[4231:4224];
        layer2[16][39:32] = buffer_data_4[4239:4232];
        layer2[16][47:40] = buffer_data_4[4247:4240];
        layer2[16][55:48] = buffer_data_4[4255:4248];
        layer3[16][7:0] = buffer_data_3[4207:4200];
        layer3[16][15:8] = buffer_data_3[4215:4208];
        layer3[16][23:16] = buffer_data_3[4223:4216];
        layer3[16][31:24] = buffer_data_3[4231:4224];
        layer3[16][39:32] = buffer_data_3[4239:4232];
        layer3[16][47:40] = buffer_data_3[4247:4240];
        layer3[16][55:48] = buffer_data_3[4255:4248];
        layer4[16][7:0] = buffer_data_2[4207:4200];
        layer4[16][15:8] = buffer_data_2[4215:4208];
        layer4[16][23:16] = buffer_data_2[4223:4216];
        layer4[16][31:24] = buffer_data_2[4231:4224];
        layer4[16][39:32] = buffer_data_2[4239:4232];
        layer4[16][47:40] = buffer_data_2[4247:4240];
        layer4[16][55:48] = buffer_data_2[4255:4248];
        layer5[16][7:0] = buffer_data_1[4207:4200];
        layer5[16][15:8] = buffer_data_1[4215:4208];
        layer5[16][23:16] = buffer_data_1[4223:4216];
        layer5[16][31:24] = buffer_data_1[4231:4224];
        layer5[16][39:32] = buffer_data_1[4239:4232];
        layer5[16][47:40] = buffer_data_1[4247:4240];
        layer5[16][55:48] = buffer_data_1[4255:4248];
        layer6[16][7:0] = buffer_data_0[4207:4200];
        layer6[16][15:8] = buffer_data_0[4215:4208];
        layer6[16][23:16] = buffer_data_0[4223:4216];
        layer6[16][31:24] = buffer_data_0[4231:4224];
        layer6[16][39:32] = buffer_data_0[4239:4232];
        layer6[16][47:40] = buffer_data_0[4247:4240];
        layer6[16][55:48] = buffer_data_0[4255:4248];
        layer0[17][7:0] = buffer_data_6[4215:4208];
        layer0[17][15:8] = buffer_data_6[4223:4216];
        layer0[17][23:16] = buffer_data_6[4231:4224];
        layer0[17][31:24] = buffer_data_6[4239:4232];
        layer0[17][39:32] = buffer_data_6[4247:4240];
        layer0[17][47:40] = buffer_data_6[4255:4248];
        layer0[17][55:48] = buffer_data_6[4263:4256];
        layer1[17][7:0] = buffer_data_5[4215:4208];
        layer1[17][15:8] = buffer_data_5[4223:4216];
        layer1[17][23:16] = buffer_data_5[4231:4224];
        layer1[17][31:24] = buffer_data_5[4239:4232];
        layer1[17][39:32] = buffer_data_5[4247:4240];
        layer1[17][47:40] = buffer_data_5[4255:4248];
        layer1[17][55:48] = buffer_data_5[4263:4256];
        layer2[17][7:0] = buffer_data_4[4215:4208];
        layer2[17][15:8] = buffer_data_4[4223:4216];
        layer2[17][23:16] = buffer_data_4[4231:4224];
        layer2[17][31:24] = buffer_data_4[4239:4232];
        layer2[17][39:32] = buffer_data_4[4247:4240];
        layer2[17][47:40] = buffer_data_4[4255:4248];
        layer2[17][55:48] = buffer_data_4[4263:4256];
        layer3[17][7:0] = buffer_data_3[4215:4208];
        layer3[17][15:8] = buffer_data_3[4223:4216];
        layer3[17][23:16] = buffer_data_3[4231:4224];
        layer3[17][31:24] = buffer_data_3[4239:4232];
        layer3[17][39:32] = buffer_data_3[4247:4240];
        layer3[17][47:40] = buffer_data_3[4255:4248];
        layer3[17][55:48] = buffer_data_3[4263:4256];
        layer4[17][7:0] = buffer_data_2[4215:4208];
        layer4[17][15:8] = buffer_data_2[4223:4216];
        layer4[17][23:16] = buffer_data_2[4231:4224];
        layer4[17][31:24] = buffer_data_2[4239:4232];
        layer4[17][39:32] = buffer_data_2[4247:4240];
        layer4[17][47:40] = buffer_data_2[4255:4248];
        layer4[17][55:48] = buffer_data_2[4263:4256];
        layer5[17][7:0] = buffer_data_1[4215:4208];
        layer5[17][15:8] = buffer_data_1[4223:4216];
        layer5[17][23:16] = buffer_data_1[4231:4224];
        layer5[17][31:24] = buffer_data_1[4239:4232];
        layer5[17][39:32] = buffer_data_1[4247:4240];
        layer5[17][47:40] = buffer_data_1[4255:4248];
        layer5[17][55:48] = buffer_data_1[4263:4256];
        layer6[17][7:0] = buffer_data_0[4215:4208];
        layer6[17][15:8] = buffer_data_0[4223:4216];
        layer6[17][23:16] = buffer_data_0[4231:4224];
        layer6[17][31:24] = buffer_data_0[4239:4232];
        layer6[17][39:32] = buffer_data_0[4247:4240];
        layer6[17][47:40] = buffer_data_0[4255:4248];
        layer6[17][55:48] = buffer_data_0[4263:4256];
        layer0[18][7:0] = buffer_data_6[4223:4216];
        layer0[18][15:8] = buffer_data_6[4231:4224];
        layer0[18][23:16] = buffer_data_6[4239:4232];
        layer0[18][31:24] = buffer_data_6[4247:4240];
        layer0[18][39:32] = buffer_data_6[4255:4248];
        layer0[18][47:40] = buffer_data_6[4263:4256];
        layer0[18][55:48] = buffer_data_6[4271:4264];
        layer1[18][7:0] = buffer_data_5[4223:4216];
        layer1[18][15:8] = buffer_data_5[4231:4224];
        layer1[18][23:16] = buffer_data_5[4239:4232];
        layer1[18][31:24] = buffer_data_5[4247:4240];
        layer1[18][39:32] = buffer_data_5[4255:4248];
        layer1[18][47:40] = buffer_data_5[4263:4256];
        layer1[18][55:48] = buffer_data_5[4271:4264];
        layer2[18][7:0] = buffer_data_4[4223:4216];
        layer2[18][15:8] = buffer_data_4[4231:4224];
        layer2[18][23:16] = buffer_data_4[4239:4232];
        layer2[18][31:24] = buffer_data_4[4247:4240];
        layer2[18][39:32] = buffer_data_4[4255:4248];
        layer2[18][47:40] = buffer_data_4[4263:4256];
        layer2[18][55:48] = buffer_data_4[4271:4264];
        layer3[18][7:0] = buffer_data_3[4223:4216];
        layer3[18][15:8] = buffer_data_3[4231:4224];
        layer3[18][23:16] = buffer_data_3[4239:4232];
        layer3[18][31:24] = buffer_data_3[4247:4240];
        layer3[18][39:32] = buffer_data_3[4255:4248];
        layer3[18][47:40] = buffer_data_3[4263:4256];
        layer3[18][55:48] = buffer_data_3[4271:4264];
        layer4[18][7:0] = buffer_data_2[4223:4216];
        layer4[18][15:8] = buffer_data_2[4231:4224];
        layer4[18][23:16] = buffer_data_2[4239:4232];
        layer4[18][31:24] = buffer_data_2[4247:4240];
        layer4[18][39:32] = buffer_data_2[4255:4248];
        layer4[18][47:40] = buffer_data_2[4263:4256];
        layer4[18][55:48] = buffer_data_2[4271:4264];
        layer5[18][7:0] = buffer_data_1[4223:4216];
        layer5[18][15:8] = buffer_data_1[4231:4224];
        layer5[18][23:16] = buffer_data_1[4239:4232];
        layer5[18][31:24] = buffer_data_1[4247:4240];
        layer5[18][39:32] = buffer_data_1[4255:4248];
        layer5[18][47:40] = buffer_data_1[4263:4256];
        layer5[18][55:48] = buffer_data_1[4271:4264];
        layer6[18][7:0] = buffer_data_0[4223:4216];
        layer6[18][15:8] = buffer_data_0[4231:4224];
        layer6[18][23:16] = buffer_data_0[4239:4232];
        layer6[18][31:24] = buffer_data_0[4247:4240];
        layer6[18][39:32] = buffer_data_0[4255:4248];
        layer6[18][47:40] = buffer_data_0[4263:4256];
        layer6[18][55:48] = buffer_data_0[4271:4264];
        layer0[19][7:0] = buffer_data_6[4231:4224];
        layer0[19][15:8] = buffer_data_6[4239:4232];
        layer0[19][23:16] = buffer_data_6[4247:4240];
        layer0[19][31:24] = buffer_data_6[4255:4248];
        layer0[19][39:32] = buffer_data_6[4263:4256];
        layer0[19][47:40] = buffer_data_6[4271:4264];
        layer0[19][55:48] = buffer_data_6[4279:4272];
        layer1[19][7:0] = buffer_data_5[4231:4224];
        layer1[19][15:8] = buffer_data_5[4239:4232];
        layer1[19][23:16] = buffer_data_5[4247:4240];
        layer1[19][31:24] = buffer_data_5[4255:4248];
        layer1[19][39:32] = buffer_data_5[4263:4256];
        layer1[19][47:40] = buffer_data_5[4271:4264];
        layer1[19][55:48] = buffer_data_5[4279:4272];
        layer2[19][7:0] = buffer_data_4[4231:4224];
        layer2[19][15:8] = buffer_data_4[4239:4232];
        layer2[19][23:16] = buffer_data_4[4247:4240];
        layer2[19][31:24] = buffer_data_4[4255:4248];
        layer2[19][39:32] = buffer_data_4[4263:4256];
        layer2[19][47:40] = buffer_data_4[4271:4264];
        layer2[19][55:48] = buffer_data_4[4279:4272];
        layer3[19][7:0] = buffer_data_3[4231:4224];
        layer3[19][15:8] = buffer_data_3[4239:4232];
        layer3[19][23:16] = buffer_data_3[4247:4240];
        layer3[19][31:24] = buffer_data_3[4255:4248];
        layer3[19][39:32] = buffer_data_3[4263:4256];
        layer3[19][47:40] = buffer_data_3[4271:4264];
        layer3[19][55:48] = buffer_data_3[4279:4272];
        layer4[19][7:0] = buffer_data_2[4231:4224];
        layer4[19][15:8] = buffer_data_2[4239:4232];
        layer4[19][23:16] = buffer_data_2[4247:4240];
        layer4[19][31:24] = buffer_data_2[4255:4248];
        layer4[19][39:32] = buffer_data_2[4263:4256];
        layer4[19][47:40] = buffer_data_2[4271:4264];
        layer4[19][55:48] = buffer_data_2[4279:4272];
        layer5[19][7:0] = buffer_data_1[4231:4224];
        layer5[19][15:8] = buffer_data_1[4239:4232];
        layer5[19][23:16] = buffer_data_1[4247:4240];
        layer5[19][31:24] = buffer_data_1[4255:4248];
        layer5[19][39:32] = buffer_data_1[4263:4256];
        layer5[19][47:40] = buffer_data_1[4271:4264];
        layer5[19][55:48] = buffer_data_1[4279:4272];
        layer6[19][7:0] = buffer_data_0[4231:4224];
        layer6[19][15:8] = buffer_data_0[4239:4232];
        layer6[19][23:16] = buffer_data_0[4247:4240];
        layer6[19][31:24] = buffer_data_0[4255:4248];
        layer6[19][39:32] = buffer_data_0[4263:4256];
        layer6[19][47:40] = buffer_data_0[4271:4264];
        layer6[19][55:48] = buffer_data_0[4279:4272];
        layer0[20][7:0] = buffer_data_6[4239:4232];
        layer0[20][15:8] = buffer_data_6[4247:4240];
        layer0[20][23:16] = buffer_data_6[4255:4248];
        layer0[20][31:24] = buffer_data_6[4263:4256];
        layer0[20][39:32] = buffer_data_6[4271:4264];
        layer0[20][47:40] = buffer_data_6[4279:4272];
        layer0[20][55:48] = buffer_data_6[4287:4280];
        layer1[20][7:0] = buffer_data_5[4239:4232];
        layer1[20][15:8] = buffer_data_5[4247:4240];
        layer1[20][23:16] = buffer_data_5[4255:4248];
        layer1[20][31:24] = buffer_data_5[4263:4256];
        layer1[20][39:32] = buffer_data_5[4271:4264];
        layer1[20][47:40] = buffer_data_5[4279:4272];
        layer1[20][55:48] = buffer_data_5[4287:4280];
        layer2[20][7:0] = buffer_data_4[4239:4232];
        layer2[20][15:8] = buffer_data_4[4247:4240];
        layer2[20][23:16] = buffer_data_4[4255:4248];
        layer2[20][31:24] = buffer_data_4[4263:4256];
        layer2[20][39:32] = buffer_data_4[4271:4264];
        layer2[20][47:40] = buffer_data_4[4279:4272];
        layer2[20][55:48] = buffer_data_4[4287:4280];
        layer3[20][7:0] = buffer_data_3[4239:4232];
        layer3[20][15:8] = buffer_data_3[4247:4240];
        layer3[20][23:16] = buffer_data_3[4255:4248];
        layer3[20][31:24] = buffer_data_3[4263:4256];
        layer3[20][39:32] = buffer_data_3[4271:4264];
        layer3[20][47:40] = buffer_data_3[4279:4272];
        layer3[20][55:48] = buffer_data_3[4287:4280];
        layer4[20][7:0] = buffer_data_2[4239:4232];
        layer4[20][15:8] = buffer_data_2[4247:4240];
        layer4[20][23:16] = buffer_data_2[4255:4248];
        layer4[20][31:24] = buffer_data_2[4263:4256];
        layer4[20][39:32] = buffer_data_2[4271:4264];
        layer4[20][47:40] = buffer_data_2[4279:4272];
        layer4[20][55:48] = buffer_data_2[4287:4280];
        layer5[20][7:0] = buffer_data_1[4239:4232];
        layer5[20][15:8] = buffer_data_1[4247:4240];
        layer5[20][23:16] = buffer_data_1[4255:4248];
        layer5[20][31:24] = buffer_data_1[4263:4256];
        layer5[20][39:32] = buffer_data_1[4271:4264];
        layer5[20][47:40] = buffer_data_1[4279:4272];
        layer5[20][55:48] = buffer_data_1[4287:4280];
        layer6[20][7:0] = buffer_data_0[4239:4232];
        layer6[20][15:8] = buffer_data_0[4247:4240];
        layer6[20][23:16] = buffer_data_0[4255:4248];
        layer6[20][31:24] = buffer_data_0[4263:4256];
        layer6[20][39:32] = buffer_data_0[4271:4264];
        layer6[20][47:40] = buffer_data_0[4279:4272];
        layer6[20][55:48] = buffer_data_0[4287:4280];
        layer0[21][7:0] = buffer_data_6[4247:4240];
        layer0[21][15:8] = buffer_data_6[4255:4248];
        layer0[21][23:16] = buffer_data_6[4263:4256];
        layer0[21][31:24] = buffer_data_6[4271:4264];
        layer0[21][39:32] = buffer_data_6[4279:4272];
        layer0[21][47:40] = buffer_data_6[4287:4280];
        layer0[21][55:48] = buffer_data_6[4295:4288];
        layer1[21][7:0] = buffer_data_5[4247:4240];
        layer1[21][15:8] = buffer_data_5[4255:4248];
        layer1[21][23:16] = buffer_data_5[4263:4256];
        layer1[21][31:24] = buffer_data_5[4271:4264];
        layer1[21][39:32] = buffer_data_5[4279:4272];
        layer1[21][47:40] = buffer_data_5[4287:4280];
        layer1[21][55:48] = buffer_data_5[4295:4288];
        layer2[21][7:0] = buffer_data_4[4247:4240];
        layer2[21][15:8] = buffer_data_4[4255:4248];
        layer2[21][23:16] = buffer_data_4[4263:4256];
        layer2[21][31:24] = buffer_data_4[4271:4264];
        layer2[21][39:32] = buffer_data_4[4279:4272];
        layer2[21][47:40] = buffer_data_4[4287:4280];
        layer2[21][55:48] = buffer_data_4[4295:4288];
        layer3[21][7:0] = buffer_data_3[4247:4240];
        layer3[21][15:8] = buffer_data_3[4255:4248];
        layer3[21][23:16] = buffer_data_3[4263:4256];
        layer3[21][31:24] = buffer_data_3[4271:4264];
        layer3[21][39:32] = buffer_data_3[4279:4272];
        layer3[21][47:40] = buffer_data_3[4287:4280];
        layer3[21][55:48] = buffer_data_3[4295:4288];
        layer4[21][7:0] = buffer_data_2[4247:4240];
        layer4[21][15:8] = buffer_data_2[4255:4248];
        layer4[21][23:16] = buffer_data_2[4263:4256];
        layer4[21][31:24] = buffer_data_2[4271:4264];
        layer4[21][39:32] = buffer_data_2[4279:4272];
        layer4[21][47:40] = buffer_data_2[4287:4280];
        layer4[21][55:48] = buffer_data_2[4295:4288];
        layer5[21][7:0] = buffer_data_1[4247:4240];
        layer5[21][15:8] = buffer_data_1[4255:4248];
        layer5[21][23:16] = buffer_data_1[4263:4256];
        layer5[21][31:24] = buffer_data_1[4271:4264];
        layer5[21][39:32] = buffer_data_1[4279:4272];
        layer5[21][47:40] = buffer_data_1[4287:4280];
        layer5[21][55:48] = buffer_data_1[4295:4288];
        layer6[21][7:0] = buffer_data_0[4247:4240];
        layer6[21][15:8] = buffer_data_0[4255:4248];
        layer6[21][23:16] = buffer_data_0[4263:4256];
        layer6[21][31:24] = buffer_data_0[4271:4264];
        layer6[21][39:32] = buffer_data_0[4279:4272];
        layer6[21][47:40] = buffer_data_0[4287:4280];
        layer6[21][55:48] = buffer_data_0[4295:4288];
        layer0[22][7:0] = buffer_data_6[4255:4248];
        layer0[22][15:8] = buffer_data_6[4263:4256];
        layer0[22][23:16] = buffer_data_6[4271:4264];
        layer0[22][31:24] = buffer_data_6[4279:4272];
        layer0[22][39:32] = buffer_data_6[4287:4280];
        layer0[22][47:40] = buffer_data_6[4295:4288];
        layer0[22][55:48] = buffer_data_6[4303:4296];
        layer1[22][7:0] = buffer_data_5[4255:4248];
        layer1[22][15:8] = buffer_data_5[4263:4256];
        layer1[22][23:16] = buffer_data_5[4271:4264];
        layer1[22][31:24] = buffer_data_5[4279:4272];
        layer1[22][39:32] = buffer_data_5[4287:4280];
        layer1[22][47:40] = buffer_data_5[4295:4288];
        layer1[22][55:48] = buffer_data_5[4303:4296];
        layer2[22][7:0] = buffer_data_4[4255:4248];
        layer2[22][15:8] = buffer_data_4[4263:4256];
        layer2[22][23:16] = buffer_data_4[4271:4264];
        layer2[22][31:24] = buffer_data_4[4279:4272];
        layer2[22][39:32] = buffer_data_4[4287:4280];
        layer2[22][47:40] = buffer_data_4[4295:4288];
        layer2[22][55:48] = buffer_data_4[4303:4296];
        layer3[22][7:0] = buffer_data_3[4255:4248];
        layer3[22][15:8] = buffer_data_3[4263:4256];
        layer3[22][23:16] = buffer_data_3[4271:4264];
        layer3[22][31:24] = buffer_data_3[4279:4272];
        layer3[22][39:32] = buffer_data_3[4287:4280];
        layer3[22][47:40] = buffer_data_3[4295:4288];
        layer3[22][55:48] = buffer_data_3[4303:4296];
        layer4[22][7:0] = buffer_data_2[4255:4248];
        layer4[22][15:8] = buffer_data_2[4263:4256];
        layer4[22][23:16] = buffer_data_2[4271:4264];
        layer4[22][31:24] = buffer_data_2[4279:4272];
        layer4[22][39:32] = buffer_data_2[4287:4280];
        layer4[22][47:40] = buffer_data_2[4295:4288];
        layer4[22][55:48] = buffer_data_2[4303:4296];
        layer5[22][7:0] = buffer_data_1[4255:4248];
        layer5[22][15:8] = buffer_data_1[4263:4256];
        layer5[22][23:16] = buffer_data_1[4271:4264];
        layer5[22][31:24] = buffer_data_1[4279:4272];
        layer5[22][39:32] = buffer_data_1[4287:4280];
        layer5[22][47:40] = buffer_data_1[4295:4288];
        layer5[22][55:48] = buffer_data_1[4303:4296];
        layer6[22][7:0] = buffer_data_0[4255:4248];
        layer6[22][15:8] = buffer_data_0[4263:4256];
        layer6[22][23:16] = buffer_data_0[4271:4264];
        layer6[22][31:24] = buffer_data_0[4279:4272];
        layer6[22][39:32] = buffer_data_0[4287:4280];
        layer6[22][47:40] = buffer_data_0[4295:4288];
        layer6[22][55:48] = buffer_data_0[4303:4296];
        layer0[23][7:0] = buffer_data_6[4263:4256];
        layer0[23][15:8] = buffer_data_6[4271:4264];
        layer0[23][23:16] = buffer_data_6[4279:4272];
        layer0[23][31:24] = buffer_data_6[4287:4280];
        layer0[23][39:32] = buffer_data_6[4295:4288];
        layer0[23][47:40] = buffer_data_6[4303:4296];
        layer0[23][55:48] = buffer_data_6[4311:4304];
        layer1[23][7:0] = buffer_data_5[4263:4256];
        layer1[23][15:8] = buffer_data_5[4271:4264];
        layer1[23][23:16] = buffer_data_5[4279:4272];
        layer1[23][31:24] = buffer_data_5[4287:4280];
        layer1[23][39:32] = buffer_data_5[4295:4288];
        layer1[23][47:40] = buffer_data_5[4303:4296];
        layer1[23][55:48] = buffer_data_5[4311:4304];
        layer2[23][7:0] = buffer_data_4[4263:4256];
        layer2[23][15:8] = buffer_data_4[4271:4264];
        layer2[23][23:16] = buffer_data_4[4279:4272];
        layer2[23][31:24] = buffer_data_4[4287:4280];
        layer2[23][39:32] = buffer_data_4[4295:4288];
        layer2[23][47:40] = buffer_data_4[4303:4296];
        layer2[23][55:48] = buffer_data_4[4311:4304];
        layer3[23][7:0] = buffer_data_3[4263:4256];
        layer3[23][15:8] = buffer_data_3[4271:4264];
        layer3[23][23:16] = buffer_data_3[4279:4272];
        layer3[23][31:24] = buffer_data_3[4287:4280];
        layer3[23][39:32] = buffer_data_3[4295:4288];
        layer3[23][47:40] = buffer_data_3[4303:4296];
        layer3[23][55:48] = buffer_data_3[4311:4304];
        layer4[23][7:0] = buffer_data_2[4263:4256];
        layer4[23][15:8] = buffer_data_2[4271:4264];
        layer4[23][23:16] = buffer_data_2[4279:4272];
        layer4[23][31:24] = buffer_data_2[4287:4280];
        layer4[23][39:32] = buffer_data_2[4295:4288];
        layer4[23][47:40] = buffer_data_2[4303:4296];
        layer4[23][55:48] = buffer_data_2[4311:4304];
        layer5[23][7:0] = buffer_data_1[4263:4256];
        layer5[23][15:8] = buffer_data_1[4271:4264];
        layer5[23][23:16] = buffer_data_1[4279:4272];
        layer5[23][31:24] = buffer_data_1[4287:4280];
        layer5[23][39:32] = buffer_data_1[4295:4288];
        layer5[23][47:40] = buffer_data_1[4303:4296];
        layer5[23][55:48] = buffer_data_1[4311:4304];
        layer6[23][7:0] = buffer_data_0[4263:4256];
        layer6[23][15:8] = buffer_data_0[4271:4264];
        layer6[23][23:16] = buffer_data_0[4279:4272];
        layer6[23][31:24] = buffer_data_0[4287:4280];
        layer6[23][39:32] = buffer_data_0[4295:4288];
        layer6[23][47:40] = buffer_data_0[4303:4296];
        layer6[23][55:48] = buffer_data_0[4311:4304];
        layer0[24][7:0] = buffer_data_6[4271:4264];
        layer0[24][15:8] = buffer_data_6[4279:4272];
        layer0[24][23:16] = buffer_data_6[4287:4280];
        layer0[24][31:24] = buffer_data_6[4295:4288];
        layer0[24][39:32] = buffer_data_6[4303:4296];
        layer0[24][47:40] = buffer_data_6[4311:4304];
        layer0[24][55:48] = buffer_data_6[4319:4312];
        layer1[24][7:0] = buffer_data_5[4271:4264];
        layer1[24][15:8] = buffer_data_5[4279:4272];
        layer1[24][23:16] = buffer_data_5[4287:4280];
        layer1[24][31:24] = buffer_data_5[4295:4288];
        layer1[24][39:32] = buffer_data_5[4303:4296];
        layer1[24][47:40] = buffer_data_5[4311:4304];
        layer1[24][55:48] = buffer_data_5[4319:4312];
        layer2[24][7:0] = buffer_data_4[4271:4264];
        layer2[24][15:8] = buffer_data_4[4279:4272];
        layer2[24][23:16] = buffer_data_4[4287:4280];
        layer2[24][31:24] = buffer_data_4[4295:4288];
        layer2[24][39:32] = buffer_data_4[4303:4296];
        layer2[24][47:40] = buffer_data_4[4311:4304];
        layer2[24][55:48] = buffer_data_4[4319:4312];
        layer3[24][7:0] = buffer_data_3[4271:4264];
        layer3[24][15:8] = buffer_data_3[4279:4272];
        layer3[24][23:16] = buffer_data_3[4287:4280];
        layer3[24][31:24] = buffer_data_3[4295:4288];
        layer3[24][39:32] = buffer_data_3[4303:4296];
        layer3[24][47:40] = buffer_data_3[4311:4304];
        layer3[24][55:48] = buffer_data_3[4319:4312];
        layer4[24][7:0] = buffer_data_2[4271:4264];
        layer4[24][15:8] = buffer_data_2[4279:4272];
        layer4[24][23:16] = buffer_data_2[4287:4280];
        layer4[24][31:24] = buffer_data_2[4295:4288];
        layer4[24][39:32] = buffer_data_2[4303:4296];
        layer4[24][47:40] = buffer_data_2[4311:4304];
        layer4[24][55:48] = buffer_data_2[4319:4312];
        layer5[24][7:0] = buffer_data_1[4271:4264];
        layer5[24][15:8] = buffer_data_1[4279:4272];
        layer5[24][23:16] = buffer_data_1[4287:4280];
        layer5[24][31:24] = buffer_data_1[4295:4288];
        layer5[24][39:32] = buffer_data_1[4303:4296];
        layer5[24][47:40] = buffer_data_1[4311:4304];
        layer5[24][55:48] = buffer_data_1[4319:4312];
        layer6[24][7:0] = buffer_data_0[4271:4264];
        layer6[24][15:8] = buffer_data_0[4279:4272];
        layer6[24][23:16] = buffer_data_0[4287:4280];
        layer6[24][31:24] = buffer_data_0[4295:4288];
        layer6[24][39:32] = buffer_data_0[4303:4296];
        layer6[24][47:40] = buffer_data_0[4311:4304];
        layer6[24][55:48] = buffer_data_0[4319:4312];
        layer0[25][7:0] = buffer_data_6[4279:4272];
        layer0[25][15:8] = buffer_data_6[4287:4280];
        layer0[25][23:16] = buffer_data_6[4295:4288];
        layer0[25][31:24] = buffer_data_6[4303:4296];
        layer0[25][39:32] = buffer_data_6[4311:4304];
        layer0[25][47:40] = buffer_data_6[4319:4312];
        layer0[25][55:48] = buffer_data_6[4327:4320];
        layer1[25][7:0] = buffer_data_5[4279:4272];
        layer1[25][15:8] = buffer_data_5[4287:4280];
        layer1[25][23:16] = buffer_data_5[4295:4288];
        layer1[25][31:24] = buffer_data_5[4303:4296];
        layer1[25][39:32] = buffer_data_5[4311:4304];
        layer1[25][47:40] = buffer_data_5[4319:4312];
        layer1[25][55:48] = buffer_data_5[4327:4320];
        layer2[25][7:0] = buffer_data_4[4279:4272];
        layer2[25][15:8] = buffer_data_4[4287:4280];
        layer2[25][23:16] = buffer_data_4[4295:4288];
        layer2[25][31:24] = buffer_data_4[4303:4296];
        layer2[25][39:32] = buffer_data_4[4311:4304];
        layer2[25][47:40] = buffer_data_4[4319:4312];
        layer2[25][55:48] = buffer_data_4[4327:4320];
        layer3[25][7:0] = buffer_data_3[4279:4272];
        layer3[25][15:8] = buffer_data_3[4287:4280];
        layer3[25][23:16] = buffer_data_3[4295:4288];
        layer3[25][31:24] = buffer_data_3[4303:4296];
        layer3[25][39:32] = buffer_data_3[4311:4304];
        layer3[25][47:40] = buffer_data_3[4319:4312];
        layer3[25][55:48] = buffer_data_3[4327:4320];
        layer4[25][7:0] = buffer_data_2[4279:4272];
        layer4[25][15:8] = buffer_data_2[4287:4280];
        layer4[25][23:16] = buffer_data_2[4295:4288];
        layer4[25][31:24] = buffer_data_2[4303:4296];
        layer4[25][39:32] = buffer_data_2[4311:4304];
        layer4[25][47:40] = buffer_data_2[4319:4312];
        layer4[25][55:48] = buffer_data_2[4327:4320];
        layer5[25][7:0] = buffer_data_1[4279:4272];
        layer5[25][15:8] = buffer_data_1[4287:4280];
        layer5[25][23:16] = buffer_data_1[4295:4288];
        layer5[25][31:24] = buffer_data_1[4303:4296];
        layer5[25][39:32] = buffer_data_1[4311:4304];
        layer5[25][47:40] = buffer_data_1[4319:4312];
        layer5[25][55:48] = buffer_data_1[4327:4320];
        layer6[25][7:0] = buffer_data_0[4279:4272];
        layer6[25][15:8] = buffer_data_0[4287:4280];
        layer6[25][23:16] = buffer_data_0[4295:4288];
        layer6[25][31:24] = buffer_data_0[4303:4296];
        layer6[25][39:32] = buffer_data_0[4311:4304];
        layer6[25][47:40] = buffer_data_0[4319:4312];
        layer6[25][55:48] = buffer_data_0[4327:4320];
        layer0[26][7:0] = buffer_data_6[4287:4280];
        layer0[26][15:8] = buffer_data_6[4295:4288];
        layer0[26][23:16] = buffer_data_6[4303:4296];
        layer0[26][31:24] = buffer_data_6[4311:4304];
        layer0[26][39:32] = buffer_data_6[4319:4312];
        layer0[26][47:40] = buffer_data_6[4327:4320];
        layer0[26][55:48] = buffer_data_6[4335:4328];
        layer1[26][7:0] = buffer_data_5[4287:4280];
        layer1[26][15:8] = buffer_data_5[4295:4288];
        layer1[26][23:16] = buffer_data_5[4303:4296];
        layer1[26][31:24] = buffer_data_5[4311:4304];
        layer1[26][39:32] = buffer_data_5[4319:4312];
        layer1[26][47:40] = buffer_data_5[4327:4320];
        layer1[26][55:48] = buffer_data_5[4335:4328];
        layer2[26][7:0] = buffer_data_4[4287:4280];
        layer2[26][15:8] = buffer_data_4[4295:4288];
        layer2[26][23:16] = buffer_data_4[4303:4296];
        layer2[26][31:24] = buffer_data_4[4311:4304];
        layer2[26][39:32] = buffer_data_4[4319:4312];
        layer2[26][47:40] = buffer_data_4[4327:4320];
        layer2[26][55:48] = buffer_data_4[4335:4328];
        layer3[26][7:0] = buffer_data_3[4287:4280];
        layer3[26][15:8] = buffer_data_3[4295:4288];
        layer3[26][23:16] = buffer_data_3[4303:4296];
        layer3[26][31:24] = buffer_data_3[4311:4304];
        layer3[26][39:32] = buffer_data_3[4319:4312];
        layer3[26][47:40] = buffer_data_3[4327:4320];
        layer3[26][55:48] = buffer_data_3[4335:4328];
        layer4[26][7:0] = buffer_data_2[4287:4280];
        layer4[26][15:8] = buffer_data_2[4295:4288];
        layer4[26][23:16] = buffer_data_2[4303:4296];
        layer4[26][31:24] = buffer_data_2[4311:4304];
        layer4[26][39:32] = buffer_data_2[4319:4312];
        layer4[26][47:40] = buffer_data_2[4327:4320];
        layer4[26][55:48] = buffer_data_2[4335:4328];
        layer5[26][7:0] = buffer_data_1[4287:4280];
        layer5[26][15:8] = buffer_data_1[4295:4288];
        layer5[26][23:16] = buffer_data_1[4303:4296];
        layer5[26][31:24] = buffer_data_1[4311:4304];
        layer5[26][39:32] = buffer_data_1[4319:4312];
        layer5[26][47:40] = buffer_data_1[4327:4320];
        layer5[26][55:48] = buffer_data_1[4335:4328];
        layer6[26][7:0] = buffer_data_0[4287:4280];
        layer6[26][15:8] = buffer_data_0[4295:4288];
        layer6[26][23:16] = buffer_data_0[4303:4296];
        layer6[26][31:24] = buffer_data_0[4311:4304];
        layer6[26][39:32] = buffer_data_0[4319:4312];
        layer6[26][47:40] = buffer_data_0[4327:4320];
        layer6[26][55:48] = buffer_data_0[4335:4328];
        layer0[27][7:0] = buffer_data_6[4295:4288];
        layer0[27][15:8] = buffer_data_6[4303:4296];
        layer0[27][23:16] = buffer_data_6[4311:4304];
        layer0[27][31:24] = buffer_data_6[4319:4312];
        layer0[27][39:32] = buffer_data_6[4327:4320];
        layer0[27][47:40] = buffer_data_6[4335:4328];
        layer0[27][55:48] = buffer_data_6[4343:4336];
        layer1[27][7:0] = buffer_data_5[4295:4288];
        layer1[27][15:8] = buffer_data_5[4303:4296];
        layer1[27][23:16] = buffer_data_5[4311:4304];
        layer1[27][31:24] = buffer_data_5[4319:4312];
        layer1[27][39:32] = buffer_data_5[4327:4320];
        layer1[27][47:40] = buffer_data_5[4335:4328];
        layer1[27][55:48] = buffer_data_5[4343:4336];
        layer2[27][7:0] = buffer_data_4[4295:4288];
        layer2[27][15:8] = buffer_data_4[4303:4296];
        layer2[27][23:16] = buffer_data_4[4311:4304];
        layer2[27][31:24] = buffer_data_4[4319:4312];
        layer2[27][39:32] = buffer_data_4[4327:4320];
        layer2[27][47:40] = buffer_data_4[4335:4328];
        layer2[27][55:48] = buffer_data_4[4343:4336];
        layer3[27][7:0] = buffer_data_3[4295:4288];
        layer3[27][15:8] = buffer_data_3[4303:4296];
        layer3[27][23:16] = buffer_data_3[4311:4304];
        layer3[27][31:24] = buffer_data_3[4319:4312];
        layer3[27][39:32] = buffer_data_3[4327:4320];
        layer3[27][47:40] = buffer_data_3[4335:4328];
        layer3[27][55:48] = buffer_data_3[4343:4336];
        layer4[27][7:0] = buffer_data_2[4295:4288];
        layer4[27][15:8] = buffer_data_2[4303:4296];
        layer4[27][23:16] = buffer_data_2[4311:4304];
        layer4[27][31:24] = buffer_data_2[4319:4312];
        layer4[27][39:32] = buffer_data_2[4327:4320];
        layer4[27][47:40] = buffer_data_2[4335:4328];
        layer4[27][55:48] = buffer_data_2[4343:4336];
        layer5[27][7:0] = buffer_data_1[4295:4288];
        layer5[27][15:8] = buffer_data_1[4303:4296];
        layer5[27][23:16] = buffer_data_1[4311:4304];
        layer5[27][31:24] = buffer_data_1[4319:4312];
        layer5[27][39:32] = buffer_data_1[4327:4320];
        layer5[27][47:40] = buffer_data_1[4335:4328];
        layer5[27][55:48] = buffer_data_1[4343:4336];
        layer6[27][7:0] = buffer_data_0[4295:4288];
        layer6[27][15:8] = buffer_data_0[4303:4296];
        layer6[27][23:16] = buffer_data_0[4311:4304];
        layer6[27][31:24] = buffer_data_0[4319:4312];
        layer6[27][39:32] = buffer_data_0[4327:4320];
        layer6[27][47:40] = buffer_data_0[4335:4328];
        layer6[27][55:48] = buffer_data_0[4343:4336];
        layer0[28][7:0] = buffer_data_6[4303:4296];
        layer0[28][15:8] = buffer_data_6[4311:4304];
        layer0[28][23:16] = buffer_data_6[4319:4312];
        layer0[28][31:24] = buffer_data_6[4327:4320];
        layer0[28][39:32] = buffer_data_6[4335:4328];
        layer0[28][47:40] = buffer_data_6[4343:4336];
        layer0[28][55:48] = buffer_data_6[4351:4344];
        layer1[28][7:0] = buffer_data_5[4303:4296];
        layer1[28][15:8] = buffer_data_5[4311:4304];
        layer1[28][23:16] = buffer_data_5[4319:4312];
        layer1[28][31:24] = buffer_data_5[4327:4320];
        layer1[28][39:32] = buffer_data_5[4335:4328];
        layer1[28][47:40] = buffer_data_5[4343:4336];
        layer1[28][55:48] = buffer_data_5[4351:4344];
        layer2[28][7:0] = buffer_data_4[4303:4296];
        layer2[28][15:8] = buffer_data_4[4311:4304];
        layer2[28][23:16] = buffer_data_4[4319:4312];
        layer2[28][31:24] = buffer_data_4[4327:4320];
        layer2[28][39:32] = buffer_data_4[4335:4328];
        layer2[28][47:40] = buffer_data_4[4343:4336];
        layer2[28][55:48] = buffer_data_4[4351:4344];
        layer3[28][7:0] = buffer_data_3[4303:4296];
        layer3[28][15:8] = buffer_data_3[4311:4304];
        layer3[28][23:16] = buffer_data_3[4319:4312];
        layer3[28][31:24] = buffer_data_3[4327:4320];
        layer3[28][39:32] = buffer_data_3[4335:4328];
        layer3[28][47:40] = buffer_data_3[4343:4336];
        layer3[28][55:48] = buffer_data_3[4351:4344];
        layer4[28][7:0] = buffer_data_2[4303:4296];
        layer4[28][15:8] = buffer_data_2[4311:4304];
        layer4[28][23:16] = buffer_data_2[4319:4312];
        layer4[28][31:24] = buffer_data_2[4327:4320];
        layer4[28][39:32] = buffer_data_2[4335:4328];
        layer4[28][47:40] = buffer_data_2[4343:4336];
        layer4[28][55:48] = buffer_data_2[4351:4344];
        layer5[28][7:0] = buffer_data_1[4303:4296];
        layer5[28][15:8] = buffer_data_1[4311:4304];
        layer5[28][23:16] = buffer_data_1[4319:4312];
        layer5[28][31:24] = buffer_data_1[4327:4320];
        layer5[28][39:32] = buffer_data_1[4335:4328];
        layer5[28][47:40] = buffer_data_1[4343:4336];
        layer5[28][55:48] = buffer_data_1[4351:4344];
        layer6[28][7:0] = buffer_data_0[4303:4296];
        layer6[28][15:8] = buffer_data_0[4311:4304];
        layer6[28][23:16] = buffer_data_0[4319:4312];
        layer6[28][31:24] = buffer_data_0[4327:4320];
        layer6[28][39:32] = buffer_data_0[4335:4328];
        layer6[28][47:40] = buffer_data_0[4343:4336];
        layer6[28][55:48] = buffer_data_0[4351:4344];
        layer0[29][7:0] = buffer_data_6[4311:4304];
        layer0[29][15:8] = buffer_data_6[4319:4312];
        layer0[29][23:16] = buffer_data_6[4327:4320];
        layer0[29][31:24] = buffer_data_6[4335:4328];
        layer0[29][39:32] = buffer_data_6[4343:4336];
        layer0[29][47:40] = buffer_data_6[4351:4344];
        layer0[29][55:48] = buffer_data_6[4359:4352];
        layer1[29][7:0] = buffer_data_5[4311:4304];
        layer1[29][15:8] = buffer_data_5[4319:4312];
        layer1[29][23:16] = buffer_data_5[4327:4320];
        layer1[29][31:24] = buffer_data_5[4335:4328];
        layer1[29][39:32] = buffer_data_5[4343:4336];
        layer1[29][47:40] = buffer_data_5[4351:4344];
        layer1[29][55:48] = buffer_data_5[4359:4352];
        layer2[29][7:0] = buffer_data_4[4311:4304];
        layer2[29][15:8] = buffer_data_4[4319:4312];
        layer2[29][23:16] = buffer_data_4[4327:4320];
        layer2[29][31:24] = buffer_data_4[4335:4328];
        layer2[29][39:32] = buffer_data_4[4343:4336];
        layer2[29][47:40] = buffer_data_4[4351:4344];
        layer2[29][55:48] = buffer_data_4[4359:4352];
        layer3[29][7:0] = buffer_data_3[4311:4304];
        layer3[29][15:8] = buffer_data_3[4319:4312];
        layer3[29][23:16] = buffer_data_3[4327:4320];
        layer3[29][31:24] = buffer_data_3[4335:4328];
        layer3[29][39:32] = buffer_data_3[4343:4336];
        layer3[29][47:40] = buffer_data_3[4351:4344];
        layer3[29][55:48] = buffer_data_3[4359:4352];
        layer4[29][7:0] = buffer_data_2[4311:4304];
        layer4[29][15:8] = buffer_data_2[4319:4312];
        layer4[29][23:16] = buffer_data_2[4327:4320];
        layer4[29][31:24] = buffer_data_2[4335:4328];
        layer4[29][39:32] = buffer_data_2[4343:4336];
        layer4[29][47:40] = buffer_data_2[4351:4344];
        layer4[29][55:48] = buffer_data_2[4359:4352];
        layer5[29][7:0] = buffer_data_1[4311:4304];
        layer5[29][15:8] = buffer_data_1[4319:4312];
        layer5[29][23:16] = buffer_data_1[4327:4320];
        layer5[29][31:24] = buffer_data_1[4335:4328];
        layer5[29][39:32] = buffer_data_1[4343:4336];
        layer5[29][47:40] = buffer_data_1[4351:4344];
        layer5[29][55:48] = buffer_data_1[4359:4352];
        layer6[29][7:0] = buffer_data_0[4311:4304];
        layer6[29][15:8] = buffer_data_0[4319:4312];
        layer6[29][23:16] = buffer_data_0[4327:4320];
        layer6[29][31:24] = buffer_data_0[4335:4328];
        layer6[29][39:32] = buffer_data_0[4343:4336];
        layer6[29][47:40] = buffer_data_0[4351:4344];
        layer6[29][55:48] = buffer_data_0[4359:4352];
        layer0[30][7:0] = buffer_data_6[4319:4312];
        layer0[30][15:8] = buffer_data_6[4327:4320];
        layer0[30][23:16] = buffer_data_6[4335:4328];
        layer0[30][31:24] = buffer_data_6[4343:4336];
        layer0[30][39:32] = buffer_data_6[4351:4344];
        layer0[30][47:40] = buffer_data_6[4359:4352];
        layer0[30][55:48] = buffer_data_6[4367:4360];
        layer1[30][7:0] = buffer_data_5[4319:4312];
        layer1[30][15:8] = buffer_data_5[4327:4320];
        layer1[30][23:16] = buffer_data_5[4335:4328];
        layer1[30][31:24] = buffer_data_5[4343:4336];
        layer1[30][39:32] = buffer_data_5[4351:4344];
        layer1[30][47:40] = buffer_data_5[4359:4352];
        layer1[30][55:48] = buffer_data_5[4367:4360];
        layer2[30][7:0] = buffer_data_4[4319:4312];
        layer2[30][15:8] = buffer_data_4[4327:4320];
        layer2[30][23:16] = buffer_data_4[4335:4328];
        layer2[30][31:24] = buffer_data_4[4343:4336];
        layer2[30][39:32] = buffer_data_4[4351:4344];
        layer2[30][47:40] = buffer_data_4[4359:4352];
        layer2[30][55:48] = buffer_data_4[4367:4360];
        layer3[30][7:0] = buffer_data_3[4319:4312];
        layer3[30][15:8] = buffer_data_3[4327:4320];
        layer3[30][23:16] = buffer_data_3[4335:4328];
        layer3[30][31:24] = buffer_data_3[4343:4336];
        layer3[30][39:32] = buffer_data_3[4351:4344];
        layer3[30][47:40] = buffer_data_3[4359:4352];
        layer3[30][55:48] = buffer_data_3[4367:4360];
        layer4[30][7:0] = buffer_data_2[4319:4312];
        layer4[30][15:8] = buffer_data_2[4327:4320];
        layer4[30][23:16] = buffer_data_2[4335:4328];
        layer4[30][31:24] = buffer_data_2[4343:4336];
        layer4[30][39:32] = buffer_data_2[4351:4344];
        layer4[30][47:40] = buffer_data_2[4359:4352];
        layer4[30][55:48] = buffer_data_2[4367:4360];
        layer5[30][7:0] = buffer_data_1[4319:4312];
        layer5[30][15:8] = buffer_data_1[4327:4320];
        layer5[30][23:16] = buffer_data_1[4335:4328];
        layer5[30][31:24] = buffer_data_1[4343:4336];
        layer5[30][39:32] = buffer_data_1[4351:4344];
        layer5[30][47:40] = buffer_data_1[4359:4352];
        layer5[30][55:48] = buffer_data_1[4367:4360];
        layer6[30][7:0] = buffer_data_0[4319:4312];
        layer6[30][15:8] = buffer_data_0[4327:4320];
        layer6[30][23:16] = buffer_data_0[4335:4328];
        layer6[30][31:24] = buffer_data_0[4343:4336];
        layer6[30][39:32] = buffer_data_0[4351:4344];
        layer6[30][47:40] = buffer_data_0[4359:4352];
        layer6[30][55:48] = buffer_data_0[4367:4360];
        layer0[31][7:0] = buffer_data_6[4327:4320];
        layer0[31][15:8] = buffer_data_6[4335:4328];
        layer0[31][23:16] = buffer_data_6[4343:4336];
        layer0[31][31:24] = buffer_data_6[4351:4344];
        layer0[31][39:32] = buffer_data_6[4359:4352];
        layer0[31][47:40] = buffer_data_6[4367:4360];
        layer0[31][55:48] = buffer_data_6[4375:4368];
        layer1[31][7:0] = buffer_data_5[4327:4320];
        layer1[31][15:8] = buffer_data_5[4335:4328];
        layer1[31][23:16] = buffer_data_5[4343:4336];
        layer1[31][31:24] = buffer_data_5[4351:4344];
        layer1[31][39:32] = buffer_data_5[4359:4352];
        layer1[31][47:40] = buffer_data_5[4367:4360];
        layer1[31][55:48] = buffer_data_5[4375:4368];
        layer2[31][7:0] = buffer_data_4[4327:4320];
        layer2[31][15:8] = buffer_data_4[4335:4328];
        layer2[31][23:16] = buffer_data_4[4343:4336];
        layer2[31][31:24] = buffer_data_4[4351:4344];
        layer2[31][39:32] = buffer_data_4[4359:4352];
        layer2[31][47:40] = buffer_data_4[4367:4360];
        layer2[31][55:48] = buffer_data_4[4375:4368];
        layer3[31][7:0] = buffer_data_3[4327:4320];
        layer3[31][15:8] = buffer_data_3[4335:4328];
        layer3[31][23:16] = buffer_data_3[4343:4336];
        layer3[31][31:24] = buffer_data_3[4351:4344];
        layer3[31][39:32] = buffer_data_3[4359:4352];
        layer3[31][47:40] = buffer_data_3[4367:4360];
        layer3[31][55:48] = buffer_data_3[4375:4368];
        layer4[31][7:0] = buffer_data_2[4327:4320];
        layer4[31][15:8] = buffer_data_2[4335:4328];
        layer4[31][23:16] = buffer_data_2[4343:4336];
        layer4[31][31:24] = buffer_data_2[4351:4344];
        layer4[31][39:32] = buffer_data_2[4359:4352];
        layer4[31][47:40] = buffer_data_2[4367:4360];
        layer4[31][55:48] = buffer_data_2[4375:4368];
        layer5[31][7:0] = buffer_data_1[4327:4320];
        layer5[31][15:8] = buffer_data_1[4335:4328];
        layer5[31][23:16] = buffer_data_1[4343:4336];
        layer5[31][31:24] = buffer_data_1[4351:4344];
        layer5[31][39:32] = buffer_data_1[4359:4352];
        layer5[31][47:40] = buffer_data_1[4367:4360];
        layer5[31][55:48] = buffer_data_1[4375:4368];
        layer6[31][7:0] = buffer_data_0[4327:4320];
        layer6[31][15:8] = buffer_data_0[4335:4328];
        layer6[31][23:16] = buffer_data_0[4343:4336];
        layer6[31][31:24] = buffer_data_0[4351:4344];
        layer6[31][39:32] = buffer_data_0[4359:4352];
        layer6[31][47:40] = buffer_data_0[4367:4360];
        layer6[31][55:48] = buffer_data_0[4375:4368];
        layer0[32][7:0] = buffer_data_6[4335:4328];
        layer0[32][15:8] = buffer_data_6[4343:4336];
        layer0[32][23:16] = buffer_data_6[4351:4344];
        layer0[32][31:24] = buffer_data_6[4359:4352];
        layer0[32][39:32] = buffer_data_6[4367:4360];
        layer0[32][47:40] = buffer_data_6[4375:4368];
        layer0[32][55:48] = buffer_data_6[4383:4376];
        layer1[32][7:0] = buffer_data_5[4335:4328];
        layer1[32][15:8] = buffer_data_5[4343:4336];
        layer1[32][23:16] = buffer_data_5[4351:4344];
        layer1[32][31:24] = buffer_data_5[4359:4352];
        layer1[32][39:32] = buffer_data_5[4367:4360];
        layer1[32][47:40] = buffer_data_5[4375:4368];
        layer1[32][55:48] = buffer_data_5[4383:4376];
        layer2[32][7:0] = buffer_data_4[4335:4328];
        layer2[32][15:8] = buffer_data_4[4343:4336];
        layer2[32][23:16] = buffer_data_4[4351:4344];
        layer2[32][31:24] = buffer_data_4[4359:4352];
        layer2[32][39:32] = buffer_data_4[4367:4360];
        layer2[32][47:40] = buffer_data_4[4375:4368];
        layer2[32][55:48] = buffer_data_4[4383:4376];
        layer3[32][7:0] = buffer_data_3[4335:4328];
        layer3[32][15:8] = buffer_data_3[4343:4336];
        layer3[32][23:16] = buffer_data_3[4351:4344];
        layer3[32][31:24] = buffer_data_3[4359:4352];
        layer3[32][39:32] = buffer_data_3[4367:4360];
        layer3[32][47:40] = buffer_data_3[4375:4368];
        layer3[32][55:48] = buffer_data_3[4383:4376];
        layer4[32][7:0] = buffer_data_2[4335:4328];
        layer4[32][15:8] = buffer_data_2[4343:4336];
        layer4[32][23:16] = buffer_data_2[4351:4344];
        layer4[32][31:24] = buffer_data_2[4359:4352];
        layer4[32][39:32] = buffer_data_2[4367:4360];
        layer4[32][47:40] = buffer_data_2[4375:4368];
        layer4[32][55:48] = buffer_data_2[4383:4376];
        layer5[32][7:0] = buffer_data_1[4335:4328];
        layer5[32][15:8] = buffer_data_1[4343:4336];
        layer5[32][23:16] = buffer_data_1[4351:4344];
        layer5[32][31:24] = buffer_data_1[4359:4352];
        layer5[32][39:32] = buffer_data_1[4367:4360];
        layer5[32][47:40] = buffer_data_1[4375:4368];
        layer5[32][55:48] = buffer_data_1[4383:4376];
        layer6[32][7:0] = buffer_data_0[4335:4328];
        layer6[32][15:8] = buffer_data_0[4343:4336];
        layer6[32][23:16] = buffer_data_0[4351:4344];
        layer6[32][31:24] = buffer_data_0[4359:4352];
        layer6[32][39:32] = buffer_data_0[4367:4360];
        layer6[32][47:40] = buffer_data_0[4375:4368];
        layer6[32][55:48] = buffer_data_0[4383:4376];
        layer0[33][7:0] = buffer_data_6[4343:4336];
        layer0[33][15:8] = buffer_data_6[4351:4344];
        layer0[33][23:16] = buffer_data_6[4359:4352];
        layer0[33][31:24] = buffer_data_6[4367:4360];
        layer0[33][39:32] = buffer_data_6[4375:4368];
        layer0[33][47:40] = buffer_data_6[4383:4376];
        layer0[33][55:48] = buffer_data_6[4391:4384];
        layer1[33][7:0] = buffer_data_5[4343:4336];
        layer1[33][15:8] = buffer_data_5[4351:4344];
        layer1[33][23:16] = buffer_data_5[4359:4352];
        layer1[33][31:24] = buffer_data_5[4367:4360];
        layer1[33][39:32] = buffer_data_5[4375:4368];
        layer1[33][47:40] = buffer_data_5[4383:4376];
        layer1[33][55:48] = buffer_data_5[4391:4384];
        layer2[33][7:0] = buffer_data_4[4343:4336];
        layer2[33][15:8] = buffer_data_4[4351:4344];
        layer2[33][23:16] = buffer_data_4[4359:4352];
        layer2[33][31:24] = buffer_data_4[4367:4360];
        layer2[33][39:32] = buffer_data_4[4375:4368];
        layer2[33][47:40] = buffer_data_4[4383:4376];
        layer2[33][55:48] = buffer_data_4[4391:4384];
        layer3[33][7:0] = buffer_data_3[4343:4336];
        layer3[33][15:8] = buffer_data_3[4351:4344];
        layer3[33][23:16] = buffer_data_3[4359:4352];
        layer3[33][31:24] = buffer_data_3[4367:4360];
        layer3[33][39:32] = buffer_data_3[4375:4368];
        layer3[33][47:40] = buffer_data_3[4383:4376];
        layer3[33][55:48] = buffer_data_3[4391:4384];
        layer4[33][7:0] = buffer_data_2[4343:4336];
        layer4[33][15:8] = buffer_data_2[4351:4344];
        layer4[33][23:16] = buffer_data_2[4359:4352];
        layer4[33][31:24] = buffer_data_2[4367:4360];
        layer4[33][39:32] = buffer_data_2[4375:4368];
        layer4[33][47:40] = buffer_data_2[4383:4376];
        layer4[33][55:48] = buffer_data_2[4391:4384];
        layer5[33][7:0] = buffer_data_1[4343:4336];
        layer5[33][15:8] = buffer_data_1[4351:4344];
        layer5[33][23:16] = buffer_data_1[4359:4352];
        layer5[33][31:24] = buffer_data_1[4367:4360];
        layer5[33][39:32] = buffer_data_1[4375:4368];
        layer5[33][47:40] = buffer_data_1[4383:4376];
        layer5[33][55:48] = buffer_data_1[4391:4384];
        layer6[33][7:0] = buffer_data_0[4343:4336];
        layer6[33][15:8] = buffer_data_0[4351:4344];
        layer6[33][23:16] = buffer_data_0[4359:4352];
        layer6[33][31:24] = buffer_data_0[4367:4360];
        layer6[33][39:32] = buffer_data_0[4375:4368];
        layer6[33][47:40] = buffer_data_0[4383:4376];
        layer6[33][55:48] = buffer_data_0[4391:4384];
        layer0[34][7:0] = buffer_data_6[4351:4344];
        layer0[34][15:8] = buffer_data_6[4359:4352];
        layer0[34][23:16] = buffer_data_6[4367:4360];
        layer0[34][31:24] = buffer_data_6[4375:4368];
        layer0[34][39:32] = buffer_data_6[4383:4376];
        layer0[34][47:40] = buffer_data_6[4391:4384];
        layer0[34][55:48] = buffer_data_6[4399:4392];
        layer1[34][7:0] = buffer_data_5[4351:4344];
        layer1[34][15:8] = buffer_data_5[4359:4352];
        layer1[34][23:16] = buffer_data_5[4367:4360];
        layer1[34][31:24] = buffer_data_5[4375:4368];
        layer1[34][39:32] = buffer_data_5[4383:4376];
        layer1[34][47:40] = buffer_data_5[4391:4384];
        layer1[34][55:48] = buffer_data_5[4399:4392];
        layer2[34][7:0] = buffer_data_4[4351:4344];
        layer2[34][15:8] = buffer_data_4[4359:4352];
        layer2[34][23:16] = buffer_data_4[4367:4360];
        layer2[34][31:24] = buffer_data_4[4375:4368];
        layer2[34][39:32] = buffer_data_4[4383:4376];
        layer2[34][47:40] = buffer_data_4[4391:4384];
        layer2[34][55:48] = buffer_data_4[4399:4392];
        layer3[34][7:0] = buffer_data_3[4351:4344];
        layer3[34][15:8] = buffer_data_3[4359:4352];
        layer3[34][23:16] = buffer_data_3[4367:4360];
        layer3[34][31:24] = buffer_data_3[4375:4368];
        layer3[34][39:32] = buffer_data_3[4383:4376];
        layer3[34][47:40] = buffer_data_3[4391:4384];
        layer3[34][55:48] = buffer_data_3[4399:4392];
        layer4[34][7:0] = buffer_data_2[4351:4344];
        layer4[34][15:8] = buffer_data_2[4359:4352];
        layer4[34][23:16] = buffer_data_2[4367:4360];
        layer4[34][31:24] = buffer_data_2[4375:4368];
        layer4[34][39:32] = buffer_data_2[4383:4376];
        layer4[34][47:40] = buffer_data_2[4391:4384];
        layer4[34][55:48] = buffer_data_2[4399:4392];
        layer5[34][7:0] = buffer_data_1[4351:4344];
        layer5[34][15:8] = buffer_data_1[4359:4352];
        layer5[34][23:16] = buffer_data_1[4367:4360];
        layer5[34][31:24] = buffer_data_1[4375:4368];
        layer5[34][39:32] = buffer_data_1[4383:4376];
        layer5[34][47:40] = buffer_data_1[4391:4384];
        layer5[34][55:48] = buffer_data_1[4399:4392];
        layer6[34][7:0] = buffer_data_0[4351:4344];
        layer6[34][15:8] = buffer_data_0[4359:4352];
        layer6[34][23:16] = buffer_data_0[4367:4360];
        layer6[34][31:24] = buffer_data_0[4375:4368];
        layer6[34][39:32] = buffer_data_0[4383:4376];
        layer6[34][47:40] = buffer_data_0[4391:4384];
        layer6[34][55:48] = buffer_data_0[4399:4392];
        layer0[35][7:0] = buffer_data_6[4359:4352];
        layer0[35][15:8] = buffer_data_6[4367:4360];
        layer0[35][23:16] = buffer_data_6[4375:4368];
        layer0[35][31:24] = buffer_data_6[4383:4376];
        layer0[35][39:32] = buffer_data_6[4391:4384];
        layer0[35][47:40] = buffer_data_6[4399:4392];
        layer0[35][55:48] = buffer_data_6[4407:4400];
        layer1[35][7:0] = buffer_data_5[4359:4352];
        layer1[35][15:8] = buffer_data_5[4367:4360];
        layer1[35][23:16] = buffer_data_5[4375:4368];
        layer1[35][31:24] = buffer_data_5[4383:4376];
        layer1[35][39:32] = buffer_data_5[4391:4384];
        layer1[35][47:40] = buffer_data_5[4399:4392];
        layer1[35][55:48] = buffer_data_5[4407:4400];
        layer2[35][7:0] = buffer_data_4[4359:4352];
        layer2[35][15:8] = buffer_data_4[4367:4360];
        layer2[35][23:16] = buffer_data_4[4375:4368];
        layer2[35][31:24] = buffer_data_4[4383:4376];
        layer2[35][39:32] = buffer_data_4[4391:4384];
        layer2[35][47:40] = buffer_data_4[4399:4392];
        layer2[35][55:48] = buffer_data_4[4407:4400];
        layer3[35][7:0] = buffer_data_3[4359:4352];
        layer3[35][15:8] = buffer_data_3[4367:4360];
        layer3[35][23:16] = buffer_data_3[4375:4368];
        layer3[35][31:24] = buffer_data_3[4383:4376];
        layer3[35][39:32] = buffer_data_3[4391:4384];
        layer3[35][47:40] = buffer_data_3[4399:4392];
        layer3[35][55:48] = buffer_data_3[4407:4400];
        layer4[35][7:0] = buffer_data_2[4359:4352];
        layer4[35][15:8] = buffer_data_2[4367:4360];
        layer4[35][23:16] = buffer_data_2[4375:4368];
        layer4[35][31:24] = buffer_data_2[4383:4376];
        layer4[35][39:32] = buffer_data_2[4391:4384];
        layer4[35][47:40] = buffer_data_2[4399:4392];
        layer4[35][55:48] = buffer_data_2[4407:4400];
        layer5[35][7:0] = buffer_data_1[4359:4352];
        layer5[35][15:8] = buffer_data_1[4367:4360];
        layer5[35][23:16] = buffer_data_1[4375:4368];
        layer5[35][31:24] = buffer_data_1[4383:4376];
        layer5[35][39:32] = buffer_data_1[4391:4384];
        layer5[35][47:40] = buffer_data_1[4399:4392];
        layer5[35][55:48] = buffer_data_1[4407:4400];
        layer6[35][7:0] = buffer_data_0[4359:4352];
        layer6[35][15:8] = buffer_data_0[4367:4360];
        layer6[35][23:16] = buffer_data_0[4375:4368];
        layer6[35][31:24] = buffer_data_0[4383:4376];
        layer6[35][39:32] = buffer_data_0[4391:4384];
        layer6[35][47:40] = buffer_data_0[4399:4392];
        layer6[35][55:48] = buffer_data_0[4407:4400];
        layer0[36][7:0] = buffer_data_6[4367:4360];
        layer0[36][15:8] = buffer_data_6[4375:4368];
        layer0[36][23:16] = buffer_data_6[4383:4376];
        layer0[36][31:24] = buffer_data_6[4391:4384];
        layer0[36][39:32] = buffer_data_6[4399:4392];
        layer0[36][47:40] = buffer_data_6[4407:4400];
        layer0[36][55:48] = buffer_data_6[4415:4408];
        layer1[36][7:0] = buffer_data_5[4367:4360];
        layer1[36][15:8] = buffer_data_5[4375:4368];
        layer1[36][23:16] = buffer_data_5[4383:4376];
        layer1[36][31:24] = buffer_data_5[4391:4384];
        layer1[36][39:32] = buffer_data_5[4399:4392];
        layer1[36][47:40] = buffer_data_5[4407:4400];
        layer1[36][55:48] = buffer_data_5[4415:4408];
        layer2[36][7:0] = buffer_data_4[4367:4360];
        layer2[36][15:8] = buffer_data_4[4375:4368];
        layer2[36][23:16] = buffer_data_4[4383:4376];
        layer2[36][31:24] = buffer_data_4[4391:4384];
        layer2[36][39:32] = buffer_data_4[4399:4392];
        layer2[36][47:40] = buffer_data_4[4407:4400];
        layer2[36][55:48] = buffer_data_4[4415:4408];
        layer3[36][7:0] = buffer_data_3[4367:4360];
        layer3[36][15:8] = buffer_data_3[4375:4368];
        layer3[36][23:16] = buffer_data_3[4383:4376];
        layer3[36][31:24] = buffer_data_3[4391:4384];
        layer3[36][39:32] = buffer_data_3[4399:4392];
        layer3[36][47:40] = buffer_data_3[4407:4400];
        layer3[36][55:48] = buffer_data_3[4415:4408];
        layer4[36][7:0] = buffer_data_2[4367:4360];
        layer4[36][15:8] = buffer_data_2[4375:4368];
        layer4[36][23:16] = buffer_data_2[4383:4376];
        layer4[36][31:24] = buffer_data_2[4391:4384];
        layer4[36][39:32] = buffer_data_2[4399:4392];
        layer4[36][47:40] = buffer_data_2[4407:4400];
        layer4[36][55:48] = buffer_data_2[4415:4408];
        layer5[36][7:0] = buffer_data_1[4367:4360];
        layer5[36][15:8] = buffer_data_1[4375:4368];
        layer5[36][23:16] = buffer_data_1[4383:4376];
        layer5[36][31:24] = buffer_data_1[4391:4384];
        layer5[36][39:32] = buffer_data_1[4399:4392];
        layer5[36][47:40] = buffer_data_1[4407:4400];
        layer5[36][55:48] = buffer_data_1[4415:4408];
        layer6[36][7:0] = buffer_data_0[4367:4360];
        layer6[36][15:8] = buffer_data_0[4375:4368];
        layer6[36][23:16] = buffer_data_0[4383:4376];
        layer6[36][31:24] = buffer_data_0[4391:4384];
        layer6[36][39:32] = buffer_data_0[4399:4392];
        layer6[36][47:40] = buffer_data_0[4407:4400];
        layer6[36][55:48] = buffer_data_0[4415:4408];
        layer0[37][7:0] = buffer_data_6[4375:4368];
        layer0[37][15:8] = buffer_data_6[4383:4376];
        layer0[37][23:16] = buffer_data_6[4391:4384];
        layer0[37][31:24] = buffer_data_6[4399:4392];
        layer0[37][39:32] = buffer_data_6[4407:4400];
        layer0[37][47:40] = buffer_data_6[4415:4408];
        layer0[37][55:48] = buffer_data_6[4423:4416];
        layer1[37][7:0] = buffer_data_5[4375:4368];
        layer1[37][15:8] = buffer_data_5[4383:4376];
        layer1[37][23:16] = buffer_data_5[4391:4384];
        layer1[37][31:24] = buffer_data_5[4399:4392];
        layer1[37][39:32] = buffer_data_5[4407:4400];
        layer1[37][47:40] = buffer_data_5[4415:4408];
        layer1[37][55:48] = buffer_data_5[4423:4416];
        layer2[37][7:0] = buffer_data_4[4375:4368];
        layer2[37][15:8] = buffer_data_4[4383:4376];
        layer2[37][23:16] = buffer_data_4[4391:4384];
        layer2[37][31:24] = buffer_data_4[4399:4392];
        layer2[37][39:32] = buffer_data_4[4407:4400];
        layer2[37][47:40] = buffer_data_4[4415:4408];
        layer2[37][55:48] = buffer_data_4[4423:4416];
        layer3[37][7:0] = buffer_data_3[4375:4368];
        layer3[37][15:8] = buffer_data_3[4383:4376];
        layer3[37][23:16] = buffer_data_3[4391:4384];
        layer3[37][31:24] = buffer_data_3[4399:4392];
        layer3[37][39:32] = buffer_data_3[4407:4400];
        layer3[37][47:40] = buffer_data_3[4415:4408];
        layer3[37][55:48] = buffer_data_3[4423:4416];
        layer4[37][7:0] = buffer_data_2[4375:4368];
        layer4[37][15:8] = buffer_data_2[4383:4376];
        layer4[37][23:16] = buffer_data_2[4391:4384];
        layer4[37][31:24] = buffer_data_2[4399:4392];
        layer4[37][39:32] = buffer_data_2[4407:4400];
        layer4[37][47:40] = buffer_data_2[4415:4408];
        layer4[37][55:48] = buffer_data_2[4423:4416];
        layer5[37][7:0] = buffer_data_1[4375:4368];
        layer5[37][15:8] = buffer_data_1[4383:4376];
        layer5[37][23:16] = buffer_data_1[4391:4384];
        layer5[37][31:24] = buffer_data_1[4399:4392];
        layer5[37][39:32] = buffer_data_1[4407:4400];
        layer5[37][47:40] = buffer_data_1[4415:4408];
        layer5[37][55:48] = buffer_data_1[4423:4416];
        layer6[37][7:0] = buffer_data_0[4375:4368];
        layer6[37][15:8] = buffer_data_0[4383:4376];
        layer6[37][23:16] = buffer_data_0[4391:4384];
        layer6[37][31:24] = buffer_data_0[4399:4392];
        layer6[37][39:32] = buffer_data_0[4407:4400];
        layer6[37][47:40] = buffer_data_0[4415:4408];
        layer6[37][55:48] = buffer_data_0[4423:4416];
        layer0[38][7:0] = buffer_data_6[4383:4376];
        layer0[38][15:8] = buffer_data_6[4391:4384];
        layer0[38][23:16] = buffer_data_6[4399:4392];
        layer0[38][31:24] = buffer_data_6[4407:4400];
        layer0[38][39:32] = buffer_data_6[4415:4408];
        layer0[38][47:40] = buffer_data_6[4423:4416];
        layer0[38][55:48] = buffer_data_6[4431:4424];
        layer1[38][7:0] = buffer_data_5[4383:4376];
        layer1[38][15:8] = buffer_data_5[4391:4384];
        layer1[38][23:16] = buffer_data_5[4399:4392];
        layer1[38][31:24] = buffer_data_5[4407:4400];
        layer1[38][39:32] = buffer_data_5[4415:4408];
        layer1[38][47:40] = buffer_data_5[4423:4416];
        layer1[38][55:48] = buffer_data_5[4431:4424];
        layer2[38][7:0] = buffer_data_4[4383:4376];
        layer2[38][15:8] = buffer_data_4[4391:4384];
        layer2[38][23:16] = buffer_data_4[4399:4392];
        layer2[38][31:24] = buffer_data_4[4407:4400];
        layer2[38][39:32] = buffer_data_4[4415:4408];
        layer2[38][47:40] = buffer_data_4[4423:4416];
        layer2[38][55:48] = buffer_data_4[4431:4424];
        layer3[38][7:0] = buffer_data_3[4383:4376];
        layer3[38][15:8] = buffer_data_3[4391:4384];
        layer3[38][23:16] = buffer_data_3[4399:4392];
        layer3[38][31:24] = buffer_data_3[4407:4400];
        layer3[38][39:32] = buffer_data_3[4415:4408];
        layer3[38][47:40] = buffer_data_3[4423:4416];
        layer3[38][55:48] = buffer_data_3[4431:4424];
        layer4[38][7:0] = buffer_data_2[4383:4376];
        layer4[38][15:8] = buffer_data_2[4391:4384];
        layer4[38][23:16] = buffer_data_2[4399:4392];
        layer4[38][31:24] = buffer_data_2[4407:4400];
        layer4[38][39:32] = buffer_data_2[4415:4408];
        layer4[38][47:40] = buffer_data_2[4423:4416];
        layer4[38][55:48] = buffer_data_2[4431:4424];
        layer5[38][7:0] = buffer_data_1[4383:4376];
        layer5[38][15:8] = buffer_data_1[4391:4384];
        layer5[38][23:16] = buffer_data_1[4399:4392];
        layer5[38][31:24] = buffer_data_1[4407:4400];
        layer5[38][39:32] = buffer_data_1[4415:4408];
        layer5[38][47:40] = buffer_data_1[4423:4416];
        layer5[38][55:48] = buffer_data_1[4431:4424];
        layer6[38][7:0] = buffer_data_0[4383:4376];
        layer6[38][15:8] = buffer_data_0[4391:4384];
        layer6[38][23:16] = buffer_data_0[4399:4392];
        layer6[38][31:24] = buffer_data_0[4407:4400];
        layer6[38][39:32] = buffer_data_0[4415:4408];
        layer6[38][47:40] = buffer_data_0[4423:4416];
        layer6[38][55:48] = buffer_data_0[4431:4424];
        layer0[39][7:0] = buffer_data_6[4391:4384];
        layer0[39][15:8] = buffer_data_6[4399:4392];
        layer0[39][23:16] = buffer_data_6[4407:4400];
        layer0[39][31:24] = buffer_data_6[4415:4408];
        layer0[39][39:32] = buffer_data_6[4423:4416];
        layer0[39][47:40] = buffer_data_6[4431:4424];
        layer0[39][55:48] = buffer_data_6[4439:4432];
        layer1[39][7:0] = buffer_data_5[4391:4384];
        layer1[39][15:8] = buffer_data_5[4399:4392];
        layer1[39][23:16] = buffer_data_5[4407:4400];
        layer1[39][31:24] = buffer_data_5[4415:4408];
        layer1[39][39:32] = buffer_data_5[4423:4416];
        layer1[39][47:40] = buffer_data_5[4431:4424];
        layer1[39][55:48] = buffer_data_5[4439:4432];
        layer2[39][7:0] = buffer_data_4[4391:4384];
        layer2[39][15:8] = buffer_data_4[4399:4392];
        layer2[39][23:16] = buffer_data_4[4407:4400];
        layer2[39][31:24] = buffer_data_4[4415:4408];
        layer2[39][39:32] = buffer_data_4[4423:4416];
        layer2[39][47:40] = buffer_data_4[4431:4424];
        layer2[39][55:48] = buffer_data_4[4439:4432];
        layer3[39][7:0] = buffer_data_3[4391:4384];
        layer3[39][15:8] = buffer_data_3[4399:4392];
        layer3[39][23:16] = buffer_data_3[4407:4400];
        layer3[39][31:24] = buffer_data_3[4415:4408];
        layer3[39][39:32] = buffer_data_3[4423:4416];
        layer3[39][47:40] = buffer_data_3[4431:4424];
        layer3[39][55:48] = buffer_data_3[4439:4432];
        layer4[39][7:0] = buffer_data_2[4391:4384];
        layer4[39][15:8] = buffer_data_2[4399:4392];
        layer4[39][23:16] = buffer_data_2[4407:4400];
        layer4[39][31:24] = buffer_data_2[4415:4408];
        layer4[39][39:32] = buffer_data_2[4423:4416];
        layer4[39][47:40] = buffer_data_2[4431:4424];
        layer4[39][55:48] = buffer_data_2[4439:4432];
        layer5[39][7:0] = buffer_data_1[4391:4384];
        layer5[39][15:8] = buffer_data_1[4399:4392];
        layer5[39][23:16] = buffer_data_1[4407:4400];
        layer5[39][31:24] = buffer_data_1[4415:4408];
        layer5[39][39:32] = buffer_data_1[4423:4416];
        layer5[39][47:40] = buffer_data_1[4431:4424];
        layer5[39][55:48] = buffer_data_1[4439:4432];
        layer6[39][7:0] = buffer_data_0[4391:4384];
        layer6[39][15:8] = buffer_data_0[4399:4392];
        layer6[39][23:16] = buffer_data_0[4407:4400];
        layer6[39][31:24] = buffer_data_0[4415:4408];
        layer6[39][39:32] = buffer_data_0[4423:4416];
        layer6[39][47:40] = buffer_data_0[4431:4424];
        layer6[39][55:48] = buffer_data_0[4439:4432];
        layer0[40][7:0] = buffer_data_6[4399:4392];
        layer0[40][15:8] = buffer_data_6[4407:4400];
        layer0[40][23:16] = buffer_data_6[4415:4408];
        layer0[40][31:24] = buffer_data_6[4423:4416];
        layer0[40][39:32] = buffer_data_6[4431:4424];
        layer0[40][47:40] = buffer_data_6[4439:4432];
        layer0[40][55:48] = buffer_data_6[4447:4440];
        layer1[40][7:0] = buffer_data_5[4399:4392];
        layer1[40][15:8] = buffer_data_5[4407:4400];
        layer1[40][23:16] = buffer_data_5[4415:4408];
        layer1[40][31:24] = buffer_data_5[4423:4416];
        layer1[40][39:32] = buffer_data_5[4431:4424];
        layer1[40][47:40] = buffer_data_5[4439:4432];
        layer1[40][55:48] = buffer_data_5[4447:4440];
        layer2[40][7:0] = buffer_data_4[4399:4392];
        layer2[40][15:8] = buffer_data_4[4407:4400];
        layer2[40][23:16] = buffer_data_4[4415:4408];
        layer2[40][31:24] = buffer_data_4[4423:4416];
        layer2[40][39:32] = buffer_data_4[4431:4424];
        layer2[40][47:40] = buffer_data_4[4439:4432];
        layer2[40][55:48] = buffer_data_4[4447:4440];
        layer3[40][7:0] = buffer_data_3[4399:4392];
        layer3[40][15:8] = buffer_data_3[4407:4400];
        layer3[40][23:16] = buffer_data_3[4415:4408];
        layer3[40][31:24] = buffer_data_3[4423:4416];
        layer3[40][39:32] = buffer_data_3[4431:4424];
        layer3[40][47:40] = buffer_data_3[4439:4432];
        layer3[40][55:48] = buffer_data_3[4447:4440];
        layer4[40][7:0] = buffer_data_2[4399:4392];
        layer4[40][15:8] = buffer_data_2[4407:4400];
        layer4[40][23:16] = buffer_data_2[4415:4408];
        layer4[40][31:24] = buffer_data_2[4423:4416];
        layer4[40][39:32] = buffer_data_2[4431:4424];
        layer4[40][47:40] = buffer_data_2[4439:4432];
        layer4[40][55:48] = buffer_data_2[4447:4440];
        layer5[40][7:0] = buffer_data_1[4399:4392];
        layer5[40][15:8] = buffer_data_1[4407:4400];
        layer5[40][23:16] = buffer_data_1[4415:4408];
        layer5[40][31:24] = buffer_data_1[4423:4416];
        layer5[40][39:32] = buffer_data_1[4431:4424];
        layer5[40][47:40] = buffer_data_1[4439:4432];
        layer5[40][55:48] = buffer_data_1[4447:4440];
        layer6[40][7:0] = buffer_data_0[4399:4392];
        layer6[40][15:8] = buffer_data_0[4407:4400];
        layer6[40][23:16] = buffer_data_0[4415:4408];
        layer6[40][31:24] = buffer_data_0[4423:4416];
        layer6[40][39:32] = buffer_data_0[4431:4424];
        layer6[40][47:40] = buffer_data_0[4439:4432];
        layer6[40][55:48] = buffer_data_0[4447:4440];
        layer0[41][7:0] = buffer_data_6[4407:4400];
        layer0[41][15:8] = buffer_data_6[4415:4408];
        layer0[41][23:16] = buffer_data_6[4423:4416];
        layer0[41][31:24] = buffer_data_6[4431:4424];
        layer0[41][39:32] = buffer_data_6[4439:4432];
        layer0[41][47:40] = buffer_data_6[4447:4440];
        layer0[41][55:48] = buffer_data_6[4455:4448];
        layer1[41][7:0] = buffer_data_5[4407:4400];
        layer1[41][15:8] = buffer_data_5[4415:4408];
        layer1[41][23:16] = buffer_data_5[4423:4416];
        layer1[41][31:24] = buffer_data_5[4431:4424];
        layer1[41][39:32] = buffer_data_5[4439:4432];
        layer1[41][47:40] = buffer_data_5[4447:4440];
        layer1[41][55:48] = buffer_data_5[4455:4448];
        layer2[41][7:0] = buffer_data_4[4407:4400];
        layer2[41][15:8] = buffer_data_4[4415:4408];
        layer2[41][23:16] = buffer_data_4[4423:4416];
        layer2[41][31:24] = buffer_data_4[4431:4424];
        layer2[41][39:32] = buffer_data_4[4439:4432];
        layer2[41][47:40] = buffer_data_4[4447:4440];
        layer2[41][55:48] = buffer_data_4[4455:4448];
        layer3[41][7:0] = buffer_data_3[4407:4400];
        layer3[41][15:8] = buffer_data_3[4415:4408];
        layer3[41][23:16] = buffer_data_3[4423:4416];
        layer3[41][31:24] = buffer_data_3[4431:4424];
        layer3[41][39:32] = buffer_data_3[4439:4432];
        layer3[41][47:40] = buffer_data_3[4447:4440];
        layer3[41][55:48] = buffer_data_3[4455:4448];
        layer4[41][7:0] = buffer_data_2[4407:4400];
        layer4[41][15:8] = buffer_data_2[4415:4408];
        layer4[41][23:16] = buffer_data_2[4423:4416];
        layer4[41][31:24] = buffer_data_2[4431:4424];
        layer4[41][39:32] = buffer_data_2[4439:4432];
        layer4[41][47:40] = buffer_data_2[4447:4440];
        layer4[41][55:48] = buffer_data_2[4455:4448];
        layer5[41][7:0] = buffer_data_1[4407:4400];
        layer5[41][15:8] = buffer_data_1[4415:4408];
        layer5[41][23:16] = buffer_data_1[4423:4416];
        layer5[41][31:24] = buffer_data_1[4431:4424];
        layer5[41][39:32] = buffer_data_1[4439:4432];
        layer5[41][47:40] = buffer_data_1[4447:4440];
        layer5[41][55:48] = buffer_data_1[4455:4448];
        layer6[41][7:0] = buffer_data_0[4407:4400];
        layer6[41][15:8] = buffer_data_0[4415:4408];
        layer6[41][23:16] = buffer_data_0[4423:4416];
        layer6[41][31:24] = buffer_data_0[4431:4424];
        layer6[41][39:32] = buffer_data_0[4439:4432];
        layer6[41][47:40] = buffer_data_0[4447:4440];
        layer6[41][55:48] = buffer_data_0[4455:4448];
        layer0[42][7:0] = buffer_data_6[4415:4408];
        layer0[42][15:8] = buffer_data_6[4423:4416];
        layer0[42][23:16] = buffer_data_6[4431:4424];
        layer0[42][31:24] = buffer_data_6[4439:4432];
        layer0[42][39:32] = buffer_data_6[4447:4440];
        layer0[42][47:40] = buffer_data_6[4455:4448];
        layer0[42][55:48] = buffer_data_6[4463:4456];
        layer1[42][7:0] = buffer_data_5[4415:4408];
        layer1[42][15:8] = buffer_data_5[4423:4416];
        layer1[42][23:16] = buffer_data_5[4431:4424];
        layer1[42][31:24] = buffer_data_5[4439:4432];
        layer1[42][39:32] = buffer_data_5[4447:4440];
        layer1[42][47:40] = buffer_data_5[4455:4448];
        layer1[42][55:48] = buffer_data_5[4463:4456];
        layer2[42][7:0] = buffer_data_4[4415:4408];
        layer2[42][15:8] = buffer_data_4[4423:4416];
        layer2[42][23:16] = buffer_data_4[4431:4424];
        layer2[42][31:24] = buffer_data_4[4439:4432];
        layer2[42][39:32] = buffer_data_4[4447:4440];
        layer2[42][47:40] = buffer_data_4[4455:4448];
        layer2[42][55:48] = buffer_data_4[4463:4456];
        layer3[42][7:0] = buffer_data_3[4415:4408];
        layer3[42][15:8] = buffer_data_3[4423:4416];
        layer3[42][23:16] = buffer_data_3[4431:4424];
        layer3[42][31:24] = buffer_data_3[4439:4432];
        layer3[42][39:32] = buffer_data_3[4447:4440];
        layer3[42][47:40] = buffer_data_3[4455:4448];
        layer3[42][55:48] = buffer_data_3[4463:4456];
        layer4[42][7:0] = buffer_data_2[4415:4408];
        layer4[42][15:8] = buffer_data_2[4423:4416];
        layer4[42][23:16] = buffer_data_2[4431:4424];
        layer4[42][31:24] = buffer_data_2[4439:4432];
        layer4[42][39:32] = buffer_data_2[4447:4440];
        layer4[42][47:40] = buffer_data_2[4455:4448];
        layer4[42][55:48] = buffer_data_2[4463:4456];
        layer5[42][7:0] = buffer_data_1[4415:4408];
        layer5[42][15:8] = buffer_data_1[4423:4416];
        layer5[42][23:16] = buffer_data_1[4431:4424];
        layer5[42][31:24] = buffer_data_1[4439:4432];
        layer5[42][39:32] = buffer_data_1[4447:4440];
        layer5[42][47:40] = buffer_data_1[4455:4448];
        layer5[42][55:48] = buffer_data_1[4463:4456];
        layer6[42][7:0] = buffer_data_0[4415:4408];
        layer6[42][15:8] = buffer_data_0[4423:4416];
        layer6[42][23:16] = buffer_data_0[4431:4424];
        layer6[42][31:24] = buffer_data_0[4439:4432];
        layer6[42][39:32] = buffer_data_0[4447:4440];
        layer6[42][47:40] = buffer_data_0[4455:4448];
        layer6[42][55:48] = buffer_data_0[4463:4456];
        layer0[43][7:0] = buffer_data_6[4423:4416];
        layer0[43][15:8] = buffer_data_6[4431:4424];
        layer0[43][23:16] = buffer_data_6[4439:4432];
        layer0[43][31:24] = buffer_data_6[4447:4440];
        layer0[43][39:32] = buffer_data_6[4455:4448];
        layer0[43][47:40] = buffer_data_6[4463:4456];
        layer0[43][55:48] = buffer_data_6[4471:4464];
        layer1[43][7:0] = buffer_data_5[4423:4416];
        layer1[43][15:8] = buffer_data_5[4431:4424];
        layer1[43][23:16] = buffer_data_5[4439:4432];
        layer1[43][31:24] = buffer_data_5[4447:4440];
        layer1[43][39:32] = buffer_data_5[4455:4448];
        layer1[43][47:40] = buffer_data_5[4463:4456];
        layer1[43][55:48] = buffer_data_5[4471:4464];
        layer2[43][7:0] = buffer_data_4[4423:4416];
        layer2[43][15:8] = buffer_data_4[4431:4424];
        layer2[43][23:16] = buffer_data_4[4439:4432];
        layer2[43][31:24] = buffer_data_4[4447:4440];
        layer2[43][39:32] = buffer_data_4[4455:4448];
        layer2[43][47:40] = buffer_data_4[4463:4456];
        layer2[43][55:48] = buffer_data_4[4471:4464];
        layer3[43][7:0] = buffer_data_3[4423:4416];
        layer3[43][15:8] = buffer_data_3[4431:4424];
        layer3[43][23:16] = buffer_data_3[4439:4432];
        layer3[43][31:24] = buffer_data_3[4447:4440];
        layer3[43][39:32] = buffer_data_3[4455:4448];
        layer3[43][47:40] = buffer_data_3[4463:4456];
        layer3[43][55:48] = buffer_data_3[4471:4464];
        layer4[43][7:0] = buffer_data_2[4423:4416];
        layer4[43][15:8] = buffer_data_2[4431:4424];
        layer4[43][23:16] = buffer_data_2[4439:4432];
        layer4[43][31:24] = buffer_data_2[4447:4440];
        layer4[43][39:32] = buffer_data_2[4455:4448];
        layer4[43][47:40] = buffer_data_2[4463:4456];
        layer4[43][55:48] = buffer_data_2[4471:4464];
        layer5[43][7:0] = buffer_data_1[4423:4416];
        layer5[43][15:8] = buffer_data_1[4431:4424];
        layer5[43][23:16] = buffer_data_1[4439:4432];
        layer5[43][31:24] = buffer_data_1[4447:4440];
        layer5[43][39:32] = buffer_data_1[4455:4448];
        layer5[43][47:40] = buffer_data_1[4463:4456];
        layer5[43][55:48] = buffer_data_1[4471:4464];
        layer6[43][7:0] = buffer_data_0[4423:4416];
        layer6[43][15:8] = buffer_data_0[4431:4424];
        layer6[43][23:16] = buffer_data_0[4439:4432];
        layer6[43][31:24] = buffer_data_0[4447:4440];
        layer6[43][39:32] = buffer_data_0[4455:4448];
        layer6[43][47:40] = buffer_data_0[4463:4456];
        layer6[43][55:48] = buffer_data_0[4471:4464];
        layer0[44][7:0] = buffer_data_6[4431:4424];
        layer0[44][15:8] = buffer_data_6[4439:4432];
        layer0[44][23:16] = buffer_data_6[4447:4440];
        layer0[44][31:24] = buffer_data_6[4455:4448];
        layer0[44][39:32] = buffer_data_6[4463:4456];
        layer0[44][47:40] = buffer_data_6[4471:4464];
        layer0[44][55:48] = buffer_data_6[4479:4472];
        layer1[44][7:0] = buffer_data_5[4431:4424];
        layer1[44][15:8] = buffer_data_5[4439:4432];
        layer1[44][23:16] = buffer_data_5[4447:4440];
        layer1[44][31:24] = buffer_data_5[4455:4448];
        layer1[44][39:32] = buffer_data_5[4463:4456];
        layer1[44][47:40] = buffer_data_5[4471:4464];
        layer1[44][55:48] = buffer_data_5[4479:4472];
        layer2[44][7:0] = buffer_data_4[4431:4424];
        layer2[44][15:8] = buffer_data_4[4439:4432];
        layer2[44][23:16] = buffer_data_4[4447:4440];
        layer2[44][31:24] = buffer_data_4[4455:4448];
        layer2[44][39:32] = buffer_data_4[4463:4456];
        layer2[44][47:40] = buffer_data_4[4471:4464];
        layer2[44][55:48] = buffer_data_4[4479:4472];
        layer3[44][7:0] = buffer_data_3[4431:4424];
        layer3[44][15:8] = buffer_data_3[4439:4432];
        layer3[44][23:16] = buffer_data_3[4447:4440];
        layer3[44][31:24] = buffer_data_3[4455:4448];
        layer3[44][39:32] = buffer_data_3[4463:4456];
        layer3[44][47:40] = buffer_data_3[4471:4464];
        layer3[44][55:48] = buffer_data_3[4479:4472];
        layer4[44][7:0] = buffer_data_2[4431:4424];
        layer4[44][15:8] = buffer_data_2[4439:4432];
        layer4[44][23:16] = buffer_data_2[4447:4440];
        layer4[44][31:24] = buffer_data_2[4455:4448];
        layer4[44][39:32] = buffer_data_2[4463:4456];
        layer4[44][47:40] = buffer_data_2[4471:4464];
        layer4[44][55:48] = buffer_data_2[4479:4472];
        layer5[44][7:0] = buffer_data_1[4431:4424];
        layer5[44][15:8] = buffer_data_1[4439:4432];
        layer5[44][23:16] = buffer_data_1[4447:4440];
        layer5[44][31:24] = buffer_data_1[4455:4448];
        layer5[44][39:32] = buffer_data_1[4463:4456];
        layer5[44][47:40] = buffer_data_1[4471:4464];
        layer5[44][55:48] = buffer_data_1[4479:4472];
        layer6[44][7:0] = buffer_data_0[4431:4424];
        layer6[44][15:8] = buffer_data_0[4439:4432];
        layer6[44][23:16] = buffer_data_0[4447:4440];
        layer6[44][31:24] = buffer_data_0[4455:4448];
        layer6[44][39:32] = buffer_data_0[4463:4456];
        layer6[44][47:40] = buffer_data_0[4471:4464];
        layer6[44][55:48] = buffer_data_0[4479:4472];
        layer0[45][7:0] = buffer_data_6[4439:4432];
        layer0[45][15:8] = buffer_data_6[4447:4440];
        layer0[45][23:16] = buffer_data_6[4455:4448];
        layer0[45][31:24] = buffer_data_6[4463:4456];
        layer0[45][39:32] = buffer_data_6[4471:4464];
        layer0[45][47:40] = buffer_data_6[4479:4472];
        layer0[45][55:48] = buffer_data_6[4487:4480];
        layer1[45][7:0] = buffer_data_5[4439:4432];
        layer1[45][15:8] = buffer_data_5[4447:4440];
        layer1[45][23:16] = buffer_data_5[4455:4448];
        layer1[45][31:24] = buffer_data_5[4463:4456];
        layer1[45][39:32] = buffer_data_5[4471:4464];
        layer1[45][47:40] = buffer_data_5[4479:4472];
        layer1[45][55:48] = buffer_data_5[4487:4480];
        layer2[45][7:0] = buffer_data_4[4439:4432];
        layer2[45][15:8] = buffer_data_4[4447:4440];
        layer2[45][23:16] = buffer_data_4[4455:4448];
        layer2[45][31:24] = buffer_data_4[4463:4456];
        layer2[45][39:32] = buffer_data_4[4471:4464];
        layer2[45][47:40] = buffer_data_4[4479:4472];
        layer2[45][55:48] = buffer_data_4[4487:4480];
        layer3[45][7:0] = buffer_data_3[4439:4432];
        layer3[45][15:8] = buffer_data_3[4447:4440];
        layer3[45][23:16] = buffer_data_3[4455:4448];
        layer3[45][31:24] = buffer_data_3[4463:4456];
        layer3[45][39:32] = buffer_data_3[4471:4464];
        layer3[45][47:40] = buffer_data_3[4479:4472];
        layer3[45][55:48] = buffer_data_3[4487:4480];
        layer4[45][7:0] = buffer_data_2[4439:4432];
        layer4[45][15:8] = buffer_data_2[4447:4440];
        layer4[45][23:16] = buffer_data_2[4455:4448];
        layer4[45][31:24] = buffer_data_2[4463:4456];
        layer4[45][39:32] = buffer_data_2[4471:4464];
        layer4[45][47:40] = buffer_data_2[4479:4472];
        layer4[45][55:48] = buffer_data_2[4487:4480];
        layer5[45][7:0] = buffer_data_1[4439:4432];
        layer5[45][15:8] = buffer_data_1[4447:4440];
        layer5[45][23:16] = buffer_data_1[4455:4448];
        layer5[45][31:24] = buffer_data_1[4463:4456];
        layer5[45][39:32] = buffer_data_1[4471:4464];
        layer5[45][47:40] = buffer_data_1[4479:4472];
        layer5[45][55:48] = buffer_data_1[4487:4480];
        layer6[45][7:0] = buffer_data_0[4439:4432];
        layer6[45][15:8] = buffer_data_0[4447:4440];
        layer6[45][23:16] = buffer_data_0[4455:4448];
        layer6[45][31:24] = buffer_data_0[4463:4456];
        layer6[45][39:32] = buffer_data_0[4471:4464];
        layer6[45][47:40] = buffer_data_0[4479:4472];
        layer6[45][55:48] = buffer_data_0[4487:4480];
        layer0[46][7:0] = buffer_data_6[4447:4440];
        layer0[46][15:8] = buffer_data_6[4455:4448];
        layer0[46][23:16] = buffer_data_6[4463:4456];
        layer0[46][31:24] = buffer_data_6[4471:4464];
        layer0[46][39:32] = buffer_data_6[4479:4472];
        layer0[46][47:40] = buffer_data_6[4487:4480];
        layer0[46][55:48] = buffer_data_6[4495:4488];
        layer1[46][7:0] = buffer_data_5[4447:4440];
        layer1[46][15:8] = buffer_data_5[4455:4448];
        layer1[46][23:16] = buffer_data_5[4463:4456];
        layer1[46][31:24] = buffer_data_5[4471:4464];
        layer1[46][39:32] = buffer_data_5[4479:4472];
        layer1[46][47:40] = buffer_data_5[4487:4480];
        layer1[46][55:48] = buffer_data_5[4495:4488];
        layer2[46][7:0] = buffer_data_4[4447:4440];
        layer2[46][15:8] = buffer_data_4[4455:4448];
        layer2[46][23:16] = buffer_data_4[4463:4456];
        layer2[46][31:24] = buffer_data_4[4471:4464];
        layer2[46][39:32] = buffer_data_4[4479:4472];
        layer2[46][47:40] = buffer_data_4[4487:4480];
        layer2[46][55:48] = buffer_data_4[4495:4488];
        layer3[46][7:0] = buffer_data_3[4447:4440];
        layer3[46][15:8] = buffer_data_3[4455:4448];
        layer3[46][23:16] = buffer_data_3[4463:4456];
        layer3[46][31:24] = buffer_data_3[4471:4464];
        layer3[46][39:32] = buffer_data_3[4479:4472];
        layer3[46][47:40] = buffer_data_3[4487:4480];
        layer3[46][55:48] = buffer_data_3[4495:4488];
        layer4[46][7:0] = buffer_data_2[4447:4440];
        layer4[46][15:8] = buffer_data_2[4455:4448];
        layer4[46][23:16] = buffer_data_2[4463:4456];
        layer4[46][31:24] = buffer_data_2[4471:4464];
        layer4[46][39:32] = buffer_data_2[4479:4472];
        layer4[46][47:40] = buffer_data_2[4487:4480];
        layer4[46][55:48] = buffer_data_2[4495:4488];
        layer5[46][7:0] = buffer_data_1[4447:4440];
        layer5[46][15:8] = buffer_data_1[4455:4448];
        layer5[46][23:16] = buffer_data_1[4463:4456];
        layer5[46][31:24] = buffer_data_1[4471:4464];
        layer5[46][39:32] = buffer_data_1[4479:4472];
        layer5[46][47:40] = buffer_data_1[4487:4480];
        layer5[46][55:48] = buffer_data_1[4495:4488];
        layer6[46][7:0] = buffer_data_0[4447:4440];
        layer6[46][15:8] = buffer_data_0[4455:4448];
        layer6[46][23:16] = buffer_data_0[4463:4456];
        layer6[46][31:24] = buffer_data_0[4471:4464];
        layer6[46][39:32] = buffer_data_0[4479:4472];
        layer6[46][47:40] = buffer_data_0[4487:4480];
        layer6[46][55:48] = buffer_data_0[4495:4488];
        layer0[47][7:0] = buffer_data_6[4455:4448];
        layer0[47][15:8] = buffer_data_6[4463:4456];
        layer0[47][23:16] = buffer_data_6[4471:4464];
        layer0[47][31:24] = buffer_data_6[4479:4472];
        layer0[47][39:32] = buffer_data_6[4487:4480];
        layer0[47][47:40] = buffer_data_6[4495:4488];
        layer0[47][55:48] = buffer_data_6[4503:4496];
        layer1[47][7:0] = buffer_data_5[4455:4448];
        layer1[47][15:8] = buffer_data_5[4463:4456];
        layer1[47][23:16] = buffer_data_5[4471:4464];
        layer1[47][31:24] = buffer_data_5[4479:4472];
        layer1[47][39:32] = buffer_data_5[4487:4480];
        layer1[47][47:40] = buffer_data_5[4495:4488];
        layer1[47][55:48] = buffer_data_5[4503:4496];
        layer2[47][7:0] = buffer_data_4[4455:4448];
        layer2[47][15:8] = buffer_data_4[4463:4456];
        layer2[47][23:16] = buffer_data_4[4471:4464];
        layer2[47][31:24] = buffer_data_4[4479:4472];
        layer2[47][39:32] = buffer_data_4[4487:4480];
        layer2[47][47:40] = buffer_data_4[4495:4488];
        layer2[47][55:48] = buffer_data_4[4503:4496];
        layer3[47][7:0] = buffer_data_3[4455:4448];
        layer3[47][15:8] = buffer_data_3[4463:4456];
        layer3[47][23:16] = buffer_data_3[4471:4464];
        layer3[47][31:24] = buffer_data_3[4479:4472];
        layer3[47][39:32] = buffer_data_3[4487:4480];
        layer3[47][47:40] = buffer_data_3[4495:4488];
        layer3[47][55:48] = buffer_data_3[4503:4496];
        layer4[47][7:0] = buffer_data_2[4455:4448];
        layer4[47][15:8] = buffer_data_2[4463:4456];
        layer4[47][23:16] = buffer_data_2[4471:4464];
        layer4[47][31:24] = buffer_data_2[4479:4472];
        layer4[47][39:32] = buffer_data_2[4487:4480];
        layer4[47][47:40] = buffer_data_2[4495:4488];
        layer4[47][55:48] = buffer_data_2[4503:4496];
        layer5[47][7:0] = buffer_data_1[4455:4448];
        layer5[47][15:8] = buffer_data_1[4463:4456];
        layer5[47][23:16] = buffer_data_1[4471:4464];
        layer5[47][31:24] = buffer_data_1[4479:4472];
        layer5[47][39:32] = buffer_data_1[4487:4480];
        layer5[47][47:40] = buffer_data_1[4495:4488];
        layer5[47][55:48] = buffer_data_1[4503:4496];
        layer6[47][7:0] = buffer_data_0[4455:4448];
        layer6[47][15:8] = buffer_data_0[4463:4456];
        layer6[47][23:16] = buffer_data_0[4471:4464];
        layer6[47][31:24] = buffer_data_0[4479:4472];
        layer6[47][39:32] = buffer_data_0[4487:4480];
        layer6[47][47:40] = buffer_data_0[4495:4488];
        layer6[47][55:48] = buffer_data_0[4503:4496];
        layer0[48][7:0] = buffer_data_6[4463:4456];
        layer0[48][15:8] = buffer_data_6[4471:4464];
        layer0[48][23:16] = buffer_data_6[4479:4472];
        layer0[48][31:24] = buffer_data_6[4487:4480];
        layer0[48][39:32] = buffer_data_6[4495:4488];
        layer0[48][47:40] = buffer_data_6[4503:4496];
        layer0[48][55:48] = buffer_data_6[4511:4504];
        layer1[48][7:0] = buffer_data_5[4463:4456];
        layer1[48][15:8] = buffer_data_5[4471:4464];
        layer1[48][23:16] = buffer_data_5[4479:4472];
        layer1[48][31:24] = buffer_data_5[4487:4480];
        layer1[48][39:32] = buffer_data_5[4495:4488];
        layer1[48][47:40] = buffer_data_5[4503:4496];
        layer1[48][55:48] = buffer_data_5[4511:4504];
        layer2[48][7:0] = buffer_data_4[4463:4456];
        layer2[48][15:8] = buffer_data_4[4471:4464];
        layer2[48][23:16] = buffer_data_4[4479:4472];
        layer2[48][31:24] = buffer_data_4[4487:4480];
        layer2[48][39:32] = buffer_data_4[4495:4488];
        layer2[48][47:40] = buffer_data_4[4503:4496];
        layer2[48][55:48] = buffer_data_4[4511:4504];
        layer3[48][7:0] = buffer_data_3[4463:4456];
        layer3[48][15:8] = buffer_data_3[4471:4464];
        layer3[48][23:16] = buffer_data_3[4479:4472];
        layer3[48][31:24] = buffer_data_3[4487:4480];
        layer3[48][39:32] = buffer_data_3[4495:4488];
        layer3[48][47:40] = buffer_data_3[4503:4496];
        layer3[48][55:48] = buffer_data_3[4511:4504];
        layer4[48][7:0] = buffer_data_2[4463:4456];
        layer4[48][15:8] = buffer_data_2[4471:4464];
        layer4[48][23:16] = buffer_data_2[4479:4472];
        layer4[48][31:24] = buffer_data_2[4487:4480];
        layer4[48][39:32] = buffer_data_2[4495:4488];
        layer4[48][47:40] = buffer_data_2[4503:4496];
        layer4[48][55:48] = buffer_data_2[4511:4504];
        layer5[48][7:0] = buffer_data_1[4463:4456];
        layer5[48][15:8] = buffer_data_1[4471:4464];
        layer5[48][23:16] = buffer_data_1[4479:4472];
        layer5[48][31:24] = buffer_data_1[4487:4480];
        layer5[48][39:32] = buffer_data_1[4495:4488];
        layer5[48][47:40] = buffer_data_1[4503:4496];
        layer5[48][55:48] = buffer_data_1[4511:4504];
        layer6[48][7:0] = buffer_data_0[4463:4456];
        layer6[48][15:8] = buffer_data_0[4471:4464];
        layer6[48][23:16] = buffer_data_0[4479:4472];
        layer6[48][31:24] = buffer_data_0[4487:4480];
        layer6[48][39:32] = buffer_data_0[4495:4488];
        layer6[48][47:40] = buffer_data_0[4503:4496];
        layer6[48][55:48] = buffer_data_0[4511:4504];
        layer0[49][7:0] = buffer_data_6[4471:4464];
        layer0[49][15:8] = buffer_data_6[4479:4472];
        layer0[49][23:16] = buffer_data_6[4487:4480];
        layer0[49][31:24] = buffer_data_6[4495:4488];
        layer0[49][39:32] = buffer_data_6[4503:4496];
        layer0[49][47:40] = buffer_data_6[4511:4504];
        layer0[49][55:48] = buffer_data_6[4519:4512];
        layer1[49][7:0] = buffer_data_5[4471:4464];
        layer1[49][15:8] = buffer_data_5[4479:4472];
        layer1[49][23:16] = buffer_data_5[4487:4480];
        layer1[49][31:24] = buffer_data_5[4495:4488];
        layer1[49][39:32] = buffer_data_5[4503:4496];
        layer1[49][47:40] = buffer_data_5[4511:4504];
        layer1[49][55:48] = buffer_data_5[4519:4512];
        layer2[49][7:0] = buffer_data_4[4471:4464];
        layer2[49][15:8] = buffer_data_4[4479:4472];
        layer2[49][23:16] = buffer_data_4[4487:4480];
        layer2[49][31:24] = buffer_data_4[4495:4488];
        layer2[49][39:32] = buffer_data_4[4503:4496];
        layer2[49][47:40] = buffer_data_4[4511:4504];
        layer2[49][55:48] = buffer_data_4[4519:4512];
        layer3[49][7:0] = buffer_data_3[4471:4464];
        layer3[49][15:8] = buffer_data_3[4479:4472];
        layer3[49][23:16] = buffer_data_3[4487:4480];
        layer3[49][31:24] = buffer_data_3[4495:4488];
        layer3[49][39:32] = buffer_data_3[4503:4496];
        layer3[49][47:40] = buffer_data_3[4511:4504];
        layer3[49][55:48] = buffer_data_3[4519:4512];
        layer4[49][7:0] = buffer_data_2[4471:4464];
        layer4[49][15:8] = buffer_data_2[4479:4472];
        layer4[49][23:16] = buffer_data_2[4487:4480];
        layer4[49][31:24] = buffer_data_2[4495:4488];
        layer4[49][39:32] = buffer_data_2[4503:4496];
        layer4[49][47:40] = buffer_data_2[4511:4504];
        layer4[49][55:48] = buffer_data_2[4519:4512];
        layer5[49][7:0] = buffer_data_1[4471:4464];
        layer5[49][15:8] = buffer_data_1[4479:4472];
        layer5[49][23:16] = buffer_data_1[4487:4480];
        layer5[49][31:24] = buffer_data_1[4495:4488];
        layer5[49][39:32] = buffer_data_1[4503:4496];
        layer5[49][47:40] = buffer_data_1[4511:4504];
        layer5[49][55:48] = buffer_data_1[4519:4512];
        layer6[49][7:0] = buffer_data_0[4471:4464];
        layer6[49][15:8] = buffer_data_0[4479:4472];
        layer6[49][23:16] = buffer_data_0[4487:4480];
        layer6[49][31:24] = buffer_data_0[4495:4488];
        layer6[49][39:32] = buffer_data_0[4503:4496];
        layer6[49][47:40] = buffer_data_0[4511:4504];
        layer6[49][55:48] = buffer_data_0[4519:4512];
        layer0[50][7:0] = buffer_data_6[4479:4472];
        layer0[50][15:8] = buffer_data_6[4487:4480];
        layer0[50][23:16] = buffer_data_6[4495:4488];
        layer0[50][31:24] = buffer_data_6[4503:4496];
        layer0[50][39:32] = buffer_data_6[4511:4504];
        layer0[50][47:40] = buffer_data_6[4519:4512];
        layer0[50][55:48] = buffer_data_6[4527:4520];
        layer1[50][7:0] = buffer_data_5[4479:4472];
        layer1[50][15:8] = buffer_data_5[4487:4480];
        layer1[50][23:16] = buffer_data_5[4495:4488];
        layer1[50][31:24] = buffer_data_5[4503:4496];
        layer1[50][39:32] = buffer_data_5[4511:4504];
        layer1[50][47:40] = buffer_data_5[4519:4512];
        layer1[50][55:48] = buffer_data_5[4527:4520];
        layer2[50][7:0] = buffer_data_4[4479:4472];
        layer2[50][15:8] = buffer_data_4[4487:4480];
        layer2[50][23:16] = buffer_data_4[4495:4488];
        layer2[50][31:24] = buffer_data_4[4503:4496];
        layer2[50][39:32] = buffer_data_4[4511:4504];
        layer2[50][47:40] = buffer_data_4[4519:4512];
        layer2[50][55:48] = buffer_data_4[4527:4520];
        layer3[50][7:0] = buffer_data_3[4479:4472];
        layer3[50][15:8] = buffer_data_3[4487:4480];
        layer3[50][23:16] = buffer_data_3[4495:4488];
        layer3[50][31:24] = buffer_data_3[4503:4496];
        layer3[50][39:32] = buffer_data_3[4511:4504];
        layer3[50][47:40] = buffer_data_3[4519:4512];
        layer3[50][55:48] = buffer_data_3[4527:4520];
        layer4[50][7:0] = buffer_data_2[4479:4472];
        layer4[50][15:8] = buffer_data_2[4487:4480];
        layer4[50][23:16] = buffer_data_2[4495:4488];
        layer4[50][31:24] = buffer_data_2[4503:4496];
        layer4[50][39:32] = buffer_data_2[4511:4504];
        layer4[50][47:40] = buffer_data_2[4519:4512];
        layer4[50][55:48] = buffer_data_2[4527:4520];
        layer5[50][7:0] = buffer_data_1[4479:4472];
        layer5[50][15:8] = buffer_data_1[4487:4480];
        layer5[50][23:16] = buffer_data_1[4495:4488];
        layer5[50][31:24] = buffer_data_1[4503:4496];
        layer5[50][39:32] = buffer_data_1[4511:4504];
        layer5[50][47:40] = buffer_data_1[4519:4512];
        layer5[50][55:48] = buffer_data_1[4527:4520];
        layer6[50][7:0] = buffer_data_0[4479:4472];
        layer6[50][15:8] = buffer_data_0[4487:4480];
        layer6[50][23:16] = buffer_data_0[4495:4488];
        layer6[50][31:24] = buffer_data_0[4503:4496];
        layer6[50][39:32] = buffer_data_0[4511:4504];
        layer6[50][47:40] = buffer_data_0[4519:4512];
        layer6[50][55:48] = buffer_data_0[4527:4520];
        layer0[51][7:0] = buffer_data_6[4487:4480];
        layer0[51][15:8] = buffer_data_6[4495:4488];
        layer0[51][23:16] = buffer_data_6[4503:4496];
        layer0[51][31:24] = buffer_data_6[4511:4504];
        layer0[51][39:32] = buffer_data_6[4519:4512];
        layer0[51][47:40] = buffer_data_6[4527:4520];
        layer0[51][55:48] = buffer_data_6[4535:4528];
        layer1[51][7:0] = buffer_data_5[4487:4480];
        layer1[51][15:8] = buffer_data_5[4495:4488];
        layer1[51][23:16] = buffer_data_5[4503:4496];
        layer1[51][31:24] = buffer_data_5[4511:4504];
        layer1[51][39:32] = buffer_data_5[4519:4512];
        layer1[51][47:40] = buffer_data_5[4527:4520];
        layer1[51][55:48] = buffer_data_5[4535:4528];
        layer2[51][7:0] = buffer_data_4[4487:4480];
        layer2[51][15:8] = buffer_data_4[4495:4488];
        layer2[51][23:16] = buffer_data_4[4503:4496];
        layer2[51][31:24] = buffer_data_4[4511:4504];
        layer2[51][39:32] = buffer_data_4[4519:4512];
        layer2[51][47:40] = buffer_data_4[4527:4520];
        layer2[51][55:48] = buffer_data_4[4535:4528];
        layer3[51][7:0] = buffer_data_3[4487:4480];
        layer3[51][15:8] = buffer_data_3[4495:4488];
        layer3[51][23:16] = buffer_data_3[4503:4496];
        layer3[51][31:24] = buffer_data_3[4511:4504];
        layer3[51][39:32] = buffer_data_3[4519:4512];
        layer3[51][47:40] = buffer_data_3[4527:4520];
        layer3[51][55:48] = buffer_data_3[4535:4528];
        layer4[51][7:0] = buffer_data_2[4487:4480];
        layer4[51][15:8] = buffer_data_2[4495:4488];
        layer4[51][23:16] = buffer_data_2[4503:4496];
        layer4[51][31:24] = buffer_data_2[4511:4504];
        layer4[51][39:32] = buffer_data_2[4519:4512];
        layer4[51][47:40] = buffer_data_2[4527:4520];
        layer4[51][55:48] = buffer_data_2[4535:4528];
        layer5[51][7:0] = buffer_data_1[4487:4480];
        layer5[51][15:8] = buffer_data_1[4495:4488];
        layer5[51][23:16] = buffer_data_1[4503:4496];
        layer5[51][31:24] = buffer_data_1[4511:4504];
        layer5[51][39:32] = buffer_data_1[4519:4512];
        layer5[51][47:40] = buffer_data_1[4527:4520];
        layer5[51][55:48] = buffer_data_1[4535:4528];
        layer6[51][7:0] = buffer_data_0[4487:4480];
        layer6[51][15:8] = buffer_data_0[4495:4488];
        layer6[51][23:16] = buffer_data_0[4503:4496];
        layer6[51][31:24] = buffer_data_0[4511:4504];
        layer6[51][39:32] = buffer_data_0[4519:4512];
        layer6[51][47:40] = buffer_data_0[4527:4520];
        layer6[51][55:48] = buffer_data_0[4535:4528];
        layer0[52][7:0] = buffer_data_6[4495:4488];
        layer0[52][15:8] = buffer_data_6[4503:4496];
        layer0[52][23:16] = buffer_data_6[4511:4504];
        layer0[52][31:24] = buffer_data_6[4519:4512];
        layer0[52][39:32] = buffer_data_6[4527:4520];
        layer0[52][47:40] = buffer_data_6[4535:4528];
        layer0[52][55:48] = buffer_data_6[4543:4536];
        layer1[52][7:0] = buffer_data_5[4495:4488];
        layer1[52][15:8] = buffer_data_5[4503:4496];
        layer1[52][23:16] = buffer_data_5[4511:4504];
        layer1[52][31:24] = buffer_data_5[4519:4512];
        layer1[52][39:32] = buffer_data_5[4527:4520];
        layer1[52][47:40] = buffer_data_5[4535:4528];
        layer1[52][55:48] = buffer_data_5[4543:4536];
        layer2[52][7:0] = buffer_data_4[4495:4488];
        layer2[52][15:8] = buffer_data_4[4503:4496];
        layer2[52][23:16] = buffer_data_4[4511:4504];
        layer2[52][31:24] = buffer_data_4[4519:4512];
        layer2[52][39:32] = buffer_data_4[4527:4520];
        layer2[52][47:40] = buffer_data_4[4535:4528];
        layer2[52][55:48] = buffer_data_4[4543:4536];
        layer3[52][7:0] = buffer_data_3[4495:4488];
        layer3[52][15:8] = buffer_data_3[4503:4496];
        layer3[52][23:16] = buffer_data_3[4511:4504];
        layer3[52][31:24] = buffer_data_3[4519:4512];
        layer3[52][39:32] = buffer_data_3[4527:4520];
        layer3[52][47:40] = buffer_data_3[4535:4528];
        layer3[52][55:48] = buffer_data_3[4543:4536];
        layer4[52][7:0] = buffer_data_2[4495:4488];
        layer4[52][15:8] = buffer_data_2[4503:4496];
        layer4[52][23:16] = buffer_data_2[4511:4504];
        layer4[52][31:24] = buffer_data_2[4519:4512];
        layer4[52][39:32] = buffer_data_2[4527:4520];
        layer4[52][47:40] = buffer_data_2[4535:4528];
        layer4[52][55:48] = buffer_data_2[4543:4536];
        layer5[52][7:0] = buffer_data_1[4495:4488];
        layer5[52][15:8] = buffer_data_1[4503:4496];
        layer5[52][23:16] = buffer_data_1[4511:4504];
        layer5[52][31:24] = buffer_data_1[4519:4512];
        layer5[52][39:32] = buffer_data_1[4527:4520];
        layer5[52][47:40] = buffer_data_1[4535:4528];
        layer5[52][55:48] = buffer_data_1[4543:4536];
        layer6[52][7:0] = buffer_data_0[4495:4488];
        layer6[52][15:8] = buffer_data_0[4503:4496];
        layer6[52][23:16] = buffer_data_0[4511:4504];
        layer6[52][31:24] = buffer_data_0[4519:4512];
        layer6[52][39:32] = buffer_data_0[4527:4520];
        layer6[52][47:40] = buffer_data_0[4535:4528];
        layer6[52][55:48] = buffer_data_0[4543:4536];
        layer0[53][7:0] = buffer_data_6[4503:4496];
        layer0[53][15:8] = buffer_data_6[4511:4504];
        layer0[53][23:16] = buffer_data_6[4519:4512];
        layer0[53][31:24] = buffer_data_6[4527:4520];
        layer0[53][39:32] = buffer_data_6[4535:4528];
        layer0[53][47:40] = buffer_data_6[4543:4536];
        layer0[53][55:48] = buffer_data_6[4551:4544];
        layer1[53][7:0] = buffer_data_5[4503:4496];
        layer1[53][15:8] = buffer_data_5[4511:4504];
        layer1[53][23:16] = buffer_data_5[4519:4512];
        layer1[53][31:24] = buffer_data_5[4527:4520];
        layer1[53][39:32] = buffer_data_5[4535:4528];
        layer1[53][47:40] = buffer_data_5[4543:4536];
        layer1[53][55:48] = buffer_data_5[4551:4544];
        layer2[53][7:0] = buffer_data_4[4503:4496];
        layer2[53][15:8] = buffer_data_4[4511:4504];
        layer2[53][23:16] = buffer_data_4[4519:4512];
        layer2[53][31:24] = buffer_data_4[4527:4520];
        layer2[53][39:32] = buffer_data_4[4535:4528];
        layer2[53][47:40] = buffer_data_4[4543:4536];
        layer2[53][55:48] = buffer_data_4[4551:4544];
        layer3[53][7:0] = buffer_data_3[4503:4496];
        layer3[53][15:8] = buffer_data_3[4511:4504];
        layer3[53][23:16] = buffer_data_3[4519:4512];
        layer3[53][31:24] = buffer_data_3[4527:4520];
        layer3[53][39:32] = buffer_data_3[4535:4528];
        layer3[53][47:40] = buffer_data_3[4543:4536];
        layer3[53][55:48] = buffer_data_3[4551:4544];
        layer4[53][7:0] = buffer_data_2[4503:4496];
        layer4[53][15:8] = buffer_data_2[4511:4504];
        layer4[53][23:16] = buffer_data_2[4519:4512];
        layer4[53][31:24] = buffer_data_2[4527:4520];
        layer4[53][39:32] = buffer_data_2[4535:4528];
        layer4[53][47:40] = buffer_data_2[4543:4536];
        layer4[53][55:48] = buffer_data_2[4551:4544];
        layer5[53][7:0] = buffer_data_1[4503:4496];
        layer5[53][15:8] = buffer_data_1[4511:4504];
        layer5[53][23:16] = buffer_data_1[4519:4512];
        layer5[53][31:24] = buffer_data_1[4527:4520];
        layer5[53][39:32] = buffer_data_1[4535:4528];
        layer5[53][47:40] = buffer_data_1[4543:4536];
        layer5[53][55:48] = buffer_data_1[4551:4544];
        layer6[53][7:0] = buffer_data_0[4503:4496];
        layer6[53][15:8] = buffer_data_0[4511:4504];
        layer6[53][23:16] = buffer_data_0[4519:4512];
        layer6[53][31:24] = buffer_data_0[4527:4520];
        layer6[53][39:32] = buffer_data_0[4535:4528];
        layer6[53][47:40] = buffer_data_0[4543:4536];
        layer6[53][55:48] = buffer_data_0[4551:4544];
        layer0[54][7:0] = buffer_data_6[4511:4504];
        layer0[54][15:8] = buffer_data_6[4519:4512];
        layer0[54][23:16] = buffer_data_6[4527:4520];
        layer0[54][31:24] = buffer_data_6[4535:4528];
        layer0[54][39:32] = buffer_data_6[4543:4536];
        layer0[54][47:40] = buffer_data_6[4551:4544];
        layer0[54][55:48] = buffer_data_6[4559:4552];
        layer1[54][7:0] = buffer_data_5[4511:4504];
        layer1[54][15:8] = buffer_data_5[4519:4512];
        layer1[54][23:16] = buffer_data_5[4527:4520];
        layer1[54][31:24] = buffer_data_5[4535:4528];
        layer1[54][39:32] = buffer_data_5[4543:4536];
        layer1[54][47:40] = buffer_data_5[4551:4544];
        layer1[54][55:48] = buffer_data_5[4559:4552];
        layer2[54][7:0] = buffer_data_4[4511:4504];
        layer2[54][15:8] = buffer_data_4[4519:4512];
        layer2[54][23:16] = buffer_data_4[4527:4520];
        layer2[54][31:24] = buffer_data_4[4535:4528];
        layer2[54][39:32] = buffer_data_4[4543:4536];
        layer2[54][47:40] = buffer_data_4[4551:4544];
        layer2[54][55:48] = buffer_data_4[4559:4552];
        layer3[54][7:0] = buffer_data_3[4511:4504];
        layer3[54][15:8] = buffer_data_3[4519:4512];
        layer3[54][23:16] = buffer_data_3[4527:4520];
        layer3[54][31:24] = buffer_data_3[4535:4528];
        layer3[54][39:32] = buffer_data_3[4543:4536];
        layer3[54][47:40] = buffer_data_3[4551:4544];
        layer3[54][55:48] = buffer_data_3[4559:4552];
        layer4[54][7:0] = buffer_data_2[4511:4504];
        layer4[54][15:8] = buffer_data_2[4519:4512];
        layer4[54][23:16] = buffer_data_2[4527:4520];
        layer4[54][31:24] = buffer_data_2[4535:4528];
        layer4[54][39:32] = buffer_data_2[4543:4536];
        layer4[54][47:40] = buffer_data_2[4551:4544];
        layer4[54][55:48] = buffer_data_2[4559:4552];
        layer5[54][7:0] = buffer_data_1[4511:4504];
        layer5[54][15:8] = buffer_data_1[4519:4512];
        layer5[54][23:16] = buffer_data_1[4527:4520];
        layer5[54][31:24] = buffer_data_1[4535:4528];
        layer5[54][39:32] = buffer_data_1[4543:4536];
        layer5[54][47:40] = buffer_data_1[4551:4544];
        layer5[54][55:48] = buffer_data_1[4559:4552];
        layer6[54][7:0] = buffer_data_0[4511:4504];
        layer6[54][15:8] = buffer_data_0[4519:4512];
        layer6[54][23:16] = buffer_data_0[4527:4520];
        layer6[54][31:24] = buffer_data_0[4535:4528];
        layer6[54][39:32] = buffer_data_0[4543:4536];
        layer6[54][47:40] = buffer_data_0[4551:4544];
        layer6[54][55:48] = buffer_data_0[4559:4552];
        layer0[55][7:0] = buffer_data_6[4519:4512];
        layer0[55][15:8] = buffer_data_6[4527:4520];
        layer0[55][23:16] = buffer_data_6[4535:4528];
        layer0[55][31:24] = buffer_data_6[4543:4536];
        layer0[55][39:32] = buffer_data_6[4551:4544];
        layer0[55][47:40] = buffer_data_6[4559:4552];
        layer0[55][55:48] = buffer_data_6[4567:4560];
        layer1[55][7:0] = buffer_data_5[4519:4512];
        layer1[55][15:8] = buffer_data_5[4527:4520];
        layer1[55][23:16] = buffer_data_5[4535:4528];
        layer1[55][31:24] = buffer_data_5[4543:4536];
        layer1[55][39:32] = buffer_data_5[4551:4544];
        layer1[55][47:40] = buffer_data_5[4559:4552];
        layer1[55][55:48] = buffer_data_5[4567:4560];
        layer2[55][7:0] = buffer_data_4[4519:4512];
        layer2[55][15:8] = buffer_data_4[4527:4520];
        layer2[55][23:16] = buffer_data_4[4535:4528];
        layer2[55][31:24] = buffer_data_4[4543:4536];
        layer2[55][39:32] = buffer_data_4[4551:4544];
        layer2[55][47:40] = buffer_data_4[4559:4552];
        layer2[55][55:48] = buffer_data_4[4567:4560];
        layer3[55][7:0] = buffer_data_3[4519:4512];
        layer3[55][15:8] = buffer_data_3[4527:4520];
        layer3[55][23:16] = buffer_data_3[4535:4528];
        layer3[55][31:24] = buffer_data_3[4543:4536];
        layer3[55][39:32] = buffer_data_3[4551:4544];
        layer3[55][47:40] = buffer_data_3[4559:4552];
        layer3[55][55:48] = buffer_data_3[4567:4560];
        layer4[55][7:0] = buffer_data_2[4519:4512];
        layer4[55][15:8] = buffer_data_2[4527:4520];
        layer4[55][23:16] = buffer_data_2[4535:4528];
        layer4[55][31:24] = buffer_data_2[4543:4536];
        layer4[55][39:32] = buffer_data_2[4551:4544];
        layer4[55][47:40] = buffer_data_2[4559:4552];
        layer4[55][55:48] = buffer_data_2[4567:4560];
        layer5[55][7:0] = buffer_data_1[4519:4512];
        layer5[55][15:8] = buffer_data_1[4527:4520];
        layer5[55][23:16] = buffer_data_1[4535:4528];
        layer5[55][31:24] = buffer_data_1[4543:4536];
        layer5[55][39:32] = buffer_data_1[4551:4544];
        layer5[55][47:40] = buffer_data_1[4559:4552];
        layer5[55][55:48] = buffer_data_1[4567:4560];
        layer6[55][7:0] = buffer_data_0[4519:4512];
        layer6[55][15:8] = buffer_data_0[4527:4520];
        layer6[55][23:16] = buffer_data_0[4535:4528];
        layer6[55][31:24] = buffer_data_0[4543:4536];
        layer6[55][39:32] = buffer_data_0[4551:4544];
        layer6[55][47:40] = buffer_data_0[4559:4552];
        layer6[55][55:48] = buffer_data_0[4567:4560];
        layer0[56][7:0] = buffer_data_6[4527:4520];
        layer0[56][15:8] = buffer_data_6[4535:4528];
        layer0[56][23:16] = buffer_data_6[4543:4536];
        layer0[56][31:24] = buffer_data_6[4551:4544];
        layer0[56][39:32] = buffer_data_6[4559:4552];
        layer0[56][47:40] = buffer_data_6[4567:4560];
        layer0[56][55:48] = buffer_data_6[4575:4568];
        layer1[56][7:0] = buffer_data_5[4527:4520];
        layer1[56][15:8] = buffer_data_5[4535:4528];
        layer1[56][23:16] = buffer_data_5[4543:4536];
        layer1[56][31:24] = buffer_data_5[4551:4544];
        layer1[56][39:32] = buffer_data_5[4559:4552];
        layer1[56][47:40] = buffer_data_5[4567:4560];
        layer1[56][55:48] = buffer_data_5[4575:4568];
        layer2[56][7:0] = buffer_data_4[4527:4520];
        layer2[56][15:8] = buffer_data_4[4535:4528];
        layer2[56][23:16] = buffer_data_4[4543:4536];
        layer2[56][31:24] = buffer_data_4[4551:4544];
        layer2[56][39:32] = buffer_data_4[4559:4552];
        layer2[56][47:40] = buffer_data_4[4567:4560];
        layer2[56][55:48] = buffer_data_4[4575:4568];
        layer3[56][7:0] = buffer_data_3[4527:4520];
        layer3[56][15:8] = buffer_data_3[4535:4528];
        layer3[56][23:16] = buffer_data_3[4543:4536];
        layer3[56][31:24] = buffer_data_3[4551:4544];
        layer3[56][39:32] = buffer_data_3[4559:4552];
        layer3[56][47:40] = buffer_data_3[4567:4560];
        layer3[56][55:48] = buffer_data_3[4575:4568];
        layer4[56][7:0] = buffer_data_2[4527:4520];
        layer4[56][15:8] = buffer_data_2[4535:4528];
        layer4[56][23:16] = buffer_data_2[4543:4536];
        layer4[56][31:24] = buffer_data_2[4551:4544];
        layer4[56][39:32] = buffer_data_2[4559:4552];
        layer4[56][47:40] = buffer_data_2[4567:4560];
        layer4[56][55:48] = buffer_data_2[4575:4568];
        layer5[56][7:0] = buffer_data_1[4527:4520];
        layer5[56][15:8] = buffer_data_1[4535:4528];
        layer5[56][23:16] = buffer_data_1[4543:4536];
        layer5[56][31:24] = buffer_data_1[4551:4544];
        layer5[56][39:32] = buffer_data_1[4559:4552];
        layer5[56][47:40] = buffer_data_1[4567:4560];
        layer5[56][55:48] = buffer_data_1[4575:4568];
        layer6[56][7:0] = buffer_data_0[4527:4520];
        layer6[56][15:8] = buffer_data_0[4535:4528];
        layer6[56][23:16] = buffer_data_0[4543:4536];
        layer6[56][31:24] = buffer_data_0[4551:4544];
        layer6[56][39:32] = buffer_data_0[4559:4552];
        layer6[56][47:40] = buffer_data_0[4567:4560];
        layer6[56][55:48] = buffer_data_0[4575:4568];
        layer0[57][7:0] = buffer_data_6[4535:4528];
        layer0[57][15:8] = buffer_data_6[4543:4536];
        layer0[57][23:16] = buffer_data_6[4551:4544];
        layer0[57][31:24] = buffer_data_6[4559:4552];
        layer0[57][39:32] = buffer_data_6[4567:4560];
        layer0[57][47:40] = buffer_data_6[4575:4568];
        layer0[57][55:48] = buffer_data_6[4583:4576];
        layer1[57][7:0] = buffer_data_5[4535:4528];
        layer1[57][15:8] = buffer_data_5[4543:4536];
        layer1[57][23:16] = buffer_data_5[4551:4544];
        layer1[57][31:24] = buffer_data_5[4559:4552];
        layer1[57][39:32] = buffer_data_5[4567:4560];
        layer1[57][47:40] = buffer_data_5[4575:4568];
        layer1[57][55:48] = buffer_data_5[4583:4576];
        layer2[57][7:0] = buffer_data_4[4535:4528];
        layer2[57][15:8] = buffer_data_4[4543:4536];
        layer2[57][23:16] = buffer_data_4[4551:4544];
        layer2[57][31:24] = buffer_data_4[4559:4552];
        layer2[57][39:32] = buffer_data_4[4567:4560];
        layer2[57][47:40] = buffer_data_4[4575:4568];
        layer2[57][55:48] = buffer_data_4[4583:4576];
        layer3[57][7:0] = buffer_data_3[4535:4528];
        layer3[57][15:8] = buffer_data_3[4543:4536];
        layer3[57][23:16] = buffer_data_3[4551:4544];
        layer3[57][31:24] = buffer_data_3[4559:4552];
        layer3[57][39:32] = buffer_data_3[4567:4560];
        layer3[57][47:40] = buffer_data_3[4575:4568];
        layer3[57][55:48] = buffer_data_3[4583:4576];
        layer4[57][7:0] = buffer_data_2[4535:4528];
        layer4[57][15:8] = buffer_data_2[4543:4536];
        layer4[57][23:16] = buffer_data_2[4551:4544];
        layer4[57][31:24] = buffer_data_2[4559:4552];
        layer4[57][39:32] = buffer_data_2[4567:4560];
        layer4[57][47:40] = buffer_data_2[4575:4568];
        layer4[57][55:48] = buffer_data_2[4583:4576];
        layer5[57][7:0] = buffer_data_1[4535:4528];
        layer5[57][15:8] = buffer_data_1[4543:4536];
        layer5[57][23:16] = buffer_data_1[4551:4544];
        layer5[57][31:24] = buffer_data_1[4559:4552];
        layer5[57][39:32] = buffer_data_1[4567:4560];
        layer5[57][47:40] = buffer_data_1[4575:4568];
        layer5[57][55:48] = buffer_data_1[4583:4576];
        layer6[57][7:0] = buffer_data_0[4535:4528];
        layer6[57][15:8] = buffer_data_0[4543:4536];
        layer6[57][23:16] = buffer_data_0[4551:4544];
        layer6[57][31:24] = buffer_data_0[4559:4552];
        layer6[57][39:32] = buffer_data_0[4567:4560];
        layer6[57][47:40] = buffer_data_0[4575:4568];
        layer6[57][55:48] = buffer_data_0[4583:4576];
        layer0[58][7:0] = buffer_data_6[4543:4536];
        layer0[58][15:8] = buffer_data_6[4551:4544];
        layer0[58][23:16] = buffer_data_6[4559:4552];
        layer0[58][31:24] = buffer_data_6[4567:4560];
        layer0[58][39:32] = buffer_data_6[4575:4568];
        layer0[58][47:40] = buffer_data_6[4583:4576];
        layer0[58][55:48] = buffer_data_6[4591:4584];
        layer1[58][7:0] = buffer_data_5[4543:4536];
        layer1[58][15:8] = buffer_data_5[4551:4544];
        layer1[58][23:16] = buffer_data_5[4559:4552];
        layer1[58][31:24] = buffer_data_5[4567:4560];
        layer1[58][39:32] = buffer_data_5[4575:4568];
        layer1[58][47:40] = buffer_data_5[4583:4576];
        layer1[58][55:48] = buffer_data_5[4591:4584];
        layer2[58][7:0] = buffer_data_4[4543:4536];
        layer2[58][15:8] = buffer_data_4[4551:4544];
        layer2[58][23:16] = buffer_data_4[4559:4552];
        layer2[58][31:24] = buffer_data_4[4567:4560];
        layer2[58][39:32] = buffer_data_4[4575:4568];
        layer2[58][47:40] = buffer_data_4[4583:4576];
        layer2[58][55:48] = buffer_data_4[4591:4584];
        layer3[58][7:0] = buffer_data_3[4543:4536];
        layer3[58][15:8] = buffer_data_3[4551:4544];
        layer3[58][23:16] = buffer_data_3[4559:4552];
        layer3[58][31:24] = buffer_data_3[4567:4560];
        layer3[58][39:32] = buffer_data_3[4575:4568];
        layer3[58][47:40] = buffer_data_3[4583:4576];
        layer3[58][55:48] = buffer_data_3[4591:4584];
        layer4[58][7:0] = buffer_data_2[4543:4536];
        layer4[58][15:8] = buffer_data_2[4551:4544];
        layer4[58][23:16] = buffer_data_2[4559:4552];
        layer4[58][31:24] = buffer_data_2[4567:4560];
        layer4[58][39:32] = buffer_data_2[4575:4568];
        layer4[58][47:40] = buffer_data_2[4583:4576];
        layer4[58][55:48] = buffer_data_2[4591:4584];
        layer5[58][7:0] = buffer_data_1[4543:4536];
        layer5[58][15:8] = buffer_data_1[4551:4544];
        layer5[58][23:16] = buffer_data_1[4559:4552];
        layer5[58][31:24] = buffer_data_1[4567:4560];
        layer5[58][39:32] = buffer_data_1[4575:4568];
        layer5[58][47:40] = buffer_data_1[4583:4576];
        layer5[58][55:48] = buffer_data_1[4591:4584];
        layer6[58][7:0] = buffer_data_0[4543:4536];
        layer6[58][15:8] = buffer_data_0[4551:4544];
        layer6[58][23:16] = buffer_data_0[4559:4552];
        layer6[58][31:24] = buffer_data_0[4567:4560];
        layer6[58][39:32] = buffer_data_0[4575:4568];
        layer6[58][47:40] = buffer_data_0[4583:4576];
        layer6[58][55:48] = buffer_data_0[4591:4584];
        layer0[59][7:0] = buffer_data_6[4551:4544];
        layer0[59][15:8] = buffer_data_6[4559:4552];
        layer0[59][23:16] = buffer_data_6[4567:4560];
        layer0[59][31:24] = buffer_data_6[4575:4568];
        layer0[59][39:32] = buffer_data_6[4583:4576];
        layer0[59][47:40] = buffer_data_6[4591:4584];
        layer0[59][55:48] = buffer_data_6[4599:4592];
        layer1[59][7:0] = buffer_data_5[4551:4544];
        layer1[59][15:8] = buffer_data_5[4559:4552];
        layer1[59][23:16] = buffer_data_5[4567:4560];
        layer1[59][31:24] = buffer_data_5[4575:4568];
        layer1[59][39:32] = buffer_data_5[4583:4576];
        layer1[59][47:40] = buffer_data_5[4591:4584];
        layer1[59][55:48] = buffer_data_5[4599:4592];
        layer2[59][7:0] = buffer_data_4[4551:4544];
        layer2[59][15:8] = buffer_data_4[4559:4552];
        layer2[59][23:16] = buffer_data_4[4567:4560];
        layer2[59][31:24] = buffer_data_4[4575:4568];
        layer2[59][39:32] = buffer_data_4[4583:4576];
        layer2[59][47:40] = buffer_data_4[4591:4584];
        layer2[59][55:48] = buffer_data_4[4599:4592];
        layer3[59][7:0] = buffer_data_3[4551:4544];
        layer3[59][15:8] = buffer_data_3[4559:4552];
        layer3[59][23:16] = buffer_data_3[4567:4560];
        layer3[59][31:24] = buffer_data_3[4575:4568];
        layer3[59][39:32] = buffer_data_3[4583:4576];
        layer3[59][47:40] = buffer_data_3[4591:4584];
        layer3[59][55:48] = buffer_data_3[4599:4592];
        layer4[59][7:0] = buffer_data_2[4551:4544];
        layer4[59][15:8] = buffer_data_2[4559:4552];
        layer4[59][23:16] = buffer_data_2[4567:4560];
        layer4[59][31:24] = buffer_data_2[4575:4568];
        layer4[59][39:32] = buffer_data_2[4583:4576];
        layer4[59][47:40] = buffer_data_2[4591:4584];
        layer4[59][55:48] = buffer_data_2[4599:4592];
        layer5[59][7:0] = buffer_data_1[4551:4544];
        layer5[59][15:8] = buffer_data_1[4559:4552];
        layer5[59][23:16] = buffer_data_1[4567:4560];
        layer5[59][31:24] = buffer_data_1[4575:4568];
        layer5[59][39:32] = buffer_data_1[4583:4576];
        layer5[59][47:40] = buffer_data_1[4591:4584];
        layer5[59][55:48] = buffer_data_1[4599:4592];
        layer6[59][7:0] = buffer_data_0[4551:4544];
        layer6[59][15:8] = buffer_data_0[4559:4552];
        layer6[59][23:16] = buffer_data_0[4567:4560];
        layer6[59][31:24] = buffer_data_0[4575:4568];
        layer6[59][39:32] = buffer_data_0[4583:4576];
        layer6[59][47:40] = buffer_data_0[4591:4584];
        layer6[59][55:48] = buffer_data_0[4599:4592];
        layer0[60][7:0] = buffer_data_6[4559:4552];
        layer0[60][15:8] = buffer_data_6[4567:4560];
        layer0[60][23:16] = buffer_data_6[4575:4568];
        layer0[60][31:24] = buffer_data_6[4583:4576];
        layer0[60][39:32] = buffer_data_6[4591:4584];
        layer0[60][47:40] = buffer_data_6[4599:4592];
        layer0[60][55:48] = buffer_data_6[4607:4600];
        layer1[60][7:0] = buffer_data_5[4559:4552];
        layer1[60][15:8] = buffer_data_5[4567:4560];
        layer1[60][23:16] = buffer_data_5[4575:4568];
        layer1[60][31:24] = buffer_data_5[4583:4576];
        layer1[60][39:32] = buffer_data_5[4591:4584];
        layer1[60][47:40] = buffer_data_5[4599:4592];
        layer1[60][55:48] = buffer_data_5[4607:4600];
        layer2[60][7:0] = buffer_data_4[4559:4552];
        layer2[60][15:8] = buffer_data_4[4567:4560];
        layer2[60][23:16] = buffer_data_4[4575:4568];
        layer2[60][31:24] = buffer_data_4[4583:4576];
        layer2[60][39:32] = buffer_data_4[4591:4584];
        layer2[60][47:40] = buffer_data_4[4599:4592];
        layer2[60][55:48] = buffer_data_4[4607:4600];
        layer3[60][7:0] = buffer_data_3[4559:4552];
        layer3[60][15:8] = buffer_data_3[4567:4560];
        layer3[60][23:16] = buffer_data_3[4575:4568];
        layer3[60][31:24] = buffer_data_3[4583:4576];
        layer3[60][39:32] = buffer_data_3[4591:4584];
        layer3[60][47:40] = buffer_data_3[4599:4592];
        layer3[60][55:48] = buffer_data_3[4607:4600];
        layer4[60][7:0] = buffer_data_2[4559:4552];
        layer4[60][15:8] = buffer_data_2[4567:4560];
        layer4[60][23:16] = buffer_data_2[4575:4568];
        layer4[60][31:24] = buffer_data_2[4583:4576];
        layer4[60][39:32] = buffer_data_2[4591:4584];
        layer4[60][47:40] = buffer_data_2[4599:4592];
        layer4[60][55:48] = buffer_data_2[4607:4600];
        layer5[60][7:0] = buffer_data_1[4559:4552];
        layer5[60][15:8] = buffer_data_1[4567:4560];
        layer5[60][23:16] = buffer_data_1[4575:4568];
        layer5[60][31:24] = buffer_data_1[4583:4576];
        layer5[60][39:32] = buffer_data_1[4591:4584];
        layer5[60][47:40] = buffer_data_1[4599:4592];
        layer5[60][55:48] = buffer_data_1[4607:4600];
        layer6[60][7:0] = buffer_data_0[4559:4552];
        layer6[60][15:8] = buffer_data_0[4567:4560];
        layer6[60][23:16] = buffer_data_0[4575:4568];
        layer6[60][31:24] = buffer_data_0[4583:4576];
        layer6[60][39:32] = buffer_data_0[4591:4584];
        layer6[60][47:40] = buffer_data_0[4599:4592];
        layer6[60][55:48] = buffer_data_0[4607:4600];
        layer0[61][7:0] = buffer_data_6[4567:4560];
        layer0[61][15:8] = buffer_data_6[4575:4568];
        layer0[61][23:16] = buffer_data_6[4583:4576];
        layer0[61][31:24] = buffer_data_6[4591:4584];
        layer0[61][39:32] = buffer_data_6[4599:4592];
        layer0[61][47:40] = buffer_data_6[4607:4600];
        layer0[61][55:48] = buffer_data_6[4615:4608];
        layer1[61][7:0] = buffer_data_5[4567:4560];
        layer1[61][15:8] = buffer_data_5[4575:4568];
        layer1[61][23:16] = buffer_data_5[4583:4576];
        layer1[61][31:24] = buffer_data_5[4591:4584];
        layer1[61][39:32] = buffer_data_5[4599:4592];
        layer1[61][47:40] = buffer_data_5[4607:4600];
        layer1[61][55:48] = buffer_data_5[4615:4608];
        layer2[61][7:0] = buffer_data_4[4567:4560];
        layer2[61][15:8] = buffer_data_4[4575:4568];
        layer2[61][23:16] = buffer_data_4[4583:4576];
        layer2[61][31:24] = buffer_data_4[4591:4584];
        layer2[61][39:32] = buffer_data_4[4599:4592];
        layer2[61][47:40] = buffer_data_4[4607:4600];
        layer2[61][55:48] = buffer_data_4[4615:4608];
        layer3[61][7:0] = buffer_data_3[4567:4560];
        layer3[61][15:8] = buffer_data_3[4575:4568];
        layer3[61][23:16] = buffer_data_3[4583:4576];
        layer3[61][31:24] = buffer_data_3[4591:4584];
        layer3[61][39:32] = buffer_data_3[4599:4592];
        layer3[61][47:40] = buffer_data_3[4607:4600];
        layer3[61][55:48] = buffer_data_3[4615:4608];
        layer4[61][7:0] = buffer_data_2[4567:4560];
        layer4[61][15:8] = buffer_data_2[4575:4568];
        layer4[61][23:16] = buffer_data_2[4583:4576];
        layer4[61][31:24] = buffer_data_2[4591:4584];
        layer4[61][39:32] = buffer_data_2[4599:4592];
        layer4[61][47:40] = buffer_data_2[4607:4600];
        layer4[61][55:48] = buffer_data_2[4615:4608];
        layer5[61][7:0] = buffer_data_1[4567:4560];
        layer5[61][15:8] = buffer_data_1[4575:4568];
        layer5[61][23:16] = buffer_data_1[4583:4576];
        layer5[61][31:24] = buffer_data_1[4591:4584];
        layer5[61][39:32] = buffer_data_1[4599:4592];
        layer5[61][47:40] = buffer_data_1[4607:4600];
        layer5[61][55:48] = buffer_data_1[4615:4608];
        layer6[61][7:0] = buffer_data_0[4567:4560];
        layer6[61][15:8] = buffer_data_0[4575:4568];
        layer6[61][23:16] = buffer_data_0[4583:4576];
        layer6[61][31:24] = buffer_data_0[4591:4584];
        layer6[61][39:32] = buffer_data_0[4599:4592];
        layer6[61][47:40] = buffer_data_0[4607:4600];
        layer6[61][55:48] = buffer_data_0[4615:4608];
        layer0[62][7:0] = buffer_data_6[4575:4568];
        layer0[62][15:8] = buffer_data_6[4583:4576];
        layer0[62][23:16] = buffer_data_6[4591:4584];
        layer0[62][31:24] = buffer_data_6[4599:4592];
        layer0[62][39:32] = buffer_data_6[4607:4600];
        layer0[62][47:40] = buffer_data_6[4615:4608];
        layer0[62][55:48] = buffer_data_6[4623:4616];
        layer1[62][7:0] = buffer_data_5[4575:4568];
        layer1[62][15:8] = buffer_data_5[4583:4576];
        layer1[62][23:16] = buffer_data_5[4591:4584];
        layer1[62][31:24] = buffer_data_5[4599:4592];
        layer1[62][39:32] = buffer_data_5[4607:4600];
        layer1[62][47:40] = buffer_data_5[4615:4608];
        layer1[62][55:48] = buffer_data_5[4623:4616];
        layer2[62][7:0] = buffer_data_4[4575:4568];
        layer2[62][15:8] = buffer_data_4[4583:4576];
        layer2[62][23:16] = buffer_data_4[4591:4584];
        layer2[62][31:24] = buffer_data_4[4599:4592];
        layer2[62][39:32] = buffer_data_4[4607:4600];
        layer2[62][47:40] = buffer_data_4[4615:4608];
        layer2[62][55:48] = buffer_data_4[4623:4616];
        layer3[62][7:0] = buffer_data_3[4575:4568];
        layer3[62][15:8] = buffer_data_3[4583:4576];
        layer3[62][23:16] = buffer_data_3[4591:4584];
        layer3[62][31:24] = buffer_data_3[4599:4592];
        layer3[62][39:32] = buffer_data_3[4607:4600];
        layer3[62][47:40] = buffer_data_3[4615:4608];
        layer3[62][55:48] = buffer_data_3[4623:4616];
        layer4[62][7:0] = buffer_data_2[4575:4568];
        layer4[62][15:8] = buffer_data_2[4583:4576];
        layer4[62][23:16] = buffer_data_2[4591:4584];
        layer4[62][31:24] = buffer_data_2[4599:4592];
        layer4[62][39:32] = buffer_data_2[4607:4600];
        layer4[62][47:40] = buffer_data_2[4615:4608];
        layer4[62][55:48] = buffer_data_2[4623:4616];
        layer5[62][7:0] = buffer_data_1[4575:4568];
        layer5[62][15:8] = buffer_data_1[4583:4576];
        layer5[62][23:16] = buffer_data_1[4591:4584];
        layer5[62][31:24] = buffer_data_1[4599:4592];
        layer5[62][39:32] = buffer_data_1[4607:4600];
        layer5[62][47:40] = buffer_data_1[4615:4608];
        layer5[62][55:48] = buffer_data_1[4623:4616];
        layer6[62][7:0] = buffer_data_0[4575:4568];
        layer6[62][15:8] = buffer_data_0[4583:4576];
        layer6[62][23:16] = buffer_data_0[4591:4584];
        layer6[62][31:24] = buffer_data_0[4599:4592];
        layer6[62][39:32] = buffer_data_0[4607:4600];
        layer6[62][47:40] = buffer_data_0[4615:4608];
        layer6[62][55:48] = buffer_data_0[4623:4616];
        layer0[63][7:0] = buffer_data_6[4583:4576];
        layer0[63][15:8] = buffer_data_6[4591:4584];
        layer0[63][23:16] = buffer_data_6[4599:4592];
        layer0[63][31:24] = buffer_data_6[4607:4600];
        layer0[63][39:32] = buffer_data_6[4615:4608];
        layer0[63][47:40] = buffer_data_6[4623:4616];
        layer0[63][55:48] = buffer_data_6[4631:4624];
        layer1[63][7:0] = buffer_data_5[4583:4576];
        layer1[63][15:8] = buffer_data_5[4591:4584];
        layer1[63][23:16] = buffer_data_5[4599:4592];
        layer1[63][31:24] = buffer_data_5[4607:4600];
        layer1[63][39:32] = buffer_data_5[4615:4608];
        layer1[63][47:40] = buffer_data_5[4623:4616];
        layer1[63][55:48] = buffer_data_5[4631:4624];
        layer2[63][7:0] = buffer_data_4[4583:4576];
        layer2[63][15:8] = buffer_data_4[4591:4584];
        layer2[63][23:16] = buffer_data_4[4599:4592];
        layer2[63][31:24] = buffer_data_4[4607:4600];
        layer2[63][39:32] = buffer_data_4[4615:4608];
        layer2[63][47:40] = buffer_data_4[4623:4616];
        layer2[63][55:48] = buffer_data_4[4631:4624];
        layer3[63][7:0] = buffer_data_3[4583:4576];
        layer3[63][15:8] = buffer_data_3[4591:4584];
        layer3[63][23:16] = buffer_data_3[4599:4592];
        layer3[63][31:24] = buffer_data_3[4607:4600];
        layer3[63][39:32] = buffer_data_3[4615:4608];
        layer3[63][47:40] = buffer_data_3[4623:4616];
        layer3[63][55:48] = buffer_data_3[4631:4624];
        layer4[63][7:0] = buffer_data_2[4583:4576];
        layer4[63][15:8] = buffer_data_2[4591:4584];
        layer4[63][23:16] = buffer_data_2[4599:4592];
        layer4[63][31:24] = buffer_data_2[4607:4600];
        layer4[63][39:32] = buffer_data_2[4615:4608];
        layer4[63][47:40] = buffer_data_2[4623:4616];
        layer4[63][55:48] = buffer_data_2[4631:4624];
        layer5[63][7:0] = buffer_data_1[4583:4576];
        layer5[63][15:8] = buffer_data_1[4591:4584];
        layer5[63][23:16] = buffer_data_1[4599:4592];
        layer5[63][31:24] = buffer_data_1[4607:4600];
        layer5[63][39:32] = buffer_data_1[4615:4608];
        layer5[63][47:40] = buffer_data_1[4623:4616];
        layer5[63][55:48] = buffer_data_1[4631:4624];
        layer6[63][7:0] = buffer_data_0[4583:4576];
        layer6[63][15:8] = buffer_data_0[4591:4584];
        layer6[63][23:16] = buffer_data_0[4599:4592];
        layer6[63][31:24] = buffer_data_0[4607:4600];
        layer6[63][39:32] = buffer_data_0[4615:4608];
        layer6[63][47:40] = buffer_data_0[4623:4616];
        layer6[63][55:48] = buffer_data_0[4631:4624];
    end
    ST_GAUSSIAN_9: begin
        layer0[0][7:0] = buffer_data_6[4591:4584];
        layer0[0][15:8] = buffer_data_6[4599:4592];
        layer0[0][23:16] = buffer_data_6[4607:4600];
        layer0[0][31:24] = buffer_data_6[4615:4608];
        layer0[0][39:32] = buffer_data_6[4623:4616];
        layer0[0][47:40] = buffer_data_6[4631:4624];
        layer0[0][55:48] = buffer_data_6[4639:4632];
        layer1[0][7:0] = buffer_data_5[4591:4584];
        layer1[0][15:8] = buffer_data_5[4599:4592];
        layer1[0][23:16] = buffer_data_5[4607:4600];
        layer1[0][31:24] = buffer_data_5[4615:4608];
        layer1[0][39:32] = buffer_data_5[4623:4616];
        layer1[0][47:40] = buffer_data_5[4631:4624];
        layer1[0][55:48] = buffer_data_5[4639:4632];
        layer2[0][7:0] = buffer_data_4[4591:4584];
        layer2[0][15:8] = buffer_data_4[4599:4592];
        layer2[0][23:16] = buffer_data_4[4607:4600];
        layer2[0][31:24] = buffer_data_4[4615:4608];
        layer2[0][39:32] = buffer_data_4[4623:4616];
        layer2[0][47:40] = buffer_data_4[4631:4624];
        layer2[0][55:48] = buffer_data_4[4639:4632];
        layer3[0][7:0] = buffer_data_3[4591:4584];
        layer3[0][15:8] = buffer_data_3[4599:4592];
        layer3[0][23:16] = buffer_data_3[4607:4600];
        layer3[0][31:24] = buffer_data_3[4615:4608];
        layer3[0][39:32] = buffer_data_3[4623:4616];
        layer3[0][47:40] = buffer_data_3[4631:4624];
        layer3[0][55:48] = buffer_data_3[4639:4632];
        layer4[0][7:0] = buffer_data_2[4591:4584];
        layer4[0][15:8] = buffer_data_2[4599:4592];
        layer4[0][23:16] = buffer_data_2[4607:4600];
        layer4[0][31:24] = buffer_data_2[4615:4608];
        layer4[0][39:32] = buffer_data_2[4623:4616];
        layer4[0][47:40] = buffer_data_2[4631:4624];
        layer4[0][55:48] = buffer_data_2[4639:4632];
        layer5[0][7:0] = buffer_data_1[4591:4584];
        layer5[0][15:8] = buffer_data_1[4599:4592];
        layer5[0][23:16] = buffer_data_1[4607:4600];
        layer5[0][31:24] = buffer_data_1[4615:4608];
        layer5[0][39:32] = buffer_data_1[4623:4616];
        layer5[0][47:40] = buffer_data_1[4631:4624];
        layer5[0][55:48] = buffer_data_1[4639:4632];
        layer6[0][7:0] = buffer_data_0[4591:4584];
        layer6[0][15:8] = buffer_data_0[4599:4592];
        layer6[0][23:16] = buffer_data_0[4607:4600];
        layer6[0][31:24] = buffer_data_0[4615:4608];
        layer6[0][39:32] = buffer_data_0[4623:4616];
        layer6[0][47:40] = buffer_data_0[4631:4624];
        layer6[0][55:48] = buffer_data_0[4639:4632];
        layer0[1][7:0] = buffer_data_6[4599:4592];
        layer0[1][15:8] = buffer_data_6[4607:4600];
        layer0[1][23:16] = buffer_data_6[4615:4608];
        layer0[1][31:24] = buffer_data_6[4623:4616];
        layer0[1][39:32] = buffer_data_6[4631:4624];
        layer0[1][47:40] = buffer_data_6[4639:4632];
        layer0[1][55:48] = buffer_data_6[4647:4640];
        layer1[1][7:0] = buffer_data_5[4599:4592];
        layer1[1][15:8] = buffer_data_5[4607:4600];
        layer1[1][23:16] = buffer_data_5[4615:4608];
        layer1[1][31:24] = buffer_data_5[4623:4616];
        layer1[1][39:32] = buffer_data_5[4631:4624];
        layer1[1][47:40] = buffer_data_5[4639:4632];
        layer1[1][55:48] = buffer_data_5[4647:4640];
        layer2[1][7:0] = buffer_data_4[4599:4592];
        layer2[1][15:8] = buffer_data_4[4607:4600];
        layer2[1][23:16] = buffer_data_4[4615:4608];
        layer2[1][31:24] = buffer_data_4[4623:4616];
        layer2[1][39:32] = buffer_data_4[4631:4624];
        layer2[1][47:40] = buffer_data_4[4639:4632];
        layer2[1][55:48] = buffer_data_4[4647:4640];
        layer3[1][7:0] = buffer_data_3[4599:4592];
        layer3[1][15:8] = buffer_data_3[4607:4600];
        layer3[1][23:16] = buffer_data_3[4615:4608];
        layer3[1][31:24] = buffer_data_3[4623:4616];
        layer3[1][39:32] = buffer_data_3[4631:4624];
        layer3[1][47:40] = buffer_data_3[4639:4632];
        layer3[1][55:48] = buffer_data_3[4647:4640];
        layer4[1][7:0] = buffer_data_2[4599:4592];
        layer4[1][15:8] = buffer_data_2[4607:4600];
        layer4[1][23:16] = buffer_data_2[4615:4608];
        layer4[1][31:24] = buffer_data_2[4623:4616];
        layer4[1][39:32] = buffer_data_2[4631:4624];
        layer4[1][47:40] = buffer_data_2[4639:4632];
        layer4[1][55:48] = buffer_data_2[4647:4640];
        layer5[1][7:0] = buffer_data_1[4599:4592];
        layer5[1][15:8] = buffer_data_1[4607:4600];
        layer5[1][23:16] = buffer_data_1[4615:4608];
        layer5[1][31:24] = buffer_data_1[4623:4616];
        layer5[1][39:32] = buffer_data_1[4631:4624];
        layer5[1][47:40] = buffer_data_1[4639:4632];
        layer5[1][55:48] = buffer_data_1[4647:4640];
        layer6[1][7:0] = buffer_data_0[4599:4592];
        layer6[1][15:8] = buffer_data_0[4607:4600];
        layer6[1][23:16] = buffer_data_0[4615:4608];
        layer6[1][31:24] = buffer_data_0[4623:4616];
        layer6[1][39:32] = buffer_data_0[4631:4624];
        layer6[1][47:40] = buffer_data_0[4639:4632];
        layer6[1][55:48] = buffer_data_0[4647:4640];
        layer0[2][7:0] = buffer_data_6[4607:4600];
        layer0[2][15:8] = buffer_data_6[4615:4608];
        layer0[2][23:16] = buffer_data_6[4623:4616];
        layer0[2][31:24] = buffer_data_6[4631:4624];
        layer0[2][39:32] = buffer_data_6[4639:4632];
        layer0[2][47:40] = buffer_data_6[4647:4640];
        layer0[2][55:48] = buffer_data_6[4655:4648];
        layer1[2][7:0] = buffer_data_5[4607:4600];
        layer1[2][15:8] = buffer_data_5[4615:4608];
        layer1[2][23:16] = buffer_data_5[4623:4616];
        layer1[2][31:24] = buffer_data_5[4631:4624];
        layer1[2][39:32] = buffer_data_5[4639:4632];
        layer1[2][47:40] = buffer_data_5[4647:4640];
        layer1[2][55:48] = buffer_data_5[4655:4648];
        layer2[2][7:0] = buffer_data_4[4607:4600];
        layer2[2][15:8] = buffer_data_4[4615:4608];
        layer2[2][23:16] = buffer_data_4[4623:4616];
        layer2[2][31:24] = buffer_data_4[4631:4624];
        layer2[2][39:32] = buffer_data_4[4639:4632];
        layer2[2][47:40] = buffer_data_4[4647:4640];
        layer2[2][55:48] = buffer_data_4[4655:4648];
        layer3[2][7:0] = buffer_data_3[4607:4600];
        layer3[2][15:8] = buffer_data_3[4615:4608];
        layer3[2][23:16] = buffer_data_3[4623:4616];
        layer3[2][31:24] = buffer_data_3[4631:4624];
        layer3[2][39:32] = buffer_data_3[4639:4632];
        layer3[2][47:40] = buffer_data_3[4647:4640];
        layer3[2][55:48] = buffer_data_3[4655:4648];
        layer4[2][7:0] = buffer_data_2[4607:4600];
        layer4[2][15:8] = buffer_data_2[4615:4608];
        layer4[2][23:16] = buffer_data_2[4623:4616];
        layer4[2][31:24] = buffer_data_2[4631:4624];
        layer4[2][39:32] = buffer_data_2[4639:4632];
        layer4[2][47:40] = buffer_data_2[4647:4640];
        layer4[2][55:48] = buffer_data_2[4655:4648];
        layer5[2][7:0] = buffer_data_1[4607:4600];
        layer5[2][15:8] = buffer_data_1[4615:4608];
        layer5[2][23:16] = buffer_data_1[4623:4616];
        layer5[2][31:24] = buffer_data_1[4631:4624];
        layer5[2][39:32] = buffer_data_1[4639:4632];
        layer5[2][47:40] = buffer_data_1[4647:4640];
        layer5[2][55:48] = buffer_data_1[4655:4648];
        layer6[2][7:0] = buffer_data_0[4607:4600];
        layer6[2][15:8] = buffer_data_0[4615:4608];
        layer6[2][23:16] = buffer_data_0[4623:4616];
        layer6[2][31:24] = buffer_data_0[4631:4624];
        layer6[2][39:32] = buffer_data_0[4639:4632];
        layer6[2][47:40] = buffer_data_0[4647:4640];
        layer6[2][55:48] = buffer_data_0[4655:4648];
        layer0[3][7:0] = buffer_data_6[4615:4608];
        layer0[3][15:8] = buffer_data_6[4623:4616];
        layer0[3][23:16] = buffer_data_6[4631:4624];
        layer0[3][31:24] = buffer_data_6[4639:4632];
        layer0[3][39:32] = buffer_data_6[4647:4640];
        layer0[3][47:40] = buffer_data_6[4655:4648];
        layer0[3][55:48] = buffer_data_6[4663:4656];
        layer1[3][7:0] = buffer_data_5[4615:4608];
        layer1[3][15:8] = buffer_data_5[4623:4616];
        layer1[3][23:16] = buffer_data_5[4631:4624];
        layer1[3][31:24] = buffer_data_5[4639:4632];
        layer1[3][39:32] = buffer_data_5[4647:4640];
        layer1[3][47:40] = buffer_data_5[4655:4648];
        layer1[3][55:48] = buffer_data_5[4663:4656];
        layer2[3][7:0] = buffer_data_4[4615:4608];
        layer2[3][15:8] = buffer_data_4[4623:4616];
        layer2[3][23:16] = buffer_data_4[4631:4624];
        layer2[3][31:24] = buffer_data_4[4639:4632];
        layer2[3][39:32] = buffer_data_4[4647:4640];
        layer2[3][47:40] = buffer_data_4[4655:4648];
        layer2[3][55:48] = buffer_data_4[4663:4656];
        layer3[3][7:0] = buffer_data_3[4615:4608];
        layer3[3][15:8] = buffer_data_3[4623:4616];
        layer3[3][23:16] = buffer_data_3[4631:4624];
        layer3[3][31:24] = buffer_data_3[4639:4632];
        layer3[3][39:32] = buffer_data_3[4647:4640];
        layer3[3][47:40] = buffer_data_3[4655:4648];
        layer3[3][55:48] = buffer_data_3[4663:4656];
        layer4[3][7:0] = buffer_data_2[4615:4608];
        layer4[3][15:8] = buffer_data_2[4623:4616];
        layer4[3][23:16] = buffer_data_2[4631:4624];
        layer4[3][31:24] = buffer_data_2[4639:4632];
        layer4[3][39:32] = buffer_data_2[4647:4640];
        layer4[3][47:40] = buffer_data_2[4655:4648];
        layer4[3][55:48] = buffer_data_2[4663:4656];
        layer5[3][7:0] = buffer_data_1[4615:4608];
        layer5[3][15:8] = buffer_data_1[4623:4616];
        layer5[3][23:16] = buffer_data_1[4631:4624];
        layer5[3][31:24] = buffer_data_1[4639:4632];
        layer5[3][39:32] = buffer_data_1[4647:4640];
        layer5[3][47:40] = buffer_data_1[4655:4648];
        layer5[3][55:48] = buffer_data_1[4663:4656];
        layer6[3][7:0] = buffer_data_0[4615:4608];
        layer6[3][15:8] = buffer_data_0[4623:4616];
        layer6[3][23:16] = buffer_data_0[4631:4624];
        layer6[3][31:24] = buffer_data_0[4639:4632];
        layer6[3][39:32] = buffer_data_0[4647:4640];
        layer6[3][47:40] = buffer_data_0[4655:4648];
        layer6[3][55:48] = buffer_data_0[4663:4656];
        layer0[4][7:0] = buffer_data_6[4623:4616];
        layer0[4][15:8] = buffer_data_6[4631:4624];
        layer0[4][23:16] = buffer_data_6[4639:4632];
        layer0[4][31:24] = buffer_data_6[4647:4640];
        layer0[4][39:32] = buffer_data_6[4655:4648];
        layer0[4][47:40] = buffer_data_6[4663:4656];
        layer0[4][55:48] = buffer_data_6[4671:4664];
        layer1[4][7:0] = buffer_data_5[4623:4616];
        layer1[4][15:8] = buffer_data_5[4631:4624];
        layer1[4][23:16] = buffer_data_5[4639:4632];
        layer1[4][31:24] = buffer_data_5[4647:4640];
        layer1[4][39:32] = buffer_data_5[4655:4648];
        layer1[4][47:40] = buffer_data_5[4663:4656];
        layer1[4][55:48] = buffer_data_5[4671:4664];
        layer2[4][7:0] = buffer_data_4[4623:4616];
        layer2[4][15:8] = buffer_data_4[4631:4624];
        layer2[4][23:16] = buffer_data_4[4639:4632];
        layer2[4][31:24] = buffer_data_4[4647:4640];
        layer2[4][39:32] = buffer_data_4[4655:4648];
        layer2[4][47:40] = buffer_data_4[4663:4656];
        layer2[4][55:48] = buffer_data_4[4671:4664];
        layer3[4][7:0] = buffer_data_3[4623:4616];
        layer3[4][15:8] = buffer_data_3[4631:4624];
        layer3[4][23:16] = buffer_data_3[4639:4632];
        layer3[4][31:24] = buffer_data_3[4647:4640];
        layer3[4][39:32] = buffer_data_3[4655:4648];
        layer3[4][47:40] = buffer_data_3[4663:4656];
        layer3[4][55:48] = buffer_data_3[4671:4664];
        layer4[4][7:0] = buffer_data_2[4623:4616];
        layer4[4][15:8] = buffer_data_2[4631:4624];
        layer4[4][23:16] = buffer_data_2[4639:4632];
        layer4[4][31:24] = buffer_data_2[4647:4640];
        layer4[4][39:32] = buffer_data_2[4655:4648];
        layer4[4][47:40] = buffer_data_2[4663:4656];
        layer4[4][55:48] = buffer_data_2[4671:4664];
        layer5[4][7:0] = buffer_data_1[4623:4616];
        layer5[4][15:8] = buffer_data_1[4631:4624];
        layer5[4][23:16] = buffer_data_1[4639:4632];
        layer5[4][31:24] = buffer_data_1[4647:4640];
        layer5[4][39:32] = buffer_data_1[4655:4648];
        layer5[4][47:40] = buffer_data_1[4663:4656];
        layer5[4][55:48] = buffer_data_1[4671:4664];
        layer6[4][7:0] = buffer_data_0[4623:4616];
        layer6[4][15:8] = buffer_data_0[4631:4624];
        layer6[4][23:16] = buffer_data_0[4639:4632];
        layer6[4][31:24] = buffer_data_0[4647:4640];
        layer6[4][39:32] = buffer_data_0[4655:4648];
        layer6[4][47:40] = buffer_data_0[4663:4656];
        layer6[4][55:48] = buffer_data_0[4671:4664];
        layer0[5][7:0] = buffer_data_6[4631:4624];
        layer0[5][15:8] = buffer_data_6[4639:4632];
        layer0[5][23:16] = buffer_data_6[4647:4640];
        layer0[5][31:24] = buffer_data_6[4655:4648];
        layer0[5][39:32] = buffer_data_6[4663:4656];
        layer0[5][47:40] = buffer_data_6[4671:4664];
        layer0[5][55:48] = buffer_data_6[4679:4672];
        layer1[5][7:0] = buffer_data_5[4631:4624];
        layer1[5][15:8] = buffer_data_5[4639:4632];
        layer1[5][23:16] = buffer_data_5[4647:4640];
        layer1[5][31:24] = buffer_data_5[4655:4648];
        layer1[5][39:32] = buffer_data_5[4663:4656];
        layer1[5][47:40] = buffer_data_5[4671:4664];
        layer1[5][55:48] = buffer_data_5[4679:4672];
        layer2[5][7:0] = buffer_data_4[4631:4624];
        layer2[5][15:8] = buffer_data_4[4639:4632];
        layer2[5][23:16] = buffer_data_4[4647:4640];
        layer2[5][31:24] = buffer_data_4[4655:4648];
        layer2[5][39:32] = buffer_data_4[4663:4656];
        layer2[5][47:40] = buffer_data_4[4671:4664];
        layer2[5][55:48] = buffer_data_4[4679:4672];
        layer3[5][7:0] = buffer_data_3[4631:4624];
        layer3[5][15:8] = buffer_data_3[4639:4632];
        layer3[5][23:16] = buffer_data_3[4647:4640];
        layer3[5][31:24] = buffer_data_3[4655:4648];
        layer3[5][39:32] = buffer_data_3[4663:4656];
        layer3[5][47:40] = buffer_data_3[4671:4664];
        layer3[5][55:48] = buffer_data_3[4679:4672];
        layer4[5][7:0] = buffer_data_2[4631:4624];
        layer4[5][15:8] = buffer_data_2[4639:4632];
        layer4[5][23:16] = buffer_data_2[4647:4640];
        layer4[5][31:24] = buffer_data_2[4655:4648];
        layer4[5][39:32] = buffer_data_2[4663:4656];
        layer4[5][47:40] = buffer_data_2[4671:4664];
        layer4[5][55:48] = buffer_data_2[4679:4672];
        layer5[5][7:0] = buffer_data_1[4631:4624];
        layer5[5][15:8] = buffer_data_1[4639:4632];
        layer5[5][23:16] = buffer_data_1[4647:4640];
        layer5[5][31:24] = buffer_data_1[4655:4648];
        layer5[5][39:32] = buffer_data_1[4663:4656];
        layer5[5][47:40] = buffer_data_1[4671:4664];
        layer5[5][55:48] = buffer_data_1[4679:4672];
        layer6[5][7:0] = buffer_data_0[4631:4624];
        layer6[5][15:8] = buffer_data_0[4639:4632];
        layer6[5][23:16] = buffer_data_0[4647:4640];
        layer6[5][31:24] = buffer_data_0[4655:4648];
        layer6[5][39:32] = buffer_data_0[4663:4656];
        layer6[5][47:40] = buffer_data_0[4671:4664];
        layer6[5][55:48] = buffer_data_0[4679:4672];
        layer0[6][7:0] = buffer_data_6[4639:4632];
        layer0[6][15:8] = buffer_data_6[4647:4640];
        layer0[6][23:16] = buffer_data_6[4655:4648];
        layer0[6][31:24] = buffer_data_6[4663:4656];
        layer0[6][39:32] = buffer_data_6[4671:4664];
        layer0[6][47:40] = buffer_data_6[4679:4672];
        layer0[6][55:48] = buffer_data_6[4687:4680];
        layer1[6][7:0] = buffer_data_5[4639:4632];
        layer1[6][15:8] = buffer_data_5[4647:4640];
        layer1[6][23:16] = buffer_data_5[4655:4648];
        layer1[6][31:24] = buffer_data_5[4663:4656];
        layer1[6][39:32] = buffer_data_5[4671:4664];
        layer1[6][47:40] = buffer_data_5[4679:4672];
        layer1[6][55:48] = buffer_data_5[4687:4680];
        layer2[6][7:0] = buffer_data_4[4639:4632];
        layer2[6][15:8] = buffer_data_4[4647:4640];
        layer2[6][23:16] = buffer_data_4[4655:4648];
        layer2[6][31:24] = buffer_data_4[4663:4656];
        layer2[6][39:32] = buffer_data_4[4671:4664];
        layer2[6][47:40] = buffer_data_4[4679:4672];
        layer2[6][55:48] = buffer_data_4[4687:4680];
        layer3[6][7:0] = buffer_data_3[4639:4632];
        layer3[6][15:8] = buffer_data_3[4647:4640];
        layer3[6][23:16] = buffer_data_3[4655:4648];
        layer3[6][31:24] = buffer_data_3[4663:4656];
        layer3[6][39:32] = buffer_data_3[4671:4664];
        layer3[6][47:40] = buffer_data_3[4679:4672];
        layer3[6][55:48] = buffer_data_3[4687:4680];
        layer4[6][7:0] = buffer_data_2[4639:4632];
        layer4[6][15:8] = buffer_data_2[4647:4640];
        layer4[6][23:16] = buffer_data_2[4655:4648];
        layer4[6][31:24] = buffer_data_2[4663:4656];
        layer4[6][39:32] = buffer_data_2[4671:4664];
        layer4[6][47:40] = buffer_data_2[4679:4672];
        layer4[6][55:48] = buffer_data_2[4687:4680];
        layer5[6][7:0] = buffer_data_1[4639:4632];
        layer5[6][15:8] = buffer_data_1[4647:4640];
        layer5[6][23:16] = buffer_data_1[4655:4648];
        layer5[6][31:24] = buffer_data_1[4663:4656];
        layer5[6][39:32] = buffer_data_1[4671:4664];
        layer5[6][47:40] = buffer_data_1[4679:4672];
        layer5[6][55:48] = buffer_data_1[4687:4680];
        layer6[6][7:0] = buffer_data_0[4639:4632];
        layer6[6][15:8] = buffer_data_0[4647:4640];
        layer6[6][23:16] = buffer_data_0[4655:4648];
        layer6[6][31:24] = buffer_data_0[4663:4656];
        layer6[6][39:32] = buffer_data_0[4671:4664];
        layer6[6][47:40] = buffer_data_0[4679:4672];
        layer6[6][55:48] = buffer_data_0[4687:4680];
        layer0[7][7:0] = buffer_data_6[4647:4640];
        layer0[7][15:8] = buffer_data_6[4655:4648];
        layer0[7][23:16] = buffer_data_6[4663:4656];
        layer0[7][31:24] = buffer_data_6[4671:4664];
        layer0[7][39:32] = buffer_data_6[4679:4672];
        layer0[7][47:40] = buffer_data_6[4687:4680];
        layer0[7][55:48] = buffer_data_6[4695:4688];
        layer1[7][7:0] = buffer_data_5[4647:4640];
        layer1[7][15:8] = buffer_data_5[4655:4648];
        layer1[7][23:16] = buffer_data_5[4663:4656];
        layer1[7][31:24] = buffer_data_5[4671:4664];
        layer1[7][39:32] = buffer_data_5[4679:4672];
        layer1[7][47:40] = buffer_data_5[4687:4680];
        layer1[7][55:48] = buffer_data_5[4695:4688];
        layer2[7][7:0] = buffer_data_4[4647:4640];
        layer2[7][15:8] = buffer_data_4[4655:4648];
        layer2[7][23:16] = buffer_data_4[4663:4656];
        layer2[7][31:24] = buffer_data_4[4671:4664];
        layer2[7][39:32] = buffer_data_4[4679:4672];
        layer2[7][47:40] = buffer_data_4[4687:4680];
        layer2[7][55:48] = buffer_data_4[4695:4688];
        layer3[7][7:0] = buffer_data_3[4647:4640];
        layer3[7][15:8] = buffer_data_3[4655:4648];
        layer3[7][23:16] = buffer_data_3[4663:4656];
        layer3[7][31:24] = buffer_data_3[4671:4664];
        layer3[7][39:32] = buffer_data_3[4679:4672];
        layer3[7][47:40] = buffer_data_3[4687:4680];
        layer3[7][55:48] = buffer_data_3[4695:4688];
        layer4[7][7:0] = buffer_data_2[4647:4640];
        layer4[7][15:8] = buffer_data_2[4655:4648];
        layer4[7][23:16] = buffer_data_2[4663:4656];
        layer4[7][31:24] = buffer_data_2[4671:4664];
        layer4[7][39:32] = buffer_data_2[4679:4672];
        layer4[7][47:40] = buffer_data_2[4687:4680];
        layer4[7][55:48] = buffer_data_2[4695:4688];
        layer5[7][7:0] = buffer_data_1[4647:4640];
        layer5[7][15:8] = buffer_data_1[4655:4648];
        layer5[7][23:16] = buffer_data_1[4663:4656];
        layer5[7][31:24] = buffer_data_1[4671:4664];
        layer5[7][39:32] = buffer_data_1[4679:4672];
        layer5[7][47:40] = buffer_data_1[4687:4680];
        layer5[7][55:48] = buffer_data_1[4695:4688];
        layer6[7][7:0] = buffer_data_0[4647:4640];
        layer6[7][15:8] = buffer_data_0[4655:4648];
        layer6[7][23:16] = buffer_data_0[4663:4656];
        layer6[7][31:24] = buffer_data_0[4671:4664];
        layer6[7][39:32] = buffer_data_0[4679:4672];
        layer6[7][47:40] = buffer_data_0[4687:4680];
        layer6[7][55:48] = buffer_data_0[4695:4688];
        layer0[8][7:0] = buffer_data_6[4655:4648];
        layer0[8][15:8] = buffer_data_6[4663:4656];
        layer0[8][23:16] = buffer_data_6[4671:4664];
        layer0[8][31:24] = buffer_data_6[4679:4672];
        layer0[8][39:32] = buffer_data_6[4687:4680];
        layer0[8][47:40] = buffer_data_6[4695:4688];
        layer0[8][55:48] = buffer_data_6[4703:4696];
        layer1[8][7:0] = buffer_data_5[4655:4648];
        layer1[8][15:8] = buffer_data_5[4663:4656];
        layer1[8][23:16] = buffer_data_5[4671:4664];
        layer1[8][31:24] = buffer_data_5[4679:4672];
        layer1[8][39:32] = buffer_data_5[4687:4680];
        layer1[8][47:40] = buffer_data_5[4695:4688];
        layer1[8][55:48] = buffer_data_5[4703:4696];
        layer2[8][7:0] = buffer_data_4[4655:4648];
        layer2[8][15:8] = buffer_data_4[4663:4656];
        layer2[8][23:16] = buffer_data_4[4671:4664];
        layer2[8][31:24] = buffer_data_4[4679:4672];
        layer2[8][39:32] = buffer_data_4[4687:4680];
        layer2[8][47:40] = buffer_data_4[4695:4688];
        layer2[8][55:48] = buffer_data_4[4703:4696];
        layer3[8][7:0] = buffer_data_3[4655:4648];
        layer3[8][15:8] = buffer_data_3[4663:4656];
        layer3[8][23:16] = buffer_data_3[4671:4664];
        layer3[8][31:24] = buffer_data_3[4679:4672];
        layer3[8][39:32] = buffer_data_3[4687:4680];
        layer3[8][47:40] = buffer_data_3[4695:4688];
        layer3[8][55:48] = buffer_data_3[4703:4696];
        layer4[8][7:0] = buffer_data_2[4655:4648];
        layer4[8][15:8] = buffer_data_2[4663:4656];
        layer4[8][23:16] = buffer_data_2[4671:4664];
        layer4[8][31:24] = buffer_data_2[4679:4672];
        layer4[8][39:32] = buffer_data_2[4687:4680];
        layer4[8][47:40] = buffer_data_2[4695:4688];
        layer4[8][55:48] = buffer_data_2[4703:4696];
        layer5[8][7:0] = buffer_data_1[4655:4648];
        layer5[8][15:8] = buffer_data_1[4663:4656];
        layer5[8][23:16] = buffer_data_1[4671:4664];
        layer5[8][31:24] = buffer_data_1[4679:4672];
        layer5[8][39:32] = buffer_data_1[4687:4680];
        layer5[8][47:40] = buffer_data_1[4695:4688];
        layer5[8][55:48] = buffer_data_1[4703:4696];
        layer6[8][7:0] = buffer_data_0[4655:4648];
        layer6[8][15:8] = buffer_data_0[4663:4656];
        layer6[8][23:16] = buffer_data_0[4671:4664];
        layer6[8][31:24] = buffer_data_0[4679:4672];
        layer6[8][39:32] = buffer_data_0[4687:4680];
        layer6[8][47:40] = buffer_data_0[4695:4688];
        layer6[8][55:48] = buffer_data_0[4703:4696];
        layer0[9][7:0] = buffer_data_6[4663:4656];
        layer0[9][15:8] = buffer_data_6[4671:4664];
        layer0[9][23:16] = buffer_data_6[4679:4672];
        layer0[9][31:24] = buffer_data_6[4687:4680];
        layer0[9][39:32] = buffer_data_6[4695:4688];
        layer0[9][47:40] = buffer_data_6[4703:4696];
        layer0[9][55:48] = buffer_data_6[4711:4704];
        layer1[9][7:0] = buffer_data_5[4663:4656];
        layer1[9][15:8] = buffer_data_5[4671:4664];
        layer1[9][23:16] = buffer_data_5[4679:4672];
        layer1[9][31:24] = buffer_data_5[4687:4680];
        layer1[9][39:32] = buffer_data_5[4695:4688];
        layer1[9][47:40] = buffer_data_5[4703:4696];
        layer1[9][55:48] = buffer_data_5[4711:4704];
        layer2[9][7:0] = buffer_data_4[4663:4656];
        layer2[9][15:8] = buffer_data_4[4671:4664];
        layer2[9][23:16] = buffer_data_4[4679:4672];
        layer2[9][31:24] = buffer_data_4[4687:4680];
        layer2[9][39:32] = buffer_data_4[4695:4688];
        layer2[9][47:40] = buffer_data_4[4703:4696];
        layer2[9][55:48] = buffer_data_4[4711:4704];
        layer3[9][7:0] = buffer_data_3[4663:4656];
        layer3[9][15:8] = buffer_data_3[4671:4664];
        layer3[9][23:16] = buffer_data_3[4679:4672];
        layer3[9][31:24] = buffer_data_3[4687:4680];
        layer3[9][39:32] = buffer_data_3[4695:4688];
        layer3[9][47:40] = buffer_data_3[4703:4696];
        layer3[9][55:48] = buffer_data_3[4711:4704];
        layer4[9][7:0] = buffer_data_2[4663:4656];
        layer4[9][15:8] = buffer_data_2[4671:4664];
        layer4[9][23:16] = buffer_data_2[4679:4672];
        layer4[9][31:24] = buffer_data_2[4687:4680];
        layer4[9][39:32] = buffer_data_2[4695:4688];
        layer4[9][47:40] = buffer_data_2[4703:4696];
        layer4[9][55:48] = buffer_data_2[4711:4704];
        layer5[9][7:0] = buffer_data_1[4663:4656];
        layer5[9][15:8] = buffer_data_1[4671:4664];
        layer5[9][23:16] = buffer_data_1[4679:4672];
        layer5[9][31:24] = buffer_data_1[4687:4680];
        layer5[9][39:32] = buffer_data_1[4695:4688];
        layer5[9][47:40] = buffer_data_1[4703:4696];
        layer5[9][55:48] = buffer_data_1[4711:4704];
        layer6[9][7:0] = buffer_data_0[4663:4656];
        layer6[9][15:8] = buffer_data_0[4671:4664];
        layer6[9][23:16] = buffer_data_0[4679:4672];
        layer6[9][31:24] = buffer_data_0[4687:4680];
        layer6[9][39:32] = buffer_data_0[4695:4688];
        layer6[9][47:40] = buffer_data_0[4703:4696];
        layer6[9][55:48] = buffer_data_0[4711:4704];
        layer0[10][7:0] = buffer_data_6[4671:4664];
        layer0[10][15:8] = buffer_data_6[4679:4672];
        layer0[10][23:16] = buffer_data_6[4687:4680];
        layer0[10][31:24] = buffer_data_6[4695:4688];
        layer0[10][39:32] = buffer_data_6[4703:4696];
        layer0[10][47:40] = buffer_data_6[4711:4704];
        layer0[10][55:48] = buffer_data_6[4719:4712];
        layer1[10][7:0] = buffer_data_5[4671:4664];
        layer1[10][15:8] = buffer_data_5[4679:4672];
        layer1[10][23:16] = buffer_data_5[4687:4680];
        layer1[10][31:24] = buffer_data_5[4695:4688];
        layer1[10][39:32] = buffer_data_5[4703:4696];
        layer1[10][47:40] = buffer_data_5[4711:4704];
        layer1[10][55:48] = buffer_data_5[4719:4712];
        layer2[10][7:0] = buffer_data_4[4671:4664];
        layer2[10][15:8] = buffer_data_4[4679:4672];
        layer2[10][23:16] = buffer_data_4[4687:4680];
        layer2[10][31:24] = buffer_data_4[4695:4688];
        layer2[10][39:32] = buffer_data_4[4703:4696];
        layer2[10][47:40] = buffer_data_4[4711:4704];
        layer2[10][55:48] = buffer_data_4[4719:4712];
        layer3[10][7:0] = buffer_data_3[4671:4664];
        layer3[10][15:8] = buffer_data_3[4679:4672];
        layer3[10][23:16] = buffer_data_3[4687:4680];
        layer3[10][31:24] = buffer_data_3[4695:4688];
        layer3[10][39:32] = buffer_data_3[4703:4696];
        layer3[10][47:40] = buffer_data_3[4711:4704];
        layer3[10][55:48] = buffer_data_3[4719:4712];
        layer4[10][7:0] = buffer_data_2[4671:4664];
        layer4[10][15:8] = buffer_data_2[4679:4672];
        layer4[10][23:16] = buffer_data_2[4687:4680];
        layer4[10][31:24] = buffer_data_2[4695:4688];
        layer4[10][39:32] = buffer_data_2[4703:4696];
        layer4[10][47:40] = buffer_data_2[4711:4704];
        layer4[10][55:48] = buffer_data_2[4719:4712];
        layer5[10][7:0] = buffer_data_1[4671:4664];
        layer5[10][15:8] = buffer_data_1[4679:4672];
        layer5[10][23:16] = buffer_data_1[4687:4680];
        layer5[10][31:24] = buffer_data_1[4695:4688];
        layer5[10][39:32] = buffer_data_1[4703:4696];
        layer5[10][47:40] = buffer_data_1[4711:4704];
        layer5[10][55:48] = buffer_data_1[4719:4712];
        layer6[10][7:0] = buffer_data_0[4671:4664];
        layer6[10][15:8] = buffer_data_0[4679:4672];
        layer6[10][23:16] = buffer_data_0[4687:4680];
        layer6[10][31:24] = buffer_data_0[4695:4688];
        layer6[10][39:32] = buffer_data_0[4703:4696];
        layer6[10][47:40] = buffer_data_0[4711:4704];
        layer6[10][55:48] = buffer_data_0[4719:4712];
        layer0[11][7:0] = buffer_data_6[4679:4672];
        layer0[11][15:8] = buffer_data_6[4687:4680];
        layer0[11][23:16] = buffer_data_6[4695:4688];
        layer0[11][31:24] = buffer_data_6[4703:4696];
        layer0[11][39:32] = buffer_data_6[4711:4704];
        layer0[11][47:40] = buffer_data_6[4719:4712];
        layer0[11][55:48] = buffer_data_6[4727:4720];
        layer1[11][7:0] = buffer_data_5[4679:4672];
        layer1[11][15:8] = buffer_data_5[4687:4680];
        layer1[11][23:16] = buffer_data_5[4695:4688];
        layer1[11][31:24] = buffer_data_5[4703:4696];
        layer1[11][39:32] = buffer_data_5[4711:4704];
        layer1[11][47:40] = buffer_data_5[4719:4712];
        layer1[11][55:48] = buffer_data_5[4727:4720];
        layer2[11][7:0] = buffer_data_4[4679:4672];
        layer2[11][15:8] = buffer_data_4[4687:4680];
        layer2[11][23:16] = buffer_data_4[4695:4688];
        layer2[11][31:24] = buffer_data_4[4703:4696];
        layer2[11][39:32] = buffer_data_4[4711:4704];
        layer2[11][47:40] = buffer_data_4[4719:4712];
        layer2[11][55:48] = buffer_data_4[4727:4720];
        layer3[11][7:0] = buffer_data_3[4679:4672];
        layer3[11][15:8] = buffer_data_3[4687:4680];
        layer3[11][23:16] = buffer_data_3[4695:4688];
        layer3[11][31:24] = buffer_data_3[4703:4696];
        layer3[11][39:32] = buffer_data_3[4711:4704];
        layer3[11][47:40] = buffer_data_3[4719:4712];
        layer3[11][55:48] = buffer_data_3[4727:4720];
        layer4[11][7:0] = buffer_data_2[4679:4672];
        layer4[11][15:8] = buffer_data_2[4687:4680];
        layer4[11][23:16] = buffer_data_2[4695:4688];
        layer4[11][31:24] = buffer_data_2[4703:4696];
        layer4[11][39:32] = buffer_data_2[4711:4704];
        layer4[11][47:40] = buffer_data_2[4719:4712];
        layer4[11][55:48] = buffer_data_2[4727:4720];
        layer5[11][7:0] = buffer_data_1[4679:4672];
        layer5[11][15:8] = buffer_data_1[4687:4680];
        layer5[11][23:16] = buffer_data_1[4695:4688];
        layer5[11][31:24] = buffer_data_1[4703:4696];
        layer5[11][39:32] = buffer_data_1[4711:4704];
        layer5[11][47:40] = buffer_data_1[4719:4712];
        layer5[11][55:48] = buffer_data_1[4727:4720];
        layer6[11][7:0] = buffer_data_0[4679:4672];
        layer6[11][15:8] = buffer_data_0[4687:4680];
        layer6[11][23:16] = buffer_data_0[4695:4688];
        layer6[11][31:24] = buffer_data_0[4703:4696];
        layer6[11][39:32] = buffer_data_0[4711:4704];
        layer6[11][47:40] = buffer_data_0[4719:4712];
        layer6[11][55:48] = buffer_data_0[4727:4720];
        layer0[12][7:0] = buffer_data_6[4687:4680];
        layer0[12][15:8] = buffer_data_6[4695:4688];
        layer0[12][23:16] = buffer_data_6[4703:4696];
        layer0[12][31:24] = buffer_data_6[4711:4704];
        layer0[12][39:32] = buffer_data_6[4719:4712];
        layer0[12][47:40] = buffer_data_6[4727:4720];
        layer0[12][55:48] = buffer_data_6[4735:4728];
        layer1[12][7:0] = buffer_data_5[4687:4680];
        layer1[12][15:8] = buffer_data_5[4695:4688];
        layer1[12][23:16] = buffer_data_5[4703:4696];
        layer1[12][31:24] = buffer_data_5[4711:4704];
        layer1[12][39:32] = buffer_data_5[4719:4712];
        layer1[12][47:40] = buffer_data_5[4727:4720];
        layer1[12][55:48] = buffer_data_5[4735:4728];
        layer2[12][7:0] = buffer_data_4[4687:4680];
        layer2[12][15:8] = buffer_data_4[4695:4688];
        layer2[12][23:16] = buffer_data_4[4703:4696];
        layer2[12][31:24] = buffer_data_4[4711:4704];
        layer2[12][39:32] = buffer_data_4[4719:4712];
        layer2[12][47:40] = buffer_data_4[4727:4720];
        layer2[12][55:48] = buffer_data_4[4735:4728];
        layer3[12][7:0] = buffer_data_3[4687:4680];
        layer3[12][15:8] = buffer_data_3[4695:4688];
        layer3[12][23:16] = buffer_data_3[4703:4696];
        layer3[12][31:24] = buffer_data_3[4711:4704];
        layer3[12][39:32] = buffer_data_3[4719:4712];
        layer3[12][47:40] = buffer_data_3[4727:4720];
        layer3[12][55:48] = buffer_data_3[4735:4728];
        layer4[12][7:0] = buffer_data_2[4687:4680];
        layer4[12][15:8] = buffer_data_2[4695:4688];
        layer4[12][23:16] = buffer_data_2[4703:4696];
        layer4[12][31:24] = buffer_data_2[4711:4704];
        layer4[12][39:32] = buffer_data_2[4719:4712];
        layer4[12][47:40] = buffer_data_2[4727:4720];
        layer4[12][55:48] = buffer_data_2[4735:4728];
        layer5[12][7:0] = buffer_data_1[4687:4680];
        layer5[12][15:8] = buffer_data_1[4695:4688];
        layer5[12][23:16] = buffer_data_1[4703:4696];
        layer5[12][31:24] = buffer_data_1[4711:4704];
        layer5[12][39:32] = buffer_data_1[4719:4712];
        layer5[12][47:40] = buffer_data_1[4727:4720];
        layer5[12][55:48] = buffer_data_1[4735:4728];
        layer6[12][7:0] = buffer_data_0[4687:4680];
        layer6[12][15:8] = buffer_data_0[4695:4688];
        layer6[12][23:16] = buffer_data_0[4703:4696];
        layer6[12][31:24] = buffer_data_0[4711:4704];
        layer6[12][39:32] = buffer_data_0[4719:4712];
        layer6[12][47:40] = buffer_data_0[4727:4720];
        layer6[12][55:48] = buffer_data_0[4735:4728];
        layer0[13][7:0] = buffer_data_6[4695:4688];
        layer0[13][15:8] = buffer_data_6[4703:4696];
        layer0[13][23:16] = buffer_data_6[4711:4704];
        layer0[13][31:24] = buffer_data_6[4719:4712];
        layer0[13][39:32] = buffer_data_6[4727:4720];
        layer0[13][47:40] = buffer_data_6[4735:4728];
        layer0[13][55:48] = buffer_data_6[4743:4736];
        layer1[13][7:0] = buffer_data_5[4695:4688];
        layer1[13][15:8] = buffer_data_5[4703:4696];
        layer1[13][23:16] = buffer_data_5[4711:4704];
        layer1[13][31:24] = buffer_data_5[4719:4712];
        layer1[13][39:32] = buffer_data_5[4727:4720];
        layer1[13][47:40] = buffer_data_5[4735:4728];
        layer1[13][55:48] = buffer_data_5[4743:4736];
        layer2[13][7:0] = buffer_data_4[4695:4688];
        layer2[13][15:8] = buffer_data_4[4703:4696];
        layer2[13][23:16] = buffer_data_4[4711:4704];
        layer2[13][31:24] = buffer_data_4[4719:4712];
        layer2[13][39:32] = buffer_data_4[4727:4720];
        layer2[13][47:40] = buffer_data_4[4735:4728];
        layer2[13][55:48] = buffer_data_4[4743:4736];
        layer3[13][7:0] = buffer_data_3[4695:4688];
        layer3[13][15:8] = buffer_data_3[4703:4696];
        layer3[13][23:16] = buffer_data_3[4711:4704];
        layer3[13][31:24] = buffer_data_3[4719:4712];
        layer3[13][39:32] = buffer_data_3[4727:4720];
        layer3[13][47:40] = buffer_data_3[4735:4728];
        layer3[13][55:48] = buffer_data_3[4743:4736];
        layer4[13][7:0] = buffer_data_2[4695:4688];
        layer4[13][15:8] = buffer_data_2[4703:4696];
        layer4[13][23:16] = buffer_data_2[4711:4704];
        layer4[13][31:24] = buffer_data_2[4719:4712];
        layer4[13][39:32] = buffer_data_2[4727:4720];
        layer4[13][47:40] = buffer_data_2[4735:4728];
        layer4[13][55:48] = buffer_data_2[4743:4736];
        layer5[13][7:0] = buffer_data_1[4695:4688];
        layer5[13][15:8] = buffer_data_1[4703:4696];
        layer5[13][23:16] = buffer_data_1[4711:4704];
        layer5[13][31:24] = buffer_data_1[4719:4712];
        layer5[13][39:32] = buffer_data_1[4727:4720];
        layer5[13][47:40] = buffer_data_1[4735:4728];
        layer5[13][55:48] = buffer_data_1[4743:4736];
        layer6[13][7:0] = buffer_data_0[4695:4688];
        layer6[13][15:8] = buffer_data_0[4703:4696];
        layer6[13][23:16] = buffer_data_0[4711:4704];
        layer6[13][31:24] = buffer_data_0[4719:4712];
        layer6[13][39:32] = buffer_data_0[4727:4720];
        layer6[13][47:40] = buffer_data_0[4735:4728];
        layer6[13][55:48] = buffer_data_0[4743:4736];
        layer0[14][7:0] = buffer_data_6[4703:4696];
        layer0[14][15:8] = buffer_data_6[4711:4704];
        layer0[14][23:16] = buffer_data_6[4719:4712];
        layer0[14][31:24] = buffer_data_6[4727:4720];
        layer0[14][39:32] = buffer_data_6[4735:4728];
        layer0[14][47:40] = buffer_data_6[4743:4736];
        layer0[14][55:48] = buffer_data_6[4751:4744];
        layer1[14][7:0] = buffer_data_5[4703:4696];
        layer1[14][15:8] = buffer_data_5[4711:4704];
        layer1[14][23:16] = buffer_data_5[4719:4712];
        layer1[14][31:24] = buffer_data_5[4727:4720];
        layer1[14][39:32] = buffer_data_5[4735:4728];
        layer1[14][47:40] = buffer_data_5[4743:4736];
        layer1[14][55:48] = buffer_data_5[4751:4744];
        layer2[14][7:0] = buffer_data_4[4703:4696];
        layer2[14][15:8] = buffer_data_4[4711:4704];
        layer2[14][23:16] = buffer_data_4[4719:4712];
        layer2[14][31:24] = buffer_data_4[4727:4720];
        layer2[14][39:32] = buffer_data_4[4735:4728];
        layer2[14][47:40] = buffer_data_4[4743:4736];
        layer2[14][55:48] = buffer_data_4[4751:4744];
        layer3[14][7:0] = buffer_data_3[4703:4696];
        layer3[14][15:8] = buffer_data_3[4711:4704];
        layer3[14][23:16] = buffer_data_3[4719:4712];
        layer3[14][31:24] = buffer_data_3[4727:4720];
        layer3[14][39:32] = buffer_data_3[4735:4728];
        layer3[14][47:40] = buffer_data_3[4743:4736];
        layer3[14][55:48] = buffer_data_3[4751:4744];
        layer4[14][7:0] = buffer_data_2[4703:4696];
        layer4[14][15:8] = buffer_data_2[4711:4704];
        layer4[14][23:16] = buffer_data_2[4719:4712];
        layer4[14][31:24] = buffer_data_2[4727:4720];
        layer4[14][39:32] = buffer_data_2[4735:4728];
        layer4[14][47:40] = buffer_data_2[4743:4736];
        layer4[14][55:48] = buffer_data_2[4751:4744];
        layer5[14][7:0] = buffer_data_1[4703:4696];
        layer5[14][15:8] = buffer_data_1[4711:4704];
        layer5[14][23:16] = buffer_data_1[4719:4712];
        layer5[14][31:24] = buffer_data_1[4727:4720];
        layer5[14][39:32] = buffer_data_1[4735:4728];
        layer5[14][47:40] = buffer_data_1[4743:4736];
        layer5[14][55:48] = buffer_data_1[4751:4744];
        layer6[14][7:0] = buffer_data_0[4703:4696];
        layer6[14][15:8] = buffer_data_0[4711:4704];
        layer6[14][23:16] = buffer_data_0[4719:4712];
        layer6[14][31:24] = buffer_data_0[4727:4720];
        layer6[14][39:32] = buffer_data_0[4735:4728];
        layer6[14][47:40] = buffer_data_0[4743:4736];
        layer6[14][55:48] = buffer_data_0[4751:4744];
        layer0[15][7:0] = buffer_data_6[4711:4704];
        layer0[15][15:8] = buffer_data_6[4719:4712];
        layer0[15][23:16] = buffer_data_6[4727:4720];
        layer0[15][31:24] = buffer_data_6[4735:4728];
        layer0[15][39:32] = buffer_data_6[4743:4736];
        layer0[15][47:40] = buffer_data_6[4751:4744];
        layer0[15][55:48] = buffer_data_6[4759:4752];
        layer1[15][7:0] = buffer_data_5[4711:4704];
        layer1[15][15:8] = buffer_data_5[4719:4712];
        layer1[15][23:16] = buffer_data_5[4727:4720];
        layer1[15][31:24] = buffer_data_5[4735:4728];
        layer1[15][39:32] = buffer_data_5[4743:4736];
        layer1[15][47:40] = buffer_data_5[4751:4744];
        layer1[15][55:48] = buffer_data_5[4759:4752];
        layer2[15][7:0] = buffer_data_4[4711:4704];
        layer2[15][15:8] = buffer_data_4[4719:4712];
        layer2[15][23:16] = buffer_data_4[4727:4720];
        layer2[15][31:24] = buffer_data_4[4735:4728];
        layer2[15][39:32] = buffer_data_4[4743:4736];
        layer2[15][47:40] = buffer_data_4[4751:4744];
        layer2[15][55:48] = buffer_data_4[4759:4752];
        layer3[15][7:0] = buffer_data_3[4711:4704];
        layer3[15][15:8] = buffer_data_3[4719:4712];
        layer3[15][23:16] = buffer_data_3[4727:4720];
        layer3[15][31:24] = buffer_data_3[4735:4728];
        layer3[15][39:32] = buffer_data_3[4743:4736];
        layer3[15][47:40] = buffer_data_3[4751:4744];
        layer3[15][55:48] = buffer_data_3[4759:4752];
        layer4[15][7:0] = buffer_data_2[4711:4704];
        layer4[15][15:8] = buffer_data_2[4719:4712];
        layer4[15][23:16] = buffer_data_2[4727:4720];
        layer4[15][31:24] = buffer_data_2[4735:4728];
        layer4[15][39:32] = buffer_data_2[4743:4736];
        layer4[15][47:40] = buffer_data_2[4751:4744];
        layer4[15][55:48] = buffer_data_2[4759:4752];
        layer5[15][7:0] = buffer_data_1[4711:4704];
        layer5[15][15:8] = buffer_data_1[4719:4712];
        layer5[15][23:16] = buffer_data_1[4727:4720];
        layer5[15][31:24] = buffer_data_1[4735:4728];
        layer5[15][39:32] = buffer_data_1[4743:4736];
        layer5[15][47:40] = buffer_data_1[4751:4744];
        layer5[15][55:48] = buffer_data_1[4759:4752];
        layer6[15][7:0] = buffer_data_0[4711:4704];
        layer6[15][15:8] = buffer_data_0[4719:4712];
        layer6[15][23:16] = buffer_data_0[4727:4720];
        layer6[15][31:24] = buffer_data_0[4735:4728];
        layer6[15][39:32] = buffer_data_0[4743:4736];
        layer6[15][47:40] = buffer_data_0[4751:4744];
        layer6[15][55:48] = buffer_data_0[4759:4752];
        layer0[16][7:0] = buffer_data_6[4719:4712];
        layer0[16][15:8] = buffer_data_6[4727:4720];
        layer0[16][23:16] = buffer_data_6[4735:4728];
        layer0[16][31:24] = buffer_data_6[4743:4736];
        layer0[16][39:32] = buffer_data_6[4751:4744];
        layer0[16][47:40] = buffer_data_6[4759:4752];
        layer0[16][55:48] = buffer_data_6[4767:4760];
        layer1[16][7:0] = buffer_data_5[4719:4712];
        layer1[16][15:8] = buffer_data_5[4727:4720];
        layer1[16][23:16] = buffer_data_5[4735:4728];
        layer1[16][31:24] = buffer_data_5[4743:4736];
        layer1[16][39:32] = buffer_data_5[4751:4744];
        layer1[16][47:40] = buffer_data_5[4759:4752];
        layer1[16][55:48] = buffer_data_5[4767:4760];
        layer2[16][7:0] = buffer_data_4[4719:4712];
        layer2[16][15:8] = buffer_data_4[4727:4720];
        layer2[16][23:16] = buffer_data_4[4735:4728];
        layer2[16][31:24] = buffer_data_4[4743:4736];
        layer2[16][39:32] = buffer_data_4[4751:4744];
        layer2[16][47:40] = buffer_data_4[4759:4752];
        layer2[16][55:48] = buffer_data_4[4767:4760];
        layer3[16][7:0] = buffer_data_3[4719:4712];
        layer3[16][15:8] = buffer_data_3[4727:4720];
        layer3[16][23:16] = buffer_data_3[4735:4728];
        layer3[16][31:24] = buffer_data_3[4743:4736];
        layer3[16][39:32] = buffer_data_3[4751:4744];
        layer3[16][47:40] = buffer_data_3[4759:4752];
        layer3[16][55:48] = buffer_data_3[4767:4760];
        layer4[16][7:0] = buffer_data_2[4719:4712];
        layer4[16][15:8] = buffer_data_2[4727:4720];
        layer4[16][23:16] = buffer_data_2[4735:4728];
        layer4[16][31:24] = buffer_data_2[4743:4736];
        layer4[16][39:32] = buffer_data_2[4751:4744];
        layer4[16][47:40] = buffer_data_2[4759:4752];
        layer4[16][55:48] = buffer_data_2[4767:4760];
        layer5[16][7:0] = buffer_data_1[4719:4712];
        layer5[16][15:8] = buffer_data_1[4727:4720];
        layer5[16][23:16] = buffer_data_1[4735:4728];
        layer5[16][31:24] = buffer_data_1[4743:4736];
        layer5[16][39:32] = buffer_data_1[4751:4744];
        layer5[16][47:40] = buffer_data_1[4759:4752];
        layer5[16][55:48] = buffer_data_1[4767:4760];
        layer6[16][7:0] = buffer_data_0[4719:4712];
        layer6[16][15:8] = buffer_data_0[4727:4720];
        layer6[16][23:16] = buffer_data_0[4735:4728];
        layer6[16][31:24] = buffer_data_0[4743:4736];
        layer6[16][39:32] = buffer_data_0[4751:4744];
        layer6[16][47:40] = buffer_data_0[4759:4752];
        layer6[16][55:48] = buffer_data_0[4767:4760];
        layer0[17][7:0] = buffer_data_6[4727:4720];
        layer0[17][15:8] = buffer_data_6[4735:4728];
        layer0[17][23:16] = buffer_data_6[4743:4736];
        layer0[17][31:24] = buffer_data_6[4751:4744];
        layer0[17][39:32] = buffer_data_6[4759:4752];
        layer0[17][47:40] = buffer_data_6[4767:4760];
        layer0[17][55:48] = buffer_data_6[4775:4768];
        layer1[17][7:0] = buffer_data_5[4727:4720];
        layer1[17][15:8] = buffer_data_5[4735:4728];
        layer1[17][23:16] = buffer_data_5[4743:4736];
        layer1[17][31:24] = buffer_data_5[4751:4744];
        layer1[17][39:32] = buffer_data_5[4759:4752];
        layer1[17][47:40] = buffer_data_5[4767:4760];
        layer1[17][55:48] = buffer_data_5[4775:4768];
        layer2[17][7:0] = buffer_data_4[4727:4720];
        layer2[17][15:8] = buffer_data_4[4735:4728];
        layer2[17][23:16] = buffer_data_4[4743:4736];
        layer2[17][31:24] = buffer_data_4[4751:4744];
        layer2[17][39:32] = buffer_data_4[4759:4752];
        layer2[17][47:40] = buffer_data_4[4767:4760];
        layer2[17][55:48] = buffer_data_4[4775:4768];
        layer3[17][7:0] = buffer_data_3[4727:4720];
        layer3[17][15:8] = buffer_data_3[4735:4728];
        layer3[17][23:16] = buffer_data_3[4743:4736];
        layer3[17][31:24] = buffer_data_3[4751:4744];
        layer3[17][39:32] = buffer_data_3[4759:4752];
        layer3[17][47:40] = buffer_data_3[4767:4760];
        layer3[17][55:48] = buffer_data_3[4775:4768];
        layer4[17][7:0] = buffer_data_2[4727:4720];
        layer4[17][15:8] = buffer_data_2[4735:4728];
        layer4[17][23:16] = buffer_data_2[4743:4736];
        layer4[17][31:24] = buffer_data_2[4751:4744];
        layer4[17][39:32] = buffer_data_2[4759:4752];
        layer4[17][47:40] = buffer_data_2[4767:4760];
        layer4[17][55:48] = buffer_data_2[4775:4768];
        layer5[17][7:0] = buffer_data_1[4727:4720];
        layer5[17][15:8] = buffer_data_1[4735:4728];
        layer5[17][23:16] = buffer_data_1[4743:4736];
        layer5[17][31:24] = buffer_data_1[4751:4744];
        layer5[17][39:32] = buffer_data_1[4759:4752];
        layer5[17][47:40] = buffer_data_1[4767:4760];
        layer5[17][55:48] = buffer_data_1[4775:4768];
        layer6[17][7:0] = buffer_data_0[4727:4720];
        layer6[17][15:8] = buffer_data_0[4735:4728];
        layer6[17][23:16] = buffer_data_0[4743:4736];
        layer6[17][31:24] = buffer_data_0[4751:4744];
        layer6[17][39:32] = buffer_data_0[4759:4752];
        layer6[17][47:40] = buffer_data_0[4767:4760];
        layer6[17][55:48] = buffer_data_0[4775:4768];
        layer0[18][7:0] = buffer_data_6[4735:4728];
        layer0[18][15:8] = buffer_data_6[4743:4736];
        layer0[18][23:16] = buffer_data_6[4751:4744];
        layer0[18][31:24] = buffer_data_6[4759:4752];
        layer0[18][39:32] = buffer_data_6[4767:4760];
        layer0[18][47:40] = buffer_data_6[4775:4768];
        layer0[18][55:48] = buffer_data_6[4783:4776];
        layer1[18][7:0] = buffer_data_5[4735:4728];
        layer1[18][15:8] = buffer_data_5[4743:4736];
        layer1[18][23:16] = buffer_data_5[4751:4744];
        layer1[18][31:24] = buffer_data_5[4759:4752];
        layer1[18][39:32] = buffer_data_5[4767:4760];
        layer1[18][47:40] = buffer_data_5[4775:4768];
        layer1[18][55:48] = buffer_data_5[4783:4776];
        layer2[18][7:0] = buffer_data_4[4735:4728];
        layer2[18][15:8] = buffer_data_4[4743:4736];
        layer2[18][23:16] = buffer_data_4[4751:4744];
        layer2[18][31:24] = buffer_data_4[4759:4752];
        layer2[18][39:32] = buffer_data_4[4767:4760];
        layer2[18][47:40] = buffer_data_4[4775:4768];
        layer2[18][55:48] = buffer_data_4[4783:4776];
        layer3[18][7:0] = buffer_data_3[4735:4728];
        layer3[18][15:8] = buffer_data_3[4743:4736];
        layer3[18][23:16] = buffer_data_3[4751:4744];
        layer3[18][31:24] = buffer_data_3[4759:4752];
        layer3[18][39:32] = buffer_data_3[4767:4760];
        layer3[18][47:40] = buffer_data_3[4775:4768];
        layer3[18][55:48] = buffer_data_3[4783:4776];
        layer4[18][7:0] = buffer_data_2[4735:4728];
        layer4[18][15:8] = buffer_data_2[4743:4736];
        layer4[18][23:16] = buffer_data_2[4751:4744];
        layer4[18][31:24] = buffer_data_2[4759:4752];
        layer4[18][39:32] = buffer_data_2[4767:4760];
        layer4[18][47:40] = buffer_data_2[4775:4768];
        layer4[18][55:48] = buffer_data_2[4783:4776];
        layer5[18][7:0] = buffer_data_1[4735:4728];
        layer5[18][15:8] = buffer_data_1[4743:4736];
        layer5[18][23:16] = buffer_data_1[4751:4744];
        layer5[18][31:24] = buffer_data_1[4759:4752];
        layer5[18][39:32] = buffer_data_1[4767:4760];
        layer5[18][47:40] = buffer_data_1[4775:4768];
        layer5[18][55:48] = buffer_data_1[4783:4776];
        layer6[18][7:0] = buffer_data_0[4735:4728];
        layer6[18][15:8] = buffer_data_0[4743:4736];
        layer6[18][23:16] = buffer_data_0[4751:4744];
        layer6[18][31:24] = buffer_data_0[4759:4752];
        layer6[18][39:32] = buffer_data_0[4767:4760];
        layer6[18][47:40] = buffer_data_0[4775:4768];
        layer6[18][55:48] = buffer_data_0[4783:4776];
        layer0[19][7:0] = buffer_data_6[4743:4736];
        layer0[19][15:8] = buffer_data_6[4751:4744];
        layer0[19][23:16] = buffer_data_6[4759:4752];
        layer0[19][31:24] = buffer_data_6[4767:4760];
        layer0[19][39:32] = buffer_data_6[4775:4768];
        layer0[19][47:40] = buffer_data_6[4783:4776];
        layer0[19][55:48] = buffer_data_6[4791:4784];
        layer1[19][7:0] = buffer_data_5[4743:4736];
        layer1[19][15:8] = buffer_data_5[4751:4744];
        layer1[19][23:16] = buffer_data_5[4759:4752];
        layer1[19][31:24] = buffer_data_5[4767:4760];
        layer1[19][39:32] = buffer_data_5[4775:4768];
        layer1[19][47:40] = buffer_data_5[4783:4776];
        layer1[19][55:48] = buffer_data_5[4791:4784];
        layer2[19][7:0] = buffer_data_4[4743:4736];
        layer2[19][15:8] = buffer_data_4[4751:4744];
        layer2[19][23:16] = buffer_data_4[4759:4752];
        layer2[19][31:24] = buffer_data_4[4767:4760];
        layer2[19][39:32] = buffer_data_4[4775:4768];
        layer2[19][47:40] = buffer_data_4[4783:4776];
        layer2[19][55:48] = buffer_data_4[4791:4784];
        layer3[19][7:0] = buffer_data_3[4743:4736];
        layer3[19][15:8] = buffer_data_3[4751:4744];
        layer3[19][23:16] = buffer_data_3[4759:4752];
        layer3[19][31:24] = buffer_data_3[4767:4760];
        layer3[19][39:32] = buffer_data_3[4775:4768];
        layer3[19][47:40] = buffer_data_3[4783:4776];
        layer3[19][55:48] = buffer_data_3[4791:4784];
        layer4[19][7:0] = buffer_data_2[4743:4736];
        layer4[19][15:8] = buffer_data_2[4751:4744];
        layer4[19][23:16] = buffer_data_2[4759:4752];
        layer4[19][31:24] = buffer_data_2[4767:4760];
        layer4[19][39:32] = buffer_data_2[4775:4768];
        layer4[19][47:40] = buffer_data_2[4783:4776];
        layer4[19][55:48] = buffer_data_2[4791:4784];
        layer5[19][7:0] = buffer_data_1[4743:4736];
        layer5[19][15:8] = buffer_data_1[4751:4744];
        layer5[19][23:16] = buffer_data_1[4759:4752];
        layer5[19][31:24] = buffer_data_1[4767:4760];
        layer5[19][39:32] = buffer_data_1[4775:4768];
        layer5[19][47:40] = buffer_data_1[4783:4776];
        layer5[19][55:48] = buffer_data_1[4791:4784];
        layer6[19][7:0] = buffer_data_0[4743:4736];
        layer6[19][15:8] = buffer_data_0[4751:4744];
        layer6[19][23:16] = buffer_data_0[4759:4752];
        layer6[19][31:24] = buffer_data_0[4767:4760];
        layer6[19][39:32] = buffer_data_0[4775:4768];
        layer6[19][47:40] = buffer_data_0[4783:4776];
        layer6[19][55:48] = buffer_data_0[4791:4784];
        layer0[20][7:0] = buffer_data_6[4751:4744];
        layer0[20][15:8] = buffer_data_6[4759:4752];
        layer0[20][23:16] = buffer_data_6[4767:4760];
        layer0[20][31:24] = buffer_data_6[4775:4768];
        layer0[20][39:32] = buffer_data_6[4783:4776];
        layer0[20][47:40] = buffer_data_6[4791:4784];
        layer0[20][55:48] = buffer_data_6[4799:4792];
        layer1[20][7:0] = buffer_data_5[4751:4744];
        layer1[20][15:8] = buffer_data_5[4759:4752];
        layer1[20][23:16] = buffer_data_5[4767:4760];
        layer1[20][31:24] = buffer_data_5[4775:4768];
        layer1[20][39:32] = buffer_data_5[4783:4776];
        layer1[20][47:40] = buffer_data_5[4791:4784];
        layer1[20][55:48] = buffer_data_5[4799:4792];
        layer2[20][7:0] = buffer_data_4[4751:4744];
        layer2[20][15:8] = buffer_data_4[4759:4752];
        layer2[20][23:16] = buffer_data_4[4767:4760];
        layer2[20][31:24] = buffer_data_4[4775:4768];
        layer2[20][39:32] = buffer_data_4[4783:4776];
        layer2[20][47:40] = buffer_data_4[4791:4784];
        layer2[20][55:48] = buffer_data_4[4799:4792];
        layer3[20][7:0] = buffer_data_3[4751:4744];
        layer3[20][15:8] = buffer_data_3[4759:4752];
        layer3[20][23:16] = buffer_data_3[4767:4760];
        layer3[20][31:24] = buffer_data_3[4775:4768];
        layer3[20][39:32] = buffer_data_3[4783:4776];
        layer3[20][47:40] = buffer_data_3[4791:4784];
        layer3[20][55:48] = buffer_data_3[4799:4792];
        layer4[20][7:0] = buffer_data_2[4751:4744];
        layer4[20][15:8] = buffer_data_2[4759:4752];
        layer4[20][23:16] = buffer_data_2[4767:4760];
        layer4[20][31:24] = buffer_data_2[4775:4768];
        layer4[20][39:32] = buffer_data_2[4783:4776];
        layer4[20][47:40] = buffer_data_2[4791:4784];
        layer4[20][55:48] = buffer_data_2[4799:4792];
        layer5[20][7:0] = buffer_data_1[4751:4744];
        layer5[20][15:8] = buffer_data_1[4759:4752];
        layer5[20][23:16] = buffer_data_1[4767:4760];
        layer5[20][31:24] = buffer_data_1[4775:4768];
        layer5[20][39:32] = buffer_data_1[4783:4776];
        layer5[20][47:40] = buffer_data_1[4791:4784];
        layer5[20][55:48] = buffer_data_1[4799:4792];
        layer6[20][7:0] = buffer_data_0[4751:4744];
        layer6[20][15:8] = buffer_data_0[4759:4752];
        layer6[20][23:16] = buffer_data_0[4767:4760];
        layer6[20][31:24] = buffer_data_0[4775:4768];
        layer6[20][39:32] = buffer_data_0[4783:4776];
        layer6[20][47:40] = buffer_data_0[4791:4784];
        layer6[20][55:48] = buffer_data_0[4799:4792];
        layer0[21][7:0] = buffer_data_6[4759:4752];
        layer0[21][15:8] = buffer_data_6[4767:4760];
        layer0[21][23:16] = buffer_data_6[4775:4768];
        layer0[21][31:24] = buffer_data_6[4783:4776];
        layer0[21][39:32] = buffer_data_6[4791:4784];
        layer0[21][47:40] = buffer_data_6[4799:4792];
        layer0[21][55:48] = buffer_data_6[4807:4800];
        layer1[21][7:0] = buffer_data_5[4759:4752];
        layer1[21][15:8] = buffer_data_5[4767:4760];
        layer1[21][23:16] = buffer_data_5[4775:4768];
        layer1[21][31:24] = buffer_data_5[4783:4776];
        layer1[21][39:32] = buffer_data_5[4791:4784];
        layer1[21][47:40] = buffer_data_5[4799:4792];
        layer1[21][55:48] = buffer_data_5[4807:4800];
        layer2[21][7:0] = buffer_data_4[4759:4752];
        layer2[21][15:8] = buffer_data_4[4767:4760];
        layer2[21][23:16] = buffer_data_4[4775:4768];
        layer2[21][31:24] = buffer_data_4[4783:4776];
        layer2[21][39:32] = buffer_data_4[4791:4784];
        layer2[21][47:40] = buffer_data_4[4799:4792];
        layer2[21][55:48] = buffer_data_4[4807:4800];
        layer3[21][7:0] = buffer_data_3[4759:4752];
        layer3[21][15:8] = buffer_data_3[4767:4760];
        layer3[21][23:16] = buffer_data_3[4775:4768];
        layer3[21][31:24] = buffer_data_3[4783:4776];
        layer3[21][39:32] = buffer_data_3[4791:4784];
        layer3[21][47:40] = buffer_data_3[4799:4792];
        layer3[21][55:48] = buffer_data_3[4807:4800];
        layer4[21][7:0] = buffer_data_2[4759:4752];
        layer4[21][15:8] = buffer_data_2[4767:4760];
        layer4[21][23:16] = buffer_data_2[4775:4768];
        layer4[21][31:24] = buffer_data_2[4783:4776];
        layer4[21][39:32] = buffer_data_2[4791:4784];
        layer4[21][47:40] = buffer_data_2[4799:4792];
        layer4[21][55:48] = buffer_data_2[4807:4800];
        layer5[21][7:0] = buffer_data_1[4759:4752];
        layer5[21][15:8] = buffer_data_1[4767:4760];
        layer5[21][23:16] = buffer_data_1[4775:4768];
        layer5[21][31:24] = buffer_data_1[4783:4776];
        layer5[21][39:32] = buffer_data_1[4791:4784];
        layer5[21][47:40] = buffer_data_1[4799:4792];
        layer5[21][55:48] = buffer_data_1[4807:4800];
        layer6[21][7:0] = buffer_data_0[4759:4752];
        layer6[21][15:8] = buffer_data_0[4767:4760];
        layer6[21][23:16] = buffer_data_0[4775:4768];
        layer6[21][31:24] = buffer_data_0[4783:4776];
        layer6[21][39:32] = buffer_data_0[4791:4784];
        layer6[21][47:40] = buffer_data_0[4799:4792];
        layer6[21][55:48] = buffer_data_0[4807:4800];
        layer0[22][7:0] = buffer_data_6[4767:4760];
        layer0[22][15:8] = buffer_data_6[4775:4768];
        layer0[22][23:16] = buffer_data_6[4783:4776];
        layer0[22][31:24] = buffer_data_6[4791:4784];
        layer0[22][39:32] = buffer_data_6[4799:4792];
        layer0[22][47:40] = buffer_data_6[4807:4800];
        layer0[22][55:48] = buffer_data_6[4815:4808];
        layer1[22][7:0] = buffer_data_5[4767:4760];
        layer1[22][15:8] = buffer_data_5[4775:4768];
        layer1[22][23:16] = buffer_data_5[4783:4776];
        layer1[22][31:24] = buffer_data_5[4791:4784];
        layer1[22][39:32] = buffer_data_5[4799:4792];
        layer1[22][47:40] = buffer_data_5[4807:4800];
        layer1[22][55:48] = buffer_data_5[4815:4808];
        layer2[22][7:0] = buffer_data_4[4767:4760];
        layer2[22][15:8] = buffer_data_4[4775:4768];
        layer2[22][23:16] = buffer_data_4[4783:4776];
        layer2[22][31:24] = buffer_data_4[4791:4784];
        layer2[22][39:32] = buffer_data_4[4799:4792];
        layer2[22][47:40] = buffer_data_4[4807:4800];
        layer2[22][55:48] = buffer_data_4[4815:4808];
        layer3[22][7:0] = buffer_data_3[4767:4760];
        layer3[22][15:8] = buffer_data_3[4775:4768];
        layer3[22][23:16] = buffer_data_3[4783:4776];
        layer3[22][31:24] = buffer_data_3[4791:4784];
        layer3[22][39:32] = buffer_data_3[4799:4792];
        layer3[22][47:40] = buffer_data_3[4807:4800];
        layer3[22][55:48] = buffer_data_3[4815:4808];
        layer4[22][7:0] = buffer_data_2[4767:4760];
        layer4[22][15:8] = buffer_data_2[4775:4768];
        layer4[22][23:16] = buffer_data_2[4783:4776];
        layer4[22][31:24] = buffer_data_2[4791:4784];
        layer4[22][39:32] = buffer_data_2[4799:4792];
        layer4[22][47:40] = buffer_data_2[4807:4800];
        layer4[22][55:48] = buffer_data_2[4815:4808];
        layer5[22][7:0] = buffer_data_1[4767:4760];
        layer5[22][15:8] = buffer_data_1[4775:4768];
        layer5[22][23:16] = buffer_data_1[4783:4776];
        layer5[22][31:24] = buffer_data_1[4791:4784];
        layer5[22][39:32] = buffer_data_1[4799:4792];
        layer5[22][47:40] = buffer_data_1[4807:4800];
        layer5[22][55:48] = buffer_data_1[4815:4808];
        layer6[22][7:0] = buffer_data_0[4767:4760];
        layer6[22][15:8] = buffer_data_0[4775:4768];
        layer6[22][23:16] = buffer_data_0[4783:4776];
        layer6[22][31:24] = buffer_data_0[4791:4784];
        layer6[22][39:32] = buffer_data_0[4799:4792];
        layer6[22][47:40] = buffer_data_0[4807:4800];
        layer6[22][55:48] = buffer_data_0[4815:4808];
        layer0[23][7:0] = buffer_data_6[4775:4768];
        layer0[23][15:8] = buffer_data_6[4783:4776];
        layer0[23][23:16] = buffer_data_6[4791:4784];
        layer0[23][31:24] = buffer_data_6[4799:4792];
        layer0[23][39:32] = buffer_data_6[4807:4800];
        layer0[23][47:40] = buffer_data_6[4815:4808];
        layer0[23][55:48] = buffer_data_6[4823:4816];
        layer1[23][7:0] = buffer_data_5[4775:4768];
        layer1[23][15:8] = buffer_data_5[4783:4776];
        layer1[23][23:16] = buffer_data_5[4791:4784];
        layer1[23][31:24] = buffer_data_5[4799:4792];
        layer1[23][39:32] = buffer_data_5[4807:4800];
        layer1[23][47:40] = buffer_data_5[4815:4808];
        layer1[23][55:48] = buffer_data_5[4823:4816];
        layer2[23][7:0] = buffer_data_4[4775:4768];
        layer2[23][15:8] = buffer_data_4[4783:4776];
        layer2[23][23:16] = buffer_data_4[4791:4784];
        layer2[23][31:24] = buffer_data_4[4799:4792];
        layer2[23][39:32] = buffer_data_4[4807:4800];
        layer2[23][47:40] = buffer_data_4[4815:4808];
        layer2[23][55:48] = buffer_data_4[4823:4816];
        layer3[23][7:0] = buffer_data_3[4775:4768];
        layer3[23][15:8] = buffer_data_3[4783:4776];
        layer3[23][23:16] = buffer_data_3[4791:4784];
        layer3[23][31:24] = buffer_data_3[4799:4792];
        layer3[23][39:32] = buffer_data_3[4807:4800];
        layer3[23][47:40] = buffer_data_3[4815:4808];
        layer3[23][55:48] = buffer_data_3[4823:4816];
        layer4[23][7:0] = buffer_data_2[4775:4768];
        layer4[23][15:8] = buffer_data_2[4783:4776];
        layer4[23][23:16] = buffer_data_2[4791:4784];
        layer4[23][31:24] = buffer_data_2[4799:4792];
        layer4[23][39:32] = buffer_data_2[4807:4800];
        layer4[23][47:40] = buffer_data_2[4815:4808];
        layer4[23][55:48] = buffer_data_2[4823:4816];
        layer5[23][7:0] = buffer_data_1[4775:4768];
        layer5[23][15:8] = buffer_data_1[4783:4776];
        layer5[23][23:16] = buffer_data_1[4791:4784];
        layer5[23][31:24] = buffer_data_1[4799:4792];
        layer5[23][39:32] = buffer_data_1[4807:4800];
        layer5[23][47:40] = buffer_data_1[4815:4808];
        layer5[23][55:48] = buffer_data_1[4823:4816];
        layer6[23][7:0] = buffer_data_0[4775:4768];
        layer6[23][15:8] = buffer_data_0[4783:4776];
        layer6[23][23:16] = buffer_data_0[4791:4784];
        layer6[23][31:24] = buffer_data_0[4799:4792];
        layer6[23][39:32] = buffer_data_0[4807:4800];
        layer6[23][47:40] = buffer_data_0[4815:4808];
        layer6[23][55:48] = buffer_data_0[4823:4816];
        layer0[24][7:0] = buffer_data_6[4783:4776];
        layer0[24][15:8] = buffer_data_6[4791:4784];
        layer0[24][23:16] = buffer_data_6[4799:4792];
        layer0[24][31:24] = buffer_data_6[4807:4800];
        layer0[24][39:32] = buffer_data_6[4815:4808];
        layer0[24][47:40] = buffer_data_6[4823:4816];
        layer0[24][55:48] = buffer_data_6[4831:4824];
        layer1[24][7:0] = buffer_data_5[4783:4776];
        layer1[24][15:8] = buffer_data_5[4791:4784];
        layer1[24][23:16] = buffer_data_5[4799:4792];
        layer1[24][31:24] = buffer_data_5[4807:4800];
        layer1[24][39:32] = buffer_data_5[4815:4808];
        layer1[24][47:40] = buffer_data_5[4823:4816];
        layer1[24][55:48] = buffer_data_5[4831:4824];
        layer2[24][7:0] = buffer_data_4[4783:4776];
        layer2[24][15:8] = buffer_data_4[4791:4784];
        layer2[24][23:16] = buffer_data_4[4799:4792];
        layer2[24][31:24] = buffer_data_4[4807:4800];
        layer2[24][39:32] = buffer_data_4[4815:4808];
        layer2[24][47:40] = buffer_data_4[4823:4816];
        layer2[24][55:48] = buffer_data_4[4831:4824];
        layer3[24][7:0] = buffer_data_3[4783:4776];
        layer3[24][15:8] = buffer_data_3[4791:4784];
        layer3[24][23:16] = buffer_data_3[4799:4792];
        layer3[24][31:24] = buffer_data_3[4807:4800];
        layer3[24][39:32] = buffer_data_3[4815:4808];
        layer3[24][47:40] = buffer_data_3[4823:4816];
        layer3[24][55:48] = buffer_data_3[4831:4824];
        layer4[24][7:0] = buffer_data_2[4783:4776];
        layer4[24][15:8] = buffer_data_2[4791:4784];
        layer4[24][23:16] = buffer_data_2[4799:4792];
        layer4[24][31:24] = buffer_data_2[4807:4800];
        layer4[24][39:32] = buffer_data_2[4815:4808];
        layer4[24][47:40] = buffer_data_2[4823:4816];
        layer4[24][55:48] = buffer_data_2[4831:4824];
        layer5[24][7:0] = buffer_data_1[4783:4776];
        layer5[24][15:8] = buffer_data_1[4791:4784];
        layer5[24][23:16] = buffer_data_1[4799:4792];
        layer5[24][31:24] = buffer_data_1[4807:4800];
        layer5[24][39:32] = buffer_data_1[4815:4808];
        layer5[24][47:40] = buffer_data_1[4823:4816];
        layer5[24][55:48] = buffer_data_1[4831:4824];
        layer6[24][7:0] = buffer_data_0[4783:4776];
        layer6[24][15:8] = buffer_data_0[4791:4784];
        layer6[24][23:16] = buffer_data_0[4799:4792];
        layer6[24][31:24] = buffer_data_0[4807:4800];
        layer6[24][39:32] = buffer_data_0[4815:4808];
        layer6[24][47:40] = buffer_data_0[4823:4816];
        layer6[24][55:48] = buffer_data_0[4831:4824];
        layer0[25][7:0] = buffer_data_6[4791:4784];
        layer0[25][15:8] = buffer_data_6[4799:4792];
        layer0[25][23:16] = buffer_data_6[4807:4800];
        layer0[25][31:24] = buffer_data_6[4815:4808];
        layer0[25][39:32] = buffer_data_6[4823:4816];
        layer0[25][47:40] = buffer_data_6[4831:4824];
        layer0[25][55:48] = buffer_data_6[4839:4832];
        layer1[25][7:0] = buffer_data_5[4791:4784];
        layer1[25][15:8] = buffer_data_5[4799:4792];
        layer1[25][23:16] = buffer_data_5[4807:4800];
        layer1[25][31:24] = buffer_data_5[4815:4808];
        layer1[25][39:32] = buffer_data_5[4823:4816];
        layer1[25][47:40] = buffer_data_5[4831:4824];
        layer1[25][55:48] = buffer_data_5[4839:4832];
        layer2[25][7:0] = buffer_data_4[4791:4784];
        layer2[25][15:8] = buffer_data_4[4799:4792];
        layer2[25][23:16] = buffer_data_4[4807:4800];
        layer2[25][31:24] = buffer_data_4[4815:4808];
        layer2[25][39:32] = buffer_data_4[4823:4816];
        layer2[25][47:40] = buffer_data_4[4831:4824];
        layer2[25][55:48] = buffer_data_4[4839:4832];
        layer3[25][7:0] = buffer_data_3[4791:4784];
        layer3[25][15:8] = buffer_data_3[4799:4792];
        layer3[25][23:16] = buffer_data_3[4807:4800];
        layer3[25][31:24] = buffer_data_3[4815:4808];
        layer3[25][39:32] = buffer_data_3[4823:4816];
        layer3[25][47:40] = buffer_data_3[4831:4824];
        layer3[25][55:48] = buffer_data_3[4839:4832];
        layer4[25][7:0] = buffer_data_2[4791:4784];
        layer4[25][15:8] = buffer_data_2[4799:4792];
        layer4[25][23:16] = buffer_data_2[4807:4800];
        layer4[25][31:24] = buffer_data_2[4815:4808];
        layer4[25][39:32] = buffer_data_2[4823:4816];
        layer4[25][47:40] = buffer_data_2[4831:4824];
        layer4[25][55:48] = buffer_data_2[4839:4832];
        layer5[25][7:0] = buffer_data_1[4791:4784];
        layer5[25][15:8] = buffer_data_1[4799:4792];
        layer5[25][23:16] = buffer_data_1[4807:4800];
        layer5[25][31:24] = buffer_data_1[4815:4808];
        layer5[25][39:32] = buffer_data_1[4823:4816];
        layer5[25][47:40] = buffer_data_1[4831:4824];
        layer5[25][55:48] = buffer_data_1[4839:4832];
        layer6[25][7:0] = buffer_data_0[4791:4784];
        layer6[25][15:8] = buffer_data_0[4799:4792];
        layer6[25][23:16] = buffer_data_0[4807:4800];
        layer6[25][31:24] = buffer_data_0[4815:4808];
        layer6[25][39:32] = buffer_data_0[4823:4816];
        layer6[25][47:40] = buffer_data_0[4831:4824];
        layer6[25][55:48] = buffer_data_0[4839:4832];
        layer0[26][7:0] = buffer_data_6[4799:4792];
        layer0[26][15:8] = buffer_data_6[4807:4800];
        layer0[26][23:16] = buffer_data_6[4815:4808];
        layer0[26][31:24] = buffer_data_6[4823:4816];
        layer0[26][39:32] = buffer_data_6[4831:4824];
        layer0[26][47:40] = buffer_data_6[4839:4832];
        layer0[26][55:48] = buffer_data_6[4847:4840];
        layer1[26][7:0] = buffer_data_5[4799:4792];
        layer1[26][15:8] = buffer_data_5[4807:4800];
        layer1[26][23:16] = buffer_data_5[4815:4808];
        layer1[26][31:24] = buffer_data_5[4823:4816];
        layer1[26][39:32] = buffer_data_5[4831:4824];
        layer1[26][47:40] = buffer_data_5[4839:4832];
        layer1[26][55:48] = buffer_data_5[4847:4840];
        layer2[26][7:0] = buffer_data_4[4799:4792];
        layer2[26][15:8] = buffer_data_4[4807:4800];
        layer2[26][23:16] = buffer_data_4[4815:4808];
        layer2[26][31:24] = buffer_data_4[4823:4816];
        layer2[26][39:32] = buffer_data_4[4831:4824];
        layer2[26][47:40] = buffer_data_4[4839:4832];
        layer2[26][55:48] = buffer_data_4[4847:4840];
        layer3[26][7:0] = buffer_data_3[4799:4792];
        layer3[26][15:8] = buffer_data_3[4807:4800];
        layer3[26][23:16] = buffer_data_3[4815:4808];
        layer3[26][31:24] = buffer_data_3[4823:4816];
        layer3[26][39:32] = buffer_data_3[4831:4824];
        layer3[26][47:40] = buffer_data_3[4839:4832];
        layer3[26][55:48] = buffer_data_3[4847:4840];
        layer4[26][7:0] = buffer_data_2[4799:4792];
        layer4[26][15:8] = buffer_data_2[4807:4800];
        layer4[26][23:16] = buffer_data_2[4815:4808];
        layer4[26][31:24] = buffer_data_2[4823:4816];
        layer4[26][39:32] = buffer_data_2[4831:4824];
        layer4[26][47:40] = buffer_data_2[4839:4832];
        layer4[26][55:48] = buffer_data_2[4847:4840];
        layer5[26][7:0] = buffer_data_1[4799:4792];
        layer5[26][15:8] = buffer_data_1[4807:4800];
        layer5[26][23:16] = buffer_data_1[4815:4808];
        layer5[26][31:24] = buffer_data_1[4823:4816];
        layer5[26][39:32] = buffer_data_1[4831:4824];
        layer5[26][47:40] = buffer_data_1[4839:4832];
        layer5[26][55:48] = buffer_data_1[4847:4840];
        layer6[26][7:0] = buffer_data_0[4799:4792];
        layer6[26][15:8] = buffer_data_0[4807:4800];
        layer6[26][23:16] = buffer_data_0[4815:4808];
        layer6[26][31:24] = buffer_data_0[4823:4816];
        layer6[26][39:32] = buffer_data_0[4831:4824];
        layer6[26][47:40] = buffer_data_0[4839:4832];
        layer6[26][55:48] = buffer_data_0[4847:4840];
        layer0[27][7:0] = buffer_data_6[4807:4800];
        layer0[27][15:8] = buffer_data_6[4815:4808];
        layer0[27][23:16] = buffer_data_6[4823:4816];
        layer0[27][31:24] = buffer_data_6[4831:4824];
        layer0[27][39:32] = buffer_data_6[4839:4832];
        layer0[27][47:40] = buffer_data_6[4847:4840];
        layer0[27][55:48] = buffer_data_6[4855:4848];
        layer1[27][7:0] = buffer_data_5[4807:4800];
        layer1[27][15:8] = buffer_data_5[4815:4808];
        layer1[27][23:16] = buffer_data_5[4823:4816];
        layer1[27][31:24] = buffer_data_5[4831:4824];
        layer1[27][39:32] = buffer_data_5[4839:4832];
        layer1[27][47:40] = buffer_data_5[4847:4840];
        layer1[27][55:48] = buffer_data_5[4855:4848];
        layer2[27][7:0] = buffer_data_4[4807:4800];
        layer2[27][15:8] = buffer_data_4[4815:4808];
        layer2[27][23:16] = buffer_data_4[4823:4816];
        layer2[27][31:24] = buffer_data_4[4831:4824];
        layer2[27][39:32] = buffer_data_4[4839:4832];
        layer2[27][47:40] = buffer_data_4[4847:4840];
        layer2[27][55:48] = buffer_data_4[4855:4848];
        layer3[27][7:0] = buffer_data_3[4807:4800];
        layer3[27][15:8] = buffer_data_3[4815:4808];
        layer3[27][23:16] = buffer_data_3[4823:4816];
        layer3[27][31:24] = buffer_data_3[4831:4824];
        layer3[27][39:32] = buffer_data_3[4839:4832];
        layer3[27][47:40] = buffer_data_3[4847:4840];
        layer3[27][55:48] = buffer_data_3[4855:4848];
        layer4[27][7:0] = buffer_data_2[4807:4800];
        layer4[27][15:8] = buffer_data_2[4815:4808];
        layer4[27][23:16] = buffer_data_2[4823:4816];
        layer4[27][31:24] = buffer_data_2[4831:4824];
        layer4[27][39:32] = buffer_data_2[4839:4832];
        layer4[27][47:40] = buffer_data_2[4847:4840];
        layer4[27][55:48] = buffer_data_2[4855:4848];
        layer5[27][7:0] = buffer_data_1[4807:4800];
        layer5[27][15:8] = buffer_data_1[4815:4808];
        layer5[27][23:16] = buffer_data_1[4823:4816];
        layer5[27][31:24] = buffer_data_1[4831:4824];
        layer5[27][39:32] = buffer_data_1[4839:4832];
        layer5[27][47:40] = buffer_data_1[4847:4840];
        layer5[27][55:48] = buffer_data_1[4855:4848];
        layer6[27][7:0] = buffer_data_0[4807:4800];
        layer6[27][15:8] = buffer_data_0[4815:4808];
        layer6[27][23:16] = buffer_data_0[4823:4816];
        layer6[27][31:24] = buffer_data_0[4831:4824];
        layer6[27][39:32] = buffer_data_0[4839:4832];
        layer6[27][47:40] = buffer_data_0[4847:4840];
        layer6[27][55:48] = buffer_data_0[4855:4848];
        layer0[28][7:0] = buffer_data_6[4815:4808];
        layer0[28][15:8] = buffer_data_6[4823:4816];
        layer0[28][23:16] = buffer_data_6[4831:4824];
        layer0[28][31:24] = buffer_data_6[4839:4832];
        layer0[28][39:32] = buffer_data_6[4847:4840];
        layer0[28][47:40] = buffer_data_6[4855:4848];
        layer0[28][55:48] = buffer_data_6[4863:4856];
        layer1[28][7:0] = buffer_data_5[4815:4808];
        layer1[28][15:8] = buffer_data_5[4823:4816];
        layer1[28][23:16] = buffer_data_5[4831:4824];
        layer1[28][31:24] = buffer_data_5[4839:4832];
        layer1[28][39:32] = buffer_data_5[4847:4840];
        layer1[28][47:40] = buffer_data_5[4855:4848];
        layer1[28][55:48] = buffer_data_5[4863:4856];
        layer2[28][7:0] = buffer_data_4[4815:4808];
        layer2[28][15:8] = buffer_data_4[4823:4816];
        layer2[28][23:16] = buffer_data_4[4831:4824];
        layer2[28][31:24] = buffer_data_4[4839:4832];
        layer2[28][39:32] = buffer_data_4[4847:4840];
        layer2[28][47:40] = buffer_data_4[4855:4848];
        layer2[28][55:48] = buffer_data_4[4863:4856];
        layer3[28][7:0] = buffer_data_3[4815:4808];
        layer3[28][15:8] = buffer_data_3[4823:4816];
        layer3[28][23:16] = buffer_data_3[4831:4824];
        layer3[28][31:24] = buffer_data_3[4839:4832];
        layer3[28][39:32] = buffer_data_3[4847:4840];
        layer3[28][47:40] = buffer_data_3[4855:4848];
        layer3[28][55:48] = buffer_data_3[4863:4856];
        layer4[28][7:0] = buffer_data_2[4815:4808];
        layer4[28][15:8] = buffer_data_2[4823:4816];
        layer4[28][23:16] = buffer_data_2[4831:4824];
        layer4[28][31:24] = buffer_data_2[4839:4832];
        layer4[28][39:32] = buffer_data_2[4847:4840];
        layer4[28][47:40] = buffer_data_2[4855:4848];
        layer4[28][55:48] = buffer_data_2[4863:4856];
        layer5[28][7:0] = buffer_data_1[4815:4808];
        layer5[28][15:8] = buffer_data_1[4823:4816];
        layer5[28][23:16] = buffer_data_1[4831:4824];
        layer5[28][31:24] = buffer_data_1[4839:4832];
        layer5[28][39:32] = buffer_data_1[4847:4840];
        layer5[28][47:40] = buffer_data_1[4855:4848];
        layer5[28][55:48] = buffer_data_1[4863:4856];
        layer6[28][7:0] = buffer_data_0[4815:4808];
        layer6[28][15:8] = buffer_data_0[4823:4816];
        layer6[28][23:16] = buffer_data_0[4831:4824];
        layer6[28][31:24] = buffer_data_0[4839:4832];
        layer6[28][39:32] = buffer_data_0[4847:4840];
        layer6[28][47:40] = buffer_data_0[4855:4848];
        layer6[28][55:48] = buffer_data_0[4863:4856];
        layer0[29][7:0] = buffer_data_6[4823:4816];
        layer0[29][15:8] = buffer_data_6[4831:4824];
        layer0[29][23:16] = buffer_data_6[4839:4832];
        layer0[29][31:24] = buffer_data_6[4847:4840];
        layer0[29][39:32] = buffer_data_6[4855:4848];
        layer0[29][47:40] = buffer_data_6[4863:4856];
        layer0[29][55:48] = buffer_data_6[4871:4864];
        layer1[29][7:0] = buffer_data_5[4823:4816];
        layer1[29][15:8] = buffer_data_5[4831:4824];
        layer1[29][23:16] = buffer_data_5[4839:4832];
        layer1[29][31:24] = buffer_data_5[4847:4840];
        layer1[29][39:32] = buffer_data_5[4855:4848];
        layer1[29][47:40] = buffer_data_5[4863:4856];
        layer1[29][55:48] = buffer_data_5[4871:4864];
        layer2[29][7:0] = buffer_data_4[4823:4816];
        layer2[29][15:8] = buffer_data_4[4831:4824];
        layer2[29][23:16] = buffer_data_4[4839:4832];
        layer2[29][31:24] = buffer_data_4[4847:4840];
        layer2[29][39:32] = buffer_data_4[4855:4848];
        layer2[29][47:40] = buffer_data_4[4863:4856];
        layer2[29][55:48] = buffer_data_4[4871:4864];
        layer3[29][7:0] = buffer_data_3[4823:4816];
        layer3[29][15:8] = buffer_data_3[4831:4824];
        layer3[29][23:16] = buffer_data_3[4839:4832];
        layer3[29][31:24] = buffer_data_3[4847:4840];
        layer3[29][39:32] = buffer_data_3[4855:4848];
        layer3[29][47:40] = buffer_data_3[4863:4856];
        layer3[29][55:48] = buffer_data_3[4871:4864];
        layer4[29][7:0] = buffer_data_2[4823:4816];
        layer4[29][15:8] = buffer_data_2[4831:4824];
        layer4[29][23:16] = buffer_data_2[4839:4832];
        layer4[29][31:24] = buffer_data_2[4847:4840];
        layer4[29][39:32] = buffer_data_2[4855:4848];
        layer4[29][47:40] = buffer_data_2[4863:4856];
        layer4[29][55:48] = buffer_data_2[4871:4864];
        layer5[29][7:0] = buffer_data_1[4823:4816];
        layer5[29][15:8] = buffer_data_1[4831:4824];
        layer5[29][23:16] = buffer_data_1[4839:4832];
        layer5[29][31:24] = buffer_data_1[4847:4840];
        layer5[29][39:32] = buffer_data_1[4855:4848];
        layer5[29][47:40] = buffer_data_1[4863:4856];
        layer5[29][55:48] = buffer_data_1[4871:4864];
        layer6[29][7:0] = buffer_data_0[4823:4816];
        layer6[29][15:8] = buffer_data_0[4831:4824];
        layer6[29][23:16] = buffer_data_0[4839:4832];
        layer6[29][31:24] = buffer_data_0[4847:4840];
        layer6[29][39:32] = buffer_data_0[4855:4848];
        layer6[29][47:40] = buffer_data_0[4863:4856];
        layer6[29][55:48] = buffer_data_0[4871:4864];
        layer0[30][7:0] = buffer_data_6[4831:4824];
        layer0[30][15:8] = buffer_data_6[4839:4832];
        layer0[30][23:16] = buffer_data_6[4847:4840];
        layer0[30][31:24] = buffer_data_6[4855:4848];
        layer0[30][39:32] = buffer_data_6[4863:4856];
        layer0[30][47:40] = buffer_data_6[4871:4864];
        layer0[30][55:48] = buffer_data_6[4879:4872];
        layer1[30][7:0] = buffer_data_5[4831:4824];
        layer1[30][15:8] = buffer_data_5[4839:4832];
        layer1[30][23:16] = buffer_data_5[4847:4840];
        layer1[30][31:24] = buffer_data_5[4855:4848];
        layer1[30][39:32] = buffer_data_5[4863:4856];
        layer1[30][47:40] = buffer_data_5[4871:4864];
        layer1[30][55:48] = buffer_data_5[4879:4872];
        layer2[30][7:0] = buffer_data_4[4831:4824];
        layer2[30][15:8] = buffer_data_4[4839:4832];
        layer2[30][23:16] = buffer_data_4[4847:4840];
        layer2[30][31:24] = buffer_data_4[4855:4848];
        layer2[30][39:32] = buffer_data_4[4863:4856];
        layer2[30][47:40] = buffer_data_4[4871:4864];
        layer2[30][55:48] = buffer_data_4[4879:4872];
        layer3[30][7:0] = buffer_data_3[4831:4824];
        layer3[30][15:8] = buffer_data_3[4839:4832];
        layer3[30][23:16] = buffer_data_3[4847:4840];
        layer3[30][31:24] = buffer_data_3[4855:4848];
        layer3[30][39:32] = buffer_data_3[4863:4856];
        layer3[30][47:40] = buffer_data_3[4871:4864];
        layer3[30][55:48] = buffer_data_3[4879:4872];
        layer4[30][7:0] = buffer_data_2[4831:4824];
        layer4[30][15:8] = buffer_data_2[4839:4832];
        layer4[30][23:16] = buffer_data_2[4847:4840];
        layer4[30][31:24] = buffer_data_2[4855:4848];
        layer4[30][39:32] = buffer_data_2[4863:4856];
        layer4[30][47:40] = buffer_data_2[4871:4864];
        layer4[30][55:48] = buffer_data_2[4879:4872];
        layer5[30][7:0] = buffer_data_1[4831:4824];
        layer5[30][15:8] = buffer_data_1[4839:4832];
        layer5[30][23:16] = buffer_data_1[4847:4840];
        layer5[30][31:24] = buffer_data_1[4855:4848];
        layer5[30][39:32] = buffer_data_1[4863:4856];
        layer5[30][47:40] = buffer_data_1[4871:4864];
        layer5[30][55:48] = buffer_data_1[4879:4872];
        layer6[30][7:0] = buffer_data_0[4831:4824];
        layer6[30][15:8] = buffer_data_0[4839:4832];
        layer6[30][23:16] = buffer_data_0[4847:4840];
        layer6[30][31:24] = buffer_data_0[4855:4848];
        layer6[30][39:32] = buffer_data_0[4863:4856];
        layer6[30][47:40] = buffer_data_0[4871:4864];
        layer6[30][55:48] = buffer_data_0[4879:4872];
        layer0[31][7:0] = buffer_data_6[4839:4832];
        layer0[31][15:8] = buffer_data_6[4847:4840];
        layer0[31][23:16] = buffer_data_6[4855:4848];
        layer0[31][31:24] = buffer_data_6[4863:4856];
        layer0[31][39:32] = buffer_data_6[4871:4864];
        layer0[31][47:40] = buffer_data_6[4879:4872];
        layer0[31][55:48] = buffer_data_6[4887:4880];
        layer1[31][7:0] = buffer_data_5[4839:4832];
        layer1[31][15:8] = buffer_data_5[4847:4840];
        layer1[31][23:16] = buffer_data_5[4855:4848];
        layer1[31][31:24] = buffer_data_5[4863:4856];
        layer1[31][39:32] = buffer_data_5[4871:4864];
        layer1[31][47:40] = buffer_data_5[4879:4872];
        layer1[31][55:48] = buffer_data_5[4887:4880];
        layer2[31][7:0] = buffer_data_4[4839:4832];
        layer2[31][15:8] = buffer_data_4[4847:4840];
        layer2[31][23:16] = buffer_data_4[4855:4848];
        layer2[31][31:24] = buffer_data_4[4863:4856];
        layer2[31][39:32] = buffer_data_4[4871:4864];
        layer2[31][47:40] = buffer_data_4[4879:4872];
        layer2[31][55:48] = buffer_data_4[4887:4880];
        layer3[31][7:0] = buffer_data_3[4839:4832];
        layer3[31][15:8] = buffer_data_3[4847:4840];
        layer3[31][23:16] = buffer_data_3[4855:4848];
        layer3[31][31:24] = buffer_data_3[4863:4856];
        layer3[31][39:32] = buffer_data_3[4871:4864];
        layer3[31][47:40] = buffer_data_3[4879:4872];
        layer3[31][55:48] = buffer_data_3[4887:4880];
        layer4[31][7:0] = buffer_data_2[4839:4832];
        layer4[31][15:8] = buffer_data_2[4847:4840];
        layer4[31][23:16] = buffer_data_2[4855:4848];
        layer4[31][31:24] = buffer_data_2[4863:4856];
        layer4[31][39:32] = buffer_data_2[4871:4864];
        layer4[31][47:40] = buffer_data_2[4879:4872];
        layer4[31][55:48] = buffer_data_2[4887:4880];
        layer5[31][7:0] = buffer_data_1[4839:4832];
        layer5[31][15:8] = buffer_data_1[4847:4840];
        layer5[31][23:16] = buffer_data_1[4855:4848];
        layer5[31][31:24] = buffer_data_1[4863:4856];
        layer5[31][39:32] = buffer_data_1[4871:4864];
        layer5[31][47:40] = buffer_data_1[4879:4872];
        layer5[31][55:48] = buffer_data_1[4887:4880];
        layer6[31][7:0] = buffer_data_0[4839:4832];
        layer6[31][15:8] = buffer_data_0[4847:4840];
        layer6[31][23:16] = buffer_data_0[4855:4848];
        layer6[31][31:24] = buffer_data_0[4863:4856];
        layer6[31][39:32] = buffer_data_0[4871:4864];
        layer6[31][47:40] = buffer_data_0[4879:4872];
        layer6[31][55:48] = buffer_data_0[4887:4880];
        layer0[32][7:0] = buffer_data_6[4847:4840];
        layer0[32][15:8] = buffer_data_6[4855:4848];
        layer0[32][23:16] = buffer_data_6[4863:4856];
        layer0[32][31:24] = buffer_data_6[4871:4864];
        layer0[32][39:32] = buffer_data_6[4879:4872];
        layer0[32][47:40] = buffer_data_6[4887:4880];
        layer0[32][55:48] = buffer_data_6[4895:4888];
        layer1[32][7:0] = buffer_data_5[4847:4840];
        layer1[32][15:8] = buffer_data_5[4855:4848];
        layer1[32][23:16] = buffer_data_5[4863:4856];
        layer1[32][31:24] = buffer_data_5[4871:4864];
        layer1[32][39:32] = buffer_data_5[4879:4872];
        layer1[32][47:40] = buffer_data_5[4887:4880];
        layer1[32][55:48] = buffer_data_5[4895:4888];
        layer2[32][7:0] = buffer_data_4[4847:4840];
        layer2[32][15:8] = buffer_data_4[4855:4848];
        layer2[32][23:16] = buffer_data_4[4863:4856];
        layer2[32][31:24] = buffer_data_4[4871:4864];
        layer2[32][39:32] = buffer_data_4[4879:4872];
        layer2[32][47:40] = buffer_data_4[4887:4880];
        layer2[32][55:48] = buffer_data_4[4895:4888];
        layer3[32][7:0] = buffer_data_3[4847:4840];
        layer3[32][15:8] = buffer_data_3[4855:4848];
        layer3[32][23:16] = buffer_data_3[4863:4856];
        layer3[32][31:24] = buffer_data_3[4871:4864];
        layer3[32][39:32] = buffer_data_3[4879:4872];
        layer3[32][47:40] = buffer_data_3[4887:4880];
        layer3[32][55:48] = buffer_data_3[4895:4888];
        layer4[32][7:0] = buffer_data_2[4847:4840];
        layer4[32][15:8] = buffer_data_2[4855:4848];
        layer4[32][23:16] = buffer_data_2[4863:4856];
        layer4[32][31:24] = buffer_data_2[4871:4864];
        layer4[32][39:32] = buffer_data_2[4879:4872];
        layer4[32][47:40] = buffer_data_2[4887:4880];
        layer4[32][55:48] = buffer_data_2[4895:4888];
        layer5[32][7:0] = buffer_data_1[4847:4840];
        layer5[32][15:8] = buffer_data_1[4855:4848];
        layer5[32][23:16] = buffer_data_1[4863:4856];
        layer5[32][31:24] = buffer_data_1[4871:4864];
        layer5[32][39:32] = buffer_data_1[4879:4872];
        layer5[32][47:40] = buffer_data_1[4887:4880];
        layer5[32][55:48] = buffer_data_1[4895:4888];
        layer6[32][7:0] = buffer_data_0[4847:4840];
        layer6[32][15:8] = buffer_data_0[4855:4848];
        layer6[32][23:16] = buffer_data_0[4863:4856];
        layer6[32][31:24] = buffer_data_0[4871:4864];
        layer6[32][39:32] = buffer_data_0[4879:4872];
        layer6[32][47:40] = buffer_data_0[4887:4880];
        layer6[32][55:48] = buffer_data_0[4895:4888];
        layer0[33][7:0] = buffer_data_6[4855:4848];
        layer0[33][15:8] = buffer_data_6[4863:4856];
        layer0[33][23:16] = buffer_data_6[4871:4864];
        layer0[33][31:24] = buffer_data_6[4879:4872];
        layer0[33][39:32] = buffer_data_6[4887:4880];
        layer0[33][47:40] = buffer_data_6[4895:4888];
        layer0[33][55:48] = buffer_data_6[4903:4896];
        layer1[33][7:0] = buffer_data_5[4855:4848];
        layer1[33][15:8] = buffer_data_5[4863:4856];
        layer1[33][23:16] = buffer_data_5[4871:4864];
        layer1[33][31:24] = buffer_data_5[4879:4872];
        layer1[33][39:32] = buffer_data_5[4887:4880];
        layer1[33][47:40] = buffer_data_5[4895:4888];
        layer1[33][55:48] = buffer_data_5[4903:4896];
        layer2[33][7:0] = buffer_data_4[4855:4848];
        layer2[33][15:8] = buffer_data_4[4863:4856];
        layer2[33][23:16] = buffer_data_4[4871:4864];
        layer2[33][31:24] = buffer_data_4[4879:4872];
        layer2[33][39:32] = buffer_data_4[4887:4880];
        layer2[33][47:40] = buffer_data_4[4895:4888];
        layer2[33][55:48] = buffer_data_4[4903:4896];
        layer3[33][7:0] = buffer_data_3[4855:4848];
        layer3[33][15:8] = buffer_data_3[4863:4856];
        layer3[33][23:16] = buffer_data_3[4871:4864];
        layer3[33][31:24] = buffer_data_3[4879:4872];
        layer3[33][39:32] = buffer_data_3[4887:4880];
        layer3[33][47:40] = buffer_data_3[4895:4888];
        layer3[33][55:48] = buffer_data_3[4903:4896];
        layer4[33][7:0] = buffer_data_2[4855:4848];
        layer4[33][15:8] = buffer_data_2[4863:4856];
        layer4[33][23:16] = buffer_data_2[4871:4864];
        layer4[33][31:24] = buffer_data_2[4879:4872];
        layer4[33][39:32] = buffer_data_2[4887:4880];
        layer4[33][47:40] = buffer_data_2[4895:4888];
        layer4[33][55:48] = buffer_data_2[4903:4896];
        layer5[33][7:0] = buffer_data_1[4855:4848];
        layer5[33][15:8] = buffer_data_1[4863:4856];
        layer5[33][23:16] = buffer_data_1[4871:4864];
        layer5[33][31:24] = buffer_data_1[4879:4872];
        layer5[33][39:32] = buffer_data_1[4887:4880];
        layer5[33][47:40] = buffer_data_1[4895:4888];
        layer5[33][55:48] = buffer_data_1[4903:4896];
        layer6[33][7:0] = buffer_data_0[4855:4848];
        layer6[33][15:8] = buffer_data_0[4863:4856];
        layer6[33][23:16] = buffer_data_0[4871:4864];
        layer6[33][31:24] = buffer_data_0[4879:4872];
        layer6[33][39:32] = buffer_data_0[4887:4880];
        layer6[33][47:40] = buffer_data_0[4895:4888];
        layer6[33][55:48] = buffer_data_0[4903:4896];
        layer0[34][7:0] = buffer_data_6[4863:4856];
        layer0[34][15:8] = buffer_data_6[4871:4864];
        layer0[34][23:16] = buffer_data_6[4879:4872];
        layer0[34][31:24] = buffer_data_6[4887:4880];
        layer0[34][39:32] = buffer_data_6[4895:4888];
        layer0[34][47:40] = buffer_data_6[4903:4896];
        layer0[34][55:48] = buffer_data_6[4911:4904];
        layer1[34][7:0] = buffer_data_5[4863:4856];
        layer1[34][15:8] = buffer_data_5[4871:4864];
        layer1[34][23:16] = buffer_data_5[4879:4872];
        layer1[34][31:24] = buffer_data_5[4887:4880];
        layer1[34][39:32] = buffer_data_5[4895:4888];
        layer1[34][47:40] = buffer_data_5[4903:4896];
        layer1[34][55:48] = buffer_data_5[4911:4904];
        layer2[34][7:0] = buffer_data_4[4863:4856];
        layer2[34][15:8] = buffer_data_4[4871:4864];
        layer2[34][23:16] = buffer_data_4[4879:4872];
        layer2[34][31:24] = buffer_data_4[4887:4880];
        layer2[34][39:32] = buffer_data_4[4895:4888];
        layer2[34][47:40] = buffer_data_4[4903:4896];
        layer2[34][55:48] = buffer_data_4[4911:4904];
        layer3[34][7:0] = buffer_data_3[4863:4856];
        layer3[34][15:8] = buffer_data_3[4871:4864];
        layer3[34][23:16] = buffer_data_3[4879:4872];
        layer3[34][31:24] = buffer_data_3[4887:4880];
        layer3[34][39:32] = buffer_data_3[4895:4888];
        layer3[34][47:40] = buffer_data_3[4903:4896];
        layer3[34][55:48] = buffer_data_3[4911:4904];
        layer4[34][7:0] = buffer_data_2[4863:4856];
        layer4[34][15:8] = buffer_data_2[4871:4864];
        layer4[34][23:16] = buffer_data_2[4879:4872];
        layer4[34][31:24] = buffer_data_2[4887:4880];
        layer4[34][39:32] = buffer_data_2[4895:4888];
        layer4[34][47:40] = buffer_data_2[4903:4896];
        layer4[34][55:48] = buffer_data_2[4911:4904];
        layer5[34][7:0] = buffer_data_1[4863:4856];
        layer5[34][15:8] = buffer_data_1[4871:4864];
        layer5[34][23:16] = buffer_data_1[4879:4872];
        layer5[34][31:24] = buffer_data_1[4887:4880];
        layer5[34][39:32] = buffer_data_1[4895:4888];
        layer5[34][47:40] = buffer_data_1[4903:4896];
        layer5[34][55:48] = buffer_data_1[4911:4904];
        layer6[34][7:0] = buffer_data_0[4863:4856];
        layer6[34][15:8] = buffer_data_0[4871:4864];
        layer6[34][23:16] = buffer_data_0[4879:4872];
        layer6[34][31:24] = buffer_data_0[4887:4880];
        layer6[34][39:32] = buffer_data_0[4895:4888];
        layer6[34][47:40] = buffer_data_0[4903:4896];
        layer6[34][55:48] = buffer_data_0[4911:4904];
        layer0[35][7:0] = buffer_data_6[4871:4864];
        layer0[35][15:8] = buffer_data_6[4879:4872];
        layer0[35][23:16] = buffer_data_6[4887:4880];
        layer0[35][31:24] = buffer_data_6[4895:4888];
        layer0[35][39:32] = buffer_data_6[4903:4896];
        layer0[35][47:40] = buffer_data_6[4911:4904];
        layer0[35][55:48] = buffer_data_6[4919:4912];
        layer1[35][7:0] = buffer_data_5[4871:4864];
        layer1[35][15:8] = buffer_data_5[4879:4872];
        layer1[35][23:16] = buffer_data_5[4887:4880];
        layer1[35][31:24] = buffer_data_5[4895:4888];
        layer1[35][39:32] = buffer_data_5[4903:4896];
        layer1[35][47:40] = buffer_data_5[4911:4904];
        layer1[35][55:48] = buffer_data_5[4919:4912];
        layer2[35][7:0] = buffer_data_4[4871:4864];
        layer2[35][15:8] = buffer_data_4[4879:4872];
        layer2[35][23:16] = buffer_data_4[4887:4880];
        layer2[35][31:24] = buffer_data_4[4895:4888];
        layer2[35][39:32] = buffer_data_4[4903:4896];
        layer2[35][47:40] = buffer_data_4[4911:4904];
        layer2[35][55:48] = buffer_data_4[4919:4912];
        layer3[35][7:0] = buffer_data_3[4871:4864];
        layer3[35][15:8] = buffer_data_3[4879:4872];
        layer3[35][23:16] = buffer_data_3[4887:4880];
        layer3[35][31:24] = buffer_data_3[4895:4888];
        layer3[35][39:32] = buffer_data_3[4903:4896];
        layer3[35][47:40] = buffer_data_3[4911:4904];
        layer3[35][55:48] = buffer_data_3[4919:4912];
        layer4[35][7:0] = buffer_data_2[4871:4864];
        layer4[35][15:8] = buffer_data_2[4879:4872];
        layer4[35][23:16] = buffer_data_2[4887:4880];
        layer4[35][31:24] = buffer_data_2[4895:4888];
        layer4[35][39:32] = buffer_data_2[4903:4896];
        layer4[35][47:40] = buffer_data_2[4911:4904];
        layer4[35][55:48] = buffer_data_2[4919:4912];
        layer5[35][7:0] = buffer_data_1[4871:4864];
        layer5[35][15:8] = buffer_data_1[4879:4872];
        layer5[35][23:16] = buffer_data_1[4887:4880];
        layer5[35][31:24] = buffer_data_1[4895:4888];
        layer5[35][39:32] = buffer_data_1[4903:4896];
        layer5[35][47:40] = buffer_data_1[4911:4904];
        layer5[35][55:48] = buffer_data_1[4919:4912];
        layer6[35][7:0] = buffer_data_0[4871:4864];
        layer6[35][15:8] = buffer_data_0[4879:4872];
        layer6[35][23:16] = buffer_data_0[4887:4880];
        layer6[35][31:24] = buffer_data_0[4895:4888];
        layer6[35][39:32] = buffer_data_0[4903:4896];
        layer6[35][47:40] = buffer_data_0[4911:4904];
        layer6[35][55:48] = buffer_data_0[4919:4912];
        layer0[36][7:0] = buffer_data_6[4879:4872];
        layer0[36][15:8] = buffer_data_6[4887:4880];
        layer0[36][23:16] = buffer_data_6[4895:4888];
        layer0[36][31:24] = buffer_data_6[4903:4896];
        layer0[36][39:32] = buffer_data_6[4911:4904];
        layer0[36][47:40] = buffer_data_6[4919:4912];
        layer0[36][55:48] = buffer_data_6[4927:4920];
        layer1[36][7:0] = buffer_data_5[4879:4872];
        layer1[36][15:8] = buffer_data_5[4887:4880];
        layer1[36][23:16] = buffer_data_5[4895:4888];
        layer1[36][31:24] = buffer_data_5[4903:4896];
        layer1[36][39:32] = buffer_data_5[4911:4904];
        layer1[36][47:40] = buffer_data_5[4919:4912];
        layer1[36][55:48] = buffer_data_5[4927:4920];
        layer2[36][7:0] = buffer_data_4[4879:4872];
        layer2[36][15:8] = buffer_data_4[4887:4880];
        layer2[36][23:16] = buffer_data_4[4895:4888];
        layer2[36][31:24] = buffer_data_4[4903:4896];
        layer2[36][39:32] = buffer_data_4[4911:4904];
        layer2[36][47:40] = buffer_data_4[4919:4912];
        layer2[36][55:48] = buffer_data_4[4927:4920];
        layer3[36][7:0] = buffer_data_3[4879:4872];
        layer3[36][15:8] = buffer_data_3[4887:4880];
        layer3[36][23:16] = buffer_data_3[4895:4888];
        layer3[36][31:24] = buffer_data_3[4903:4896];
        layer3[36][39:32] = buffer_data_3[4911:4904];
        layer3[36][47:40] = buffer_data_3[4919:4912];
        layer3[36][55:48] = buffer_data_3[4927:4920];
        layer4[36][7:0] = buffer_data_2[4879:4872];
        layer4[36][15:8] = buffer_data_2[4887:4880];
        layer4[36][23:16] = buffer_data_2[4895:4888];
        layer4[36][31:24] = buffer_data_2[4903:4896];
        layer4[36][39:32] = buffer_data_2[4911:4904];
        layer4[36][47:40] = buffer_data_2[4919:4912];
        layer4[36][55:48] = buffer_data_2[4927:4920];
        layer5[36][7:0] = buffer_data_1[4879:4872];
        layer5[36][15:8] = buffer_data_1[4887:4880];
        layer5[36][23:16] = buffer_data_1[4895:4888];
        layer5[36][31:24] = buffer_data_1[4903:4896];
        layer5[36][39:32] = buffer_data_1[4911:4904];
        layer5[36][47:40] = buffer_data_1[4919:4912];
        layer5[36][55:48] = buffer_data_1[4927:4920];
        layer6[36][7:0] = buffer_data_0[4879:4872];
        layer6[36][15:8] = buffer_data_0[4887:4880];
        layer6[36][23:16] = buffer_data_0[4895:4888];
        layer6[36][31:24] = buffer_data_0[4903:4896];
        layer6[36][39:32] = buffer_data_0[4911:4904];
        layer6[36][47:40] = buffer_data_0[4919:4912];
        layer6[36][55:48] = buffer_data_0[4927:4920];
        layer0[37][7:0] = buffer_data_6[4887:4880];
        layer0[37][15:8] = buffer_data_6[4895:4888];
        layer0[37][23:16] = buffer_data_6[4903:4896];
        layer0[37][31:24] = buffer_data_6[4911:4904];
        layer0[37][39:32] = buffer_data_6[4919:4912];
        layer0[37][47:40] = buffer_data_6[4927:4920];
        layer0[37][55:48] = buffer_data_6[4935:4928];
        layer1[37][7:0] = buffer_data_5[4887:4880];
        layer1[37][15:8] = buffer_data_5[4895:4888];
        layer1[37][23:16] = buffer_data_5[4903:4896];
        layer1[37][31:24] = buffer_data_5[4911:4904];
        layer1[37][39:32] = buffer_data_5[4919:4912];
        layer1[37][47:40] = buffer_data_5[4927:4920];
        layer1[37][55:48] = buffer_data_5[4935:4928];
        layer2[37][7:0] = buffer_data_4[4887:4880];
        layer2[37][15:8] = buffer_data_4[4895:4888];
        layer2[37][23:16] = buffer_data_4[4903:4896];
        layer2[37][31:24] = buffer_data_4[4911:4904];
        layer2[37][39:32] = buffer_data_4[4919:4912];
        layer2[37][47:40] = buffer_data_4[4927:4920];
        layer2[37][55:48] = buffer_data_4[4935:4928];
        layer3[37][7:0] = buffer_data_3[4887:4880];
        layer3[37][15:8] = buffer_data_3[4895:4888];
        layer3[37][23:16] = buffer_data_3[4903:4896];
        layer3[37][31:24] = buffer_data_3[4911:4904];
        layer3[37][39:32] = buffer_data_3[4919:4912];
        layer3[37][47:40] = buffer_data_3[4927:4920];
        layer3[37][55:48] = buffer_data_3[4935:4928];
        layer4[37][7:0] = buffer_data_2[4887:4880];
        layer4[37][15:8] = buffer_data_2[4895:4888];
        layer4[37][23:16] = buffer_data_2[4903:4896];
        layer4[37][31:24] = buffer_data_2[4911:4904];
        layer4[37][39:32] = buffer_data_2[4919:4912];
        layer4[37][47:40] = buffer_data_2[4927:4920];
        layer4[37][55:48] = buffer_data_2[4935:4928];
        layer5[37][7:0] = buffer_data_1[4887:4880];
        layer5[37][15:8] = buffer_data_1[4895:4888];
        layer5[37][23:16] = buffer_data_1[4903:4896];
        layer5[37][31:24] = buffer_data_1[4911:4904];
        layer5[37][39:32] = buffer_data_1[4919:4912];
        layer5[37][47:40] = buffer_data_1[4927:4920];
        layer5[37][55:48] = buffer_data_1[4935:4928];
        layer6[37][7:0] = buffer_data_0[4887:4880];
        layer6[37][15:8] = buffer_data_0[4895:4888];
        layer6[37][23:16] = buffer_data_0[4903:4896];
        layer6[37][31:24] = buffer_data_0[4911:4904];
        layer6[37][39:32] = buffer_data_0[4919:4912];
        layer6[37][47:40] = buffer_data_0[4927:4920];
        layer6[37][55:48] = buffer_data_0[4935:4928];
        layer0[38][7:0] = buffer_data_6[4895:4888];
        layer0[38][15:8] = buffer_data_6[4903:4896];
        layer0[38][23:16] = buffer_data_6[4911:4904];
        layer0[38][31:24] = buffer_data_6[4919:4912];
        layer0[38][39:32] = buffer_data_6[4927:4920];
        layer0[38][47:40] = buffer_data_6[4935:4928];
        layer0[38][55:48] = buffer_data_6[4943:4936];
        layer1[38][7:0] = buffer_data_5[4895:4888];
        layer1[38][15:8] = buffer_data_5[4903:4896];
        layer1[38][23:16] = buffer_data_5[4911:4904];
        layer1[38][31:24] = buffer_data_5[4919:4912];
        layer1[38][39:32] = buffer_data_5[4927:4920];
        layer1[38][47:40] = buffer_data_5[4935:4928];
        layer1[38][55:48] = buffer_data_5[4943:4936];
        layer2[38][7:0] = buffer_data_4[4895:4888];
        layer2[38][15:8] = buffer_data_4[4903:4896];
        layer2[38][23:16] = buffer_data_4[4911:4904];
        layer2[38][31:24] = buffer_data_4[4919:4912];
        layer2[38][39:32] = buffer_data_4[4927:4920];
        layer2[38][47:40] = buffer_data_4[4935:4928];
        layer2[38][55:48] = buffer_data_4[4943:4936];
        layer3[38][7:0] = buffer_data_3[4895:4888];
        layer3[38][15:8] = buffer_data_3[4903:4896];
        layer3[38][23:16] = buffer_data_3[4911:4904];
        layer3[38][31:24] = buffer_data_3[4919:4912];
        layer3[38][39:32] = buffer_data_3[4927:4920];
        layer3[38][47:40] = buffer_data_3[4935:4928];
        layer3[38][55:48] = buffer_data_3[4943:4936];
        layer4[38][7:0] = buffer_data_2[4895:4888];
        layer4[38][15:8] = buffer_data_2[4903:4896];
        layer4[38][23:16] = buffer_data_2[4911:4904];
        layer4[38][31:24] = buffer_data_2[4919:4912];
        layer4[38][39:32] = buffer_data_2[4927:4920];
        layer4[38][47:40] = buffer_data_2[4935:4928];
        layer4[38][55:48] = buffer_data_2[4943:4936];
        layer5[38][7:0] = buffer_data_1[4895:4888];
        layer5[38][15:8] = buffer_data_1[4903:4896];
        layer5[38][23:16] = buffer_data_1[4911:4904];
        layer5[38][31:24] = buffer_data_1[4919:4912];
        layer5[38][39:32] = buffer_data_1[4927:4920];
        layer5[38][47:40] = buffer_data_1[4935:4928];
        layer5[38][55:48] = buffer_data_1[4943:4936];
        layer6[38][7:0] = buffer_data_0[4895:4888];
        layer6[38][15:8] = buffer_data_0[4903:4896];
        layer6[38][23:16] = buffer_data_0[4911:4904];
        layer6[38][31:24] = buffer_data_0[4919:4912];
        layer6[38][39:32] = buffer_data_0[4927:4920];
        layer6[38][47:40] = buffer_data_0[4935:4928];
        layer6[38][55:48] = buffer_data_0[4943:4936];
        layer0[39][7:0] = buffer_data_6[4903:4896];
        layer0[39][15:8] = buffer_data_6[4911:4904];
        layer0[39][23:16] = buffer_data_6[4919:4912];
        layer0[39][31:24] = buffer_data_6[4927:4920];
        layer0[39][39:32] = buffer_data_6[4935:4928];
        layer0[39][47:40] = buffer_data_6[4943:4936];
        layer0[39][55:48] = buffer_data_6[4951:4944];
        layer1[39][7:0] = buffer_data_5[4903:4896];
        layer1[39][15:8] = buffer_data_5[4911:4904];
        layer1[39][23:16] = buffer_data_5[4919:4912];
        layer1[39][31:24] = buffer_data_5[4927:4920];
        layer1[39][39:32] = buffer_data_5[4935:4928];
        layer1[39][47:40] = buffer_data_5[4943:4936];
        layer1[39][55:48] = buffer_data_5[4951:4944];
        layer2[39][7:0] = buffer_data_4[4903:4896];
        layer2[39][15:8] = buffer_data_4[4911:4904];
        layer2[39][23:16] = buffer_data_4[4919:4912];
        layer2[39][31:24] = buffer_data_4[4927:4920];
        layer2[39][39:32] = buffer_data_4[4935:4928];
        layer2[39][47:40] = buffer_data_4[4943:4936];
        layer2[39][55:48] = buffer_data_4[4951:4944];
        layer3[39][7:0] = buffer_data_3[4903:4896];
        layer3[39][15:8] = buffer_data_3[4911:4904];
        layer3[39][23:16] = buffer_data_3[4919:4912];
        layer3[39][31:24] = buffer_data_3[4927:4920];
        layer3[39][39:32] = buffer_data_3[4935:4928];
        layer3[39][47:40] = buffer_data_3[4943:4936];
        layer3[39][55:48] = buffer_data_3[4951:4944];
        layer4[39][7:0] = buffer_data_2[4903:4896];
        layer4[39][15:8] = buffer_data_2[4911:4904];
        layer4[39][23:16] = buffer_data_2[4919:4912];
        layer4[39][31:24] = buffer_data_2[4927:4920];
        layer4[39][39:32] = buffer_data_2[4935:4928];
        layer4[39][47:40] = buffer_data_2[4943:4936];
        layer4[39][55:48] = buffer_data_2[4951:4944];
        layer5[39][7:0] = buffer_data_1[4903:4896];
        layer5[39][15:8] = buffer_data_1[4911:4904];
        layer5[39][23:16] = buffer_data_1[4919:4912];
        layer5[39][31:24] = buffer_data_1[4927:4920];
        layer5[39][39:32] = buffer_data_1[4935:4928];
        layer5[39][47:40] = buffer_data_1[4943:4936];
        layer5[39][55:48] = buffer_data_1[4951:4944];
        layer6[39][7:0] = buffer_data_0[4903:4896];
        layer6[39][15:8] = buffer_data_0[4911:4904];
        layer6[39][23:16] = buffer_data_0[4919:4912];
        layer6[39][31:24] = buffer_data_0[4927:4920];
        layer6[39][39:32] = buffer_data_0[4935:4928];
        layer6[39][47:40] = buffer_data_0[4943:4936];
        layer6[39][55:48] = buffer_data_0[4951:4944];
        layer0[40][7:0] = buffer_data_6[4911:4904];
        layer0[40][15:8] = buffer_data_6[4919:4912];
        layer0[40][23:16] = buffer_data_6[4927:4920];
        layer0[40][31:24] = buffer_data_6[4935:4928];
        layer0[40][39:32] = buffer_data_6[4943:4936];
        layer0[40][47:40] = buffer_data_6[4951:4944];
        layer0[40][55:48] = buffer_data_6[4959:4952];
        layer1[40][7:0] = buffer_data_5[4911:4904];
        layer1[40][15:8] = buffer_data_5[4919:4912];
        layer1[40][23:16] = buffer_data_5[4927:4920];
        layer1[40][31:24] = buffer_data_5[4935:4928];
        layer1[40][39:32] = buffer_data_5[4943:4936];
        layer1[40][47:40] = buffer_data_5[4951:4944];
        layer1[40][55:48] = buffer_data_5[4959:4952];
        layer2[40][7:0] = buffer_data_4[4911:4904];
        layer2[40][15:8] = buffer_data_4[4919:4912];
        layer2[40][23:16] = buffer_data_4[4927:4920];
        layer2[40][31:24] = buffer_data_4[4935:4928];
        layer2[40][39:32] = buffer_data_4[4943:4936];
        layer2[40][47:40] = buffer_data_4[4951:4944];
        layer2[40][55:48] = buffer_data_4[4959:4952];
        layer3[40][7:0] = buffer_data_3[4911:4904];
        layer3[40][15:8] = buffer_data_3[4919:4912];
        layer3[40][23:16] = buffer_data_3[4927:4920];
        layer3[40][31:24] = buffer_data_3[4935:4928];
        layer3[40][39:32] = buffer_data_3[4943:4936];
        layer3[40][47:40] = buffer_data_3[4951:4944];
        layer3[40][55:48] = buffer_data_3[4959:4952];
        layer4[40][7:0] = buffer_data_2[4911:4904];
        layer4[40][15:8] = buffer_data_2[4919:4912];
        layer4[40][23:16] = buffer_data_2[4927:4920];
        layer4[40][31:24] = buffer_data_2[4935:4928];
        layer4[40][39:32] = buffer_data_2[4943:4936];
        layer4[40][47:40] = buffer_data_2[4951:4944];
        layer4[40][55:48] = buffer_data_2[4959:4952];
        layer5[40][7:0] = buffer_data_1[4911:4904];
        layer5[40][15:8] = buffer_data_1[4919:4912];
        layer5[40][23:16] = buffer_data_1[4927:4920];
        layer5[40][31:24] = buffer_data_1[4935:4928];
        layer5[40][39:32] = buffer_data_1[4943:4936];
        layer5[40][47:40] = buffer_data_1[4951:4944];
        layer5[40][55:48] = buffer_data_1[4959:4952];
        layer6[40][7:0] = buffer_data_0[4911:4904];
        layer6[40][15:8] = buffer_data_0[4919:4912];
        layer6[40][23:16] = buffer_data_0[4927:4920];
        layer6[40][31:24] = buffer_data_0[4935:4928];
        layer6[40][39:32] = buffer_data_0[4943:4936];
        layer6[40][47:40] = buffer_data_0[4951:4944];
        layer6[40][55:48] = buffer_data_0[4959:4952];
        layer0[41][7:0] = buffer_data_6[4919:4912];
        layer0[41][15:8] = buffer_data_6[4927:4920];
        layer0[41][23:16] = buffer_data_6[4935:4928];
        layer0[41][31:24] = buffer_data_6[4943:4936];
        layer0[41][39:32] = buffer_data_6[4951:4944];
        layer0[41][47:40] = buffer_data_6[4959:4952];
        layer0[41][55:48] = buffer_data_6[4967:4960];
        layer1[41][7:0] = buffer_data_5[4919:4912];
        layer1[41][15:8] = buffer_data_5[4927:4920];
        layer1[41][23:16] = buffer_data_5[4935:4928];
        layer1[41][31:24] = buffer_data_5[4943:4936];
        layer1[41][39:32] = buffer_data_5[4951:4944];
        layer1[41][47:40] = buffer_data_5[4959:4952];
        layer1[41][55:48] = buffer_data_5[4967:4960];
        layer2[41][7:0] = buffer_data_4[4919:4912];
        layer2[41][15:8] = buffer_data_4[4927:4920];
        layer2[41][23:16] = buffer_data_4[4935:4928];
        layer2[41][31:24] = buffer_data_4[4943:4936];
        layer2[41][39:32] = buffer_data_4[4951:4944];
        layer2[41][47:40] = buffer_data_4[4959:4952];
        layer2[41][55:48] = buffer_data_4[4967:4960];
        layer3[41][7:0] = buffer_data_3[4919:4912];
        layer3[41][15:8] = buffer_data_3[4927:4920];
        layer3[41][23:16] = buffer_data_3[4935:4928];
        layer3[41][31:24] = buffer_data_3[4943:4936];
        layer3[41][39:32] = buffer_data_3[4951:4944];
        layer3[41][47:40] = buffer_data_3[4959:4952];
        layer3[41][55:48] = buffer_data_3[4967:4960];
        layer4[41][7:0] = buffer_data_2[4919:4912];
        layer4[41][15:8] = buffer_data_2[4927:4920];
        layer4[41][23:16] = buffer_data_2[4935:4928];
        layer4[41][31:24] = buffer_data_2[4943:4936];
        layer4[41][39:32] = buffer_data_2[4951:4944];
        layer4[41][47:40] = buffer_data_2[4959:4952];
        layer4[41][55:48] = buffer_data_2[4967:4960];
        layer5[41][7:0] = buffer_data_1[4919:4912];
        layer5[41][15:8] = buffer_data_1[4927:4920];
        layer5[41][23:16] = buffer_data_1[4935:4928];
        layer5[41][31:24] = buffer_data_1[4943:4936];
        layer5[41][39:32] = buffer_data_1[4951:4944];
        layer5[41][47:40] = buffer_data_1[4959:4952];
        layer5[41][55:48] = buffer_data_1[4967:4960];
        layer6[41][7:0] = buffer_data_0[4919:4912];
        layer6[41][15:8] = buffer_data_0[4927:4920];
        layer6[41][23:16] = buffer_data_0[4935:4928];
        layer6[41][31:24] = buffer_data_0[4943:4936];
        layer6[41][39:32] = buffer_data_0[4951:4944];
        layer6[41][47:40] = buffer_data_0[4959:4952];
        layer6[41][55:48] = buffer_data_0[4967:4960];
        layer0[42][7:0] = buffer_data_6[4927:4920];
        layer0[42][15:8] = buffer_data_6[4935:4928];
        layer0[42][23:16] = buffer_data_6[4943:4936];
        layer0[42][31:24] = buffer_data_6[4951:4944];
        layer0[42][39:32] = buffer_data_6[4959:4952];
        layer0[42][47:40] = buffer_data_6[4967:4960];
        layer0[42][55:48] = buffer_data_6[4975:4968];
        layer1[42][7:0] = buffer_data_5[4927:4920];
        layer1[42][15:8] = buffer_data_5[4935:4928];
        layer1[42][23:16] = buffer_data_5[4943:4936];
        layer1[42][31:24] = buffer_data_5[4951:4944];
        layer1[42][39:32] = buffer_data_5[4959:4952];
        layer1[42][47:40] = buffer_data_5[4967:4960];
        layer1[42][55:48] = buffer_data_5[4975:4968];
        layer2[42][7:0] = buffer_data_4[4927:4920];
        layer2[42][15:8] = buffer_data_4[4935:4928];
        layer2[42][23:16] = buffer_data_4[4943:4936];
        layer2[42][31:24] = buffer_data_4[4951:4944];
        layer2[42][39:32] = buffer_data_4[4959:4952];
        layer2[42][47:40] = buffer_data_4[4967:4960];
        layer2[42][55:48] = buffer_data_4[4975:4968];
        layer3[42][7:0] = buffer_data_3[4927:4920];
        layer3[42][15:8] = buffer_data_3[4935:4928];
        layer3[42][23:16] = buffer_data_3[4943:4936];
        layer3[42][31:24] = buffer_data_3[4951:4944];
        layer3[42][39:32] = buffer_data_3[4959:4952];
        layer3[42][47:40] = buffer_data_3[4967:4960];
        layer3[42][55:48] = buffer_data_3[4975:4968];
        layer4[42][7:0] = buffer_data_2[4927:4920];
        layer4[42][15:8] = buffer_data_2[4935:4928];
        layer4[42][23:16] = buffer_data_2[4943:4936];
        layer4[42][31:24] = buffer_data_2[4951:4944];
        layer4[42][39:32] = buffer_data_2[4959:4952];
        layer4[42][47:40] = buffer_data_2[4967:4960];
        layer4[42][55:48] = buffer_data_2[4975:4968];
        layer5[42][7:0] = buffer_data_1[4927:4920];
        layer5[42][15:8] = buffer_data_1[4935:4928];
        layer5[42][23:16] = buffer_data_1[4943:4936];
        layer5[42][31:24] = buffer_data_1[4951:4944];
        layer5[42][39:32] = buffer_data_1[4959:4952];
        layer5[42][47:40] = buffer_data_1[4967:4960];
        layer5[42][55:48] = buffer_data_1[4975:4968];
        layer6[42][7:0] = buffer_data_0[4927:4920];
        layer6[42][15:8] = buffer_data_0[4935:4928];
        layer6[42][23:16] = buffer_data_0[4943:4936];
        layer6[42][31:24] = buffer_data_0[4951:4944];
        layer6[42][39:32] = buffer_data_0[4959:4952];
        layer6[42][47:40] = buffer_data_0[4967:4960];
        layer6[42][55:48] = buffer_data_0[4975:4968];
        layer0[43][7:0] = buffer_data_6[4935:4928];
        layer0[43][15:8] = buffer_data_6[4943:4936];
        layer0[43][23:16] = buffer_data_6[4951:4944];
        layer0[43][31:24] = buffer_data_6[4959:4952];
        layer0[43][39:32] = buffer_data_6[4967:4960];
        layer0[43][47:40] = buffer_data_6[4975:4968];
        layer0[43][55:48] = buffer_data_6[4983:4976];
        layer1[43][7:0] = buffer_data_5[4935:4928];
        layer1[43][15:8] = buffer_data_5[4943:4936];
        layer1[43][23:16] = buffer_data_5[4951:4944];
        layer1[43][31:24] = buffer_data_5[4959:4952];
        layer1[43][39:32] = buffer_data_5[4967:4960];
        layer1[43][47:40] = buffer_data_5[4975:4968];
        layer1[43][55:48] = buffer_data_5[4983:4976];
        layer2[43][7:0] = buffer_data_4[4935:4928];
        layer2[43][15:8] = buffer_data_4[4943:4936];
        layer2[43][23:16] = buffer_data_4[4951:4944];
        layer2[43][31:24] = buffer_data_4[4959:4952];
        layer2[43][39:32] = buffer_data_4[4967:4960];
        layer2[43][47:40] = buffer_data_4[4975:4968];
        layer2[43][55:48] = buffer_data_4[4983:4976];
        layer3[43][7:0] = buffer_data_3[4935:4928];
        layer3[43][15:8] = buffer_data_3[4943:4936];
        layer3[43][23:16] = buffer_data_3[4951:4944];
        layer3[43][31:24] = buffer_data_3[4959:4952];
        layer3[43][39:32] = buffer_data_3[4967:4960];
        layer3[43][47:40] = buffer_data_3[4975:4968];
        layer3[43][55:48] = buffer_data_3[4983:4976];
        layer4[43][7:0] = buffer_data_2[4935:4928];
        layer4[43][15:8] = buffer_data_2[4943:4936];
        layer4[43][23:16] = buffer_data_2[4951:4944];
        layer4[43][31:24] = buffer_data_2[4959:4952];
        layer4[43][39:32] = buffer_data_2[4967:4960];
        layer4[43][47:40] = buffer_data_2[4975:4968];
        layer4[43][55:48] = buffer_data_2[4983:4976];
        layer5[43][7:0] = buffer_data_1[4935:4928];
        layer5[43][15:8] = buffer_data_1[4943:4936];
        layer5[43][23:16] = buffer_data_1[4951:4944];
        layer5[43][31:24] = buffer_data_1[4959:4952];
        layer5[43][39:32] = buffer_data_1[4967:4960];
        layer5[43][47:40] = buffer_data_1[4975:4968];
        layer5[43][55:48] = buffer_data_1[4983:4976];
        layer6[43][7:0] = buffer_data_0[4935:4928];
        layer6[43][15:8] = buffer_data_0[4943:4936];
        layer6[43][23:16] = buffer_data_0[4951:4944];
        layer6[43][31:24] = buffer_data_0[4959:4952];
        layer6[43][39:32] = buffer_data_0[4967:4960];
        layer6[43][47:40] = buffer_data_0[4975:4968];
        layer6[43][55:48] = buffer_data_0[4983:4976];
        layer0[44][7:0] = buffer_data_6[4943:4936];
        layer0[44][15:8] = buffer_data_6[4951:4944];
        layer0[44][23:16] = buffer_data_6[4959:4952];
        layer0[44][31:24] = buffer_data_6[4967:4960];
        layer0[44][39:32] = buffer_data_6[4975:4968];
        layer0[44][47:40] = buffer_data_6[4983:4976];
        layer0[44][55:48] = buffer_data_6[4991:4984];
        layer1[44][7:0] = buffer_data_5[4943:4936];
        layer1[44][15:8] = buffer_data_5[4951:4944];
        layer1[44][23:16] = buffer_data_5[4959:4952];
        layer1[44][31:24] = buffer_data_5[4967:4960];
        layer1[44][39:32] = buffer_data_5[4975:4968];
        layer1[44][47:40] = buffer_data_5[4983:4976];
        layer1[44][55:48] = buffer_data_5[4991:4984];
        layer2[44][7:0] = buffer_data_4[4943:4936];
        layer2[44][15:8] = buffer_data_4[4951:4944];
        layer2[44][23:16] = buffer_data_4[4959:4952];
        layer2[44][31:24] = buffer_data_4[4967:4960];
        layer2[44][39:32] = buffer_data_4[4975:4968];
        layer2[44][47:40] = buffer_data_4[4983:4976];
        layer2[44][55:48] = buffer_data_4[4991:4984];
        layer3[44][7:0] = buffer_data_3[4943:4936];
        layer3[44][15:8] = buffer_data_3[4951:4944];
        layer3[44][23:16] = buffer_data_3[4959:4952];
        layer3[44][31:24] = buffer_data_3[4967:4960];
        layer3[44][39:32] = buffer_data_3[4975:4968];
        layer3[44][47:40] = buffer_data_3[4983:4976];
        layer3[44][55:48] = buffer_data_3[4991:4984];
        layer4[44][7:0] = buffer_data_2[4943:4936];
        layer4[44][15:8] = buffer_data_2[4951:4944];
        layer4[44][23:16] = buffer_data_2[4959:4952];
        layer4[44][31:24] = buffer_data_2[4967:4960];
        layer4[44][39:32] = buffer_data_2[4975:4968];
        layer4[44][47:40] = buffer_data_2[4983:4976];
        layer4[44][55:48] = buffer_data_2[4991:4984];
        layer5[44][7:0] = buffer_data_1[4943:4936];
        layer5[44][15:8] = buffer_data_1[4951:4944];
        layer5[44][23:16] = buffer_data_1[4959:4952];
        layer5[44][31:24] = buffer_data_1[4967:4960];
        layer5[44][39:32] = buffer_data_1[4975:4968];
        layer5[44][47:40] = buffer_data_1[4983:4976];
        layer5[44][55:48] = buffer_data_1[4991:4984];
        layer6[44][7:0] = buffer_data_0[4943:4936];
        layer6[44][15:8] = buffer_data_0[4951:4944];
        layer6[44][23:16] = buffer_data_0[4959:4952];
        layer6[44][31:24] = buffer_data_0[4967:4960];
        layer6[44][39:32] = buffer_data_0[4975:4968];
        layer6[44][47:40] = buffer_data_0[4983:4976];
        layer6[44][55:48] = buffer_data_0[4991:4984];
        layer0[45][7:0] = buffer_data_6[4951:4944];
        layer0[45][15:8] = buffer_data_6[4959:4952];
        layer0[45][23:16] = buffer_data_6[4967:4960];
        layer0[45][31:24] = buffer_data_6[4975:4968];
        layer0[45][39:32] = buffer_data_6[4983:4976];
        layer0[45][47:40] = buffer_data_6[4991:4984];
        layer0[45][55:48] = buffer_data_6[4999:4992];
        layer1[45][7:0] = buffer_data_5[4951:4944];
        layer1[45][15:8] = buffer_data_5[4959:4952];
        layer1[45][23:16] = buffer_data_5[4967:4960];
        layer1[45][31:24] = buffer_data_5[4975:4968];
        layer1[45][39:32] = buffer_data_5[4983:4976];
        layer1[45][47:40] = buffer_data_5[4991:4984];
        layer1[45][55:48] = buffer_data_5[4999:4992];
        layer2[45][7:0] = buffer_data_4[4951:4944];
        layer2[45][15:8] = buffer_data_4[4959:4952];
        layer2[45][23:16] = buffer_data_4[4967:4960];
        layer2[45][31:24] = buffer_data_4[4975:4968];
        layer2[45][39:32] = buffer_data_4[4983:4976];
        layer2[45][47:40] = buffer_data_4[4991:4984];
        layer2[45][55:48] = buffer_data_4[4999:4992];
        layer3[45][7:0] = buffer_data_3[4951:4944];
        layer3[45][15:8] = buffer_data_3[4959:4952];
        layer3[45][23:16] = buffer_data_3[4967:4960];
        layer3[45][31:24] = buffer_data_3[4975:4968];
        layer3[45][39:32] = buffer_data_3[4983:4976];
        layer3[45][47:40] = buffer_data_3[4991:4984];
        layer3[45][55:48] = buffer_data_3[4999:4992];
        layer4[45][7:0] = buffer_data_2[4951:4944];
        layer4[45][15:8] = buffer_data_2[4959:4952];
        layer4[45][23:16] = buffer_data_2[4967:4960];
        layer4[45][31:24] = buffer_data_2[4975:4968];
        layer4[45][39:32] = buffer_data_2[4983:4976];
        layer4[45][47:40] = buffer_data_2[4991:4984];
        layer4[45][55:48] = buffer_data_2[4999:4992];
        layer5[45][7:0] = buffer_data_1[4951:4944];
        layer5[45][15:8] = buffer_data_1[4959:4952];
        layer5[45][23:16] = buffer_data_1[4967:4960];
        layer5[45][31:24] = buffer_data_1[4975:4968];
        layer5[45][39:32] = buffer_data_1[4983:4976];
        layer5[45][47:40] = buffer_data_1[4991:4984];
        layer5[45][55:48] = buffer_data_1[4999:4992];
        layer6[45][7:0] = buffer_data_0[4951:4944];
        layer6[45][15:8] = buffer_data_0[4959:4952];
        layer6[45][23:16] = buffer_data_0[4967:4960];
        layer6[45][31:24] = buffer_data_0[4975:4968];
        layer6[45][39:32] = buffer_data_0[4983:4976];
        layer6[45][47:40] = buffer_data_0[4991:4984];
        layer6[45][55:48] = buffer_data_0[4999:4992];
        layer0[46][7:0] = buffer_data_6[4959:4952];
        layer0[46][15:8] = buffer_data_6[4967:4960];
        layer0[46][23:16] = buffer_data_6[4975:4968];
        layer0[46][31:24] = buffer_data_6[4983:4976];
        layer0[46][39:32] = buffer_data_6[4991:4984];
        layer0[46][47:40] = buffer_data_6[4999:4992];
        layer0[46][55:48] = buffer_data_6[5007:5000];
        layer1[46][7:0] = buffer_data_5[4959:4952];
        layer1[46][15:8] = buffer_data_5[4967:4960];
        layer1[46][23:16] = buffer_data_5[4975:4968];
        layer1[46][31:24] = buffer_data_5[4983:4976];
        layer1[46][39:32] = buffer_data_5[4991:4984];
        layer1[46][47:40] = buffer_data_5[4999:4992];
        layer1[46][55:48] = buffer_data_5[5007:5000];
        layer2[46][7:0] = buffer_data_4[4959:4952];
        layer2[46][15:8] = buffer_data_4[4967:4960];
        layer2[46][23:16] = buffer_data_4[4975:4968];
        layer2[46][31:24] = buffer_data_4[4983:4976];
        layer2[46][39:32] = buffer_data_4[4991:4984];
        layer2[46][47:40] = buffer_data_4[4999:4992];
        layer2[46][55:48] = buffer_data_4[5007:5000];
        layer3[46][7:0] = buffer_data_3[4959:4952];
        layer3[46][15:8] = buffer_data_3[4967:4960];
        layer3[46][23:16] = buffer_data_3[4975:4968];
        layer3[46][31:24] = buffer_data_3[4983:4976];
        layer3[46][39:32] = buffer_data_3[4991:4984];
        layer3[46][47:40] = buffer_data_3[4999:4992];
        layer3[46][55:48] = buffer_data_3[5007:5000];
        layer4[46][7:0] = buffer_data_2[4959:4952];
        layer4[46][15:8] = buffer_data_2[4967:4960];
        layer4[46][23:16] = buffer_data_2[4975:4968];
        layer4[46][31:24] = buffer_data_2[4983:4976];
        layer4[46][39:32] = buffer_data_2[4991:4984];
        layer4[46][47:40] = buffer_data_2[4999:4992];
        layer4[46][55:48] = buffer_data_2[5007:5000];
        layer5[46][7:0] = buffer_data_1[4959:4952];
        layer5[46][15:8] = buffer_data_1[4967:4960];
        layer5[46][23:16] = buffer_data_1[4975:4968];
        layer5[46][31:24] = buffer_data_1[4983:4976];
        layer5[46][39:32] = buffer_data_1[4991:4984];
        layer5[46][47:40] = buffer_data_1[4999:4992];
        layer5[46][55:48] = buffer_data_1[5007:5000];
        layer6[46][7:0] = buffer_data_0[4959:4952];
        layer6[46][15:8] = buffer_data_0[4967:4960];
        layer6[46][23:16] = buffer_data_0[4975:4968];
        layer6[46][31:24] = buffer_data_0[4983:4976];
        layer6[46][39:32] = buffer_data_0[4991:4984];
        layer6[46][47:40] = buffer_data_0[4999:4992];
        layer6[46][55:48] = buffer_data_0[5007:5000];
        layer0[47][7:0] = buffer_data_6[4967:4960];
        layer0[47][15:8] = buffer_data_6[4975:4968];
        layer0[47][23:16] = buffer_data_6[4983:4976];
        layer0[47][31:24] = buffer_data_6[4991:4984];
        layer0[47][39:32] = buffer_data_6[4999:4992];
        layer0[47][47:40] = buffer_data_6[5007:5000];
        layer0[47][55:48] = buffer_data_6[5015:5008];
        layer1[47][7:0] = buffer_data_5[4967:4960];
        layer1[47][15:8] = buffer_data_5[4975:4968];
        layer1[47][23:16] = buffer_data_5[4983:4976];
        layer1[47][31:24] = buffer_data_5[4991:4984];
        layer1[47][39:32] = buffer_data_5[4999:4992];
        layer1[47][47:40] = buffer_data_5[5007:5000];
        layer1[47][55:48] = buffer_data_5[5015:5008];
        layer2[47][7:0] = buffer_data_4[4967:4960];
        layer2[47][15:8] = buffer_data_4[4975:4968];
        layer2[47][23:16] = buffer_data_4[4983:4976];
        layer2[47][31:24] = buffer_data_4[4991:4984];
        layer2[47][39:32] = buffer_data_4[4999:4992];
        layer2[47][47:40] = buffer_data_4[5007:5000];
        layer2[47][55:48] = buffer_data_4[5015:5008];
        layer3[47][7:0] = buffer_data_3[4967:4960];
        layer3[47][15:8] = buffer_data_3[4975:4968];
        layer3[47][23:16] = buffer_data_3[4983:4976];
        layer3[47][31:24] = buffer_data_3[4991:4984];
        layer3[47][39:32] = buffer_data_3[4999:4992];
        layer3[47][47:40] = buffer_data_3[5007:5000];
        layer3[47][55:48] = buffer_data_3[5015:5008];
        layer4[47][7:0] = buffer_data_2[4967:4960];
        layer4[47][15:8] = buffer_data_2[4975:4968];
        layer4[47][23:16] = buffer_data_2[4983:4976];
        layer4[47][31:24] = buffer_data_2[4991:4984];
        layer4[47][39:32] = buffer_data_2[4999:4992];
        layer4[47][47:40] = buffer_data_2[5007:5000];
        layer4[47][55:48] = buffer_data_2[5015:5008];
        layer5[47][7:0] = buffer_data_1[4967:4960];
        layer5[47][15:8] = buffer_data_1[4975:4968];
        layer5[47][23:16] = buffer_data_1[4983:4976];
        layer5[47][31:24] = buffer_data_1[4991:4984];
        layer5[47][39:32] = buffer_data_1[4999:4992];
        layer5[47][47:40] = buffer_data_1[5007:5000];
        layer5[47][55:48] = buffer_data_1[5015:5008];
        layer6[47][7:0] = buffer_data_0[4967:4960];
        layer6[47][15:8] = buffer_data_0[4975:4968];
        layer6[47][23:16] = buffer_data_0[4983:4976];
        layer6[47][31:24] = buffer_data_0[4991:4984];
        layer6[47][39:32] = buffer_data_0[4999:4992];
        layer6[47][47:40] = buffer_data_0[5007:5000];
        layer6[47][55:48] = buffer_data_0[5015:5008];
        layer0[48][7:0] = buffer_data_6[4975:4968];
        layer0[48][15:8] = buffer_data_6[4983:4976];
        layer0[48][23:16] = buffer_data_6[4991:4984];
        layer0[48][31:24] = buffer_data_6[4999:4992];
        layer0[48][39:32] = buffer_data_6[5007:5000];
        layer0[48][47:40] = buffer_data_6[5015:5008];
        layer0[48][55:48] = buffer_data_6[5023:5016];
        layer1[48][7:0] = buffer_data_5[4975:4968];
        layer1[48][15:8] = buffer_data_5[4983:4976];
        layer1[48][23:16] = buffer_data_5[4991:4984];
        layer1[48][31:24] = buffer_data_5[4999:4992];
        layer1[48][39:32] = buffer_data_5[5007:5000];
        layer1[48][47:40] = buffer_data_5[5015:5008];
        layer1[48][55:48] = buffer_data_5[5023:5016];
        layer2[48][7:0] = buffer_data_4[4975:4968];
        layer2[48][15:8] = buffer_data_4[4983:4976];
        layer2[48][23:16] = buffer_data_4[4991:4984];
        layer2[48][31:24] = buffer_data_4[4999:4992];
        layer2[48][39:32] = buffer_data_4[5007:5000];
        layer2[48][47:40] = buffer_data_4[5015:5008];
        layer2[48][55:48] = buffer_data_4[5023:5016];
        layer3[48][7:0] = buffer_data_3[4975:4968];
        layer3[48][15:8] = buffer_data_3[4983:4976];
        layer3[48][23:16] = buffer_data_3[4991:4984];
        layer3[48][31:24] = buffer_data_3[4999:4992];
        layer3[48][39:32] = buffer_data_3[5007:5000];
        layer3[48][47:40] = buffer_data_3[5015:5008];
        layer3[48][55:48] = buffer_data_3[5023:5016];
        layer4[48][7:0] = buffer_data_2[4975:4968];
        layer4[48][15:8] = buffer_data_2[4983:4976];
        layer4[48][23:16] = buffer_data_2[4991:4984];
        layer4[48][31:24] = buffer_data_2[4999:4992];
        layer4[48][39:32] = buffer_data_2[5007:5000];
        layer4[48][47:40] = buffer_data_2[5015:5008];
        layer4[48][55:48] = buffer_data_2[5023:5016];
        layer5[48][7:0] = buffer_data_1[4975:4968];
        layer5[48][15:8] = buffer_data_1[4983:4976];
        layer5[48][23:16] = buffer_data_1[4991:4984];
        layer5[48][31:24] = buffer_data_1[4999:4992];
        layer5[48][39:32] = buffer_data_1[5007:5000];
        layer5[48][47:40] = buffer_data_1[5015:5008];
        layer5[48][55:48] = buffer_data_1[5023:5016];
        layer6[48][7:0] = buffer_data_0[4975:4968];
        layer6[48][15:8] = buffer_data_0[4983:4976];
        layer6[48][23:16] = buffer_data_0[4991:4984];
        layer6[48][31:24] = buffer_data_0[4999:4992];
        layer6[48][39:32] = buffer_data_0[5007:5000];
        layer6[48][47:40] = buffer_data_0[5015:5008];
        layer6[48][55:48] = buffer_data_0[5023:5016];
        layer0[49][7:0] = buffer_data_6[4983:4976];
        layer0[49][15:8] = buffer_data_6[4991:4984];
        layer0[49][23:16] = buffer_data_6[4999:4992];
        layer0[49][31:24] = buffer_data_6[5007:5000];
        layer0[49][39:32] = buffer_data_6[5015:5008];
        layer0[49][47:40] = buffer_data_6[5023:5016];
        layer0[49][55:48] = buffer_data_6[5031:5024];
        layer1[49][7:0] = buffer_data_5[4983:4976];
        layer1[49][15:8] = buffer_data_5[4991:4984];
        layer1[49][23:16] = buffer_data_5[4999:4992];
        layer1[49][31:24] = buffer_data_5[5007:5000];
        layer1[49][39:32] = buffer_data_5[5015:5008];
        layer1[49][47:40] = buffer_data_5[5023:5016];
        layer1[49][55:48] = buffer_data_5[5031:5024];
        layer2[49][7:0] = buffer_data_4[4983:4976];
        layer2[49][15:8] = buffer_data_4[4991:4984];
        layer2[49][23:16] = buffer_data_4[4999:4992];
        layer2[49][31:24] = buffer_data_4[5007:5000];
        layer2[49][39:32] = buffer_data_4[5015:5008];
        layer2[49][47:40] = buffer_data_4[5023:5016];
        layer2[49][55:48] = buffer_data_4[5031:5024];
        layer3[49][7:0] = buffer_data_3[4983:4976];
        layer3[49][15:8] = buffer_data_3[4991:4984];
        layer3[49][23:16] = buffer_data_3[4999:4992];
        layer3[49][31:24] = buffer_data_3[5007:5000];
        layer3[49][39:32] = buffer_data_3[5015:5008];
        layer3[49][47:40] = buffer_data_3[5023:5016];
        layer3[49][55:48] = buffer_data_3[5031:5024];
        layer4[49][7:0] = buffer_data_2[4983:4976];
        layer4[49][15:8] = buffer_data_2[4991:4984];
        layer4[49][23:16] = buffer_data_2[4999:4992];
        layer4[49][31:24] = buffer_data_2[5007:5000];
        layer4[49][39:32] = buffer_data_2[5015:5008];
        layer4[49][47:40] = buffer_data_2[5023:5016];
        layer4[49][55:48] = buffer_data_2[5031:5024];
        layer5[49][7:0] = buffer_data_1[4983:4976];
        layer5[49][15:8] = buffer_data_1[4991:4984];
        layer5[49][23:16] = buffer_data_1[4999:4992];
        layer5[49][31:24] = buffer_data_1[5007:5000];
        layer5[49][39:32] = buffer_data_1[5015:5008];
        layer5[49][47:40] = buffer_data_1[5023:5016];
        layer5[49][55:48] = buffer_data_1[5031:5024];
        layer6[49][7:0] = buffer_data_0[4983:4976];
        layer6[49][15:8] = buffer_data_0[4991:4984];
        layer6[49][23:16] = buffer_data_0[4999:4992];
        layer6[49][31:24] = buffer_data_0[5007:5000];
        layer6[49][39:32] = buffer_data_0[5015:5008];
        layer6[49][47:40] = buffer_data_0[5023:5016];
        layer6[49][55:48] = buffer_data_0[5031:5024];
        layer0[50][7:0] = buffer_data_6[4991:4984];
        layer0[50][15:8] = buffer_data_6[4999:4992];
        layer0[50][23:16] = buffer_data_6[5007:5000];
        layer0[50][31:24] = buffer_data_6[5015:5008];
        layer0[50][39:32] = buffer_data_6[5023:5016];
        layer0[50][47:40] = buffer_data_6[5031:5024];
        layer0[50][55:48] = buffer_data_6[5039:5032];
        layer1[50][7:0] = buffer_data_5[4991:4984];
        layer1[50][15:8] = buffer_data_5[4999:4992];
        layer1[50][23:16] = buffer_data_5[5007:5000];
        layer1[50][31:24] = buffer_data_5[5015:5008];
        layer1[50][39:32] = buffer_data_5[5023:5016];
        layer1[50][47:40] = buffer_data_5[5031:5024];
        layer1[50][55:48] = buffer_data_5[5039:5032];
        layer2[50][7:0] = buffer_data_4[4991:4984];
        layer2[50][15:8] = buffer_data_4[4999:4992];
        layer2[50][23:16] = buffer_data_4[5007:5000];
        layer2[50][31:24] = buffer_data_4[5015:5008];
        layer2[50][39:32] = buffer_data_4[5023:5016];
        layer2[50][47:40] = buffer_data_4[5031:5024];
        layer2[50][55:48] = buffer_data_4[5039:5032];
        layer3[50][7:0] = buffer_data_3[4991:4984];
        layer3[50][15:8] = buffer_data_3[4999:4992];
        layer3[50][23:16] = buffer_data_3[5007:5000];
        layer3[50][31:24] = buffer_data_3[5015:5008];
        layer3[50][39:32] = buffer_data_3[5023:5016];
        layer3[50][47:40] = buffer_data_3[5031:5024];
        layer3[50][55:48] = buffer_data_3[5039:5032];
        layer4[50][7:0] = buffer_data_2[4991:4984];
        layer4[50][15:8] = buffer_data_2[4999:4992];
        layer4[50][23:16] = buffer_data_2[5007:5000];
        layer4[50][31:24] = buffer_data_2[5015:5008];
        layer4[50][39:32] = buffer_data_2[5023:5016];
        layer4[50][47:40] = buffer_data_2[5031:5024];
        layer4[50][55:48] = buffer_data_2[5039:5032];
        layer5[50][7:0] = buffer_data_1[4991:4984];
        layer5[50][15:8] = buffer_data_1[4999:4992];
        layer5[50][23:16] = buffer_data_1[5007:5000];
        layer5[50][31:24] = buffer_data_1[5015:5008];
        layer5[50][39:32] = buffer_data_1[5023:5016];
        layer5[50][47:40] = buffer_data_1[5031:5024];
        layer5[50][55:48] = buffer_data_1[5039:5032];
        layer6[50][7:0] = buffer_data_0[4991:4984];
        layer6[50][15:8] = buffer_data_0[4999:4992];
        layer6[50][23:16] = buffer_data_0[5007:5000];
        layer6[50][31:24] = buffer_data_0[5015:5008];
        layer6[50][39:32] = buffer_data_0[5023:5016];
        layer6[50][47:40] = buffer_data_0[5031:5024];
        layer6[50][55:48] = buffer_data_0[5039:5032];
        layer0[51][7:0] = buffer_data_6[4999:4992];
        layer0[51][15:8] = buffer_data_6[5007:5000];
        layer0[51][23:16] = buffer_data_6[5015:5008];
        layer0[51][31:24] = buffer_data_6[5023:5016];
        layer0[51][39:32] = buffer_data_6[5031:5024];
        layer0[51][47:40] = buffer_data_6[5039:5032];
        layer0[51][55:48] = buffer_data_6[5047:5040];
        layer1[51][7:0] = buffer_data_5[4999:4992];
        layer1[51][15:8] = buffer_data_5[5007:5000];
        layer1[51][23:16] = buffer_data_5[5015:5008];
        layer1[51][31:24] = buffer_data_5[5023:5016];
        layer1[51][39:32] = buffer_data_5[5031:5024];
        layer1[51][47:40] = buffer_data_5[5039:5032];
        layer1[51][55:48] = buffer_data_5[5047:5040];
        layer2[51][7:0] = buffer_data_4[4999:4992];
        layer2[51][15:8] = buffer_data_4[5007:5000];
        layer2[51][23:16] = buffer_data_4[5015:5008];
        layer2[51][31:24] = buffer_data_4[5023:5016];
        layer2[51][39:32] = buffer_data_4[5031:5024];
        layer2[51][47:40] = buffer_data_4[5039:5032];
        layer2[51][55:48] = buffer_data_4[5047:5040];
        layer3[51][7:0] = buffer_data_3[4999:4992];
        layer3[51][15:8] = buffer_data_3[5007:5000];
        layer3[51][23:16] = buffer_data_3[5015:5008];
        layer3[51][31:24] = buffer_data_3[5023:5016];
        layer3[51][39:32] = buffer_data_3[5031:5024];
        layer3[51][47:40] = buffer_data_3[5039:5032];
        layer3[51][55:48] = buffer_data_3[5047:5040];
        layer4[51][7:0] = buffer_data_2[4999:4992];
        layer4[51][15:8] = buffer_data_2[5007:5000];
        layer4[51][23:16] = buffer_data_2[5015:5008];
        layer4[51][31:24] = buffer_data_2[5023:5016];
        layer4[51][39:32] = buffer_data_2[5031:5024];
        layer4[51][47:40] = buffer_data_2[5039:5032];
        layer4[51][55:48] = buffer_data_2[5047:5040];
        layer5[51][7:0] = buffer_data_1[4999:4992];
        layer5[51][15:8] = buffer_data_1[5007:5000];
        layer5[51][23:16] = buffer_data_1[5015:5008];
        layer5[51][31:24] = buffer_data_1[5023:5016];
        layer5[51][39:32] = buffer_data_1[5031:5024];
        layer5[51][47:40] = buffer_data_1[5039:5032];
        layer5[51][55:48] = buffer_data_1[5047:5040];
        layer6[51][7:0] = buffer_data_0[4999:4992];
        layer6[51][15:8] = buffer_data_0[5007:5000];
        layer6[51][23:16] = buffer_data_0[5015:5008];
        layer6[51][31:24] = buffer_data_0[5023:5016];
        layer6[51][39:32] = buffer_data_0[5031:5024];
        layer6[51][47:40] = buffer_data_0[5039:5032];
        layer6[51][55:48] = buffer_data_0[5047:5040];
        layer0[52][7:0] = buffer_data_6[5007:5000];
        layer0[52][15:8] = buffer_data_6[5015:5008];
        layer0[52][23:16] = buffer_data_6[5023:5016];
        layer0[52][31:24] = buffer_data_6[5031:5024];
        layer0[52][39:32] = buffer_data_6[5039:5032];
        layer0[52][47:40] = buffer_data_6[5047:5040];
        layer0[52][55:48] = buffer_data_6[5055:5048];
        layer1[52][7:0] = buffer_data_5[5007:5000];
        layer1[52][15:8] = buffer_data_5[5015:5008];
        layer1[52][23:16] = buffer_data_5[5023:5016];
        layer1[52][31:24] = buffer_data_5[5031:5024];
        layer1[52][39:32] = buffer_data_5[5039:5032];
        layer1[52][47:40] = buffer_data_5[5047:5040];
        layer1[52][55:48] = buffer_data_5[5055:5048];
        layer2[52][7:0] = buffer_data_4[5007:5000];
        layer2[52][15:8] = buffer_data_4[5015:5008];
        layer2[52][23:16] = buffer_data_4[5023:5016];
        layer2[52][31:24] = buffer_data_4[5031:5024];
        layer2[52][39:32] = buffer_data_4[5039:5032];
        layer2[52][47:40] = buffer_data_4[5047:5040];
        layer2[52][55:48] = buffer_data_4[5055:5048];
        layer3[52][7:0] = buffer_data_3[5007:5000];
        layer3[52][15:8] = buffer_data_3[5015:5008];
        layer3[52][23:16] = buffer_data_3[5023:5016];
        layer3[52][31:24] = buffer_data_3[5031:5024];
        layer3[52][39:32] = buffer_data_3[5039:5032];
        layer3[52][47:40] = buffer_data_3[5047:5040];
        layer3[52][55:48] = buffer_data_3[5055:5048];
        layer4[52][7:0] = buffer_data_2[5007:5000];
        layer4[52][15:8] = buffer_data_2[5015:5008];
        layer4[52][23:16] = buffer_data_2[5023:5016];
        layer4[52][31:24] = buffer_data_2[5031:5024];
        layer4[52][39:32] = buffer_data_2[5039:5032];
        layer4[52][47:40] = buffer_data_2[5047:5040];
        layer4[52][55:48] = buffer_data_2[5055:5048];
        layer5[52][7:0] = buffer_data_1[5007:5000];
        layer5[52][15:8] = buffer_data_1[5015:5008];
        layer5[52][23:16] = buffer_data_1[5023:5016];
        layer5[52][31:24] = buffer_data_1[5031:5024];
        layer5[52][39:32] = buffer_data_1[5039:5032];
        layer5[52][47:40] = buffer_data_1[5047:5040];
        layer5[52][55:48] = buffer_data_1[5055:5048];
        layer6[52][7:0] = buffer_data_0[5007:5000];
        layer6[52][15:8] = buffer_data_0[5015:5008];
        layer6[52][23:16] = buffer_data_0[5023:5016];
        layer6[52][31:24] = buffer_data_0[5031:5024];
        layer6[52][39:32] = buffer_data_0[5039:5032];
        layer6[52][47:40] = buffer_data_0[5047:5040];
        layer6[52][55:48] = buffer_data_0[5055:5048];
        layer0[53][7:0] = buffer_data_6[5015:5008];
        layer0[53][15:8] = buffer_data_6[5023:5016];
        layer0[53][23:16] = buffer_data_6[5031:5024];
        layer0[53][31:24] = buffer_data_6[5039:5032];
        layer0[53][39:32] = buffer_data_6[5047:5040];
        layer0[53][47:40] = buffer_data_6[5055:5048];
        layer0[53][55:48] = buffer_data_6[5063:5056];
        layer1[53][7:0] = buffer_data_5[5015:5008];
        layer1[53][15:8] = buffer_data_5[5023:5016];
        layer1[53][23:16] = buffer_data_5[5031:5024];
        layer1[53][31:24] = buffer_data_5[5039:5032];
        layer1[53][39:32] = buffer_data_5[5047:5040];
        layer1[53][47:40] = buffer_data_5[5055:5048];
        layer1[53][55:48] = buffer_data_5[5063:5056];
        layer2[53][7:0] = buffer_data_4[5015:5008];
        layer2[53][15:8] = buffer_data_4[5023:5016];
        layer2[53][23:16] = buffer_data_4[5031:5024];
        layer2[53][31:24] = buffer_data_4[5039:5032];
        layer2[53][39:32] = buffer_data_4[5047:5040];
        layer2[53][47:40] = buffer_data_4[5055:5048];
        layer2[53][55:48] = buffer_data_4[5063:5056];
        layer3[53][7:0] = buffer_data_3[5015:5008];
        layer3[53][15:8] = buffer_data_3[5023:5016];
        layer3[53][23:16] = buffer_data_3[5031:5024];
        layer3[53][31:24] = buffer_data_3[5039:5032];
        layer3[53][39:32] = buffer_data_3[5047:5040];
        layer3[53][47:40] = buffer_data_3[5055:5048];
        layer3[53][55:48] = buffer_data_3[5063:5056];
        layer4[53][7:0] = buffer_data_2[5015:5008];
        layer4[53][15:8] = buffer_data_2[5023:5016];
        layer4[53][23:16] = buffer_data_2[5031:5024];
        layer4[53][31:24] = buffer_data_2[5039:5032];
        layer4[53][39:32] = buffer_data_2[5047:5040];
        layer4[53][47:40] = buffer_data_2[5055:5048];
        layer4[53][55:48] = buffer_data_2[5063:5056];
        layer5[53][7:0] = buffer_data_1[5015:5008];
        layer5[53][15:8] = buffer_data_1[5023:5016];
        layer5[53][23:16] = buffer_data_1[5031:5024];
        layer5[53][31:24] = buffer_data_1[5039:5032];
        layer5[53][39:32] = buffer_data_1[5047:5040];
        layer5[53][47:40] = buffer_data_1[5055:5048];
        layer5[53][55:48] = buffer_data_1[5063:5056];
        layer6[53][7:0] = buffer_data_0[5015:5008];
        layer6[53][15:8] = buffer_data_0[5023:5016];
        layer6[53][23:16] = buffer_data_0[5031:5024];
        layer6[53][31:24] = buffer_data_0[5039:5032];
        layer6[53][39:32] = buffer_data_0[5047:5040];
        layer6[53][47:40] = buffer_data_0[5055:5048];
        layer6[53][55:48] = buffer_data_0[5063:5056];
        layer0[54][7:0] = buffer_data_6[5023:5016];
        layer0[54][15:8] = buffer_data_6[5031:5024];
        layer0[54][23:16] = buffer_data_6[5039:5032];
        layer0[54][31:24] = buffer_data_6[5047:5040];
        layer0[54][39:32] = buffer_data_6[5055:5048];
        layer0[54][47:40] = buffer_data_6[5063:5056];
        layer0[54][55:48] = buffer_data_6[5071:5064];
        layer1[54][7:0] = buffer_data_5[5023:5016];
        layer1[54][15:8] = buffer_data_5[5031:5024];
        layer1[54][23:16] = buffer_data_5[5039:5032];
        layer1[54][31:24] = buffer_data_5[5047:5040];
        layer1[54][39:32] = buffer_data_5[5055:5048];
        layer1[54][47:40] = buffer_data_5[5063:5056];
        layer1[54][55:48] = buffer_data_5[5071:5064];
        layer2[54][7:0] = buffer_data_4[5023:5016];
        layer2[54][15:8] = buffer_data_4[5031:5024];
        layer2[54][23:16] = buffer_data_4[5039:5032];
        layer2[54][31:24] = buffer_data_4[5047:5040];
        layer2[54][39:32] = buffer_data_4[5055:5048];
        layer2[54][47:40] = buffer_data_4[5063:5056];
        layer2[54][55:48] = buffer_data_4[5071:5064];
        layer3[54][7:0] = buffer_data_3[5023:5016];
        layer3[54][15:8] = buffer_data_3[5031:5024];
        layer3[54][23:16] = buffer_data_3[5039:5032];
        layer3[54][31:24] = buffer_data_3[5047:5040];
        layer3[54][39:32] = buffer_data_3[5055:5048];
        layer3[54][47:40] = buffer_data_3[5063:5056];
        layer3[54][55:48] = buffer_data_3[5071:5064];
        layer4[54][7:0] = buffer_data_2[5023:5016];
        layer4[54][15:8] = buffer_data_2[5031:5024];
        layer4[54][23:16] = buffer_data_2[5039:5032];
        layer4[54][31:24] = buffer_data_2[5047:5040];
        layer4[54][39:32] = buffer_data_2[5055:5048];
        layer4[54][47:40] = buffer_data_2[5063:5056];
        layer4[54][55:48] = buffer_data_2[5071:5064];
        layer5[54][7:0] = buffer_data_1[5023:5016];
        layer5[54][15:8] = buffer_data_1[5031:5024];
        layer5[54][23:16] = buffer_data_1[5039:5032];
        layer5[54][31:24] = buffer_data_1[5047:5040];
        layer5[54][39:32] = buffer_data_1[5055:5048];
        layer5[54][47:40] = buffer_data_1[5063:5056];
        layer5[54][55:48] = buffer_data_1[5071:5064];
        layer6[54][7:0] = buffer_data_0[5023:5016];
        layer6[54][15:8] = buffer_data_0[5031:5024];
        layer6[54][23:16] = buffer_data_0[5039:5032];
        layer6[54][31:24] = buffer_data_0[5047:5040];
        layer6[54][39:32] = buffer_data_0[5055:5048];
        layer6[54][47:40] = buffer_data_0[5063:5056];
        layer6[54][55:48] = buffer_data_0[5071:5064];
        layer0[55][7:0] = buffer_data_6[5031:5024];
        layer0[55][15:8] = buffer_data_6[5039:5032];
        layer0[55][23:16] = buffer_data_6[5047:5040];
        layer0[55][31:24] = buffer_data_6[5055:5048];
        layer0[55][39:32] = buffer_data_6[5063:5056];
        layer0[55][47:40] = buffer_data_6[5071:5064];
        layer0[55][55:48] = buffer_data_6[5079:5072];
        layer1[55][7:0] = buffer_data_5[5031:5024];
        layer1[55][15:8] = buffer_data_5[5039:5032];
        layer1[55][23:16] = buffer_data_5[5047:5040];
        layer1[55][31:24] = buffer_data_5[5055:5048];
        layer1[55][39:32] = buffer_data_5[5063:5056];
        layer1[55][47:40] = buffer_data_5[5071:5064];
        layer1[55][55:48] = buffer_data_5[5079:5072];
        layer2[55][7:0] = buffer_data_4[5031:5024];
        layer2[55][15:8] = buffer_data_4[5039:5032];
        layer2[55][23:16] = buffer_data_4[5047:5040];
        layer2[55][31:24] = buffer_data_4[5055:5048];
        layer2[55][39:32] = buffer_data_4[5063:5056];
        layer2[55][47:40] = buffer_data_4[5071:5064];
        layer2[55][55:48] = buffer_data_4[5079:5072];
        layer3[55][7:0] = buffer_data_3[5031:5024];
        layer3[55][15:8] = buffer_data_3[5039:5032];
        layer3[55][23:16] = buffer_data_3[5047:5040];
        layer3[55][31:24] = buffer_data_3[5055:5048];
        layer3[55][39:32] = buffer_data_3[5063:5056];
        layer3[55][47:40] = buffer_data_3[5071:5064];
        layer3[55][55:48] = buffer_data_3[5079:5072];
        layer4[55][7:0] = buffer_data_2[5031:5024];
        layer4[55][15:8] = buffer_data_2[5039:5032];
        layer4[55][23:16] = buffer_data_2[5047:5040];
        layer4[55][31:24] = buffer_data_2[5055:5048];
        layer4[55][39:32] = buffer_data_2[5063:5056];
        layer4[55][47:40] = buffer_data_2[5071:5064];
        layer4[55][55:48] = buffer_data_2[5079:5072];
        layer5[55][7:0] = buffer_data_1[5031:5024];
        layer5[55][15:8] = buffer_data_1[5039:5032];
        layer5[55][23:16] = buffer_data_1[5047:5040];
        layer5[55][31:24] = buffer_data_1[5055:5048];
        layer5[55][39:32] = buffer_data_1[5063:5056];
        layer5[55][47:40] = buffer_data_1[5071:5064];
        layer5[55][55:48] = buffer_data_1[5079:5072];
        layer6[55][7:0] = buffer_data_0[5031:5024];
        layer6[55][15:8] = buffer_data_0[5039:5032];
        layer6[55][23:16] = buffer_data_0[5047:5040];
        layer6[55][31:24] = buffer_data_0[5055:5048];
        layer6[55][39:32] = buffer_data_0[5063:5056];
        layer6[55][47:40] = buffer_data_0[5071:5064];
        layer6[55][55:48] = buffer_data_0[5079:5072];
        layer0[56][7:0] = buffer_data_6[5039:5032];
        layer0[56][15:8] = buffer_data_6[5047:5040];
        layer0[56][23:16] = buffer_data_6[5055:5048];
        layer0[56][31:24] = buffer_data_6[5063:5056];
        layer0[56][39:32] = buffer_data_6[5071:5064];
        layer0[56][47:40] = buffer_data_6[5079:5072];
        layer0[56][55:48] = buffer_data_6[5087:5080];
        layer1[56][7:0] = buffer_data_5[5039:5032];
        layer1[56][15:8] = buffer_data_5[5047:5040];
        layer1[56][23:16] = buffer_data_5[5055:5048];
        layer1[56][31:24] = buffer_data_5[5063:5056];
        layer1[56][39:32] = buffer_data_5[5071:5064];
        layer1[56][47:40] = buffer_data_5[5079:5072];
        layer1[56][55:48] = buffer_data_5[5087:5080];
        layer2[56][7:0] = buffer_data_4[5039:5032];
        layer2[56][15:8] = buffer_data_4[5047:5040];
        layer2[56][23:16] = buffer_data_4[5055:5048];
        layer2[56][31:24] = buffer_data_4[5063:5056];
        layer2[56][39:32] = buffer_data_4[5071:5064];
        layer2[56][47:40] = buffer_data_4[5079:5072];
        layer2[56][55:48] = buffer_data_4[5087:5080];
        layer3[56][7:0] = buffer_data_3[5039:5032];
        layer3[56][15:8] = buffer_data_3[5047:5040];
        layer3[56][23:16] = buffer_data_3[5055:5048];
        layer3[56][31:24] = buffer_data_3[5063:5056];
        layer3[56][39:32] = buffer_data_3[5071:5064];
        layer3[56][47:40] = buffer_data_3[5079:5072];
        layer3[56][55:48] = buffer_data_3[5087:5080];
        layer4[56][7:0] = buffer_data_2[5039:5032];
        layer4[56][15:8] = buffer_data_2[5047:5040];
        layer4[56][23:16] = buffer_data_2[5055:5048];
        layer4[56][31:24] = buffer_data_2[5063:5056];
        layer4[56][39:32] = buffer_data_2[5071:5064];
        layer4[56][47:40] = buffer_data_2[5079:5072];
        layer4[56][55:48] = buffer_data_2[5087:5080];
        layer5[56][7:0] = buffer_data_1[5039:5032];
        layer5[56][15:8] = buffer_data_1[5047:5040];
        layer5[56][23:16] = buffer_data_1[5055:5048];
        layer5[56][31:24] = buffer_data_1[5063:5056];
        layer5[56][39:32] = buffer_data_1[5071:5064];
        layer5[56][47:40] = buffer_data_1[5079:5072];
        layer5[56][55:48] = buffer_data_1[5087:5080];
        layer6[56][7:0] = buffer_data_0[5039:5032];
        layer6[56][15:8] = buffer_data_0[5047:5040];
        layer6[56][23:16] = buffer_data_0[5055:5048];
        layer6[56][31:24] = buffer_data_0[5063:5056];
        layer6[56][39:32] = buffer_data_0[5071:5064];
        layer6[56][47:40] = buffer_data_0[5079:5072];
        layer6[56][55:48] = buffer_data_0[5087:5080];
        layer0[57][7:0] = buffer_data_6[5047:5040];
        layer0[57][15:8] = buffer_data_6[5055:5048];
        layer0[57][23:16] = buffer_data_6[5063:5056];
        layer0[57][31:24] = buffer_data_6[5071:5064];
        layer0[57][39:32] = buffer_data_6[5079:5072];
        layer0[57][47:40] = buffer_data_6[5087:5080];
        layer0[57][55:48] = buffer_data_6[5095:5088];
        layer1[57][7:0] = buffer_data_5[5047:5040];
        layer1[57][15:8] = buffer_data_5[5055:5048];
        layer1[57][23:16] = buffer_data_5[5063:5056];
        layer1[57][31:24] = buffer_data_5[5071:5064];
        layer1[57][39:32] = buffer_data_5[5079:5072];
        layer1[57][47:40] = buffer_data_5[5087:5080];
        layer1[57][55:48] = buffer_data_5[5095:5088];
        layer2[57][7:0] = buffer_data_4[5047:5040];
        layer2[57][15:8] = buffer_data_4[5055:5048];
        layer2[57][23:16] = buffer_data_4[5063:5056];
        layer2[57][31:24] = buffer_data_4[5071:5064];
        layer2[57][39:32] = buffer_data_4[5079:5072];
        layer2[57][47:40] = buffer_data_4[5087:5080];
        layer2[57][55:48] = buffer_data_4[5095:5088];
        layer3[57][7:0] = buffer_data_3[5047:5040];
        layer3[57][15:8] = buffer_data_3[5055:5048];
        layer3[57][23:16] = buffer_data_3[5063:5056];
        layer3[57][31:24] = buffer_data_3[5071:5064];
        layer3[57][39:32] = buffer_data_3[5079:5072];
        layer3[57][47:40] = buffer_data_3[5087:5080];
        layer3[57][55:48] = buffer_data_3[5095:5088];
        layer4[57][7:0] = buffer_data_2[5047:5040];
        layer4[57][15:8] = buffer_data_2[5055:5048];
        layer4[57][23:16] = buffer_data_2[5063:5056];
        layer4[57][31:24] = buffer_data_2[5071:5064];
        layer4[57][39:32] = buffer_data_2[5079:5072];
        layer4[57][47:40] = buffer_data_2[5087:5080];
        layer4[57][55:48] = buffer_data_2[5095:5088];
        layer5[57][7:0] = buffer_data_1[5047:5040];
        layer5[57][15:8] = buffer_data_1[5055:5048];
        layer5[57][23:16] = buffer_data_1[5063:5056];
        layer5[57][31:24] = buffer_data_1[5071:5064];
        layer5[57][39:32] = buffer_data_1[5079:5072];
        layer5[57][47:40] = buffer_data_1[5087:5080];
        layer5[57][55:48] = buffer_data_1[5095:5088];
        layer6[57][7:0] = buffer_data_0[5047:5040];
        layer6[57][15:8] = buffer_data_0[5055:5048];
        layer6[57][23:16] = buffer_data_0[5063:5056];
        layer6[57][31:24] = buffer_data_0[5071:5064];
        layer6[57][39:32] = buffer_data_0[5079:5072];
        layer6[57][47:40] = buffer_data_0[5087:5080];
        layer6[57][55:48] = buffer_data_0[5095:5088];
        layer0[58][7:0] = buffer_data_6[5055:5048];
        layer0[58][15:8] = buffer_data_6[5063:5056];
        layer0[58][23:16] = buffer_data_6[5071:5064];
        layer0[58][31:24] = buffer_data_6[5079:5072];
        layer0[58][39:32] = buffer_data_6[5087:5080];
        layer0[58][47:40] = buffer_data_6[5095:5088];
        layer0[58][55:48] = buffer_data_6[5103:5096];
        layer1[58][7:0] = buffer_data_5[5055:5048];
        layer1[58][15:8] = buffer_data_5[5063:5056];
        layer1[58][23:16] = buffer_data_5[5071:5064];
        layer1[58][31:24] = buffer_data_5[5079:5072];
        layer1[58][39:32] = buffer_data_5[5087:5080];
        layer1[58][47:40] = buffer_data_5[5095:5088];
        layer1[58][55:48] = buffer_data_5[5103:5096];
        layer2[58][7:0] = buffer_data_4[5055:5048];
        layer2[58][15:8] = buffer_data_4[5063:5056];
        layer2[58][23:16] = buffer_data_4[5071:5064];
        layer2[58][31:24] = buffer_data_4[5079:5072];
        layer2[58][39:32] = buffer_data_4[5087:5080];
        layer2[58][47:40] = buffer_data_4[5095:5088];
        layer2[58][55:48] = buffer_data_4[5103:5096];
        layer3[58][7:0] = buffer_data_3[5055:5048];
        layer3[58][15:8] = buffer_data_3[5063:5056];
        layer3[58][23:16] = buffer_data_3[5071:5064];
        layer3[58][31:24] = buffer_data_3[5079:5072];
        layer3[58][39:32] = buffer_data_3[5087:5080];
        layer3[58][47:40] = buffer_data_3[5095:5088];
        layer3[58][55:48] = buffer_data_3[5103:5096];
        layer4[58][7:0] = buffer_data_2[5055:5048];
        layer4[58][15:8] = buffer_data_2[5063:5056];
        layer4[58][23:16] = buffer_data_2[5071:5064];
        layer4[58][31:24] = buffer_data_2[5079:5072];
        layer4[58][39:32] = buffer_data_2[5087:5080];
        layer4[58][47:40] = buffer_data_2[5095:5088];
        layer4[58][55:48] = buffer_data_2[5103:5096];
        layer5[58][7:0] = buffer_data_1[5055:5048];
        layer5[58][15:8] = buffer_data_1[5063:5056];
        layer5[58][23:16] = buffer_data_1[5071:5064];
        layer5[58][31:24] = buffer_data_1[5079:5072];
        layer5[58][39:32] = buffer_data_1[5087:5080];
        layer5[58][47:40] = buffer_data_1[5095:5088];
        layer5[58][55:48] = buffer_data_1[5103:5096];
        layer6[58][7:0] = buffer_data_0[5055:5048];
        layer6[58][15:8] = buffer_data_0[5063:5056];
        layer6[58][23:16] = buffer_data_0[5071:5064];
        layer6[58][31:24] = buffer_data_0[5079:5072];
        layer6[58][39:32] = buffer_data_0[5087:5080];
        layer6[58][47:40] = buffer_data_0[5095:5088];
        layer6[58][55:48] = buffer_data_0[5103:5096];
        layer0[59][7:0] = buffer_data_6[5063:5056];
        layer0[59][15:8] = buffer_data_6[5071:5064];
        layer0[59][23:16] = buffer_data_6[5079:5072];
        layer0[59][31:24] = buffer_data_6[5087:5080];
        layer0[59][39:32] = buffer_data_6[5095:5088];
        layer0[59][47:40] = buffer_data_6[5103:5096];
        layer0[59][55:48] = buffer_data_6[5111:5104];
        layer1[59][7:0] = buffer_data_5[5063:5056];
        layer1[59][15:8] = buffer_data_5[5071:5064];
        layer1[59][23:16] = buffer_data_5[5079:5072];
        layer1[59][31:24] = buffer_data_5[5087:5080];
        layer1[59][39:32] = buffer_data_5[5095:5088];
        layer1[59][47:40] = buffer_data_5[5103:5096];
        layer1[59][55:48] = buffer_data_5[5111:5104];
        layer2[59][7:0] = buffer_data_4[5063:5056];
        layer2[59][15:8] = buffer_data_4[5071:5064];
        layer2[59][23:16] = buffer_data_4[5079:5072];
        layer2[59][31:24] = buffer_data_4[5087:5080];
        layer2[59][39:32] = buffer_data_4[5095:5088];
        layer2[59][47:40] = buffer_data_4[5103:5096];
        layer2[59][55:48] = buffer_data_4[5111:5104];
        layer3[59][7:0] = buffer_data_3[5063:5056];
        layer3[59][15:8] = buffer_data_3[5071:5064];
        layer3[59][23:16] = buffer_data_3[5079:5072];
        layer3[59][31:24] = buffer_data_3[5087:5080];
        layer3[59][39:32] = buffer_data_3[5095:5088];
        layer3[59][47:40] = buffer_data_3[5103:5096];
        layer3[59][55:48] = buffer_data_3[5111:5104];
        layer4[59][7:0] = buffer_data_2[5063:5056];
        layer4[59][15:8] = buffer_data_2[5071:5064];
        layer4[59][23:16] = buffer_data_2[5079:5072];
        layer4[59][31:24] = buffer_data_2[5087:5080];
        layer4[59][39:32] = buffer_data_2[5095:5088];
        layer4[59][47:40] = buffer_data_2[5103:5096];
        layer4[59][55:48] = buffer_data_2[5111:5104];
        layer5[59][7:0] = buffer_data_1[5063:5056];
        layer5[59][15:8] = buffer_data_1[5071:5064];
        layer5[59][23:16] = buffer_data_1[5079:5072];
        layer5[59][31:24] = buffer_data_1[5087:5080];
        layer5[59][39:32] = buffer_data_1[5095:5088];
        layer5[59][47:40] = buffer_data_1[5103:5096];
        layer5[59][55:48] = buffer_data_1[5111:5104];
        layer6[59][7:0] = buffer_data_0[5063:5056];
        layer6[59][15:8] = buffer_data_0[5071:5064];
        layer6[59][23:16] = buffer_data_0[5079:5072];
        layer6[59][31:24] = buffer_data_0[5087:5080];
        layer6[59][39:32] = buffer_data_0[5095:5088];
        layer6[59][47:40] = buffer_data_0[5103:5096];
        layer6[59][55:48] = buffer_data_0[5111:5104];
        layer0[60][7:0] = buffer_data_6[5071:5064];
        layer0[60][15:8] = buffer_data_6[5079:5072];
        layer0[60][23:16] = buffer_data_6[5087:5080];
        layer0[60][31:24] = buffer_data_6[5095:5088];
        layer0[60][39:32] = buffer_data_6[5103:5096];
        layer0[60][47:40] = buffer_data_6[5111:5104];
        layer0[60][55:48] = buffer_data_6[5119:5112];
        layer1[60][7:0] = buffer_data_5[5071:5064];
        layer1[60][15:8] = buffer_data_5[5079:5072];
        layer1[60][23:16] = buffer_data_5[5087:5080];
        layer1[60][31:24] = buffer_data_5[5095:5088];
        layer1[60][39:32] = buffer_data_5[5103:5096];
        layer1[60][47:40] = buffer_data_5[5111:5104];
        layer1[60][55:48] = buffer_data_5[5119:5112];
        layer2[60][7:0] = buffer_data_4[5071:5064];
        layer2[60][15:8] = buffer_data_4[5079:5072];
        layer2[60][23:16] = buffer_data_4[5087:5080];
        layer2[60][31:24] = buffer_data_4[5095:5088];
        layer2[60][39:32] = buffer_data_4[5103:5096];
        layer2[60][47:40] = buffer_data_4[5111:5104];
        layer2[60][55:48] = buffer_data_4[5119:5112];
        layer3[60][7:0] = buffer_data_3[5071:5064];
        layer3[60][15:8] = buffer_data_3[5079:5072];
        layer3[60][23:16] = buffer_data_3[5087:5080];
        layer3[60][31:24] = buffer_data_3[5095:5088];
        layer3[60][39:32] = buffer_data_3[5103:5096];
        layer3[60][47:40] = buffer_data_3[5111:5104];
        layer3[60][55:48] = buffer_data_3[5119:5112];
        layer4[60][7:0] = buffer_data_2[5071:5064];
        layer4[60][15:8] = buffer_data_2[5079:5072];
        layer4[60][23:16] = buffer_data_2[5087:5080];
        layer4[60][31:24] = buffer_data_2[5095:5088];
        layer4[60][39:32] = buffer_data_2[5103:5096];
        layer4[60][47:40] = buffer_data_2[5111:5104];
        layer4[60][55:48] = buffer_data_2[5119:5112];
        layer5[60][7:0] = buffer_data_1[5071:5064];
        layer5[60][15:8] = buffer_data_1[5079:5072];
        layer5[60][23:16] = buffer_data_1[5087:5080];
        layer5[60][31:24] = buffer_data_1[5095:5088];
        layer5[60][39:32] = buffer_data_1[5103:5096];
        layer5[60][47:40] = buffer_data_1[5111:5104];
        layer5[60][55:48] = buffer_data_1[5119:5112];
        layer6[60][7:0] = buffer_data_0[5071:5064];
        layer6[60][15:8] = buffer_data_0[5079:5072];
        layer6[60][23:16] = buffer_data_0[5087:5080];
        layer6[60][31:24] = buffer_data_0[5095:5088];
        layer6[60][39:32] = buffer_data_0[5103:5096];
        layer6[60][47:40] = buffer_data_0[5111:5104];
        layer6[60][55:48] = buffer_data_0[5119:5112];
        layer0[61][7:0] = buffer_data_6[5079:5072];
        layer0[61][15:8] = buffer_data_6[5087:5080];
        layer0[61][23:16] = buffer_data_6[5095:5088];
        layer0[61][31:24] = buffer_data_6[5103:5096];
        layer0[61][39:32] = 0;
        layer0[61][47:40] = 0;
        layer0[61][55:48] = 0;
        layer1[61][7:0] = buffer_data_5[5079:5072];
        layer1[61][15:8] = buffer_data_5[5087:5080];
        layer1[61][23:16] = buffer_data_5[5095:5088];
        layer1[61][31:24] = buffer_data_5[5103:5096];
        layer1[61][39:32] = 0;
        layer1[61][47:40] = 0;
        layer1[61][55:48] = 0;
        layer2[61][7:0] = buffer_data_4[5079:5072];
        layer2[61][15:8] = buffer_data_4[5087:5080];
        layer2[61][23:16] = buffer_data_4[5095:5088];
        layer2[61][31:24] = buffer_data_4[5103:5096];
        layer2[61][39:32] = 0;
        layer2[61][47:40] = 0;
        layer2[61][55:48] = 0;
        layer3[61][7:0] = buffer_data_3[5079:5072];
        layer3[61][15:8] = buffer_data_3[5087:5080];
        layer3[61][23:16] = buffer_data_3[5095:5088];
        layer3[61][31:24] = buffer_data_3[5103:5096];
        layer3[61][39:32] = 0;
        layer3[61][47:40] = 0;
        layer3[61][55:48] = 0;
        layer4[61][7:0] = buffer_data_2[5079:5072];
        layer4[61][15:8] = buffer_data_2[5087:5080];
        layer4[61][23:16] = buffer_data_2[5095:5088];
        layer4[61][31:24] = buffer_data_2[5103:5096];
        layer4[61][39:32] = 0;
        layer4[61][47:40] = 0;
        layer4[61][55:48] = 0;
        layer5[61][7:0] = buffer_data_1[5079:5072];
        layer5[61][15:8] = buffer_data_1[5087:5080];
        layer5[61][23:16] = buffer_data_1[5095:5088];
        layer5[61][31:24] = buffer_data_1[5103:5096];
        layer5[61][39:32] = 0;
        layer5[61][47:40] = 0;
        layer5[61][55:48] = 0;
        layer6[61][7:0] = buffer_data_0[5079:5072];
        layer6[61][15:8] = buffer_data_0[5087:5080];
        layer6[61][23:16] = buffer_data_0[5095:5088];
        layer6[61][31:24] = buffer_data_0[5103:5096];
        layer6[61][39:32] = 0;
        layer6[61][47:40] = 0;
        layer6[61][55:48] = 0;
        layer0[62][7:0] = buffer_data_6[5087:5080];
        layer0[62][15:8] = buffer_data_6[5095:5088];
        layer0[62][23:16] = buffer_data_6[5103:5096];
        layer0[62][31:24] = 0;
        layer0[62][39:32] = 0;
        layer0[62][47:40] = 0;
        layer0[62][55:48] = 0;
        layer1[62][7:0] = buffer_data_5[5087:5080];
        layer1[62][15:8] = buffer_data_5[5095:5088];
        layer1[62][23:16] = buffer_data_5[5103:5096];
        layer1[62][31:24] = 0;
        layer1[62][39:32] = 0;
        layer1[62][47:40] = 0;
        layer1[62][55:48] = 0;
        layer2[62][7:0] = buffer_data_4[5087:5080];
        layer2[62][15:8] = buffer_data_4[5095:5088];
        layer2[62][23:16] = buffer_data_4[5103:5096];
        layer2[62][31:24] = 0;
        layer2[62][39:32] = 0;
        layer2[62][47:40] = 0;
        layer2[62][55:48] = 0;
        layer3[62][7:0] = buffer_data_3[5087:5080];
        layer3[62][15:8] = buffer_data_3[5095:5088];
        layer3[62][23:16] = buffer_data_3[5103:5096];
        layer3[62][31:24] = 0;
        layer3[62][39:32] = 0;
        layer3[62][47:40] = 0;
        layer3[62][55:48] = 0;
        layer4[62][7:0] = buffer_data_2[5087:5080];
        layer4[62][15:8] = buffer_data_2[5095:5088];
        layer4[62][23:16] = buffer_data_2[5103:5096];
        layer4[62][31:24] = 0;
        layer4[62][39:32] = 0;
        layer4[62][47:40] = 0;
        layer4[62][55:48] = 0;
        layer5[62][7:0] = buffer_data_1[5087:5080];
        layer5[62][15:8] = buffer_data_1[5095:5088];
        layer5[62][23:16] = buffer_data_1[5103:5096];
        layer5[62][31:24] = 0;
        layer5[62][39:32] = 0;
        layer5[62][47:40] = 0;
        layer5[62][55:48] = 0;
        layer6[62][7:0] = buffer_data_0[5087:5080];
        layer6[62][15:8] = buffer_data_0[5095:5088];
        layer6[62][23:16] = buffer_data_0[5103:5096];
        layer6[62][31:24] = 0;
        layer6[62][39:32] = 0;
        layer6[62][47:40] = 0;
        layer6[62][55:48] = 0;
        layer0[63][7:0] = buffer_data_6[5095:5088];
        layer0[63][15:8] = buffer_data_6[5103:5096];
        layer0[63][23:16] = 0;
        layer0[63][31:24] = 0;
        layer0[63][39:32] = 0;
        layer0[63][47:40] = 0;
        layer0[63][55:48] = 0;
        layer1[63][7:0] = buffer_data_5[5095:5088];
        layer1[63][15:8] = buffer_data_5[5103:5096];
        layer1[63][23:16] = 0;
        layer1[63][31:24] = 0;
        layer1[63][39:32] = 0;
        layer1[63][47:40] = 0;
        layer1[63][55:48] = 0;
        layer2[63][7:0] = buffer_data_4[5095:5088];
        layer2[63][15:8] = buffer_data_4[5103:5096];
        layer2[63][23:16] = 0;
        layer2[63][31:24] = 0;
        layer2[63][39:32] = 0;
        layer2[63][47:40] = 0;
        layer2[63][55:48] = 0;
        layer3[63][7:0] = buffer_data_3[5095:5088];
        layer3[63][15:8] = buffer_data_3[5103:5096];
        layer3[63][23:16] = 0;
        layer3[63][31:24] = 0;
        layer3[63][39:32] = 0;
        layer3[63][47:40] = 0;
        layer3[63][55:48] = 0;
        layer4[63][7:0] = buffer_data_2[5095:5088];
        layer4[63][15:8] = buffer_data_2[5103:5096];
        layer4[63][23:16] = 0;
        layer4[63][31:24] = 0;
        layer4[63][39:32] = 0;
        layer4[63][47:40] = 0;
        layer4[63][55:48] = 0;
        layer5[63][7:0] = buffer_data_1[5095:5088];
        layer5[63][15:8] = buffer_data_1[5103:5096];
        layer5[63][23:16] = 0;
        layer5[63][31:24] = 0;
        layer5[63][39:32] = 0;
        layer5[63][47:40] = 0;
        layer5[63][55:48] = 0;
        layer6[63][7:0] = buffer_data_0[5095:5088];
        layer6[63][15:8] = buffer_data_0[5103:5096];
        layer6[63][23:16] = 0;
        layer6[63][31:24] = 0;
        layer6[63][39:32] = 0;
        layer6[63][47:40] = 0;
        layer6[63][55:48] = 0;
    end
  endcase
end

wire  [39:0]  kernel_img_mul_0[0:48];
assign kernel_img_mul_0[0] = layer0[0][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_0[1] = layer0[0][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_0[2] = layer0[0][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_0[3] = layer0[0][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_0[4] = layer0[0][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_0[5] = layer0[0][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_0[6] = layer0[0][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_0[7] = layer1[0][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_0[8] = layer1[0][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_0[9] = layer1[0][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_0[10] = layer1[0][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_0[11] = layer1[0][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_0[12] = layer1[0][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_0[13] = layer1[0][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_0[14] = layer2[0][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_0[15] = layer2[0][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_0[16] = layer2[0][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_0[17] = layer2[0][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_0[18] = layer2[0][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_0[19] = layer2[0][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_0[20] = layer2[0][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_0[21] = layer3[0][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_0[22] = layer3[0][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_0[23] = layer3[0][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_0[24] = layer3[0][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_0[25] = layer3[0][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_0[26] = layer3[0][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_0[27] = layer3[0][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_0[28] = layer4[0][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_0[29] = layer4[0][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_0[30] = layer4[0][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_0[31] = layer4[0][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_0[32] = layer4[0][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_0[33] = layer4[0][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_0[34] = layer4[0][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_0[35] = layer5[0][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_0[36] = layer5[0][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_0[37] = layer5[0][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_0[38] = layer5[0][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_0[39] = layer5[0][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_0[40] = layer5[0][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_0[41] = layer5[0][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_0[42] = layer6[0][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_0[43] = layer6[0][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_0[44] = layer6[0][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_0[45] = layer6[0][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_0[46] = layer6[0][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_0[47] = layer6[0][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_0[48] = layer6[0][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_0 = kernel_img_mul_0[0] + kernel_img_mul_0[1] + kernel_img_mul_0[2] + 
                kernel_img_mul_0[3] + kernel_img_mul_0[4] + kernel_img_mul_0[5] + 
                kernel_img_mul_0[6] + kernel_img_mul_0[7] + kernel_img_mul_0[8] + 
                kernel_img_mul_0[9] + kernel_img_mul_0[10] + kernel_img_mul_0[11] + 
                kernel_img_mul_0[12] + kernel_img_mul_0[13] + kernel_img_mul_0[14] + 
                kernel_img_mul_0[15] + kernel_img_mul_0[16] + kernel_img_mul_0[17] + 
                kernel_img_mul_0[18] + kernel_img_mul_0[19] + kernel_img_mul_0[20] + 
                kernel_img_mul_0[21] + kernel_img_mul_0[22] + kernel_img_mul_0[23] + 
                kernel_img_mul_0[24] + kernel_img_mul_0[25] + kernel_img_mul_0[26] + 
                kernel_img_mul_0[27] + kernel_img_mul_0[28] + kernel_img_mul_0[29] + 
                kernel_img_mul_0[30] + kernel_img_mul_0[31] + kernel_img_mul_0[32] + 
                kernel_img_mul_0[33] + kernel_img_mul_0[34] + kernel_img_mul_0[35] + 
                kernel_img_mul_0[36] + kernel_img_mul_0[37] + kernel_img_mul_0[38] + 
                kernel_img_mul_0[39] + kernel_img_mul_0[40] + kernel_img_mul_0[41] + 
                kernel_img_mul_0[42] + kernel_img_mul_0[43] + kernel_img_mul_0[44] + 
                kernel_img_mul_0[45] + kernel_img_mul_0[46] + kernel_img_mul_0[47] + 
                kernel_img_mul_0[48];
wire  [39:0]  kernel_img_mul_1[0:48];
assign kernel_img_mul_1[0] = layer0[1][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_1[1] = layer0[1][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_1[2] = layer0[1][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_1[3] = layer0[1][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_1[4] = layer0[1][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_1[5] = layer0[1][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_1[6] = layer0[1][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_1[7] = layer1[1][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_1[8] = layer1[1][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_1[9] = layer1[1][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_1[10] = layer1[1][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_1[11] = layer1[1][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_1[12] = layer1[1][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_1[13] = layer1[1][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_1[14] = layer2[1][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_1[15] = layer2[1][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_1[16] = layer2[1][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_1[17] = layer2[1][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_1[18] = layer2[1][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_1[19] = layer2[1][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_1[20] = layer2[1][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_1[21] = layer3[1][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_1[22] = layer3[1][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_1[23] = layer3[1][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_1[24] = layer3[1][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_1[25] = layer3[1][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_1[26] = layer3[1][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_1[27] = layer3[1][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_1[28] = layer4[1][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_1[29] = layer4[1][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_1[30] = layer4[1][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_1[31] = layer4[1][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_1[32] = layer4[1][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_1[33] = layer4[1][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_1[34] = layer4[1][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_1[35] = layer5[1][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_1[36] = layer5[1][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_1[37] = layer5[1][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_1[38] = layer5[1][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_1[39] = layer5[1][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_1[40] = layer5[1][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_1[41] = layer5[1][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_1[42] = layer6[1][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_1[43] = layer6[1][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_1[44] = layer6[1][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_1[45] = layer6[1][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_1[46] = layer6[1][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_1[47] = layer6[1][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_1[48] = layer6[1][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_1 = kernel_img_mul_1[0] + kernel_img_mul_1[1] + kernel_img_mul_1[2] + 
                kernel_img_mul_1[3] + kernel_img_mul_1[4] + kernel_img_mul_1[5] + 
                kernel_img_mul_1[6] + kernel_img_mul_1[7] + kernel_img_mul_1[8] + 
                kernel_img_mul_1[9] + kernel_img_mul_1[10] + kernel_img_mul_1[11] + 
                kernel_img_mul_1[12] + kernel_img_mul_1[13] + kernel_img_mul_1[14] + 
                kernel_img_mul_1[15] + kernel_img_mul_1[16] + kernel_img_mul_1[17] + 
                kernel_img_mul_1[18] + kernel_img_mul_1[19] + kernel_img_mul_1[20] + 
                kernel_img_mul_1[21] + kernel_img_mul_1[22] + kernel_img_mul_1[23] + 
                kernel_img_mul_1[24] + kernel_img_mul_1[25] + kernel_img_mul_1[26] + 
                kernel_img_mul_1[27] + kernel_img_mul_1[28] + kernel_img_mul_1[29] + 
                kernel_img_mul_1[30] + kernel_img_mul_1[31] + kernel_img_mul_1[32] + 
                kernel_img_mul_1[33] + kernel_img_mul_1[34] + kernel_img_mul_1[35] + 
                kernel_img_mul_1[36] + kernel_img_mul_1[37] + kernel_img_mul_1[38] + 
                kernel_img_mul_1[39] + kernel_img_mul_1[40] + kernel_img_mul_1[41] + 
                kernel_img_mul_1[42] + kernel_img_mul_1[43] + kernel_img_mul_1[44] + 
                kernel_img_mul_1[45] + kernel_img_mul_1[46] + kernel_img_mul_1[47] + 
                kernel_img_mul_1[48];
wire  [39:0]  kernel_img_mul_2[0:48];
assign kernel_img_mul_2[0] = layer0[2][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_2[1] = layer0[2][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_2[2] = layer0[2][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_2[3] = layer0[2][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_2[4] = layer0[2][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_2[5] = layer0[2][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_2[6] = layer0[2][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_2[7] = layer1[2][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_2[8] = layer1[2][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_2[9] = layer1[2][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_2[10] = layer1[2][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_2[11] = layer1[2][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_2[12] = layer1[2][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_2[13] = layer1[2][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_2[14] = layer2[2][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_2[15] = layer2[2][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_2[16] = layer2[2][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_2[17] = layer2[2][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_2[18] = layer2[2][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_2[19] = layer2[2][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_2[20] = layer2[2][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_2[21] = layer3[2][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_2[22] = layer3[2][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_2[23] = layer3[2][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_2[24] = layer3[2][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_2[25] = layer3[2][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_2[26] = layer3[2][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_2[27] = layer3[2][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_2[28] = layer4[2][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_2[29] = layer4[2][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_2[30] = layer4[2][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_2[31] = layer4[2][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_2[32] = layer4[2][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_2[33] = layer4[2][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_2[34] = layer4[2][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_2[35] = layer5[2][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_2[36] = layer5[2][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_2[37] = layer5[2][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_2[38] = layer5[2][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_2[39] = layer5[2][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_2[40] = layer5[2][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_2[41] = layer5[2][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_2[42] = layer6[2][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_2[43] = layer6[2][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_2[44] = layer6[2][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_2[45] = layer6[2][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_2[46] = layer6[2][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_2[47] = layer6[2][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_2[48] = layer6[2][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_2 = kernel_img_mul_2[0] + kernel_img_mul_2[1] + kernel_img_mul_2[2] + 
                kernel_img_mul_2[3] + kernel_img_mul_2[4] + kernel_img_mul_2[5] + 
                kernel_img_mul_2[6] + kernel_img_mul_2[7] + kernel_img_mul_2[8] + 
                kernel_img_mul_2[9] + kernel_img_mul_2[10] + kernel_img_mul_2[11] + 
                kernel_img_mul_2[12] + kernel_img_mul_2[13] + kernel_img_mul_2[14] + 
                kernel_img_mul_2[15] + kernel_img_mul_2[16] + kernel_img_mul_2[17] + 
                kernel_img_mul_2[18] + kernel_img_mul_2[19] + kernel_img_mul_2[20] + 
                kernel_img_mul_2[21] + kernel_img_mul_2[22] + kernel_img_mul_2[23] + 
                kernel_img_mul_2[24] + kernel_img_mul_2[25] + kernel_img_mul_2[26] + 
                kernel_img_mul_2[27] + kernel_img_mul_2[28] + kernel_img_mul_2[29] + 
                kernel_img_mul_2[30] + kernel_img_mul_2[31] + kernel_img_mul_2[32] + 
                kernel_img_mul_2[33] + kernel_img_mul_2[34] + kernel_img_mul_2[35] + 
                kernel_img_mul_2[36] + kernel_img_mul_2[37] + kernel_img_mul_2[38] + 
                kernel_img_mul_2[39] + kernel_img_mul_2[40] + kernel_img_mul_2[41] + 
                kernel_img_mul_2[42] + kernel_img_mul_2[43] + kernel_img_mul_2[44] + 
                kernel_img_mul_2[45] + kernel_img_mul_2[46] + kernel_img_mul_2[47] + 
                kernel_img_mul_2[48];
wire  [39:0]  kernel_img_mul_3[0:48];
assign kernel_img_mul_3[0] = layer0[3][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_3[1] = layer0[3][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_3[2] = layer0[3][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_3[3] = layer0[3][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_3[4] = layer0[3][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_3[5] = layer0[3][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_3[6] = layer0[3][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_3[7] = layer1[3][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_3[8] = layer1[3][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_3[9] = layer1[3][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_3[10] = layer1[3][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_3[11] = layer1[3][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_3[12] = layer1[3][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_3[13] = layer1[3][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_3[14] = layer2[3][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_3[15] = layer2[3][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_3[16] = layer2[3][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_3[17] = layer2[3][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_3[18] = layer2[3][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_3[19] = layer2[3][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_3[20] = layer2[3][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_3[21] = layer3[3][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_3[22] = layer3[3][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_3[23] = layer3[3][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_3[24] = layer3[3][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_3[25] = layer3[3][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_3[26] = layer3[3][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_3[27] = layer3[3][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_3[28] = layer4[3][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_3[29] = layer4[3][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_3[30] = layer4[3][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_3[31] = layer4[3][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_3[32] = layer4[3][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_3[33] = layer4[3][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_3[34] = layer4[3][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_3[35] = layer5[3][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_3[36] = layer5[3][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_3[37] = layer5[3][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_3[38] = layer5[3][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_3[39] = layer5[3][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_3[40] = layer5[3][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_3[41] = layer5[3][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_3[42] = layer6[3][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_3[43] = layer6[3][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_3[44] = layer6[3][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_3[45] = layer6[3][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_3[46] = layer6[3][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_3[47] = layer6[3][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_3[48] = layer6[3][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_3 = kernel_img_mul_3[0] + kernel_img_mul_3[1] + kernel_img_mul_3[2] + 
                kernel_img_mul_3[3] + kernel_img_mul_3[4] + kernel_img_mul_3[5] + 
                kernel_img_mul_3[6] + kernel_img_mul_3[7] + kernel_img_mul_3[8] + 
                kernel_img_mul_3[9] + kernel_img_mul_3[10] + kernel_img_mul_3[11] + 
                kernel_img_mul_3[12] + kernel_img_mul_3[13] + kernel_img_mul_3[14] + 
                kernel_img_mul_3[15] + kernel_img_mul_3[16] + kernel_img_mul_3[17] + 
                kernel_img_mul_3[18] + kernel_img_mul_3[19] + kernel_img_mul_3[20] + 
                kernel_img_mul_3[21] + kernel_img_mul_3[22] + kernel_img_mul_3[23] + 
                kernel_img_mul_3[24] + kernel_img_mul_3[25] + kernel_img_mul_3[26] + 
                kernel_img_mul_3[27] + kernel_img_mul_3[28] + kernel_img_mul_3[29] + 
                kernel_img_mul_3[30] + kernel_img_mul_3[31] + kernel_img_mul_3[32] + 
                kernel_img_mul_3[33] + kernel_img_mul_3[34] + kernel_img_mul_3[35] + 
                kernel_img_mul_3[36] + kernel_img_mul_3[37] + kernel_img_mul_3[38] + 
                kernel_img_mul_3[39] + kernel_img_mul_3[40] + kernel_img_mul_3[41] + 
                kernel_img_mul_3[42] + kernel_img_mul_3[43] + kernel_img_mul_3[44] + 
                kernel_img_mul_3[45] + kernel_img_mul_3[46] + kernel_img_mul_3[47] + 
                kernel_img_mul_3[48];
wire  [39:0]  kernel_img_mul_4[0:48];
assign kernel_img_mul_4[0] = layer0[4][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_4[1] = layer0[4][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_4[2] = layer0[4][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_4[3] = layer0[4][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_4[4] = layer0[4][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_4[5] = layer0[4][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_4[6] = layer0[4][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_4[7] = layer1[4][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_4[8] = layer1[4][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_4[9] = layer1[4][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_4[10] = layer1[4][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_4[11] = layer1[4][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_4[12] = layer1[4][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_4[13] = layer1[4][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_4[14] = layer2[4][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_4[15] = layer2[4][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_4[16] = layer2[4][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_4[17] = layer2[4][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_4[18] = layer2[4][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_4[19] = layer2[4][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_4[20] = layer2[4][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_4[21] = layer3[4][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_4[22] = layer3[4][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_4[23] = layer3[4][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_4[24] = layer3[4][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_4[25] = layer3[4][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_4[26] = layer3[4][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_4[27] = layer3[4][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_4[28] = layer4[4][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_4[29] = layer4[4][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_4[30] = layer4[4][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_4[31] = layer4[4][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_4[32] = layer4[4][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_4[33] = layer4[4][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_4[34] = layer4[4][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_4[35] = layer5[4][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_4[36] = layer5[4][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_4[37] = layer5[4][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_4[38] = layer5[4][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_4[39] = layer5[4][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_4[40] = layer5[4][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_4[41] = layer5[4][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_4[42] = layer6[4][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_4[43] = layer6[4][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_4[44] = layer6[4][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_4[45] = layer6[4][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_4[46] = layer6[4][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_4[47] = layer6[4][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_4[48] = layer6[4][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_4 = kernel_img_mul_4[0] + kernel_img_mul_4[1] + kernel_img_mul_4[2] + 
                kernel_img_mul_4[3] + kernel_img_mul_4[4] + kernel_img_mul_4[5] + 
                kernel_img_mul_4[6] + kernel_img_mul_4[7] + kernel_img_mul_4[8] + 
                kernel_img_mul_4[9] + kernel_img_mul_4[10] + kernel_img_mul_4[11] + 
                kernel_img_mul_4[12] + kernel_img_mul_4[13] + kernel_img_mul_4[14] + 
                kernel_img_mul_4[15] + kernel_img_mul_4[16] + kernel_img_mul_4[17] + 
                kernel_img_mul_4[18] + kernel_img_mul_4[19] + kernel_img_mul_4[20] + 
                kernel_img_mul_4[21] + kernel_img_mul_4[22] + kernel_img_mul_4[23] + 
                kernel_img_mul_4[24] + kernel_img_mul_4[25] + kernel_img_mul_4[26] + 
                kernel_img_mul_4[27] + kernel_img_mul_4[28] + kernel_img_mul_4[29] + 
                kernel_img_mul_4[30] + kernel_img_mul_4[31] + kernel_img_mul_4[32] + 
                kernel_img_mul_4[33] + kernel_img_mul_4[34] + kernel_img_mul_4[35] + 
                kernel_img_mul_4[36] + kernel_img_mul_4[37] + kernel_img_mul_4[38] + 
                kernel_img_mul_4[39] + kernel_img_mul_4[40] + kernel_img_mul_4[41] + 
                kernel_img_mul_4[42] + kernel_img_mul_4[43] + kernel_img_mul_4[44] + 
                kernel_img_mul_4[45] + kernel_img_mul_4[46] + kernel_img_mul_4[47] + 
                kernel_img_mul_4[48];
wire  [39:0]  kernel_img_mul_5[0:48];
assign kernel_img_mul_5[0] = layer0[5][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_5[1] = layer0[5][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_5[2] = layer0[5][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_5[3] = layer0[5][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_5[4] = layer0[5][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_5[5] = layer0[5][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_5[6] = layer0[5][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_5[7] = layer1[5][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_5[8] = layer1[5][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_5[9] = layer1[5][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_5[10] = layer1[5][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_5[11] = layer1[5][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_5[12] = layer1[5][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_5[13] = layer1[5][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_5[14] = layer2[5][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_5[15] = layer2[5][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_5[16] = layer2[5][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_5[17] = layer2[5][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_5[18] = layer2[5][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_5[19] = layer2[5][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_5[20] = layer2[5][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_5[21] = layer3[5][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_5[22] = layer3[5][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_5[23] = layer3[5][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_5[24] = layer3[5][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_5[25] = layer3[5][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_5[26] = layer3[5][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_5[27] = layer3[5][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_5[28] = layer4[5][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_5[29] = layer4[5][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_5[30] = layer4[5][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_5[31] = layer4[5][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_5[32] = layer4[5][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_5[33] = layer4[5][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_5[34] = layer4[5][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_5[35] = layer5[5][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_5[36] = layer5[5][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_5[37] = layer5[5][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_5[38] = layer5[5][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_5[39] = layer5[5][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_5[40] = layer5[5][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_5[41] = layer5[5][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_5[42] = layer6[5][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_5[43] = layer6[5][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_5[44] = layer6[5][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_5[45] = layer6[5][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_5[46] = layer6[5][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_5[47] = layer6[5][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_5[48] = layer6[5][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_5 = kernel_img_mul_5[0] + kernel_img_mul_5[1] + kernel_img_mul_5[2] + 
                kernel_img_mul_5[3] + kernel_img_mul_5[4] + kernel_img_mul_5[5] + 
                kernel_img_mul_5[6] + kernel_img_mul_5[7] + kernel_img_mul_5[8] + 
                kernel_img_mul_5[9] + kernel_img_mul_5[10] + kernel_img_mul_5[11] + 
                kernel_img_mul_5[12] + kernel_img_mul_5[13] + kernel_img_mul_5[14] + 
                kernel_img_mul_5[15] + kernel_img_mul_5[16] + kernel_img_mul_5[17] + 
                kernel_img_mul_5[18] + kernel_img_mul_5[19] + kernel_img_mul_5[20] + 
                kernel_img_mul_5[21] + kernel_img_mul_5[22] + kernel_img_mul_5[23] + 
                kernel_img_mul_5[24] + kernel_img_mul_5[25] + kernel_img_mul_5[26] + 
                kernel_img_mul_5[27] + kernel_img_mul_5[28] + kernel_img_mul_5[29] + 
                kernel_img_mul_5[30] + kernel_img_mul_5[31] + kernel_img_mul_5[32] + 
                kernel_img_mul_5[33] + kernel_img_mul_5[34] + kernel_img_mul_5[35] + 
                kernel_img_mul_5[36] + kernel_img_mul_5[37] + kernel_img_mul_5[38] + 
                kernel_img_mul_5[39] + kernel_img_mul_5[40] + kernel_img_mul_5[41] + 
                kernel_img_mul_5[42] + kernel_img_mul_5[43] + kernel_img_mul_5[44] + 
                kernel_img_mul_5[45] + kernel_img_mul_5[46] + kernel_img_mul_5[47] + 
                kernel_img_mul_5[48];
wire  [39:0]  kernel_img_mul_6[0:48];
assign kernel_img_mul_6[0] = layer0[6][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_6[1] = layer0[6][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_6[2] = layer0[6][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_6[3] = layer0[6][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_6[4] = layer0[6][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_6[5] = layer0[6][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_6[6] = layer0[6][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_6[7] = layer1[6][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_6[8] = layer1[6][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_6[9] = layer1[6][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_6[10] = layer1[6][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_6[11] = layer1[6][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_6[12] = layer1[6][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_6[13] = layer1[6][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_6[14] = layer2[6][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_6[15] = layer2[6][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_6[16] = layer2[6][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_6[17] = layer2[6][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_6[18] = layer2[6][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_6[19] = layer2[6][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_6[20] = layer2[6][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_6[21] = layer3[6][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_6[22] = layer3[6][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_6[23] = layer3[6][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_6[24] = layer3[6][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_6[25] = layer3[6][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_6[26] = layer3[6][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_6[27] = layer3[6][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_6[28] = layer4[6][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_6[29] = layer4[6][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_6[30] = layer4[6][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_6[31] = layer4[6][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_6[32] = layer4[6][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_6[33] = layer4[6][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_6[34] = layer4[6][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_6[35] = layer5[6][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_6[36] = layer5[6][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_6[37] = layer5[6][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_6[38] = layer5[6][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_6[39] = layer5[6][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_6[40] = layer5[6][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_6[41] = layer5[6][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_6[42] = layer6[6][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_6[43] = layer6[6][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_6[44] = layer6[6][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_6[45] = layer6[6][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_6[46] = layer6[6][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_6[47] = layer6[6][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_6[48] = layer6[6][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_6 = kernel_img_mul_6[0] + kernel_img_mul_6[1] + kernel_img_mul_6[2] + 
                kernel_img_mul_6[3] + kernel_img_mul_6[4] + kernel_img_mul_6[5] + 
                kernel_img_mul_6[6] + kernel_img_mul_6[7] + kernel_img_mul_6[8] + 
                kernel_img_mul_6[9] + kernel_img_mul_6[10] + kernel_img_mul_6[11] + 
                kernel_img_mul_6[12] + kernel_img_mul_6[13] + kernel_img_mul_6[14] + 
                kernel_img_mul_6[15] + kernel_img_mul_6[16] + kernel_img_mul_6[17] + 
                kernel_img_mul_6[18] + kernel_img_mul_6[19] + kernel_img_mul_6[20] + 
                kernel_img_mul_6[21] + kernel_img_mul_6[22] + kernel_img_mul_6[23] + 
                kernel_img_mul_6[24] + kernel_img_mul_6[25] + kernel_img_mul_6[26] + 
                kernel_img_mul_6[27] + kernel_img_mul_6[28] + kernel_img_mul_6[29] + 
                kernel_img_mul_6[30] + kernel_img_mul_6[31] + kernel_img_mul_6[32] + 
                kernel_img_mul_6[33] + kernel_img_mul_6[34] + kernel_img_mul_6[35] + 
                kernel_img_mul_6[36] + kernel_img_mul_6[37] + kernel_img_mul_6[38] + 
                kernel_img_mul_6[39] + kernel_img_mul_6[40] + kernel_img_mul_6[41] + 
                kernel_img_mul_6[42] + kernel_img_mul_6[43] + kernel_img_mul_6[44] + 
                kernel_img_mul_6[45] + kernel_img_mul_6[46] + kernel_img_mul_6[47] + 
                kernel_img_mul_6[48];
wire  [39:0]  kernel_img_mul_7[0:48];
assign kernel_img_mul_7[0] = layer0[7][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_7[1] = layer0[7][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_7[2] = layer0[7][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_7[3] = layer0[7][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_7[4] = layer0[7][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_7[5] = layer0[7][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_7[6] = layer0[7][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_7[7] = layer1[7][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_7[8] = layer1[7][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_7[9] = layer1[7][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_7[10] = layer1[7][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_7[11] = layer1[7][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_7[12] = layer1[7][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_7[13] = layer1[7][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_7[14] = layer2[7][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_7[15] = layer2[7][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_7[16] = layer2[7][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_7[17] = layer2[7][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_7[18] = layer2[7][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_7[19] = layer2[7][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_7[20] = layer2[7][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_7[21] = layer3[7][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_7[22] = layer3[7][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_7[23] = layer3[7][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_7[24] = layer3[7][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_7[25] = layer3[7][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_7[26] = layer3[7][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_7[27] = layer3[7][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_7[28] = layer4[7][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_7[29] = layer4[7][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_7[30] = layer4[7][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_7[31] = layer4[7][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_7[32] = layer4[7][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_7[33] = layer4[7][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_7[34] = layer4[7][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_7[35] = layer5[7][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_7[36] = layer5[7][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_7[37] = layer5[7][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_7[38] = layer5[7][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_7[39] = layer5[7][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_7[40] = layer5[7][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_7[41] = layer5[7][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_7[42] = layer6[7][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_7[43] = layer6[7][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_7[44] = layer6[7][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_7[45] = layer6[7][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_7[46] = layer6[7][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_7[47] = layer6[7][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_7[48] = layer6[7][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_7 = kernel_img_mul_7[0] + kernel_img_mul_7[1] + kernel_img_mul_7[2] + 
                kernel_img_mul_7[3] + kernel_img_mul_7[4] + kernel_img_mul_7[5] + 
                kernel_img_mul_7[6] + kernel_img_mul_7[7] + kernel_img_mul_7[8] + 
                kernel_img_mul_7[9] + kernel_img_mul_7[10] + kernel_img_mul_7[11] + 
                kernel_img_mul_7[12] + kernel_img_mul_7[13] + kernel_img_mul_7[14] + 
                kernel_img_mul_7[15] + kernel_img_mul_7[16] + kernel_img_mul_7[17] + 
                kernel_img_mul_7[18] + kernel_img_mul_7[19] + kernel_img_mul_7[20] + 
                kernel_img_mul_7[21] + kernel_img_mul_7[22] + kernel_img_mul_7[23] + 
                kernel_img_mul_7[24] + kernel_img_mul_7[25] + kernel_img_mul_7[26] + 
                kernel_img_mul_7[27] + kernel_img_mul_7[28] + kernel_img_mul_7[29] + 
                kernel_img_mul_7[30] + kernel_img_mul_7[31] + kernel_img_mul_7[32] + 
                kernel_img_mul_7[33] + kernel_img_mul_7[34] + kernel_img_mul_7[35] + 
                kernel_img_mul_7[36] + kernel_img_mul_7[37] + kernel_img_mul_7[38] + 
                kernel_img_mul_7[39] + kernel_img_mul_7[40] + kernel_img_mul_7[41] + 
                kernel_img_mul_7[42] + kernel_img_mul_7[43] + kernel_img_mul_7[44] + 
                kernel_img_mul_7[45] + kernel_img_mul_7[46] + kernel_img_mul_7[47] + 
                kernel_img_mul_7[48];
wire  [39:0]  kernel_img_mul_8[0:48];
assign kernel_img_mul_8[0] = layer0[8][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_8[1] = layer0[8][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_8[2] = layer0[8][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_8[3] = layer0[8][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_8[4] = layer0[8][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_8[5] = layer0[8][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_8[6] = layer0[8][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_8[7] = layer1[8][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_8[8] = layer1[8][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_8[9] = layer1[8][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_8[10] = layer1[8][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_8[11] = layer1[8][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_8[12] = layer1[8][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_8[13] = layer1[8][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_8[14] = layer2[8][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_8[15] = layer2[8][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_8[16] = layer2[8][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_8[17] = layer2[8][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_8[18] = layer2[8][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_8[19] = layer2[8][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_8[20] = layer2[8][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_8[21] = layer3[8][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_8[22] = layer3[8][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_8[23] = layer3[8][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_8[24] = layer3[8][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_8[25] = layer3[8][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_8[26] = layer3[8][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_8[27] = layer3[8][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_8[28] = layer4[8][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_8[29] = layer4[8][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_8[30] = layer4[8][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_8[31] = layer4[8][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_8[32] = layer4[8][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_8[33] = layer4[8][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_8[34] = layer4[8][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_8[35] = layer5[8][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_8[36] = layer5[8][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_8[37] = layer5[8][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_8[38] = layer5[8][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_8[39] = layer5[8][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_8[40] = layer5[8][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_8[41] = layer5[8][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_8[42] = layer6[8][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_8[43] = layer6[8][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_8[44] = layer6[8][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_8[45] = layer6[8][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_8[46] = layer6[8][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_8[47] = layer6[8][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_8[48] = layer6[8][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_8 = kernel_img_mul_8[0] + kernel_img_mul_8[1] + kernel_img_mul_8[2] + 
                kernel_img_mul_8[3] + kernel_img_mul_8[4] + kernel_img_mul_8[5] + 
                kernel_img_mul_8[6] + kernel_img_mul_8[7] + kernel_img_mul_8[8] + 
                kernel_img_mul_8[9] + kernel_img_mul_8[10] + kernel_img_mul_8[11] + 
                kernel_img_mul_8[12] + kernel_img_mul_8[13] + kernel_img_mul_8[14] + 
                kernel_img_mul_8[15] + kernel_img_mul_8[16] + kernel_img_mul_8[17] + 
                kernel_img_mul_8[18] + kernel_img_mul_8[19] + kernel_img_mul_8[20] + 
                kernel_img_mul_8[21] + kernel_img_mul_8[22] + kernel_img_mul_8[23] + 
                kernel_img_mul_8[24] + kernel_img_mul_8[25] + kernel_img_mul_8[26] + 
                kernel_img_mul_8[27] + kernel_img_mul_8[28] + kernel_img_mul_8[29] + 
                kernel_img_mul_8[30] + kernel_img_mul_8[31] + kernel_img_mul_8[32] + 
                kernel_img_mul_8[33] + kernel_img_mul_8[34] + kernel_img_mul_8[35] + 
                kernel_img_mul_8[36] + kernel_img_mul_8[37] + kernel_img_mul_8[38] + 
                kernel_img_mul_8[39] + kernel_img_mul_8[40] + kernel_img_mul_8[41] + 
                kernel_img_mul_8[42] + kernel_img_mul_8[43] + kernel_img_mul_8[44] + 
                kernel_img_mul_8[45] + kernel_img_mul_8[46] + kernel_img_mul_8[47] + 
                kernel_img_mul_8[48];
wire  [39:0]  kernel_img_mul_9[0:48];
assign kernel_img_mul_9[0] = layer0[9][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_9[1] = layer0[9][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_9[2] = layer0[9][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_9[3] = layer0[9][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_9[4] = layer0[9][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_9[5] = layer0[9][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_9[6] = layer0[9][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_9[7] = layer1[9][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_9[8] = layer1[9][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_9[9] = layer1[9][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_9[10] = layer1[9][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_9[11] = layer1[9][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_9[12] = layer1[9][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_9[13] = layer1[9][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_9[14] = layer2[9][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_9[15] = layer2[9][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_9[16] = layer2[9][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_9[17] = layer2[9][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_9[18] = layer2[9][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_9[19] = layer2[9][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_9[20] = layer2[9][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_9[21] = layer3[9][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_9[22] = layer3[9][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_9[23] = layer3[9][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_9[24] = layer3[9][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_9[25] = layer3[9][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_9[26] = layer3[9][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_9[27] = layer3[9][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_9[28] = layer4[9][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_9[29] = layer4[9][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_9[30] = layer4[9][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_9[31] = layer4[9][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_9[32] = layer4[9][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_9[33] = layer4[9][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_9[34] = layer4[9][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_9[35] = layer5[9][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_9[36] = layer5[9][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_9[37] = layer5[9][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_9[38] = layer5[9][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_9[39] = layer5[9][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_9[40] = layer5[9][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_9[41] = layer5[9][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_9[42] = layer6[9][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_9[43] = layer6[9][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_9[44] = layer6[9][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_9[45] = layer6[9][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_9[46] = layer6[9][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_9[47] = layer6[9][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_9[48] = layer6[9][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_9 = kernel_img_mul_9[0] + kernel_img_mul_9[1] + kernel_img_mul_9[2] + 
                kernel_img_mul_9[3] + kernel_img_mul_9[4] + kernel_img_mul_9[5] + 
                kernel_img_mul_9[6] + kernel_img_mul_9[7] + kernel_img_mul_9[8] + 
                kernel_img_mul_9[9] + kernel_img_mul_9[10] + kernel_img_mul_9[11] + 
                kernel_img_mul_9[12] + kernel_img_mul_9[13] + kernel_img_mul_9[14] + 
                kernel_img_mul_9[15] + kernel_img_mul_9[16] + kernel_img_mul_9[17] + 
                kernel_img_mul_9[18] + kernel_img_mul_9[19] + kernel_img_mul_9[20] + 
                kernel_img_mul_9[21] + kernel_img_mul_9[22] + kernel_img_mul_9[23] + 
                kernel_img_mul_9[24] + kernel_img_mul_9[25] + kernel_img_mul_9[26] + 
                kernel_img_mul_9[27] + kernel_img_mul_9[28] + kernel_img_mul_9[29] + 
                kernel_img_mul_9[30] + kernel_img_mul_9[31] + kernel_img_mul_9[32] + 
                kernel_img_mul_9[33] + kernel_img_mul_9[34] + kernel_img_mul_9[35] + 
                kernel_img_mul_9[36] + kernel_img_mul_9[37] + kernel_img_mul_9[38] + 
                kernel_img_mul_9[39] + kernel_img_mul_9[40] + kernel_img_mul_9[41] + 
                kernel_img_mul_9[42] + kernel_img_mul_9[43] + kernel_img_mul_9[44] + 
                kernel_img_mul_9[45] + kernel_img_mul_9[46] + kernel_img_mul_9[47] + 
                kernel_img_mul_9[48];
wire  [39:0]  kernel_img_mul_10[0:48];
assign kernel_img_mul_10[0] = layer0[10][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_10[1] = layer0[10][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_10[2] = layer0[10][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_10[3] = layer0[10][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_10[4] = layer0[10][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_10[5] = layer0[10][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_10[6] = layer0[10][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_10[7] = layer1[10][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_10[8] = layer1[10][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_10[9] = layer1[10][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_10[10] = layer1[10][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_10[11] = layer1[10][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_10[12] = layer1[10][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_10[13] = layer1[10][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_10[14] = layer2[10][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_10[15] = layer2[10][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_10[16] = layer2[10][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_10[17] = layer2[10][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_10[18] = layer2[10][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_10[19] = layer2[10][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_10[20] = layer2[10][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_10[21] = layer3[10][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_10[22] = layer3[10][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_10[23] = layer3[10][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_10[24] = layer3[10][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_10[25] = layer3[10][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_10[26] = layer3[10][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_10[27] = layer3[10][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_10[28] = layer4[10][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_10[29] = layer4[10][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_10[30] = layer4[10][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_10[31] = layer4[10][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_10[32] = layer4[10][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_10[33] = layer4[10][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_10[34] = layer4[10][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_10[35] = layer5[10][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_10[36] = layer5[10][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_10[37] = layer5[10][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_10[38] = layer5[10][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_10[39] = layer5[10][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_10[40] = layer5[10][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_10[41] = layer5[10][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_10[42] = layer6[10][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_10[43] = layer6[10][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_10[44] = layer6[10][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_10[45] = layer6[10][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_10[46] = layer6[10][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_10[47] = layer6[10][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_10[48] = layer6[10][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_10 = kernel_img_mul_10[0] + kernel_img_mul_10[1] + kernel_img_mul_10[2] + 
                kernel_img_mul_10[3] + kernel_img_mul_10[4] + kernel_img_mul_10[5] + 
                kernel_img_mul_10[6] + kernel_img_mul_10[7] + kernel_img_mul_10[8] + 
                kernel_img_mul_10[9] + kernel_img_mul_10[10] + kernel_img_mul_10[11] + 
                kernel_img_mul_10[12] + kernel_img_mul_10[13] + kernel_img_mul_10[14] + 
                kernel_img_mul_10[15] + kernel_img_mul_10[16] + kernel_img_mul_10[17] + 
                kernel_img_mul_10[18] + kernel_img_mul_10[19] + kernel_img_mul_10[20] + 
                kernel_img_mul_10[21] + kernel_img_mul_10[22] + kernel_img_mul_10[23] + 
                kernel_img_mul_10[24] + kernel_img_mul_10[25] + kernel_img_mul_10[26] + 
                kernel_img_mul_10[27] + kernel_img_mul_10[28] + kernel_img_mul_10[29] + 
                kernel_img_mul_10[30] + kernel_img_mul_10[31] + kernel_img_mul_10[32] + 
                kernel_img_mul_10[33] + kernel_img_mul_10[34] + kernel_img_mul_10[35] + 
                kernel_img_mul_10[36] + kernel_img_mul_10[37] + kernel_img_mul_10[38] + 
                kernel_img_mul_10[39] + kernel_img_mul_10[40] + kernel_img_mul_10[41] + 
                kernel_img_mul_10[42] + kernel_img_mul_10[43] + kernel_img_mul_10[44] + 
                kernel_img_mul_10[45] + kernel_img_mul_10[46] + kernel_img_mul_10[47] + 
                kernel_img_mul_10[48];
wire  [39:0]  kernel_img_mul_11[0:48];
assign kernel_img_mul_11[0] = layer0[11][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_11[1] = layer0[11][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_11[2] = layer0[11][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_11[3] = layer0[11][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_11[4] = layer0[11][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_11[5] = layer0[11][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_11[6] = layer0[11][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_11[7] = layer1[11][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_11[8] = layer1[11][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_11[9] = layer1[11][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_11[10] = layer1[11][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_11[11] = layer1[11][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_11[12] = layer1[11][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_11[13] = layer1[11][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_11[14] = layer2[11][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_11[15] = layer2[11][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_11[16] = layer2[11][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_11[17] = layer2[11][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_11[18] = layer2[11][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_11[19] = layer2[11][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_11[20] = layer2[11][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_11[21] = layer3[11][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_11[22] = layer3[11][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_11[23] = layer3[11][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_11[24] = layer3[11][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_11[25] = layer3[11][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_11[26] = layer3[11][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_11[27] = layer3[11][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_11[28] = layer4[11][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_11[29] = layer4[11][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_11[30] = layer4[11][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_11[31] = layer4[11][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_11[32] = layer4[11][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_11[33] = layer4[11][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_11[34] = layer4[11][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_11[35] = layer5[11][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_11[36] = layer5[11][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_11[37] = layer5[11][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_11[38] = layer5[11][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_11[39] = layer5[11][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_11[40] = layer5[11][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_11[41] = layer5[11][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_11[42] = layer6[11][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_11[43] = layer6[11][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_11[44] = layer6[11][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_11[45] = layer6[11][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_11[46] = layer6[11][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_11[47] = layer6[11][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_11[48] = layer6[11][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_11 = kernel_img_mul_11[0] + kernel_img_mul_11[1] + kernel_img_mul_11[2] + 
                kernel_img_mul_11[3] + kernel_img_mul_11[4] + kernel_img_mul_11[5] + 
                kernel_img_mul_11[6] + kernel_img_mul_11[7] + kernel_img_mul_11[8] + 
                kernel_img_mul_11[9] + kernel_img_mul_11[10] + kernel_img_mul_11[11] + 
                kernel_img_mul_11[12] + kernel_img_mul_11[13] + kernel_img_mul_11[14] + 
                kernel_img_mul_11[15] + kernel_img_mul_11[16] + kernel_img_mul_11[17] + 
                kernel_img_mul_11[18] + kernel_img_mul_11[19] + kernel_img_mul_11[20] + 
                kernel_img_mul_11[21] + kernel_img_mul_11[22] + kernel_img_mul_11[23] + 
                kernel_img_mul_11[24] + kernel_img_mul_11[25] + kernel_img_mul_11[26] + 
                kernel_img_mul_11[27] + kernel_img_mul_11[28] + kernel_img_mul_11[29] + 
                kernel_img_mul_11[30] + kernel_img_mul_11[31] + kernel_img_mul_11[32] + 
                kernel_img_mul_11[33] + kernel_img_mul_11[34] + kernel_img_mul_11[35] + 
                kernel_img_mul_11[36] + kernel_img_mul_11[37] + kernel_img_mul_11[38] + 
                kernel_img_mul_11[39] + kernel_img_mul_11[40] + kernel_img_mul_11[41] + 
                kernel_img_mul_11[42] + kernel_img_mul_11[43] + kernel_img_mul_11[44] + 
                kernel_img_mul_11[45] + kernel_img_mul_11[46] + kernel_img_mul_11[47] + 
                kernel_img_mul_11[48];
wire  [39:0]  kernel_img_mul_12[0:48];
assign kernel_img_mul_12[0] = layer0[12][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_12[1] = layer0[12][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_12[2] = layer0[12][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_12[3] = layer0[12][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_12[4] = layer0[12][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_12[5] = layer0[12][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_12[6] = layer0[12][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_12[7] = layer1[12][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_12[8] = layer1[12][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_12[9] = layer1[12][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_12[10] = layer1[12][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_12[11] = layer1[12][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_12[12] = layer1[12][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_12[13] = layer1[12][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_12[14] = layer2[12][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_12[15] = layer2[12][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_12[16] = layer2[12][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_12[17] = layer2[12][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_12[18] = layer2[12][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_12[19] = layer2[12][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_12[20] = layer2[12][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_12[21] = layer3[12][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_12[22] = layer3[12][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_12[23] = layer3[12][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_12[24] = layer3[12][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_12[25] = layer3[12][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_12[26] = layer3[12][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_12[27] = layer3[12][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_12[28] = layer4[12][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_12[29] = layer4[12][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_12[30] = layer4[12][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_12[31] = layer4[12][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_12[32] = layer4[12][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_12[33] = layer4[12][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_12[34] = layer4[12][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_12[35] = layer5[12][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_12[36] = layer5[12][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_12[37] = layer5[12][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_12[38] = layer5[12][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_12[39] = layer5[12][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_12[40] = layer5[12][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_12[41] = layer5[12][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_12[42] = layer6[12][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_12[43] = layer6[12][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_12[44] = layer6[12][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_12[45] = layer6[12][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_12[46] = layer6[12][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_12[47] = layer6[12][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_12[48] = layer6[12][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_12 = kernel_img_mul_12[0] + kernel_img_mul_12[1] + kernel_img_mul_12[2] + 
                kernel_img_mul_12[3] + kernel_img_mul_12[4] + kernel_img_mul_12[5] + 
                kernel_img_mul_12[6] + kernel_img_mul_12[7] + kernel_img_mul_12[8] + 
                kernel_img_mul_12[9] + kernel_img_mul_12[10] + kernel_img_mul_12[11] + 
                kernel_img_mul_12[12] + kernel_img_mul_12[13] + kernel_img_mul_12[14] + 
                kernel_img_mul_12[15] + kernel_img_mul_12[16] + kernel_img_mul_12[17] + 
                kernel_img_mul_12[18] + kernel_img_mul_12[19] + kernel_img_mul_12[20] + 
                kernel_img_mul_12[21] + kernel_img_mul_12[22] + kernel_img_mul_12[23] + 
                kernel_img_mul_12[24] + kernel_img_mul_12[25] + kernel_img_mul_12[26] + 
                kernel_img_mul_12[27] + kernel_img_mul_12[28] + kernel_img_mul_12[29] + 
                kernel_img_mul_12[30] + kernel_img_mul_12[31] + kernel_img_mul_12[32] + 
                kernel_img_mul_12[33] + kernel_img_mul_12[34] + kernel_img_mul_12[35] + 
                kernel_img_mul_12[36] + kernel_img_mul_12[37] + kernel_img_mul_12[38] + 
                kernel_img_mul_12[39] + kernel_img_mul_12[40] + kernel_img_mul_12[41] + 
                kernel_img_mul_12[42] + kernel_img_mul_12[43] + kernel_img_mul_12[44] + 
                kernel_img_mul_12[45] + kernel_img_mul_12[46] + kernel_img_mul_12[47] + 
                kernel_img_mul_12[48];
wire  [39:0]  kernel_img_mul_13[0:48];
assign kernel_img_mul_13[0] = layer0[13][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_13[1] = layer0[13][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_13[2] = layer0[13][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_13[3] = layer0[13][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_13[4] = layer0[13][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_13[5] = layer0[13][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_13[6] = layer0[13][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_13[7] = layer1[13][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_13[8] = layer1[13][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_13[9] = layer1[13][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_13[10] = layer1[13][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_13[11] = layer1[13][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_13[12] = layer1[13][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_13[13] = layer1[13][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_13[14] = layer2[13][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_13[15] = layer2[13][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_13[16] = layer2[13][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_13[17] = layer2[13][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_13[18] = layer2[13][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_13[19] = layer2[13][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_13[20] = layer2[13][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_13[21] = layer3[13][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_13[22] = layer3[13][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_13[23] = layer3[13][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_13[24] = layer3[13][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_13[25] = layer3[13][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_13[26] = layer3[13][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_13[27] = layer3[13][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_13[28] = layer4[13][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_13[29] = layer4[13][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_13[30] = layer4[13][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_13[31] = layer4[13][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_13[32] = layer4[13][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_13[33] = layer4[13][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_13[34] = layer4[13][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_13[35] = layer5[13][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_13[36] = layer5[13][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_13[37] = layer5[13][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_13[38] = layer5[13][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_13[39] = layer5[13][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_13[40] = layer5[13][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_13[41] = layer5[13][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_13[42] = layer6[13][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_13[43] = layer6[13][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_13[44] = layer6[13][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_13[45] = layer6[13][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_13[46] = layer6[13][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_13[47] = layer6[13][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_13[48] = layer6[13][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_13 = kernel_img_mul_13[0] + kernel_img_mul_13[1] + kernel_img_mul_13[2] + 
                kernel_img_mul_13[3] + kernel_img_mul_13[4] + kernel_img_mul_13[5] + 
                kernel_img_mul_13[6] + kernel_img_mul_13[7] + kernel_img_mul_13[8] + 
                kernel_img_mul_13[9] + kernel_img_mul_13[10] + kernel_img_mul_13[11] + 
                kernel_img_mul_13[12] + kernel_img_mul_13[13] + kernel_img_mul_13[14] + 
                kernel_img_mul_13[15] + kernel_img_mul_13[16] + kernel_img_mul_13[17] + 
                kernel_img_mul_13[18] + kernel_img_mul_13[19] + kernel_img_mul_13[20] + 
                kernel_img_mul_13[21] + kernel_img_mul_13[22] + kernel_img_mul_13[23] + 
                kernel_img_mul_13[24] + kernel_img_mul_13[25] + kernel_img_mul_13[26] + 
                kernel_img_mul_13[27] + kernel_img_mul_13[28] + kernel_img_mul_13[29] + 
                kernel_img_mul_13[30] + kernel_img_mul_13[31] + kernel_img_mul_13[32] + 
                kernel_img_mul_13[33] + kernel_img_mul_13[34] + kernel_img_mul_13[35] + 
                kernel_img_mul_13[36] + kernel_img_mul_13[37] + kernel_img_mul_13[38] + 
                kernel_img_mul_13[39] + kernel_img_mul_13[40] + kernel_img_mul_13[41] + 
                kernel_img_mul_13[42] + kernel_img_mul_13[43] + kernel_img_mul_13[44] + 
                kernel_img_mul_13[45] + kernel_img_mul_13[46] + kernel_img_mul_13[47] + 
                kernel_img_mul_13[48];
wire  [39:0]  kernel_img_mul_14[0:48];
assign kernel_img_mul_14[0] = layer0[14][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_14[1] = layer0[14][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_14[2] = layer0[14][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_14[3] = layer0[14][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_14[4] = layer0[14][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_14[5] = layer0[14][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_14[6] = layer0[14][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_14[7] = layer1[14][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_14[8] = layer1[14][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_14[9] = layer1[14][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_14[10] = layer1[14][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_14[11] = layer1[14][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_14[12] = layer1[14][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_14[13] = layer1[14][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_14[14] = layer2[14][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_14[15] = layer2[14][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_14[16] = layer2[14][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_14[17] = layer2[14][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_14[18] = layer2[14][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_14[19] = layer2[14][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_14[20] = layer2[14][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_14[21] = layer3[14][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_14[22] = layer3[14][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_14[23] = layer3[14][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_14[24] = layer3[14][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_14[25] = layer3[14][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_14[26] = layer3[14][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_14[27] = layer3[14][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_14[28] = layer4[14][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_14[29] = layer4[14][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_14[30] = layer4[14][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_14[31] = layer4[14][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_14[32] = layer4[14][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_14[33] = layer4[14][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_14[34] = layer4[14][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_14[35] = layer5[14][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_14[36] = layer5[14][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_14[37] = layer5[14][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_14[38] = layer5[14][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_14[39] = layer5[14][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_14[40] = layer5[14][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_14[41] = layer5[14][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_14[42] = layer6[14][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_14[43] = layer6[14][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_14[44] = layer6[14][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_14[45] = layer6[14][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_14[46] = layer6[14][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_14[47] = layer6[14][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_14[48] = layer6[14][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_14 = kernel_img_mul_14[0] + kernel_img_mul_14[1] + kernel_img_mul_14[2] + 
                kernel_img_mul_14[3] + kernel_img_mul_14[4] + kernel_img_mul_14[5] + 
                kernel_img_mul_14[6] + kernel_img_mul_14[7] + kernel_img_mul_14[8] + 
                kernel_img_mul_14[9] + kernel_img_mul_14[10] + kernel_img_mul_14[11] + 
                kernel_img_mul_14[12] + kernel_img_mul_14[13] + kernel_img_mul_14[14] + 
                kernel_img_mul_14[15] + kernel_img_mul_14[16] + kernel_img_mul_14[17] + 
                kernel_img_mul_14[18] + kernel_img_mul_14[19] + kernel_img_mul_14[20] + 
                kernel_img_mul_14[21] + kernel_img_mul_14[22] + kernel_img_mul_14[23] + 
                kernel_img_mul_14[24] + kernel_img_mul_14[25] + kernel_img_mul_14[26] + 
                kernel_img_mul_14[27] + kernel_img_mul_14[28] + kernel_img_mul_14[29] + 
                kernel_img_mul_14[30] + kernel_img_mul_14[31] + kernel_img_mul_14[32] + 
                kernel_img_mul_14[33] + kernel_img_mul_14[34] + kernel_img_mul_14[35] + 
                kernel_img_mul_14[36] + kernel_img_mul_14[37] + kernel_img_mul_14[38] + 
                kernel_img_mul_14[39] + kernel_img_mul_14[40] + kernel_img_mul_14[41] + 
                kernel_img_mul_14[42] + kernel_img_mul_14[43] + kernel_img_mul_14[44] + 
                kernel_img_mul_14[45] + kernel_img_mul_14[46] + kernel_img_mul_14[47] + 
                kernel_img_mul_14[48];
wire  [39:0]  kernel_img_mul_15[0:48];
assign kernel_img_mul_15[0] = layer0[15][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_15[1] = layer0[15][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_15[2] = layer0[15][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_15[3] = layer0[15][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_15[4] = layer0[15][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_15[5] = layer0[15][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_15[6] = layer0[15][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_15[7] = layer1[15][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_15[8] = layer1[15][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_15[9] = layer1[15][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_15[10] = layer1[15][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_15[11] = layer1[15][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_15[12] = layer1[15][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_15[13] = layer1[15][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_15[14] = layer2[15][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_15[15] = layer2[15][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_15[16] = layer2[15][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_15[17] = layer2[15][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_15[18] = layer2[15][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_15[19] = layer2[15][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_15[20] = layer2[15][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_15[21] = layer3[15][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_15[22] = layer3[15][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_15[23] = layer3[15][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_15[24] = layer3[15][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_15[25] = layer3[15][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_15[26] = layer3[15][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_15[27] = layer3[15][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_15[28] = layer4[15][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_15[29] = layer4[15][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_15[30] = layer4[15][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_15[31] = layer4[15][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_15[32] = layer4[15][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_15[33] = layer4[15][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_15[34] = layer4[15][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_15[35] = layer5[15][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_15[36] = layer5[15][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_15[37] = layer5[15][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_15[38] = layer5[15][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_15[39] = layer5[15][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_15[40] = layer5[15][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_15[41] = layer5[15][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_15[42] = layer6[15][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_15[43] = layer6[15][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_15[44] = layer6[15][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_15[45] = layer6[15][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_15[46] = layer6[15][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_15[47] = layer6[15][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_15[48] = layer6[15][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_15 = kernel_img_mul_15[0] + kernel_img_mul_15[1] + kernel_img_mul_15[2] + 
                kernel_img_mul_15[3] + kernel_img_mul_15[4] + kernel_img_mul_15[5] + 
                kernel_img_mul_15[6] + kernel_img_mul_15[7] + kernel_img_mul_15[8] + 
                kernel_img_mul_15[9] + kernel_img_mul_15[10] + kernel_img_mul_15[11] + 
                kernel_img_mul_15[12] + kernel_img_mul_15[13] + kernel_img_mul_15[14] + 
                kernel_img_mul_15[15] + kernel_img_mul_15[16] + kernel_img_mul_15[17] + 
                kernel_img_mul_15[18] + kernel_img_mul_15[19] + kernel_img_mul_15[20] + 
                kernel_img_mul_15[21] + kernel_img_mul_15[22] + kernel_img_mul_15[23] + 
                kernel_img_mul_15[24] + kernel_img_mul_15[25] + kernel_img_mul_15[26] + 
                kernel_img_mul_15[27] + kernel_img_mul_15[28] + kernel_img_mul_15[29] + 
                kernel_img_mul_15[30] + kernel_img_mul_15[31] + kernel_img_mul_15[32] + 
                kernel_img_mul_15[33] + kernel_img_mul_15[34] + kernel_img_mul_15[35] + 
                kernel_img_mul_15[36] + kernel_img_mul_15[37] + kernel_img_mul_15[38] + 
                kernel_img_mul_15[39] + kernel_img_mul_15[40] + kernel_img_mul_15[41] + 
                kernel_img_mul_15[42] + kernel_img_mul_15[43] + kernel_img_mul_15[44] + 
                kernel_img_mul_15[45] + kernel_img_mul_15[46] + kernel_img_mul_15[47] + 
                kernel_img_mul_15[48];
wire  [39:0]  kernel_img_mul_16[0:48];
assign kernel_img_mul_16[0] = layer0[16][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_16[1] = layer0[16][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_16[2] = layer0[16][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_16[3] = layer0[16][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_16[4] = layer0[16][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_16[5] = layer0[16][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_16[6] = layer0[16][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_16[7] = layer1[16][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_16[8] = layer1[16][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_16[9] = layer1[16][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_16[10] = layer1[16][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_16[11] = layer1[16][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_16[12] = layer1[16][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_16[13] = layer1[16][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_16[14] = layer2[16][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_16[15] = layer2[16][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_16[16] = layer2[16][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_16[17] = layer2[16][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_16[18] = layer2[16][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_16[19] = layer2[16][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_16[20] = layer2[16][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_16[21] = layer3[16][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_16[22] = layer3[16][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_16[23] = layer3[16][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_16[24] = layer3[16][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_16[25] = layer3[16][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_16[26] = layer3[16][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_16[27] = layer3[16][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_16[28] = layer4[16][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_16[29] = layer4[16][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_16[30] = layer4[16][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_16[31] = layer4[16][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_16[32] = layer4[16][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_16[33] = layer4[16][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_16[34] = layer4[16][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_16[35] = layer5[16][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_16[36] = layer5[16][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_16[37] = layer5[16][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_16[38] = layer5[16][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_16[39] = layer5[16][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_16[40] = layer5[16][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_16[41] = layer5[16][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_16[42] = layer6[16][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_16[43] = layer6[16][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_16[44] = layer6[16][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_16[45] = layer6[16][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_16[46] = layer6[16][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_16[47] = layer6[16][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_16[48] = layer6[16][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_16 = kernel_img_mul_16[0] + kernel_img_mul_16[1] + kernel_img_mul_16[2] + 
                kernel_img_mul_16[3] + kernel_img_mul_16[4] + kernel_img_mul_16[5] + 
                kernel_img_mul_16[6] + kernel_img_mul_16[7] + kernel_img_mul_16[8] + 
                kernel_img_mul_16[9] + kernel_img_mul_16[10] + kernel_img_mul_16[11] + 
                kernel_img_mul_16[12] + kernel_img_mul_16[13] + kernel_img_mul_16[14] + 
                kernel_img_mul_16[15] + kernel_img_mul_16[16] + kernel_img_mul_16[17] + 
                kernel_img_mul_16[18] + kernel_img_mul_16[19] + kernel_img_mul_16[20] + 
                kernel_img_mul_16[21] + kernel_img_mul_16[22] + kernel_img_mul_16[23] + 
                kernel_img_mul_16[24] + kernel_img_mul_16[25] + kernel_img_mul_16[26] + 
                kernel_img_mul_16[27] + kernel_img_mul_16[28] + kernel_img_mul_16[29] + 
                kernel_img_mul_16[30] + kernel_img_mul_16[31] + kernel_img_mul_16[32] + 
                kernel_img_mul_16[33] + kernel_img_mul_16[34] + kernel_img_mul_16[35] + 
                kernel_img_mul_16[36] + kernel_img_mul_16[37] + kernel_img_mul_16[38] + 
                kernel_img_mul_16[39] + kernel_img_mul_16[40] + kernel_img_mul_16[41] + 
                kernel_img_mul_16[42] + kernel_img_mul_16[43] + kernel_img_mul_16[44] + 
                kernel_img_mul_16[45] + kernel_img_mul_16[46] + kernel_img_mul_16[47] + 
                kernel_img_mul_16[48];
wire  [39:0]  kernel_img_mul_17[0:48];
assign kernel_img_mul_17[0] = layer0[17][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_17[1] = layer0[17][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_17[2] = layer0[17][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_17[3] = layer0[17][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_17[4] = layer0[17][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_17[5] = layer0[17][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_17[6] = layer0[17][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_17[7] = layer1[17][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_17[8] = layer1[17][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_17[9] = layer1[17][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_17[10] = layer1[17][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_17[11] = layer1[17][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_17[12] = layer1[17][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_17[13] = layer1[17][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_17[14] = layer2[17][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_17[15] = layer2[17][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_17[16] = layer2[17][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_17[17] = layer2[17][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_17[18] = layer2[17][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_17[19] = layer2[17][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_17[20] = layer2[17][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_17[21] = layer3[17][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_17[22] = layer3[17][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_17[23] = layer3[17][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_17[24] = layer3[17][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_17[25] = layer3[17][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_17[26] = layer3[17][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_17[27] = layer3[17][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_17[28] = layer4[17][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_17[29] = layer4[17][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_17[30] = layer4[17][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_17[31] = layer4[17][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_17[32] = layer4[17][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_17[33] = layer4[17][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_17[34] = layer4[17][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_17[35] = layer5[17][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_17[36] = layer5[17][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_17[37] = layer5[17][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_17[38] = layer5[17][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_17[39] = layer5[17][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_17[40] = layer5[17][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_17[41] = layer5[17][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_17[42] = layer6[17][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_17[43] = layer6[17][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_17[44] = layer6[17][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_17[45] = layer6[17][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_17[46] = layer6[17][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_17[47] = layer6[17][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_17[48] = layer6[17][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_17 = kernel_img_mul_17[0] + kernel_img_mul_17[1] + kernel_img_mul_17[2] + 
                kernel_img_mul_17[3] + kernel_img_mul_17[4] + kernel_img_mul_17[5] + 
                kernel_img_mul_17[6] + kernel_img_mul_17[7] + kernel_img_mul_17[8] + 
                kernel_img_mul_17[9] + kernel_img_mul_17[10] + kernel_img_mul_17[11] + 
                kernel_img_mul_17[12] + kernel_img_mul_17[13] + kernel_img_mul_17[14] + 
                kernel_img_mul_17[15] + kernel_img_mul_17[16] + kernel_img_mul_17[17] + 
                kernel_img_mul_17[18] + kernel_img_mul_17[19] + kernel_img_mul_17[20] + 
                kernel_img_mul_17[21] + kernel_img_mul_17[22] + kernel_img_mul_17[23] + 
                kernel_img_mul_17[24] + kernel_img_mul_17[25] + kernel_img_mul_17[26] + 
                kernel_img_mul_17[27] + kernel_img_mul_17[28] + kernel_img_mul_17[29] + 
                kernel_img_mul_17[30] + kernel_img_mul_17[31] + kernel_img_mul_17[32] + 
                kernel_img_mul_17[33] + kernel_img_mul_17[34] + kernel_img_mul_17[35] + 
                kernel_img_mul_17[36] + kernel_img_mul_17[37] + kernel_img_mul_17[38] + 
                kernel_img_mul_17[39] + kernel_img_mul_17[40] + kernel_img_mul_17[41] + 
                kernel_img_mul_17[42] + kernel_img_mul_17[43] + kernel_img_mul_17[44] + 
                kernel_img_mul_17[45] + kernel_img_mul_17[46] + kernel_img_mul_17[47] + 
                kernel_img_mul_17[48];
wire  [39:0]  kernel_img_mul_18[0:48];
assign kernel_img_mul_18[0] = layer0[18][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_18[1] = layer0[18][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_18[2] = layer0[18][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_18[3] = layer0[18][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_18[4] = layer0[18][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_18[5] = layer0[18][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_18[6] = layer0[18][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_18[7] = layer1[18][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_18[8] = layer1[18][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_18[9] = layer1[18][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_18[10] = layer1[18][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_18[11] = layer1[18][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_18[12] = layer1[18][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_18[13] = layer1[18][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_18[14] = layer2[18][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_18[15] = layer2[18][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_18[16] = layer2[18][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_18[17] = layer2[18][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_18[18] = layer2[18][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_18[19] = layer2[18][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_18[20] = layer2[18][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_18[21] = layer3[18][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_18[22] = layer3[18][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_18[23] = layer3[18][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_18[24] = layer3[18][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_18[25] = layer3[18][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_18[26] = layer3[18][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_18[27] = layer3[18][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_18[28] = layer4[18][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_18[29] = layer4[18][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_18[30] = layer4[18][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_18[31] = layer4[18][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_18[32] = layer4[18][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_18[33] = layer4[18][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_18[34] = layer4[18][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_18[35] = layer5[18][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_18[36] = layer5[18][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_18[37] = layer5[18][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_18[38] = layer5[18][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_18[39] = layer5[18][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_18[40] = layer5[18][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_18[41] = layer5[18][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_18[42] = layer6[18][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_18[43] = layer6[18][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_18[44] = layer6[18][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_18[45] = layer6[18][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_18[46] = layer6[18][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_18[47] = layer6[18][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_18[48] = layer6[18][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_18 = kernel_img_mul_18[0] + kernel_img_mul_18[1] + kernel_img_mul_18[2] + 
                kernel_img_mul_18[3] + kernel_img_mul_18[4] + kernel_img_mul_18[5] + 
                kernel_img_mul_18[6] + kernel_img_mul_18[7] + kernel_img_mul_18[8] + 
                kernel_img_mul_18[9] + kernel_img_mul_18[10] + kernel_img_mul_18[11] + 
                kernel_img_mul_18[12] + kernel_img_mul_18[13] + kernel_img_mul_18[14] + 
                kernel_img_mul_18[15] + kernel_img_mul_18[16] + kernel_img_mul_18[17] + 
                kernel_img_mul_18[18] + kernel_img_mul_18[19] + kernel_img_mul_18[20] + 
                kernel_img_mul_18[21] + kernel_img_mul_18[22] + kernel_img_mul_18[23] + 
                kernel_img_mul_18[24] + kernel_img_mul_18[25] + kernel_img_mul_18[26] + 
                kernel_img_mul_18[27] + kernel_img_mul_18[28] + kernel_img_mul_18[29] + 
                kernel_img_mul_18[30] + kernel_img_mul_18[31] + kernel_img_mul_18[32] + 
                kernel_img_mul_18[33] + kernel_img_mul_18[34] + kernel_img_mul_18[35] + 
                kernel_img_mul_18[36] + kernel_img_mul_18[37] + kernel_img_mul_18[38] + 
                kernel_img_mul_18[39] + kernel_img_mul_18[40] + kernel_img_mul_18[41] + 
                kernel_img_mul_18[42] + kernel_img_mul_18[43] + kernel_img_mul_18[44] + 
                kernel_img_mul_18[45] + kernel_img_mul_18[46] + kernel_img_mul_18[47] + 
                kernel_img_mul_18[48];
wire  [39:0]  kernel_img_mul_19[0:48];
assign kernel_img_mul_19[0] = layer0[19][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_19[1] = layer0[19][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_19[2] = layer0[19][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_19[3] = layer0[19][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_19[4] = layer0[19][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_19[5] = layer0[19][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_19[6] = layer0[19][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_19[7] = layer1[19][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_19[8] = layer1[19][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_19[9] = layer1[19][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_19[10] = layer1[19][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_19[11] = layer1[19][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_19[12] = layer1[19][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_19[13] = layer1[19][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_19[14] = layer2[19][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_19[15] = layer2[19][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_19[16] = layer2[19][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_19[17] = layer2[19][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_19[18] = layer2[19][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_19[19] = layer2[19][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_19[20] = layer2[19][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_19[21] = layer3[19][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_19[22] = layer3[19][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_19[23] = layer3[19][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_19[24] = layer3[19][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_19[25] = layer3[19][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_19[26] = layer3[19][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_19[27] = layer3[19][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_19[28] = layer4[19][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_19[29] = layer4[19][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_19[30] = layer4[19][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_19[31] = layer4[19][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_19[32] = layer4[19][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_19[33] = layer4[19][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_19[34] = layer4[19][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_19[35] = layer5[19][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_19[36] = layer5[19][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_19[37] = layer5[19][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_19[38] = layer5[19][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_19[39] = layer5[19][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_19[40] = layer5[19][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_19[41] = layer5[19][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_19[42] = layer6[19][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_19[43] = layer6[19][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_19[44] = layer6[19][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_19[45] = layer6[19][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_19[46] = layer6[19][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_19[47] = layer6[19][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_19[48] = layer6[19][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_19 = kernel_img_mul_19[0] + kernel_img_mul_19[1] + kernel_img_mul_19[2] + 
                kernel_img_mul_19[3] + kernel_img_mul_19[4] + kernel_img_mul_19[5] + 
                kernel_img_mul_19[6] + kernel_img_mul_19[7] + kernel_img_mul_19[8] + 
                kernel_img_mul_19[9] + kernel_img_mul_19[10] + kernel_img_mul_19[11] + 
                kernel_img_mul_19[12] + kernel_img_mul_19[13] + kernel_img_mul_19[14] + 
                kernel_img_mul_19[15] + kernel_img_mul_19[16] + kernel_img_mul_19[17] + 
                kernel_img_mul_19[18] + kernel_img_mul_19[19] + kernel_img_mul_19[20] + 
                kernel_img_mul_19[21] + kernel_img_mul_19[22] + kernel_img_mul_19[23] + 
                kernel_img_mul_19[24] + kernel_img_mul_19[25] + kernel_img_mul_19[26] + 
                kernel_img_mul_19[27] + kernel_img_mul_19[28] + kernel_img_mul_19[29] + 
                kernel_img_mul_19[30] + kernel_img_mul_19[31] + kernel_img_mul_19[32] + 
                kernel_img_mul_19[33] + kernel_img_mul_19[34] + kernel_img_mul_19[35] + 
                kernel_img_mul_19[36] + kernel_img_mul_19[37] + kernel_img_mul_19[38] + 
                kernel_img_mul_19[39] + kernel_img_mul_19[40] + kernel_img_mul_19[41] + 
                kernel_img_mul_19[42] + kernel_img_mul_19[43] + kernel_img_mul_19[44] + 
                kernel_img_mul_19[45] + kernel_img_mul_19[46] + kernel_img_mul_19[47] + 
                kernel_img_mul_19[48];
wire  [39:0]  kernel_img_mul_20[0:48];
assign kernel_img_mul_20[0] = layer0[20][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_20[1] = layer0[20][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_20[2] = layer0[20][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_20[3] = layer0[20][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_20[4] = layer0[20][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_20[5] = layer0[20][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_20[6] = layer0[20][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_20[7] = layer1[20][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_20[8] = layer1[20][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_20[9] = layer1[20][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_20[10] = layer1[20][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_20[11] = layer1[20][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_20[12] = layer1[20][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_20[13] = layer1[20][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_20[14] = layer2[20][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_20[15] = layer2[20][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_20[16] = layer2[20][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_20[17] = layer2[20][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_20[18] = layer2[20][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_20[19] = layer2[20][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_20[20] = layer2[20][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_20[21] = layer3[20][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_20[22] = layer3[20][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_20[23] = layer3[20][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_20[24] = layer3[20][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_20[25] = layer3[20][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_20[26] = layer3[20][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_20[27] = layer3[20][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_20[28] = layer4[20][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_20[29] = layer4[20][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_20[30] = layer4[20][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_20[31] = layer4[20][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_20[32] = layer4[20][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_20[33] = layer4[20][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_20[34] = layer4[20][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_20[35] = layer5[20][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_20[36] = layer5[20][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_20[37] = layer5[20][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_20[38] = layer5[20][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_20[39] = layer5[20][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_20[40] = layer5[20][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_20[41] = layer5[20][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_20[42] = layer6[20][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_20[43] = layer6[20][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_20[44] = layer6[20][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_20[45] = layer6[20][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_20[46] = layer6[20][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_20[47] = layer6[20][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_20[48] = layer6[20][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_20 = kernel_img_mul_20[0] + kernel_img_mul_20[1] + kernel_img_mul_20[2] + 
                kernel_img_mul_20[3] + kernel_img_mul_20[4] + kernel_img_mul_20[5] + 
                kernel_img_mul_20[6] + kernel_img_mul_20[7] + kernel_img_mul_20[8] + 
                kernel_img_mul_20[9] + kernel_img_mul_20[10] + kernel_img_mul_20[11] + 
                kernel_img_mul_20[12] + kernel_img_mul_20[13] + kernel_img_mul_20[14] + 
                kernel_img_mul_20[15] + kernel_img_mul_20[16] + kernel_img_mul_20[17] + 
                kernel_img_mul_20[18] + kernel_img_mul_20[19] + kernel_img_mul_20[20] + 
                kernel_img_mul_20[21] + kernel_img_mul_20[22] + kernel_img_mul_20[23] + 
                kernel_img_mul_20[24] + kernel_img_mul_20[25] + kernel_img_mul_20[26] + 
                kernel_img_mul_20[27] + kernel_img_mul_20[28] + kernel_img_mul_20[29] + 
                kernel_img_mul_20[30] + kernel_img_mul_20[31] + kernel_img_mul_20[32] + 
                kernel_img_mul_20[33] + kernel_img_mul_20[34] + kernel_img_mul_20[35] + 
                kernel_img_mul_20[36] + kernel_img_mul_20[37] + kernel_img_mul_20[38] + 
                kernel_img_mul_20[39] + kernel_img_mul_20[40] + kernel_img_mul_20[41] + 
                kernel_img_mul_20[42] + kernel_img_mul_20[43] + kernel_img_mul_20[44] + 
                kernel_img_mul_20[45] + kernel_img_mul_20[46] + kernel_img_mul_20[47] + 
                kernel_img_mul_20[48];
wire  [39:0]  kernel_img_mul_21[0:48];
assign kernel_img_mul_21[0] = layer0[21][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_21[1] = layer0[21][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_21[2] = layer0[21][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_21[3] = layer0[21][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_21[4] = layer0[21][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_21[5] = layer0[21][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_21[6] = layer0[21][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_21[7] = layer1[21][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_21[8] = layer1[21][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_21[9] = layer1[21][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_21[10] = layer1[21][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_21[11] = layer1[21][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_21[12] = layer1[21][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_21[13] = layer1[21][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_21[14] = layer2[21][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_21[15] = layer2[21][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_21[16] = layer2[21][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_21[17] = layer2[21][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_21[18] = layer2[21][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_21[19] = layer2[21][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_21[20] = layer2[21][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_21[21] = layer3[21][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_21[22] = layer3[21][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_21[23] = layer3[21][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_21[24] = layer3[21][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_21[25] = layer3[21][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_21[26] = layer3[21][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_21[27] = layer3[21][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_21[28] = layer4[21][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_21[29] = layer4[21][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_21[30] = layer4[21][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_21[31] = layer4[21][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_21[32] = layer4[21][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_21[33] = layer4[21][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_21[34] = layer4[21][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_21[35] = layer5[21][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_21[36] = layer5[21][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_21[37] = layer5[21][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_21[38] = layer5[21][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_21[39] = layer5[21][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_21[40] = layer5[21][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_21[41] = layer5[21][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_21[42] = layer6[21][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_21[43] = layer6[21][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_21[44] = layer6[21][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_21[45] = layer6[21][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_21[46] = layer6[21][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_21[47] = layer6[21][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_21[48] = layer6[21][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_21 = kernel_img_mul_21[0] + kernel_img_mul_21[1] + kernel_img_mul_21[2] + 
                kernel_img_mul_21[3] + kernel_img_mul_21[4] + kernel_img_mul_21[5] + 
                kernel_img_mul_21[6] + kernel_img_mul_21[7] + kernel_img_mul_21[8] + 
                kernel_img_mul_21[9] + kernel_img_mul_21[10] + kernel_img_mul_21[11] + 
                kernel_img_mul_21[12] + kernel_img_mul_21[13] + kernel_img_mul_21[14] + 
                kernel_img_mul_21[15] + kernel_img_mul_21[16] + kernel_img_mul_21[17] + 
                kernel_img_mul_21[18] + kernel_img_mul_21[19] + kernel_img_mul_21[20] + 
                kernel_img_mul_21[21] + kernel_img_mul_21[22] + kernel_img_mul_21[23] + 
                kernel_img_mul_21[24] + kernel_img_mul_21[25] + kernel_img_mul_21[26] + 
                kernel_img_mul_21[27] + kernel_img_mul_21[28] + kernel_img_mul_21[29] + 
                kernel_img_mul_21[30] + kernel_img_mul_21[31] + kernel_img_mul_21[32] + 
                kernel_img_mul_21[33] + kernel_img_mul_21[34] + kernel_img_mul_21[35] + 
                kernel_img_mul_21[36] + kernel_img_mul_21[37] + kernel_img_mul_21[38] + 
                kernel_img_mul_21[39] + kernel_img_mul_21[40] + kernel_img_mul_21[41] + 
                kernel_img_mul_21[42] + kernel_img_mul_21[43] + kernel_img_mul_21[44] + 
                kernel_img_mul_21[45] + kernel_img_mul_21[46] + kernel_img_mul_21[47] + 
                kernel_img_mul_21[48];
wire  [39:0]  kernel_img_mul_22[0:48];
assign kernel_img_mul_22[0] = layer0[22][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_22[1] = layer0[22][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_22[2] = layer0[22][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_22[3] = layer0[22][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_22[4] = layer0[22][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_22[5] = layer0[22][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_22[6] = layer0[22][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_22[7] = layer1[22][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_22[8] = layer1[22][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_22[9] = layer1[22][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_22[10] = layer1[22][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_22[11] = layer1[22][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_22[12] = layer1[22][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_22[13] = layer1[22][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_22[14] = layer2[22][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_22[15] = layer2[22][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_22[16] = layer2[22][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_22[17] = layer2[22][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_22[18] = layer2[22][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_22[19] = layer2[22][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_22[20] = layer2[22][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_22[21] = layer3[22][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_22[22] = layer3[22][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_22[23] = layer3[22][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_22[24] = layer3[22][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_22[25] = layer3[22][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_22[26] = layer3[22][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_22[27] = layer3[22][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_22[28] = layer4[22][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_22[29] = layer4[22][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_22[30] = layer4[22][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_22[31] = layer4[22][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_22[32] = layer4[22][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_22[33] = layer4[22][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_22[34] = layer4[22][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_22[35] = layer5[22][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_22[36] = layer5[22][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_22[37] = layer5[22][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_22[38] = layer5[22][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_22[39] = layer5[22][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_22[40] = layer5[22][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_22[41] = layer5[22][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_22[42] = layer6[22][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_22[43] = layer6[22][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_22[44] = layer6[22][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_22[45] = layer6[22][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_22[46] = layer6[22][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_22[47] = layer6[22][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_22[48] = layer6[22][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_22 = kernel_img_mul_22[0] + kernel_img_mul_22[1] + kernel_img_mul_22[2] + 
                kernel_img_mul_22[3] + kernel_img_mul_22[4] + kernel_img_mul_22[5] + 
                kernel_img_mul_22[6] + kernel_img_mul_22[7] + kernel_img_mul_22[8] + 
                kernel_img_mul_22[9] + kernel_img_mul_22[10] + kernel_img_mul_22[11] + 
                kernel_img_mul_22[12] + kernel_img_mul_22[13] + kernel_img_mul_22[14] + 
                kernel_img_mul_22[15] + kernel_img_mul_22[16] + kernel_img_mul_22[17] + 
                kernel_img_mul_22[18] + kernel_img_mul_22[19] + kernel_img_mul_22[20] + 
                kernel_img_mul_22[21] + kernel_img_mul_22[22] + kernel_img_mul_22[23] + 
                kernel_img_mul_22[24] + kernel_img_mul_22[25] + kernel_img_mul_22[26] + 
                kernel_img_mul_22[27] + kernel_img_mul_22[28] + kernel_img_mul_22[29] + 
                kernel_img_mul_22[30] + kernel_img_mul_22[31] + kernel_img_mul_22[32] + 
                kernel_img_mul_22[33] + kernel_img_mul_22[34] + kernel_img_mul_22[35] + 
                kernel_img_mul_22[36] + kernel_img_mul_22[37] + kernel_img_mul_22[38] + 
                kernel_img_mul_22[39] + kernel_img_mul_22[40] + kernel_img_mul_22[41] + 
                kernel_img_mul_22[42] + kernel_img_mul_22[43] + kernel_img_mul_22[44] + 
                kernel_img_mul_22[45] + kernel_img_mul_22[46] + kernel_img_mul_22[47] + 
                kernel_img_mul_22[48];
wire  [39:0]  kernel_img_mul_23[0:48];
assign kernel_img_mul_23[0] = layer0[23][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_23[1] = layer0[23][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_23[2] = layer0[23][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_23[3] = layer0[23][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_23[4] = layer0[23][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_23[5] = layer0[23][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_23[6] = layer0[23][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_23[7] = layer1[23][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_23[8] = layer1[23][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_23[9] = layer1[23][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_23[10] = layer1[23][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_23[11] = layer1[23][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_23[12] = layer1[23][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_23[13] = layer1[23][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_23[14] = layer2[23][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_23[15] = layer2[23][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_23[16] = layer2[23][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_23[17] = layer2[23][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_23[18] = layer2[23][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_23[19] = layer2[23][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_23[20] = layer2[23][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_23[21] = layer3[23][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_23[22] = layer3[23][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_23[23] = layer3[23][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_23[24] = layer3[23][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_23[25] = layer3[23][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_23[26] = layer3[23][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_23[27] = layer3[23][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_23[28] = layer4[23][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_23[29] = layer4[23][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_23[30] = layer4[23][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_23[31] = layer4[23][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_23[32] = layer4[23][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_23[33] = layer4[23][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_23[34] = layer4[23][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_23[35] = layer5[23][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_23[36] = layer5[23][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_23[37] = layer5[23][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_23[38] = layer5[23][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_23[39] = layer5[23][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_23[40] = layer5[23][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_23[41] = layer5[23][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_23[42] = layer6[23][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_23[43] = layer6[23][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_23[44] = layer6[23][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_23[45] = layer6[23][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_23[46] = layer6[23][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_23[47] = layer6[23][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_23[48] = layer6[23][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_23 = kernel_img_mul_23[0] + kernel_img_mul_23[1] + kernel_img_mul_23[2] + 
                kernel_img_mul_23[3] + kernel_img_mul_23[4] + kernel_img_mul_23[5] + 
                kernel_img_mul_23[6] + kernel_img_mul_23[7] + kernel_img_mul_23[8] + 
                kernel_img_mul_23[9] + kernel_img_mul_23[10] + kernel_img_mul_23[11] + 
                kernel_img_mul_23[12] + kernel_img_mul_23[13] + kernel_img_mul_23[14] + 
                kernel_img_mul_23[15] + kernel_img_mul_23[16] + kernel_img_mul_23[17] + 
                kernel_img_mul_23[18] + kernel_img_mul_23[19] + kernel_img_mul_23[20] + 
                kernel_img_mul_23[21] + kernel_img_mul_23[22] + kernel_img_mul_23[23] + 
                kernel_img_mul_23[24] + kernel_img_mul_23[25] + kernel_img_mul_23[26] + 
                kernel_img_mul_23[27] + kernel_img_mul_23[28] + kernel_img_mul_23[29] + 
                kernel_img_mul_23[30] + kernel_img_mul_23[31] + kernel_img_mul_23[32] + 
                kernel_img_mul_23[33] + kernel_img_mul_23[34] + kernel_img_mul_23[35] + 
                kernel_img_mul_23[36] + kernel_img_mul_23[37] + kernel_img_mul_23[38] + 
                kernel_img_mul_23[39] + kernel_img_mul_23[40] + kernel_img_mul_23[41] + 
                kernel_img_mul_23[42] + kernel_img_mul_23[43] + kernel_img_mul_23[44] + 
                kernel_img_mul_23[45] + kernel_img_mul_23[46] + kernel_img_mul_23[47] + 
                kernel_img_mul_23[48];
wire  [39:0]  kernel_img_mul_24[0:48];
assign kernel_img_mul_24[0] = layer0[24][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_24[1] = layer0[24][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_24[2] = layer0[24][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_24[3] = layer0[24][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_24[4] = layer0[24][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_24[5] = layer0[24][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_24[6] = layer0[24][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_24[7] = layer1[24][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_24[8] = layer1[24][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_24[9] = layer1[24][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_24[10] = layer1[24][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_24[11] = layer1[24][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_24[12] = layer1[24][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_24[13] = layer1[24][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_24[14] = layer2[24][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_24[15] = layer2[24][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_24[16] = layer2[24][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_24[17] = layer2[24][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_24[18] = layer2[24][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_24[19] = layer2[24][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_24[20] = layer2[24][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_24[21] = layer3[24][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_24[22] = layer3[24][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_24[23] = layer3[24][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_24[24] = layer3[24][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_24[25] = layer3[24][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_24[26] = layer3[24][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_24[27] = layer3[24][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_24[28] = layer4[24][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_24[29] = layer4[24][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_24[30] = layer4[24][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_24[31] = layer4[24][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_24[32] = layer4[24][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_24[33] = layer4[24][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_24[34] = layer4[24][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_24[35] = layer5[24][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_24[36] = layer5[24][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_24[37] = layer5[24][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_24[38] = layer5[24][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_24[39] = layer5[24][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_24[40] = layer5[24][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_24[41] = layer5[24][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_24[42] = layer6[24][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_24[43] = layer6[24][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_24[44] = layer6[24][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_24[45] = layer6[24][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_24[46] = layer6[24][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_24[47] = layer6[24][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_24[48] = layer6[24][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_24 = kernel_img_mul_24[0] + kernel_img_mul_24[1] + kernel_img_mul_24[2] + 
                kernel_img_mul_24[3] + kernel_img_mul_24[4] + kernel_img_mul_24[5] + 
                kernel_img_mul_24[6] + kernel_img_mul_24[7] + kernel_img_mul_24[8] + 
                kernel_img_mul_24[9] + kernel_img_mul_24[10] + kernel_img_mul_24[11] + 
                kernel_img_mul_24[12] + kernel_img_mul_24[13] + kernel_img_mul_24[14] + 
                kernel_img_mul_24[15] + kernel_img_mul_24[16] + kernel_img_mul_24[17] + 
                kernel_img_mul_24[18] + kernel_img_mul_24[19] + kernel_img_mul_24[20] + 
                kernel_img_mul_24[21] + kernel_img_mul_24[22] + kernel_img_mul_24[23] + 
                kernel_img_mul_24[24] + kernel_img_mul_24[25] + kernel_img_mul_24[26] + 
                kernel_img_mul_24[27] + kernel_img_mul_24[28] + kernel_img_mul_24[29] + 
                kernel_img_mul_24[30] + kernel_img_mul_24[31] + kernel_img_mul_24[32] + 
                kernel_img_mul_24[33] + kernel_img_mul_24[34] + kernel_img_mul_24[35] + 
                kernel_img_mul_24[36] + kernel_img_mul_24[37] + kernel_img_mul_24[38] + 
                kernel_img_mul_24[39] + kernel_img_mul_24[40] + kernel_img_mul_24[41] + 
                kernel_img_mul_24[42] + kernel_img_mul_24[43] + kernel_img_mul_24[44] + 
                kernel_img_mul_24[45] + kernel_img_mul_24[46] + kernel_img_mul_24[47] + 
                kernel_img_mul_24[48];
wire  [39:0]  kernel_img_mul_25[0:48];
assign kernel_img_mul_25[0] = layer0[25][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_25[1] = layer0[25][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_25[2] = layer0[25][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_25[3] = layer0[25][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_25[4] = layer0[25][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_25[5] = layer0[25][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_25[6] = layer0[25][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_25[7] = layer1[25][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_25[8] = layer1[25][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_25[9] = layer1[25][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_25[10] = layer1[25][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_25[11] = layer1[25][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_25[12] = layer1[25][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_25[13] = layer1[25][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_25[14] = layer2[25][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_25[15] = layer2[25][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_25[16] = layer2[25][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_25[17] = layer2[25][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_25[18] = layer2[25][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_25[19] = layer2[25][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_25[20] = layer2[25][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_25[21] = layer3[25][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_25[22] = layer3[25][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_25[23] = layer3[25][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_25[24] = layer3[25][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_25[25] = layer3[25][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_25[26] = layer3[25][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_25[27] = layer3[25][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_25[28] = layer4[25][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_25[29] = layer4[25][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_25[30] = layer4[25][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_25[31] = layer4[25][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_25[32] = layer4[25][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_25[33] = layer4[25][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_25[34] = layer4[25][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_25[35] = layer5[25][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_25[36] = layer5[25][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_25[37] = layer5[25][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_25[38] = layer5[25][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_25[39] = layer5[25][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_25[40] = layer5[25][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_25[41] = layer5[25][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_25[42] = layer6[25][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_25[43] = layer6[25][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_25[44] = layer6[25][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_25[45] = layer6[25][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_25[46] = layer6[25][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_25[47] = layer6[25][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_25[48] = layer6[25][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_25 = kernel_img_mul_25[0] + kernel_img_mul_25[1] + kernel_img_mul_25[2] + 
                kernel_img_mul_25[3] + kernel_img_mul_25[4] + kernel_img_mul_25[5] + 
                kernel_img_mul_25[6] + kernel_img_mul_25[7] + kernel_img_mul_25[8] + 
                kernel_img_mul_25[9] + kernel_img_mul_25[10] + kernel_img_mul_25[11] + 
                kernel_img_mul_25[12] + kernel_img_mul_25[13] + kernel_img_mul_25[14] + 
                kernel_img_mul_25[15] + kernel_img_mul_25[16] + kernel_img_mul_25[17] + 
                kernel_img_mul_25[18] + kernel_img_mul_25[19] + kernel_img_mul_25[20] + 
                kernel_img_mul_25[21] + kernel_img_mul_25[22] + kernel_img_mul_25[23] + 
                kernel_img_mul_25[24] + kernel_img_mul_25[25] + kernel_img_mul_25[26] + 
                kernel_img_mul_25[27] + kernel_img_mul_25[28] + kernel_img_mul_25[29] + 
                kernel_img_mul_25[30] + kernel_img_mul_25[31] + kernel_img_mul_25[32] + 
                kernel_img_mul_25[33] + kernel_img_mul_25[34] + kernel_img_mul_25[35] + 
                kernel_img_mul_25[36] + kernel_img_mul_25[37] + kernel_img_mul_25[38] + 
                kernel_img_mul_25[39] + kernel_img_mul_25[40] + kernel_img_mul_25[41] + 
                kernel_img_mul_25[42] + kernel_img_mul_25[43] + kernel_img_mul_25[44] + 
                kernel_img_mul_25[45] + kernel_img_mul_25[46] + kernel_img_mul_25[47] + 
                kernel_img_mul_25[48];
wire  [39:0]  kernel_img_mul_26[0:48];
assign kernel_img_mul_26[0] = layer0[26][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_26[1] = layer0[26][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_26[2] = layer0[26][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_26[3] = layer0[26][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_26[4] = layer0[26][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_26[5] = layer0[26][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_26[6] = layer0[26][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_26[7] = layer1[26][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_26[8] = layer1[26][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_26[9] = layer1[26][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_26[10] = layer1[26][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_26[11] = layer1[26][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_26[12] = layer1[26][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_26[13] = layer1[26][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_26[14] = layer2[26][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_26[15] = layer2[26][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_26[16] = layer2[26][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_26[17] = layer2[26][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_26[18] = layer2[26][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_26[19] = layer2[26][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_26[20] = layer2[26][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_26[21] = layer3[26][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_26[22] = layer3[26][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_26[23] = layer3[26][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_26[24] = layer3[26][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_26[25] = layer3[26][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_26[26] = layer3[26][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_26[27] = layer3[26][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_26[28] = layer4[26][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_26[29] = layer4[26][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_26[30] = layer4[26][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_26[31] = layer4[26][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_26[32] = layer4[26][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_26[33] = layer4[26][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_26[34] = layer4[26][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_26[35] = layer5[26][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_26[36] = layer5[26][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_26[37] = layer5[26][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_26[38] = layer5[26][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_26[39] = layer5[26][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_26[40] = layer5[26][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_26[41] = layer5[26][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_26[42] = layer6[26][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_26[43] = layer6[26][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_26[44] = layer6[26][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_26[45] = layer6[26][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_26[46] = layer6[26][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_26[47] = layer6[26][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_26[48] = layer6[26][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_26 = kernel_img_mul_26[0] + kernel_img_mul_26[1] + kernel_img_mul_26[2] + 
                kernel_img_mul_26[3] + kernel_img_mul_26[4] + kernel_img_mul_26[5] + 
                kernel_img_mul_26[6] + kernel_img_mul_26[7] + kernel_img_mul_26[8] + 
                kernel_img_mul_26[9] + kernel_img_mul_26[10] + kernel_img_mul_26[11] + 
                kernel_img_mul_26[12] + kernel_img_mul_26[13] + kernel_img_mul_26[14] + 
                kernel_img_mul_26[15] + kernel_img_mul_26[16] + kernel_img_mul_26[17] + 
                kernel_img_mul_26[18] + kernel_img_mul_26[19] + kernel_img_mul_26[20] + 
                kernel_img_mul_26[21] + kernel_img_mul_26[22] + kernel_img_mul_26[23] + 
                kernel_img_mul_26[24] + kernel_img_mul_26[25] + kernel_img_mul_26[26] + 
                kernel_img_mul_26[27] + kernel_img_mul_26[28] + kernel_img_mul_26[29] + 
                kernel_img_mul_26[30] + kernel_img_mul_26[31] + kernel_img_mul_26[32] + 
                kernel_img_mul_26[33] + kernel_img_mul_26[34] + kernel_img_mul_26[35] + 
                kernel_img_mul_26[36] + kernel_img_mul_26[37] + kernel_img_mul_26[38] + 
                kernel_img_mul_26[39] + kernel_img_mul_26[40] + kernel_img_mul_26[41] + 
                kernel_img_mul_26[42] + kernel_img_mul_26[43] + kernel_img_mul_26[44] + 
                kernel_img_mul_26[45] + kernel_img_mul_26[46] + kernel_img_mul_26[47] + 
                kernel_img_mul_26[48];
wire  [39:0]  kernel_img_mul_27[0:48];
assign kernel_img_mul_27[0] = layer0[27][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_27[1] = layer0[27][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_27[2] = layer0[27][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_27[3] = layer0[27][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_27[4] = layer0[27][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_27[5] = layer0[27][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_27[6] = layer0[27][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_27[7] = layer1[27][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_27[8] = layer1[27][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_27[9] = layer1[27][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_27[10] = layer1[27][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_27[11] = layer1[27][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_27[12] = layer1[27][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_27[13] = layer1[27][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_27[14] = layer2[27][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_27[15] = layer2[27][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_27[16] = layer2[27][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_27[17] = layer2[27][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_27[18] = layer2[27][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_27[19] = layer2[27][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_27[20] = layer2[27][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_27[21] = layer3[27][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_27[22] = layer3[27][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_27[23] = layer3[27][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_27[24] = layer3[27][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_27[25] = layer3[27][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_27[26] = layer3[27][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_27[27] = layer3[27][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_27[28] = layer4[27][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_27[29] = layer4[27][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_27[30] = layer4[27][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_27[31] = layer4[27][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_27[32] = layer4[27][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_27[33] = layer4[27][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_27[34] = layer4[27][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_27[35] = layer5[27][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_27[36] = layer5[27][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_27[37] = layer5[27][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_27[38] = layer5[27][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_27[39] = layer5[27][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_27[40] = layer5[27][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_27[41] = layer5[27][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_27[42] = layer6[27][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_27[43] = layer6[27][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_27[44] = layer6[27][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_27[45] = layer6[27][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_27[46] = layer6[27][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_27[47] = layer6[27][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_27[48] = layer6[27][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_27 = kernel_img_mul_27[0] + kernel_img_mul_27[1] + kernel_img_mul_27[2] + 
                kernel_img_mul_27[3] + kernel_img_mul_27[4] + kernel_img_mul_27[5] + 
                kernel_img_mul_27[6] + kernel_img_mul_27[7] + kernel_img_mul_27[8] + 
                kernel_img_mul_27[9] + kernel_img_mul_27[10] + kernel_img_mul_27[11] + 
                kernel_img_mul_27[12] + kernel_img_mul_27[13] + kernel_img_mul_27[14] + 
                kernel_img_mul_27[15] + kernel_img_mul_27[16] + kernel_img_mul_27[17] + 
                kernel_img_mul_27[18] + kernel_img_mul_27[19] + kernel_img_mul_27[20] + 
                kernel_img_mul_27[21] + kernel_img_mul_27[22] + kernel_img_mul_27[23] + 
                kernel_img_mul_27[24] + kernel_img_mul_27[25] + kernel_img_mul_27[26] + 
                kernel_img_mul_27[27] + kernel_img_mul_27[28] + kernel_img_mul_27[29] + 
                kernel_img_mul_27[30] + kernel_img_mul_27[31] + kernel_img_mul_27[32] + 
                kernel_img_mul_27[33] + kernel_img_mul_27[34] + kernel_img_mul_27[35] + 
                kernel_img_mul_27[36] + kernel_img_mul_27[37] + kernel_img_mul_27[38] + 
                kernel_img_mul_27[39] + kernel_img_mul_27[40] + kernel_img_mul_27[41] + 
                kernel_img_mul_27[42] + kernel_img_mul_27[43] + kernel_img_mul_27[44] + 
                kernel_img_mul_27[45] + kernel_img_mul_27[46] + kernel_img_mul_27[47] + 
                kernel_img_mul_27[48];
wire  [39:0]  kernel_img_mul_28[0:48];
assign kernel_img_mul_28[0] = layer0[28][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_28[1] = layer0[28][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_28[2] = layer0[28][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_28[3] = layer0[28][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_28[4] = layer0[28][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_28[5] = layer0[28][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_28[6] = layer0[28][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_28[7] = layer1[28][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_28[8] = layer1[28][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_28[9] = layer1[28][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_28[10] = layer1[28][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_28[11] = layer1[28][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_28[12] = layer1[28][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_28[13] = layer1[28][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_28[14] = layer2[28][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_28[15] = layer2[28][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_28[16] = layer2[28][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_28[17] = layer2[28][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_28[18] = layer2[28][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_28[19] = layer2[28][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_28[20] = layer2[28][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_28[21] = layer3[28][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_28[22] = layer3[28][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_28[23] = layer3[28][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_28[24] = layer3[28][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_28[25] = layer3[28][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_28[26] = layer3[28][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_28[27] = layer3[28][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_28[28] = layer4[28][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_28[29] = layer4[28][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_28[30] = layer4[28][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_28[31] = layer4[28][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_28[32] = layer4[28][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_28[33] = layer4[28][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_28[34] = layer4[28][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_28[35] = layer5[28][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_28[36] = layer5[28][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_28[37] = layer5[28][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_28[38] = layer5[28][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_28[39] = layer5[28][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_28[40] = layer5[28][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_28[41] = layer5[28][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_28[42] = layer6[28][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_28[43] = layer6[28][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_28[44] = layer6[28][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_28[45] = layer6[28][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_28[46] = layer6[28][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_28[47] = layer6[28][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_28[48] = layer6[28][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_28 = kernel_img_mul_28[0] + kernel_img_mul_28[1] + kernel_img_mul_28[2] + 
                kernel_img_mul_28[3] + kernel_img_mul_28[4] + kernel_img_mul_28[5] + 
                kernel_img_mul_28[6] + kernel_img_mul_28[7] + kernel_img_mul_28[8] + 
                kernel_img_mul_28[9] + kernel_img_mul_28[10] + kernel_img_mul_28[11] + 
                kernel_img_mul_28[12] + kernel_img_mul_28[13] + kernel_img_mul_28[14] + 
                kernel_img_mul_28[15] + kernel_img_mul_28[16] + kernel_img_mul_28[17] + 
                kernel_img_mul_28[18] + kernel_img_mul_28[19] + kernel_img_mul_28[20] + 
                kernel_img_mul_28[21] + kernel_img_mul_28[22] + kernel_img_mul_28[23] + 
                kernel_img_mul_28[24] + kernel_img_mul_28[25] + kernel_img_mul_28[26] + 
                kernel_img_mul_28[27] + kernel_img_mul_28[28] + kernel_img_mul_28[29] + 
                kernel_img_mul_28[30] + kernel_img_mul_28[31] + kernel_img_mul_28[32] + 
                kernel_img_mul_28[33] + kernel_img_mul_28[34] + kernel_img_mul_28[35] + 
                kernel_img_mul_28[36] + kernel_img_mul_28[37] + kernel_img_mul_28[38] + 
                kernel_img_mul_28[39] + kernel_img_mul_28[40] + kernel_img_mul_28[41] + 
                kernel_img_mul_28[42] + kernel_img_mul_28[43] + kernel_img_mul_28[44] + 
                kernel_img_mul_28[45] + kernel_img_mul_28[46] + kernel_img_mul_28[47] + 
                kernel_img_mul_28[48];
wire  [39:0]  kernel_img_mul_29[0:48];
assign kernel_img_mul_29[0] = layer0[29][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_29[1] = layer0[29][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_29[2] = layer0[29][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_29[3] = layer0[29][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_29[4] = layer0[29][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_29[5] = layer0[29][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_29[6] = layer0[29][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_29[7] = layer1[29][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_29[8] = layer1[29][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_29[9] = layer1[29][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_29[10] = layer1[29][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_29[11] = layer1[29][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_29[12] = layer1[29][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_29[13] = layer1[29][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_29[14] = layer2[29][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_29[15] = layer2[29][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_29[16] = layer2[29][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_29[17] = layer2[29][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_29[18] = layer2[29][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_29[19] = layer2[29][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_29[20] = layer2[29][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_29[21] = layer3[29][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_29[22] = layer3[29][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_29[23] = layer3[29][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_29[24] = layer3[29][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_29[25] = layer3[29][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_29[26] = layer3[29][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_29[27] = layer3[29][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_29[28] = layer4[29][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_29[29] = layer4[29][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_29[30] = layer4[29][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_29[31] = layer4[29][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_29[32] = layer4[29][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_29[33] = layer4[29][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_29[34] = layer4[29][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_29[35] = layer5[29][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_29[36] = layer5[29][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_29[37] = layer5[29][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_29[38] = layer5[29][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_29[39] = layer5[29][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_29[40] = layer5[29][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_29[41] = layer5[29][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_29[42] = layer6[29][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_29[43] = layer6[29][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_29[44] = layer6[29][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_29[45] = layer6[29][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_29[46] = layer6[29][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_29[47] = layer6[29][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_29[48] = layer6[29][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_29 = kernel_img_mul_29[0] + kernel_img_mul_29[1] + kernel_img_mul_29[2] + 
                kernel_img_mul_29[3] + kernel_img_mul_29[4] + kernel_img_mul_29[5] + 
                kernel_img_mul_29[6] + kernel_img_mul_29[7] + kernel_img_mul_29[8] + 
                kernel_img_mul_29[9] + kernel_img_mul_29[10] + kernel_img_mul_29[11] + 
                kernel_img_mul_29[12] + kernel_img_mul_29[13] + kernel_img_mul_29[14] + 
                kernel_img_mul_29[15] + kernel_img_mul_29[16] + kernel_img_mul_29[17] + 
                kernel_img_mul_29[18] + kernel_img_mul_29[19] + kernel_img_mul_29[20] + 
                kernel_img_mul_29[21] + kernel_img_mul_29[22] + kernel_img_mul_29[23] + 
                kernel_img_mul_29[24] + kernel_img_mul_29[25] + kernel_img_mul_29[26] + 
                kernel_img_mul_29[27] + kernel_img_mul_29[28] + kernel_img_mul_29[29] + 
                kernel_img_mul_29[30] + kernel_img_mul_29[31] + kernel_img_mul_29[32] + 
                kernel_img_mul_29[33] + kernel_img_mul_29[34] + kernel_img_mul_29[35] + 
                kernel_img_mul_29[36] + kernel_img_mul_29[37] + kernel_img_mul_29[38] + 
                kernel_img_mul_29[39] + kernel_img_mul_29[40] + kernel_img_mul_29[41] + 
                kernel_img_mul_29[42] + kernel_img_mul_29[43] + kernel_img_mul_29[44] + 
                kernel_img_mul_29[45] + kernel_img_mul_29[46] + kernel_img_mul_29[47] + 
                kernel_img_mul_29[48];
wire  [39:0]  kernel_img_mul_30[0:48];
assign kernel_img_mul_30[0] = layer0[30][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_30[1] = layer0[30][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_30[2] = layer0[30][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_30[3] = layer0[30][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_30[4] = layer0[30][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_30[5] = layer0[30][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_30[6] = layer0[30][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_30[7] = layer1[30][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_30[8] = layer1[30][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_30[9] = layer1[30][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_30[10] = layer1[30][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_30[11] = layer1[30][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_30[12] = layer1[30][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_30[13] = layer1[30][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_30[14] = layer2[30][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_30[15] = layer2[30][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_30[16] = layer2[30][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_30[17] = layer2[30][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_30[18] = layer2[30][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_30[19] = layer2[30][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_30[20] = layer2[30][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_30[21] = layer3[30][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_30[22] = layer3[30][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_30[23] = layer3[30][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_30[24] = layer3[30][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_30[25] = layer3[30][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_30[26] = layer3[30][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_30[27] = layer3[30][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_30[28] = layer4[30][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_30[29] = layer4[30][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_30[30] = layer4[30][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_30[31] = layer4[30][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_30[32] = layer4[30][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_30[33] = layer4[30][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_30[34] = layer4[30][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_30[35] = layer5[30][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_30[36] = layer5[30][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_30[37] = layer5[30][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_30[38] = layer5[30][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_30[39] = layer5[30][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_30[40] = layer5[30][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_30[41] = layer5[30][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_30[42] = layer6[30][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_30[43] = layer6[30][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_30[44] = layer6[30][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_30[45] = layer6[30][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_30[46] = layer6[30][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_30[47] = layer6[30][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_30[48] = layer6[30][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_30 = kernel_img_mul_30[0] + kernel_img_mul_30[1] + kernel_img_mul_30[2] + 
                kernel_img_mul_30[3] + kernel_img_mul_30[4] + kernel_img_mul_30[5] + 
                kernel_img_mul_30[6] + kernel_img_mul_30[7] + kernel_img_mul_30[8] + 
                kernel_img_mul_30[9] + kernel_img_mul_30[10] + kernel_img_mul_30[11] + 
                kernel_img_mul_30[12] + kernel_img_mul_30[13] + kernel_img_mul_30[14] + 
                kernel_img_mul_30[15] + kernel_img_mul_30[16] + kernel_img_mul_30[17] + 
                kernel_img_mul_30[18] + kernel_img_mul_30[19] + kernel_img_mul_30[20] + 
                kernel_img_mul_30[21] + kernel_img_mul_30[22] + kernel_img_mul_30[23] + 
                kernel_img_mul_30[24] + kernel_img_mul_30[25] + kernel_img_mul_30[26] + 
                kernel_img_mul_30[27] + kernel_img_mul_30[28] + kernel_img_mul_30[29] + 
                kernel_img_mul_30[30] + kernel_img_mul_30[31] + kernel_img_mul_30[32] + 
                kernel_img_mul_30[33] + kernel_img_mul_30[34] + kernel_img_mul_30[35] + 
                kernel_img_mul_30[36] + kernel_img_mul_30[37] + kernel_img_mul_30[38] + 
                kernel_img_mul_30[39] + kernel_img_mul_30[40] + kernel_img_mul_30[41] + 
                kernel_img_mul_30[42] + kernel_img_mul_30[43] + kernel_img_mul_30[44] + 
                kernel_img_mul_30[45] + kernel_img_mul_30[46] + kernel_img_mul_30[47] + 
                kernel_img_mul_30[48];
wire  [39:0]  kernel_img_mul_31[0:48];
assign kernel_img_mul_31[0] = layer0[31][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_31[1] = layer0[31][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_31[2] = layer0[31][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_31[3] = layer0[31][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_31[4] = layer0[31][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_31[5] = layer0[31][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_31[6] = layer0[31][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_31[7] = layer1[31][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_31[8] = layer1[31][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_31[9] = layer1[31][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_31[10] = layer1[31][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_31[11] = layer1[31][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_31[12] = layer1[31][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_31[13] = layer1[31][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_31[14] = layer2[31][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_31[15] = layer2[31][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_31[16] = layer2[31][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_31[17] = layer2[31][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_31[18] = layer2[31][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_31[19] = layer2[31][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_31[20] = layer2[31][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_31[21] = layer3[31][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_31[22] = layer3[31][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_31[23] = layer3[31][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_31[24] = layer3[31][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_31[25] = layer3[31][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_31[26] = layer3[31][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_31[27] = layer3[31][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_31[28] = layer4[31][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_31[29] = layer4[31][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_31[30] = layer4[31][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_31[31] = layer4[31][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_31[32] = layer4[31][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_31[33] = layer4[31][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_31[34] = layer4[31][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_31[35] = layer5[31][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_31[36] = layer5[31][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_31[37] = layer5[31][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_31[38] = layer5[31][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_31[39] = layer5[31][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_31[40] = layer5[31][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_31[41] = layer5[31][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_31[42] = layer6[31][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_31[43] = layer6[31][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_31[44] = layer6[31][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_31[45] = layer6[31][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_31[46] = layer6[31][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_31[47] = layer6[31][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_31[48] = layer6[31][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_31 = kernel_img_mul_31[0] + kernel_img_mul_31[1] + kernel_img_mul_31[2] + 
                kernel_img_mul_31[3] + kernel_img_mul_31[4] + kernel_img_mul_31[5] + 
                kernel_img_mul_31[6] + kernel_img_mul_31[7] + kernel_img_mul_31[8] + 
                kernel_img_mul_31[9] + kernel_img_mul_31[10] + kernel_img_mul_31[11] + 
                kernel_img_mul_31[12] + kernel_img_mul_31[13] + kernel_img_mul_31[14] + 
                kernel_img_mul_31[15] + kernel_img_mul_31[16] + kernel_img_mul_31[17] + 
                kernel_img_mul_31[18] + kernel_img_mul_31[19] + kernel_img_mul_31[20] + 
                kernel_img_mul_31[21] + kernel_img_mul_31[22] + kernel_img_mul_31[23] + 
                kernel_img_mul_31[24] + kernel_img_mul_31[25] + kernel_img_mul_31[26] + 
                kernel_img_mul_31[27] + kernel_img_mul_31[28] + kernel_img_mul_31[29] + 
                kernel_img_mul_31[30] + kernel_img_mul_31[31] + kernel_img_mul_31[32] + 
                kernel_img_mul_31[33] + kernel_img_mul_31[34] + kernel_img_mul_31[35] + 
                kernel_img_mul_31[36] + kernel_img_mul_31[37] + kernel_img_mul_31[38] + 
                kernel_img_mul_31[39] + kernel_img_mul_31[40] + kernel_img_mul_31[41] + 
                kernel_img_mul_31[42] + kernel_img_mul_31[43] + kernel_img_mul_31[44] + 
                kernel_img_mul_31[45] + kernel_img_mul_31[46] + kernel_img_mul_31[47] + 
                kernel_img_mul_31[48];
wire  [39:0]  kernel_img_mul_32[0:48];
assign kernel_img_mul_32[0] = layer0[32][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_32[1] = layer0[32][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_32[2] = layer0[32][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_32[3] = layer0[32][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_32[4] = layer0[32][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_32[5] = layer0[32][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_32[6] = layer0[32][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_32[7] = layer1[32][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_32[8] = layer1[32][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_32[9] = layer1[32][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_32[10] = layer1[32][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_32[11] = layer1[32][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_32[12] = layer1[32][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_32[13] = layer1[32][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_32[14] = layer2[32][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_32[15] = layer2[32][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_32[16] = layer2[32][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_32[17] = layer2[32][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_32[18] = layer2[32][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_32[19] = layer2[32][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_32[20] = layer2[32][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_32[21] = layer3[32][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_32[22] = layer3[32][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_32[23] = layer3[32][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_32[24] = layer3[32][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_32[25] = layer3[32][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_32[26] = layer3[32][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_32[27] = layer3[32][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_32[28] = layer4[32][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_32[29] = layer4[32][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_32[30] = layer4[32][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_32[31] = layer4[32][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_32[32] = layer4[32][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_32[33] = layer4[32][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_32[34] = layer4[32][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_32[35] = layer5[32][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_32[36] = layer5[32][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_32[37] = layer5[32][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_32[38] = layer5[32][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_32[39] = layer5[32][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_32[40] = layer5[32][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_32[41] = layer5[32][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_32[42] = layer6[32][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_32[43] = layer6[32][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_32[44] = layer6[32][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_32[45] = layer6[32][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_32[46] = layer6[32][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_32[47] = layer6[32][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_32[48] = layer6[32][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_32 = kernel_img_mul_32[0] + kernel_img_mul_32[1] + kernel_img_mul_32[2] + 
                kernel_img_mul_32[3] + kernel_img_mul_32[4] + kernel_img_mul_32[5] + 
                kernel_img_mul_32[6] + kernel_img_mul_32[7] + kernel_img_mul_32[8] + 
                kernel_img_mul_32[9] + kernel_img_mul_32[10] + kernel_img_mul_32[11] + 
                kernel_img_mul_32[12] + kernel_img_mul_32[13] + kernel_img_mul_32[14] + 
                kernel_img_mul_32[15] + kernel_img_mul_32[16] + kernel_img_mul_32[17] + 
                kernel_img_mul_32[18] + kernel_img_mul_32[19] + kernel_img_mul_32[20] + 
                kernel_img_mul_32[21] + kernel_img_mul_32[22] + kernel_img_mul_32[23] + 
                kernel_img_mul_32[24] + kernel_img_mul_32[25] + kernel_img_mul_32[26] + 
                kernel_img_mul_32[27] + kernel_img_mul_32[28] + kernel_img_mul_32[29] + 
                kernel_img_mul_32[30] + kernel_img_mul_32[31] + kernel_img_mul_32[32] + 
                kernel_img_mul_32[33] + kernel_img_mul_32[34] + kernel_img_mul_32[35] + 
                kernel_img_mul_32[36] + kernel_img_mul_32[37] + kernel_img_mul_32[38] + 
                kernel_img_mul_32[39] + kernel_img_mul_32[40] + kernel_img_mul_32[41] + 
                kernel_img_mul_32[42] + kernel_img_mul_32[43] + kernel_img_mul_32[44] + 
                kernel_img_mul_32[45] + kernel_img_mul_32[46] + kernel_img_mul_32[47] + 
                kernel_img_mul_32[48];
wire  [39:0]  kernel_img_mul_33[0:48];
assign kernel_img_mul_33[0] = layer0[33][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_33[1] = layer0[33][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_33[2] = layer0[33][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_33[3] = layer0[33][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_33[4] = layer0[33][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_33[5] = layer0[33][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_33[6] = layer0[33][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_33[7] = layer1[33][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_33[8] = layer1[33][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_33[9] = layer1[33][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_33[10] = layer1[33][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_33[11] = layer1[33][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_33[12] = layer1[33][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_33[13] = layer1[33][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_33[14] = layer2[33][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_33[15] = layer2[33][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_33[16] = layer2[33][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_33[17] = layer2[33][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_33[18] = layer2[33][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_33[19] = layer2[33][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_33[20] = layer2[33][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_33[21] = layer3[33][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_33[22] = layer3[33][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_33[23] = layer3[33][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_33[24] = layer3[33][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_33[25] = layer3[33][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_33[26] = layer3[33][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_33[27] = layer3[33][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_33[28] = layer4[33][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_33[29] = layer4[33][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_33[30] = layer4[33][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_33[31] = layer4[33][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_33[32] = layer4[33][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_33[33] = layer4[33][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_33[34] = layer4[33][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_33[35] = layer5[33][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_33[36] = layer5[33][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_33[37] = layer5[33][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_33[38] = layer5[33][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_33[39] = layer5[33][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_33[40] = layer5[33][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_33[41] = layer5[33][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_33[42] = layer6[33][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_33[43] = layer6[33][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_33[44] = layer6[33][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_33[45] = layer6[33][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_33[46] = layer6[33][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_33[47] = layer6[33][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_33[48] = layer6[33][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_33 = kernel_img_mul_33[0] + kernel_img_mul_33[1] + kernel_img_mul_33[2] + 
                kernel_img_mul_33[3] + kernel_img_mul_33[4] + kernel_img_mul_33[5] + 
                kernel_img_mul_33[6] + kernel_img_mul_33[7] + kernel_img_mul_33[8] + 
                kernel_img_mul_33[9] + kernel_img_mul_33[10] + kernel_img_mul_33[11] + 
                kernel_img_mul_33[12] + kernel_img_mul_33[13] + kernel_img_mul_33[14] + 
                kernel_img_mul_33[15] + kernel_img_mul_33[16] + kernel_img_mul_33[17] + 
                kernel_img_mul_33[18] + kernel_img_mul_33[19] + kernel_img_mul_33[20] + 
                kernel_img_mul_33[21] + kernel_img_mul_33[22] + kernel_img_mul_33[23] + 
                kernel_img_mul_33[24] + kernel_img_mul_33[25] + kernel_img_mul_33[26] + 
                kernel_img_mul_33[27] + kernel_img_mul_33[28] + kernel_img_mul_33[29] + 
                kernel_img_mul_33[30] + kernel_img_mul_33[31] + kernel_img_mul_33[32] + 
                kernel_img_mul_33[33] + kernel_img_mul_33[34] + kernel_img_mul_33[35] + 
                kernel_img_mul_33[36] + kernel_img_mul_33[37] + kernel_img_mul_33[38] + 
                kernel_img_mul_33[39] + kernel_img_mul_33[40] + kernel_img_mul_33[41] + 
                kernel_img_mul_33[42] + kernel_img_mul_33[43] + kernel_img_mul_33[44] + 
                kernel_img_mul_33[45] + kernel_img_mul_33[46] + kernel_img_mul_33[47] + 
                kernel_img_mul_33[48];
wire  [39:0]  kernel_img_mul_34[0:48];
assign kernel_img_mul_34[0] = layer0[34][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_34[1] = layer0[34][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_34[2] = layer0[34][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_34[3] = layer0[34][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_34[4] = layer0[34][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_34[5] = layer0[34][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_34[6] = layer0[34][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_34[7] = layer1[34][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_34[8] = layer1[34][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_34[9] = layer1[34][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_34[10] = layer1[34][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_34[11] = layer1[34][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_34[12] = layer1[34][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_34[13] = layer1[34][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_34[14] = layer2[34][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_34[15] = layer2[34][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_34[16] = layer2[34][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_34[17] = layer2[34][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_34[18] = layer2[34][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_34[19] = layer2[34][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_34[20] = layer2[34][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_34[21] = layer3[34][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_34[22] = layer3[34][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_34[23] = layer3[34][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_34[24] = layer3[34][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_34[25] = layer3[34][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_34[26] = layer3[34][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_34[27] = layer3[34][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_34[28] = layer4[34][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_34[29] = layer4[34][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_34[30] = layer4[34][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_34[31] = layer4[34][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_34[32] = layer4[34][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_34[33] = layer4[34][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_34[34] = layer4[34][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_34[35] = layer5[34][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_34[36] = layer5[34][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_34[37] = layer5[34][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_34[38] = layer5[34][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_34[39] = layer5[34][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_34[40] = layer5[34][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_34[41] = layer5[34][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_34[42] = layer6[34][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_34[43] = layer6[34][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_34[44] = layer6[34][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_34[45] = layer6[34][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_34[46] = layer6[34][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_34[47] = layer6[34][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_34[48] = layer6[34][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_34 = kernel_img_mul_34[0] + kernel_img_mul_34[1] + kernel_img_mul_34[2] + 
                kernel_img_mul_34[3] + kernel_img_mul_34[4] + kernel_img_mul_34[5] + 
                kernel_img_mul_34[6] + kernel_img_mul_34[7] + kernel_img_mul_34[8] + 
                kernel_img_mul_34[9] + kernel_img_mul_34[10] + kernel_img_mul_34[11] + 
                kernel_img_mul_34[12] + kernel_img_mul_34[13] + kernel_img_mul_34[14] + 
                kernel_img_mul_34[15] + kernel_img_mul_34[16] + kernel_img_mul_34[17] + 
                kernel_img_mul_34[18] + kernel_img_mul_34[19] + kernel_img_mul_34[20] + 
                kernel_img_mul_34[21] + kernel_img_mul_34[22] + kernel_img_mul_34[23] + 
                kernel_img_mul_34[24] + kernel_img_mul_34[25] + kernel_img_mul_34[26] + 
                kernel_img_mul_34[27] + kernel_img_mul_34[28] + kernel_img_mul_34[29] + 
                kernel_img_mul_34[30] + kernel_img_mul_34[31] + kernel_img_mul_34[32] + 
                kernel_img_mul_34[33] + kernel_img_mul_34[34] + kernel_img_mul_34[35] + 
                kernel_img_mul_34[36] + kernel_img_mul_34[37] + kernel_img_mul_34[38] + 
                kernel_img_mul_34[39] + kernel_img_mul_34[40] + kernel_img_mul_34[41] + 
                kernel_img_mul_34[42] + kernel_img_mul_34[43] + kernel_img_mul_34[44] + 
                kernel_img_mul_34[45] + kernel_img_mul_34[46] + kernel_img_mul_34[47] + 
                kernel_img_mul_34[48];
wire  [39:0]  kernel_img_mul_35[0:48];
assign kernel_img_mul_35[0] = layer0[35][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_35[1] = layer0[35][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_35[2] = layer0[35][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_35[3] = layer0[35][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_35[4] = layer0[35][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_35[5] = layer0[35][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_35[6] = layer0[35][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_35[7] = layer1[35][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_35[8] = layer1[35][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_35[9] = layer1[35][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_35[10] = layer1[35][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_35[11] = layer1[35][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_35[12] = layer1[35][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_35[13] = layer1[35][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_35[14] = layer2[35][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_35[15] = layer2[35][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_35[16] = layer2[35][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_35[17] = layer2[35][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_35[18] = layer2[35][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_35[19] = layer2[35][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_35[20] = layer2[35][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_35[21] = layer3[35][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_35[22] = layer3[35][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_35[23] = layer3[35][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_35[24] = layer3[35][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_35[25] = layer3[35][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_35[26] = layer3[35][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_35[27] = layer3[35][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_35[28] = layer4[35][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_35[29] = layer4[35][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_35[30] = layer4[35][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_35[31] = layer4[35][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_35[32] = layer4[35][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_35[33] = layer4[35][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_35[34] = layer4[35][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_35[35] = layer5[35][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_35[36] = layer5[35][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_35[37] = layer5[35][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_35[38] = layer5[35][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_35[39] = layer5[35][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_35[40] = layer5[35][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_35[41] = layer5[35][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_35[42] = layer6[35][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_35[43] = layer6[35][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_35[44] = layer6[35][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_35[45] = layer6[35][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_35[46] = layer6[35][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_35[47] = layer6[35][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_35[48] = layer6[35][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_35 = kernel_img_mul_35[0] + kernel_img_mul_35[1] + kernel_img_mul_35[2] + 
                kernel_img_mul_35[3] + kernel_img_mul_35[4] + kernel_img_mul_35[5] + 
                kernel_img_mul_35[6] + kernel_img_mul_35[7] + kernel_img_mul_35[8] + 
                kernel_img_mul_35[9] + kernel_img_mul_35[10] + kernel_img_mul_35[11] + 
                kernel_img_mul_35[12] + kernel_img_mul_35[13] + kernel_img_mul_35[14] + 
                kernel_img_mul_35[15] + kernel_img_mul_35[16] + kernel_img_mul_35[17] + 
                kernel_img_mul_35[18] + kernel_img_mul_35[19] + kernel_img_mul_35[20] + 
                kernel_img_mul_35[21] + kernel_img_mul_35[22] + kernel_img_mul_35[23] + 
                kernel_img_mul_35[24] + kernel_img_mul_35[25] + kernel_img_mul_35[26] + 
                kernel_img_mul_35[27] + kernel_img_mul_35[28] + kernel_img_mul_35[29] + 
                kernel_img_mul_35[30] + kernel_img_mul_35[31] + kernel_img_mul_35[32] + 
                kernel_img_mul_35[33] + kernel_img_mul_35[34] + kernel_img_mul_35[35] + 
                kernel_img_mul_35[36] + kernel_img_mul_35[37] + kernel_img_mul_35[38] + 
                kernel_img_mul_35[39] + kernel_img_mul_35[40] + kernel_img_mul_35[41] + 
                kernel_img_mul_35[42] + kernel_img_mul_35[43] + kernel_img_mul_35[44] + 
                kernel_img_mul_35[45] + kernel_img_mul_35[46] + kernel_img_mul_35[47] + 
                kernel_img_mul_35[48];
wire  [39:0]  kernel_img_mul_36[0:48];
assign kernel_img_mul_36[0] = layer0[36][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_36[1] = layer0[36][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_36[2] = layer0[36][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_36[3] = layer0[36][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_36[4] = layer0[36][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_36[5] = layer0[36][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_36[6] = layer0[36][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_36[7] = layer1[36][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_36[8] = layer1[36][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_36[9] = layer1[36][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_36[10] = layer1[36][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_36[11] = layer1[36][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_36[12] = layer1[36][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_36[13] = layer1[36][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_36[14] = layer2[36][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_36[15] = layer2[36][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_36[16] = layer2[36][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_36[17] = layer2[36][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_36[18] = layer2[36][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_36[19] = layer2[36][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_36[20] = layer2[36][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_36[21] = layer3[36][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_36[22] = layer3[36][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_36[23] = layer3[36][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_36[24] = layer3[36][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_36[25] = layer3[36][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_36[26] = layer3[36][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_36[27] = layer3[36][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_36[28] = layer4[36][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_36[29] = layer4[36][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_36[30] = layer4[36][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_36[31] = layer4[36][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_36[32] = layer4[36][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_36[33] = layer4[36][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_36[34] = layer4[36][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_36[35] = layer5[36][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_36[36] = layer5[36][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_36[37] = layer5[36][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_36[38] = layer5[36][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_36[39] = layer5[36][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_36[40] = layer5[36][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_36[41] = layer5[36][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_36[42] = layer6[36][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_36[43] = layer6[36][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_36[44] = layer6[36][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_36[45] = layer6[36][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_36[46] = layer6[36][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_36[47] = layer6[36][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_36[48] = layer6[36][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_36 = kernel_img_mul_36[0] + kernel_img_mul_36[1] + kernel_img_mul_36[2] + 
                kernel_img_mul_36[3] + kernel_img_mul_36[4] + kernel_img_mul_36[5] + 
                kernel_img_mul_36[6] + kernel_img_mul_36[7] + kernel_img_mul_36[8] + 
                kernel_img_mul_36[9] + kernel_img_mul_36[10] + kernel_img_mul_36[11] + 
                kernel_img_mul_36[12] + kernel_img_mul_36[13] + kernel_img_mul_36[14] + 
                kernel_img_mul_36[15] + kernel_img_mul_36[16] + kernel_img_mul_36[17] + 
                kernel_img_mul_36[18] + kernel_img_mul_36[19] + kernel_img_mul_36[20] + 
                kernel_img_mul_36[21] + kernel_img_mul_36[22] + kernel_img_mul_36[23] + 
                kernel_img_mul_36[24] + kernel_img_mul_36[25] + kernel_img_mul_36[26] + 
                kernel_img_mul_36[27] + kernel_img_mul_36[28] + kernel_img_mul_36[29] + 
                kernel_img_mul_36[30] + kernel_img_mul_36[31] + kernel_img_mul_36[32] + 
                kernel_img_mul_36[33] + kernel_img_mul_36[34] + kernel_img_mul_36[35] + 
                kernel_img_mul_36[36] + kernel_img_mul_36[37] + kernel_img_mul_36[38] + 
                kernel_img_mul_36[39] + kernel_img_mul_36[40] + kernel_img_mul_36[41] + 
                kernel_img_mul_36[42] + kernel_img_mul_36[43] + kernel_img_mul_36[44] + 
                kernel_img_mul_36[45] + kernel_img_mul_36[46] + kernel_img_mul_36[47] + 
                kernel_img_mul_36[48];
wire  [39:0]  kernel_img_mul_37[0:48];
assign kernel_img_mul_37[0] = layer0[37][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_37[1] = layer0[37][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_37[2] = layer0[37][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_37[3] = layer0[37][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_37[4] = layer0[37][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_37[5] = layer0[37][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_37[6] = layer0[37][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_37[7] = layer1[37][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_37[8] = layer1[37][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_37[9] = layer1[37][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_37[10] = layer1[37][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_37[11] = layer1[37][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_37[12] = layer1[37][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_37[13] = layer1[37][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_37[14] = layer2[37][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_37[15] = layer2[37][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_37[16] = layer2[37][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_37[17] = layer2[37][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_37[18] = layer2[37][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_37[19] = layer2[37][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_37[20] = layer2[37][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_37[21] = layer3[37][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_37[22] = layer3[37][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_37[23] = layer3[37][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_37[24] = layer3[37][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_37[25] = layer3[37][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_37[26] = layer3[37][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_37[27] = layer3[37][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_37[28] = layer4[37][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_37[29] = layer4[37][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_37[30] = layer4[37][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_37[31] = layer4[37][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_37[32] = layer4[37][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_37[33] = layer4[37][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_37[34] = layer4[37][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_37[35] = layer5[37][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_37[36] = layer5[37][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_37[37] = layer5[37][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_37[38] = layer5[37][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_37[39] = layer5[37][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_37[40] = layer5[37][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_37[41] = layer5[37][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_37[42] = layer6[37][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_37[43] = layer6[37][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_37[44] = layer6[37][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_37[45] = layer6[37][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_37[46] = layer6[37][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_37[47] = layer6[37][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_37[48] = layer6[37][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_37 = kernel_img_mul_37[0] + kernel_img_mul_37[1] + kernel_img_mul_37[2] + 
                kernel_img_mul_37[3] + kernel_img_mul_37[4] + kernel_img_mul_37[5] + 
                kernel_img_mul_37[6] + kernel_img_mul_37[7] + kernel_img_mul_37[8] + 
                kernel_img_mul_37[9] + kernel_img_mul_37[10] + kernel_img_mul_37[11] + 
                kernel_img_mul_37[12] + kernel_img_mul_37[13] + kernel_img_mul_37[14] + 
                kernel_img_mul_37[15] + kernel_img_mul_37[16] + kernel_img_mul_37[17] + 
                kernel_img_mul_37[18] + kernel_img_mul_37[19] + kernel_img_mul_37[20] + 
                kernel_img_mul_37[21] + kernel_img_mul_37[22] + kernel_img_mul_37[23] + 
                kernel_img_mul_37[24] + kernel_img_mul_37[25] + kernel_img_mul_37[26] + 
                kernel_img_mul_37[27] + kernel_img_mul_37[28] + kernel_img_mul_37[29] + 
                kernel_img_mul_37[30] + kernel_img_mul_37[31] + kernel_img_mul_37[32] + 
                kernel_img_mul_37[33] + kernel_img_mul_37[34] + kernel_img_mul_37[35] + 
                kernel_img_mul_37[36] + kernel_img_mul_37[37] + kernel_img_mul_37[38] + 
                kernel_img_mul_37[39] + kernel_img_mul_37[40] + kernel_img_mul_37[41] + 
                kernel_img_mul_37[42] + kernel_img_mul_37[43] + kernel_img_mul_37[44] + 
                kernel_img_mul_37[45] + kernel_img_mul_37[46] + kernel_img_mul_37[47] + 
                kernel_img_mul_37[48];
wire  [39:0]  kernel_img_mul_38[0:48];
assign kernel_img_mul_38[0] = layer0[38][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_38[1] = layer0[38][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_38[2] = layer0[38][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_38[3] = layer0[38][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_38[4] = layer0[38][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_38[5] = layer0[38][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_38[6] = layer0[38][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_38[7] = layer1[38][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_38[8] = layer1[38][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_38[9] = layer1[38][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_38[10] = layer1[38][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_38[11] = layer1[38][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_38[12] = layer1[38][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_38[13] = layer1[38][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_38[14] = layer2[38][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_38[15] = layer2[38][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_38[16] = layer2[38][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_38[17] = layer2[38][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_38[18] = layer2[38][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_38[19] = layer2[38][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_38[20] = layer2[38][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_38[21] = layer3[38][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_38[22] = layer3[38][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_38[23] = layer3[38][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_38[24] = layer3[38][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_38[25] = layer3[38][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_38[26] = layer3[38][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_38[27] = layer3[38][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_38[28] = layer4[38][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_38[29] = layer4[38][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_38[30] = layer4[38][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_38[31] = layer4[38][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_38[32] = layer4[38][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_38[33] = layer4[38][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_38[34] = layer4[38][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_38[35] = layer5[38][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_38[36] = layer5[38][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_38[37] = layer5[38][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_38[38] = layer5[38][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_38[39] = layer5[38][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_38[40] = layer5[38][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_38[41] = layer5[38][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_38[42] = layer6[38][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_38[43] = layer6[38][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_38[44] = layer6[38][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_38[45] = layer6[38][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_38[46] = layer6[38][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_38[47] = layer6[38][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_38[48] = layer6[38][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_38 = kernel_img_mul_38[0] + kernel_img_mul_38[1] + kernel_img_mul_38[2] + 
                kernel_img_mul_38[3] + kernel_img_mul_38[4] + kernel_img_mul_38[5] + 
                kernel_img_mul_38[6] + kernel_img_mul_38[7] + kernel_img_mul_38[8] + 
                kernel_img_mul_38[9] + kernel_img_mul_38[10] + kernel_img_mul_38[11] + 
                kernel_img_mul_38[12] + kernel_img_mul_38[13] + kernel_img_mul_38[14] + 
                kernel_img_mul_38[15] + kernel_img_mul_38[16] + kernel_img_mul_38[17] + 
                kernel_img_mul_38[18] + kernel_img_mul_38[19] + kernel_img_mul_38[20] + 
                kernel_img_mul_38[21] + kernel_img_mul_38[22] + kernel_img_mul_38[23] + 
                kernel_img_mul_38[24] + kernel_img_mul_38[25] + kernel_img_mul_38[26] + 
                kernel_img_mul_38[27] + kernel_img_mul_38[28] + kernel_img_mul_38[29] + 
                kernel_img_mul_38[30] + kernel_img_mul_38[31] + kernel_img_mul_38[32] + 
                kernel_img_mul_38[33] + kernel_img_mul_38[34] + kernel_img_mul_38[35] + 
                kernel_img_mul_38[36] + kernel_img_mul_38[37] + kernel_img_mul_38[38] + 
                kernel_img_mul_38[39] + kernel_img_mul_38[40] + kernel_img_mul_38[41] + 
                kernel_img_mul_38[42] + kernel_img_mul_38[43] + kernel_img_mul_38[44] + 
                kernel_img_mul_38[45] + kernel_img_mul_38[46] + kernel_img_mul_38[47] + 
                kernel_img_mul_38[48];
wire  [39:0]  kernel_img_mul_39[0:48];
assign kernel_img_mul_39[0] = layer0[39][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_39[1] = layer0[39][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_39[2] = layer0[39][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_39[3] = layer0[39][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_39[4] = layer0[39][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_39[5] = layer0[39][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_39[6] = layer0[39][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_39[7] = layer1[39][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_39[8] = layer1[39][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_39[9] = layer1[39][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_39[10] = layer1[39][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_39[11] = layer1[39][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_39[12] = layer1[39][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_39[13] = layer1[39][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_39[14] = layer2[39][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_39[15] = layer2[39][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_39[16] = layer2[39][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_39[17] = layer2[39][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_39[18] = layer2[39][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_39[19] = layer2[39][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_39[20] = layer2[39][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_39[21] = layer3[39][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_39[22] = layer3[39][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_39[23] = layer3[39][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_39[24] = layer3[39][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_39[25] = layer3[39][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_39[26] = layer3[39][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_39[27] = layer3[39][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_39[28] = layer4[39][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_39[29] = layer4[39][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_39[30] = layer4[39][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_39[31] = layer4[39][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_39[32] = layer4[39][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_39[33] = layer4[39][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_39[34] = layer4[39][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_39[35] = layer5[39][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_39[36] = layer5[39][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_39[37] = layer5[39][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_39[38] = layer5[39][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_39[39] = layer5[39][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_39[40] = layer5[39][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_39[41] = layer5[39][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_39[42] = layer6[39][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_39[43] = layer6[39][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_39[44] = layer6[39][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_39[45] = layer6[39][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_39[46] = layer6[39][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_39[47] = layer6[39][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_39[48] = layer6[39][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_39 = kernel_img_mul_39[0] + kernel_img_mul_39[1] + kernel_img_mul_39[2] + 
                kernel_img_mul_39[3] + kernel_img_mul_39[4] + kernel_img_mul_39[5] + 
                kernel_img_mul_39[6] + kernel_img_mul_39[7] + kernel_img_mul_39[8] + 
                kernel_img_mul_39[9] + kernel_img_mul_39[10] + kernel_img_mul_39[11] + 
                kernel_img_mul_39[12] + kernel_img_mul_39[13] + kernel_img_mul_39[14] + 
                kernel_img_mul_39[15] + kernel_img_mul_39[16] + kernel_img_mul_39[17] + 
                kernel_img_mul_39[18] + kernel_img_mul_39[19] + kernel_img_mul_39[20] + 
                kernel_img_mul_39[21] + kernel_img_mul_39[22] + kernel_img_mul_39[23] + 
                kernel_img_mul_39[24] + kernel_img_mul_39[25] + kernel_img_mul_39[26] + 
                kernel_img_mul_39[27] + kernel_img_mul_39[28] + kernel_img_mul_39[29] + 
                kernel_img_mul_39[30] + kernel_img_mul_39[31] + kernel_img_mul_39[32] + 
                kernel_img_mul_39[33] + kernel_img_mul_39[34] + kernel_img_mul_39[35] + 
                kernel_img_mul_39[36] + kernel_img_mul_39[37] + kernel_img_mul_39[38] + 
                kernel_img_mul_39[39] + kernel_img_mul_39[40] + kernel_img_mul_39[41] + 
                kernel_img_mul_39[42] + kernel_img_mul_39[43] + kernel_img_mul_39[44] + 
                kernel_img_mul_39[45] + kernel_img_mul_39[46] + kernel_img_mul_39[47] + 
                kernel_img_mul_39[48];
wire  [39:0]  kernel_img_mul_40[0:48];
assign kernel_img_mul_40[0] = layer0[40][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_40[1] = layer0[40][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_40[2] = layer0[40][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_40[3] = layer0[40][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_40[4] = layer0[40][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_40[5] = layer0[40][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_40[6] = layer0[40][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_40[7] = layer1[40][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_40[8] = layer1[40][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_40[9] = layer1[40][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_40[10] = layer1[40][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_40[11] = layer1[40][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_40[12] = layer1[40][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_40[13] = layer1[40][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_40[14] = layer2[40][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_40[15] = layer2[40][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_40[16] = layer2[40][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_40[17] = layer2[40][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_40[18] = layer2[40][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_40[19] = layer2[40][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_40[20] = layer2[40][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_40[21] = layer3[40][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_40[22] = layer3[40][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_40[23] = layer3[40][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_40[24] = layer3[40][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_40[25] = layer3[40][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_40[26] = layer3[40][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_40[27] = layer3[40][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_40[28] = layer4[40][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_40[29] = layer4[40][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_40[30] = layer4[40][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_40[31] = layer4[40][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_40[32] = layer4[40][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_40[33] = layer4[40][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_40[34] = layer4[40][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_40[35] = layer5[40][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_40[36] = layer5[40][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_40[37] = layer5[40][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_40[38] = layer5[40][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_40[39] = layer5[40][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_40[40] = layer5[40][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_40[41] = layer5[40][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_40[42] = layer6[40][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_40[43] = layer6[40][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_40[44] = layer6[40][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_40[45] = layer6[40][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_40[46] = layer6[40][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_40[47] = layer6[40][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_40[48] = layer6[40][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_40 = kernel_img_mul_40[0] + kernel_img_mul_40[1] + kernel_img_mul_40[2] + 
                kernel_img_mul_40[3] + kernel_img_mul_40[4] + kernel_img_mul_40[5] + 
                kernel_img_mul_40[6] + kernel_img_mul_40[7] + kernel_img_mul_40[8] + 
                kernel_img_mul_40[9] + kernel_img_mul_40[10] + kernel_img_mul_40[11] + 
                kernel_img_mul_40[12] + kernel_img_mul_40[13] + kernel_img_mul_40[14] + 
                kernel_img_mul_40[15] + kernel_img_mul_40[16] + kernel_img_mul_40[17] + 
                kernel_img_mul_40[18] + kernel_img_mul_40[19] + kernel_img_mul_40[20] + 
                kernel_img_mul_40[21] + kernel_img_mul_40[22] + kernel_img_mul_40[23] + 
                kernel_img_mul_40[24] + kernel_img_mul_40[25] + kernel_img_mul_40[26] + 
                kernel_img_mul_40[27] + kernel_img_mul_40[28] + kernel_img_mul_40[29] + 
                kernel_img_mul_40[30] + kernel_img_mul_40[31] + kernel_img_mul_40[32] + 
                kernel_img_mul_40[33] + kernel_img_mul_40[34] + kernel_img_mul_40[35] + 
                kernel_img_mul_40[36] + kernel_img_mul_40[37] + kernel_img_mul_40[38] + 
                kernel_img_mul_40[39] + kernel_img_mul_40[40] + kernel_img_mul_40[41] + 
                kernel_img_mul_40[42] + kernel_img_mul_40[43] + kernel_img_mul_40[44] + 
                kernel_img_mul_40[45] + kernel_img_mul_40[46] + kernel_img_mul_40[47] + 
                kernel_img_mul_40[48];
wire  [39:0]  kernel_img_mul_41[0:48];
assign kernel_img_mul_41[0] = layer0[41][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_41[1] = layer0[41][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_41[2] = layer0[41][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_41[3] = layer0[41][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_41[4] = layer0[41][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_41[5] = layer0[41][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_41[6] = layer0[41][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_41[7] = layer1[41][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_41[8] = layer1[41][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_41[9] = layer1[41][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_41[10] = layer1[41][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_41[11] = layer1[41][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_41[12] = layer1[41][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_41[13] = layer1[41][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_41[14] = layer2[41][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_41[15] = layer2[41][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_41[16] = layer2[41][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_41[17] = layer2[41][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_41[18] = layer2[41][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_41[19] = layer2[41][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_41[20] = layer2[41][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_41[21] = layer3[41][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_41[22] = layer3[41][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_41[23] = layer3[41][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_41[24] = layer3[41][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_41[25] = layer3[41][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_41[26] = layer3[41][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_41[27] = layer3[41][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_41[28] = layer4[41][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_41[29] = layer4[41][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_41[30] = layer4[41][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_41[31] = layer4[41][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_41[32] = layer4[41][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_41[33] = layer4[41][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_41[34] = layer4[41][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_41[35] = layer5[41][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_41[36] = layer5[41][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_41[37] = layer5[41][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_41[38] = layer5[41][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_41[39] = layer5[41][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_41[40] = layer5[41][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_41[41] = layer5[41][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_41[42] = layer6[41][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_41[43] = layer6[41][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_41[44] = layer6[41][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_41[45] = layer6[41][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_41[46] = layer6[41][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_41[47] = layer6[41][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_41[48] = layer6[41][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_41 = kernel_img_mul_41[0] + kernel_img_mul_41[1] + kernel_img_mul_41[2] + 
                kernel_img_mul_41[3] + kernel_img_mul_41[4] + kernel_img_mul_41[5] + 
                kernel_img_mul_41[6] + kernel_img_mul_41[7] + kernel_img_mul_41[8] + 
                kernel_img_mul_41[9] + kernel_img_mul_41[10] + kernel_img_mul_41[11] + 
                kernel_img_mul_41[12] + kernel_img_mul_41[13] + kernel_img_mul_41[14] + 
                kernel_img_mul_41[15] + kernel_img_mul_41[16] + kernel_img_mul_41[17] + 
                kernel_img_mul_41[18] + kernel_img_mul_41[19] + kernel_img_mul_41[20] + 
                kernel_img_mul_41[21] + kernel_img_mul_41[22] + kernel_img_mul_41[23] + 
                kernel_img_mul_41[24] + kernel_img_mul_41[25] + kernel_img_mul_41[26] + 
                kernel_img_mul_41[27] + kernel_img_mul_41[28] + kernel_img_mul_41[29] + 
                kernel_img_mul_41[30] + kernel_img_mul_41[31] + kernel_img_mul_41[32] + 
                kernel_img_mul_41[33] + kernel_img_mul_41[34] + kernel_img_mul_41[35] + 
                kernel_img_mul_41[36] + kernel_img_mul_41[37] + kernel_img_mul_41[38] + 
                kernel_img_mul_41[39] + kernel_img_mul_41[40] + kernel_img_mul_41[41] + 
                kernel_img_mul_41[42] + kernel_img_mul_41[43] + kernel_img_mul_41[44] + 
                kernel_img_mul_41[45] + kernel_img_mul_41[46] + kernel_img_mul_41[47] + 
                kernel_img_mul_41[48];
wire  [39:0]  kernel_img_mul_42[0:48];
assign kernel_img_mul_42[0] = layer0[42][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_42[1] = layer0[42][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_42[2] = layer0[42][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_42[3] = layer0[42][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_42[4] = layer0[42][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_42[5] = layer0[42][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_42[6] = layer0[42][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_42[7] = layer1[42][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_42[8] = layer1[42][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_42[9] = layer1[42][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_42[10] = layer1[42][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_42[11] = layer1[42][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_42[12] = layer1[42][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_42[13] = layer1[42][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_42[14] = layer2[42][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_42[15] = layer2[42][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_42[16] = layer2[42][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_42[17] = layer2[42][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_42[18] = layer2[42][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_42[19] = layer2[42][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_42[20] = layer2[42][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_42[21] = layer3[42][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_42[22] = layer3[42][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_42[23] = layer3[42][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_42[24] = layer3[42][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_42[25] = layer3[42][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_42[26] = layer3[42][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_42[27] = layer3[42][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_42[28] = layer4[42][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_42[29] = layer4[42][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_42[30] = layer4[42][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_42[31] = layer4[42][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_42[32] = layer4[42][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_42[33] = layer4[42][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_42[34] = layer4[42][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_42[35] = layer5[42][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_42[36] = layer5[42][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_42[37] = layer5[42][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_42[38] = layer5[42][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_42[39] = layer5[42][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_42[40] = layer5[42][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_42[41] = layer5[42][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_42[42] = layer6[42][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_42[43] = layer6[42][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_42[44] = layer6[42][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_42[45] = layer6[42][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_42[46] = layer6[42][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_42[47] = layer6[42][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_42[48] = layer6[42][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_42 = kernel_img_mul_42[0] + kernel_img_mul_42[1] + kernel_img_mul_42[2] + 
                kernel_img_mul_42[3] + kernel_img_mul_42[4] + kernel_img_mul_42[5] + 
                kernel_img_mul_42[6] + kernel_img_mul_42[7] + kernel_img_mul_42[8] + 
                kernel_img_mul_42[9] + kernel_img_mul_42[10] + kernel_img_mul_42[11] + 
                kernel_img_mul_42[12] + kernel_img_mul_42[13] + kernel_img_mul_42[14] + 
                kernel_img_mul_42[15] + kernel_img_mul_42[16] + kernel_img_mul_42[17] + 
                kernel_img_mul_42[18] + kernel_img_mul_42[19] + kernel_img_mul_42[20] + 
                kernel_img_mul_42[21] + kernel_img_mul_42[22] + kernel_img_mul_42[23] + 
                kernel_img_mul_42[24] + kernel_img_mul_42[25] + kernel_img_mul_42[26] + 
                kernel_img_mul_42[27] + kernel_img_mul_42[28] + kernel_img_mul_42[29] + 
                kernel_img_mul_42[30] + kernel_img_mul_42[31] + kernel_img_mul_42[32] + 
                kernel_img_mul_42[33] + kernel_img_mul_42[34] + kernel_img_mul_42[35] + 
                kernel_img_mul_42[36] + kernel_img_mul_42[37] + kernel_img_mul_42[38] + 
                kernel_img_mul_42[39] + kernel_img_mul_42[40] + kernel_img_mul_42[41] + 
                kernel_img_mul_42[42] + kernel_img_mul_42[43] + kernel_img_mul_42[44] + 
                kernel_img_mul_42[45] + kernel_img_mul_42[46] + kernel_img_mul_42[47] + 
                kernel_img_mul_42[48];
wire  [39:0]  kernel_img_mul_43[0:48];
assign kernel_img_mul_43[0] = layer0[43][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_43[1] = layer0[43][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_43[2] = layer0[43][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_43[3] = layer0[43][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_43[4] = layer0[43][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_43[5] = layer0[43][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_43[6] = layer0[43][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_43[7] = layer1[43][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_43[8] = layer1[43][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_43[9] = layer1[43][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_43[10] = layer1[43][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_43[11] = layer1[43][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_43[12] = layer1[43][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_43[13] = layer1[43][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_43[14] = layer2[43][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_43[15] = layer2[43][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_43[16] = layer2[43][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_43[17] = layer2[43][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_43[18] = layer2[43][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_43[19] = layer2[43][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_43[20] = layer2[43][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_43[21] = layer3[43][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_43[22] = layer3[43][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_43[23] = layer3[43][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_43[24] = layer3[43][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_43[25] = layer3[43][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_43[26] = layer3[43][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_43[27] = layer3[43][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_43[28] = layer4[43][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_43[29] = layer4[43][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_43[30] = layer4[43][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_43[31] = layer4[43][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_43[32] = layer4[43][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_43[33] = layer4[43][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_43[34] = layer4[43][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_43[35] = layer5[43][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_43[36] = layer5[43][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_43[37] = layer5[43][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_43[38] = layer5[43][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_43[39] = layer5[43][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_43[40] = layer5[43][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_43[41] = layer5[43][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_43[42] = layer6[43][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_43[43] = layer6[43][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_43[44] = layer6[43][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_43[45] = layer6[43][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_43[46] = layer6[43][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_43[47] = layer6[43][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_43[48] = layer6[43][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_43 = kernel_img_mul_43[0] + kernel_img_mul_43[1] + kernel_img_mul_43[2] + 
                kernel_img_mul_43[3] + kernel_img_mul_43[4] + kernel_img_mul_43[5] + 
                kernel_img_mul_43[6] + kernel_img_mul_43[7] + kernel_img_mul_43[8] + 
                kernel_img_mul_43[9] + kernel_img_mul_43[10] + kernel_img_mul_43[11] + 
                kernel_img_mul_43[12] + kernel_img_mul_43[13] + kernel_img_mul_43[14] + 
                kernel_img_mul_43[15] + kernel_img_mul_43[16] + kernel_img_mul_43[17] + 
                kernel_img_mul_43[18] + kernel_img_mul_43[19] + kernel_img_mul_43[20] + 
                kernel_img_mul_43[21] + kernel_img_mul_43[22] + kernel_img_mul_43[23] + 
                kernel_img_mul_43[24] + kernel_img_mul_43[25] + kernel_img_mul_43[26] + 
                kernel_img_mul_43[27] + kernel_img_mul_43[28] + kernel_img_mul_43[29] + 
                kernel_img_mul_43[30] + kernel_img_mul_43[31] + kernel_img_mul_43[32] + 
                kernel_img_mul_43[33] + kernel_img_mul_43[34] + kernel_img_mul_43[35] + 
                kernel_img_mul_43[36] + kernel_img_mul_43[37] + kernel_img_mul_43[38] + 
                kernel_img_mul_43[39] + kernel_img_mul_43[40] + kernel_img_mul_43[41] + 
                kernel_img_mul_43[42] + kernel_img_mul_43[43] + kernel_img_mul_43[44] + 
                kernel_img_mul_43[45] + kernel_img_mul_43[46] + kernel_img_mul_43[47] + 
                kernel_img_mul_43[48];
wire  [39:0]  kernel_img_mul_44[0:48];
assign kernel_img_mul_44[0] = layer0[44][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_44[1] = layer0[44][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_44[2] = layer0[44][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_44[3] = layer0[44][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_44[4] = layer0[44][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_44[5] = layer0[44][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_44[6] = layer0[44][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_44[7] = layer1[44][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_44[8] = layer1[44][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_44[9] = layer1[44][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_44[10] = layer1[44][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_44[11] = layer1[44][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_44[12] = layer1[44][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_44[13] = layer1[44][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_44[14] = layer2[44][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_44[15] = layer2[44][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_44[16] = layer2[44][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_44[17] = layer2[44][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_44[18] = layer2[44][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_44[19] = layer2[44][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_44[20] = layer2[44][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_44[21] = layer3[44][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_44[22] = layer3[44][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_44[23] = layer3[44][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_44[24] = layer3[44][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_44[25] = layer3[44][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_44[26] = layer3[44][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_44[27] = layer3[44][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_44[28] = layer4[44][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_44[29] = layer4[44][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_44[30] = layer4[44][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_44[31] = layer4[44][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_44[32] = layer4[44][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_44[33] = layer4[44][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_44[34] = layer4[44][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_44[35] = layer5[44][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_44[36] = layer5[44][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_44[37] = layer5[44][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_44[38] = layer5[44][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_44[39] = layer5[44][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_44[40] = layer5[44][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_44[41] = layer5[44][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_44[42] = layer6[44][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_44[43] = layer6[44][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_44[44] = layer6[44][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_44[45] = layer6[44][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_44[46] = layer6[44][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_44[47] = layer6[44][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_44[48] = layer6[44][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_44 = kernel_img_mul_44[0] + kernel_img_mul_44[1] + kernel_img_mul_44[2] + 
                kernel_img_mul_44[3] + kernel_img_mul_44[4] + kernel_img_mul_44[5] + 
                kernel_img_mul_44[6] + kernel_img_mul_44[7] + kernel_img_mul_44[8] + 
                kernel_img_mul_44[9] + kernel_img_mul_44[10] + kernel_img_mul_44[11] + 
                kernel_img_mul_44[12] + kernel_img_mul_44[13] + kernel_img_mul_44[14] + 
                kernel_img_mul_44[15] + kernel_img_mul_44[16] + kernel_img_mul_44[17] + 
                kernel_img_mul_44[18] + kernel_img_mul_44[19] + kernel_img_mul_44[20] + 
                kernel_img_mul_44[21] + kernel_img_mul_44[22] + kernel_img_mul_44[23] + 
                kernel_img_mul_44[24] + kernel_img_mul_44[25] + kernel_img_mul_44[26] + 
                kernel_img_mul_44[27] + kernel_img_mul_44[28] + kernel_img_mul_44[29] + 
                kernel_img_mul_44[30] + kernel_img_mul_44[31] + kernel_img_mul_44[32] + 
                kernel_img_mul_44[33] + kernel_img_mul_44[34] + kernel_img_mul_44[35] + 
                kernel_img_mul_44[36] + kernel_img_mul_44[37] + kernel_img_mul_44[38] + 
                kernel_img_mul_44[39] + kernel_img_mul_44[40] + kernel_img_mul_44[41] + 
                kernel_img_mul_44[42] + kernel_img_mul_44[43] + kernel_img_mul_44[44] + 
                kernel_img_mul_44[45] + kernel_img_mul_44[46] + kernel_img_mul_44[47] + 
                kernel_img_mul_44[48];
wire  [39:0]  kernel_img_mul_45[0:48];
assign kernel_img_mul_45[0] = layer0[45][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_45[1] = layer0[45][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_45[2] = layer0[45][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_45[3] = layer0[45][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_45[4] = layer0[45][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_45[5] = layer0[45][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_45[6] = layer0[45][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_45[7] = layer1[45][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_45[8] = layer1[45][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_45[9] = layer1[45][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_45[10] = layer1[45][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_45[11] = layer1[45][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_45[12] = layer1[45][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_45[13] = layer1[45][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_45[14] = layer2[45][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_45[15] = layer2[45][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_45[16] = layer2[45][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_45[17] = layer2[45][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_45[18] = layer2[45][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_45[19] = layer2[45][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_45[20] = layer2[45][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_45[21] = layer3[45][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_45[22] = layer3[45][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_45[23] = layer3[45][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_45[24] = layer3[45][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_45[25] = layer3[45][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_45[26] = layer3[45][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_45[27] = layer3[45][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_45[28] = layer4[45][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_45[29] = layer4[45][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_45[30] = layer4[45][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_45[31] = layer4[45][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_45[32] = layer4[45][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_45[33] = layer4[45][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_45[34] = layer4[45][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_45[35] = layer5[45][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_45[36] = layer5[45][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_45[37] = layer5[45][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_45[38] = layer5[45][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_45[39] = layer5[45][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_45[40] = layer5[45][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_45[41] = layer5[45][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_45[42] = layer6[45][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_45[43] = layer6[45][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_45[44] = layer6[45][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_45[45] = layer6[45][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_45[46] = layer6[45][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_45[47] = layer6[45][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_45[48] = layer6[45][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_45 = kernel_img_mul_45[0] + kernel_img_mul_45[1] + kernel_img_mul_45[2] + 
                kernel_img_mul_45[3] + kernel_img_mul_45[4] + kernel_img_mul_45[5] + 
                kernel_img_mul_45[6] + kernel_img_mul_45[7] + kernel_img_mul_45[8] + 
                kernel_img_mul_45[9] + kernel_img_mul_45[10] + kernel_img_mul_45[11] + 
                kernel_img_mul_45[12] + kernel_img_mul_45[13] + kernel_img_mul_45[14] + 
                kernel_img_mul_45[15] + kernel_img_mul_45[16] + kernel_img_mul_45[17] + 
                kernel_img_mul_45[18] + kernel_img_mul_45[19] + kernel_img_mul_45[20] + 
                kernel_img_mul_45[21] + kernel_img_mul_45[22] + kernel_img_mul_45[23] + 
                kernel_img_mul_45[24] + kernel_img_mul_45[25] + kernel_img_mul_45[26] + 
                kernel_img_mul_45[27] + kernel_img_mul_45[28] + kernel_img_mul_45[29] + 
                kernel_img_mul_45[30] + kernel_img_mul_45[31] + kernel_img_mul_45[32] + 
                kernel_img_mul_45[33] + kernel_img_mul_45[34] + kernel_img_mul_45[35] + 
                kernel_img_mul_45[36] + kernel_img_mul_45[37] + kernel_img_mul_45[38] + 
                kernel_img_mul_45[39] + kernel_img_mul_45[40] + kernel_img_mul_45[41] + 
                kernel_img_mul_45[42] + kernel_img_mul_45[43] + kernel_img_mul_45[44] + 
                kernel_img_mul_45[45] + kernel_img_mul_45[46] + kernel_img_mul_45[47] + 
                kernel_img_mul_45[48];
wire  [39:0]  kernel_img_mul_46[0:48];
assign kernel_img_mul_46[0] = layer0[46][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_46[1] = layer0[46][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_46[2] = layer0[46][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_46[3] = layer0[46][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_46[4] = layer0[46][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_46[5] = layer0[46][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_46[6] = layer0[46][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_46[7] = layer1[46][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_46[8] = layer1[46][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_46[9] = layer1[46][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_46[10] = layer1[46][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_46[11] = layer1[46][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_46[12] = layer1[46][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_46[13] = layer1[46][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_46[14] = layer2[46][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_46[15] = layer2[46][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_46[16] = layer2[46][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_46[17] = layer2[46][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_46[18] = layer2[46][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_46[19] = layer2[46][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_46[20] = layer2[46][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_46[21] = layer3[46][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_46[22] = layer3[46][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_46[23] = layer3[46][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_46[24] = layer3[46][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_46[25] = layer3[46][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_46[26] = layer3[46][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_46[27] = layer3[46][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_46[28] = layer4[46][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_46[29] = layer4[46][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_46[30] = layer4[46][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_46[31] = layer4[46][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_46[32] = layer4[46][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_46[33] = layer4[46][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_46[34] = layer4[46][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_46[35] = layer5[46][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_46[36] = layer5[46][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_46[37] = layer5[46][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_46[38] = layer5[46][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_46[39] = layer5[46][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_46[40] = layer5[46][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_46[41] = layer5[46][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_46[42] = layer6[46][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_46[43] = layer6[46][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_46[44] = layer6[46][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_46[45] = layer6[46][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_46[46] = layer6[46][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_46[47] = layer6[46][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_46[48] = layer6[46][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_46 = kernel_img_mul_46[0] + kernel_img_mul_46[1] + kernel_img_mul_46[2] + 
                kernel_img_mul_46[3] + kernel_img_mul_46[4] + kernel_img_mul_46[5] + 
                kernel_img_mul_46[6] + kernel_img_mul_46[7] + kernel_img_mul_46[8] + 
                kernel_img_mul_46[9] + kernel_img_mul_46[10] + kernel_img_mul_46[11] + 
                kernel_img_mul_46[12] + kernel_img_mul_46[13] + kernel_img_mul_46[14] + 
                kernel_img_mul_46[15] + kernel_img_mul_46[16] + kernel_img_mul_46[17] + 
                kernel_img_mul_46[18] + kernel_img_mul_46[19] + kernel_img_mul_46[20] + 
                kernel_img_mul_46[21] + kernel_img_mul_46[22] + kernel_img_mul_46[23] + 
                kernel_img_mul_46[24] + kernel_img_mul_46[25] + kernel_img_mul_46[26] + 
                kernel_img_mul_46[27] + kernel_img_mul_46[28] + kernel_img_mul_46[29] + 
                kernel_img_mul_46[30] + kernel_img_mul_46[31] + kernel_img_mul_46[32] + 
                kernel_img_mul_46[33] + kernel_img_mul_46[34] + kernel_img_mul_46[35] + 
                kernel_img_mul_46[36] + kernel_img_mul_46[37] + kernel_img_mul_46[38] + 
                kernel_img_mul_46[39] + kernel_img_mul_46[40] + kernel_img_mul_46[41] + 
                kernel_img_mul_46[42] + kernel_img_mul_46[43] + kernel_img_mul_46[44] + 
                kernel_img_mul_46[45] + kernel_img_mul_46[46] + kernel_img_mul_46[47] + 
                kernel_img_mul_46[48];
wire  [39:0]  kernel_img_mul_47[0:48];
assign kernel_img_mul_47[0] = layer0[47][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_47[1] = layer0[47][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_47[2] = layer0[47][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_47[3] = layer0[47][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_47[4] = layer0[47][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_47[5] = layer0[47][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_47[6] = layer0[47][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_47[7] = layer1[47][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_47[8] = layer1[47][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_47[9] = layer1[47][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_47[10] = layer1[47][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_47[11] = layer1[47][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_47[12] = layer1[47][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_47[13] = layer1[47][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_47[14] = layer2[47][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_47[15] = layer2[47][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_47[16] = layer2[47][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_47[17] = layer2[47][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_47[18] = layer2[47][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_47[19] = layer2[47][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_47[20] = layer2[47][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_47[21] = layer3[47][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_47[22] = layer3[47][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_47[23] = layer3[47][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_47[24] = layer3[47][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_47[25] = layer3[47][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_47[26] = layer3[47][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_47[27] = layer3[47][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_47[28] = layer4[47][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_47[29] = layer4[47][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_47[30] = layer4[47][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_47[31] = layer4[47][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_47[32] = layer4[47][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_47[33] = layer4[47][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_47[34] = layer4[47][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_47[35] = layer5[47][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_47[36] = layer5[47][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_47[37] = layer5[47][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_47[38] = layer5[47][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_47[39] = layer5[47][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_47[40] = layer5[47][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_47[41] = layer5[47][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_47[42] = layer6[47][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_47[43] = layer6[47][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_47[44] = layer6[47][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_47[45] = layer6[47][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_47[46] = layer6[47][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_47[47] = layer6[47][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_47[48] = layer6[47][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_47 = kernel_img_mul_47[0] + kernel_img_mul_47[1] + kernel_img_mul_47[2] + 
                kernel_img_mul_47[3] + kernel_img_mul_47[4] + kernel_img_mul_47[5] + 
                kernel_img_mul_47[6] + kernel_img_mul_47[7] + kernel_img_mul_47[8] + 
                kernel_img_mul_47[9] + kernel_img_mul_47[10] + kernel_img_mul_47[11] + 
                kernel_img_mul_47[12] + kernel_img_mul_47[13] + kernel_img_mul_47[14] + 
                kernel_img_mul_47[15] + kernel_img_mul_47[16] + kernel_img_mul_47[17] + 
                kernel_img_mul_47[18] + kernel_img_mul_47[19] + kernel_img_mul_47[20] + 
                kernel_img_mul_47[21] + kernel_img_mul_47[22] + kernel_img_mul_47[23] + 
                kernel_img_mul_47[24] + kernel_img_mul_47[25] + kernel_img_mul_47[26] + 
                kernel_img_mul_47[27] + kernel_img_mul_47[28] + kernel_img_mul_47[29] + 
                kernel_img_mul_47[30] + kernel_img_mul_47[31] + kernel_img_mul_47[32] + 
                kernel_img_mul_47[33] + kernel_img_mul_47[34] + kernel_img_mul_47[35] + 
                kernel_img_mul_47[36] + kernel_img_mul_47[37] + kernel_img_mul_47[38] + 
                kernel_img_mul_47[39] + kernel_img_mul_47[40] + kernel_img_mul_47[41] + 
                kernel_img_mul_47[42] + kernel_img_mul_47[43] + kernel_img_mul_47[44] + 
                kernel_img_mul_47[45] + kernel_img_mul_47[46] + kernel_img_mul_47[47] + 
                kernel_img_mul_47[48];
wire  [39:0]  kernel_img_mul_48[0:48];
assign kernel_img_mul_48[0] = layer0[48][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_48[1] = layer0[48][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_48[2] = layer0[48][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_48[3] = layer0[48][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_48[4] = layer0[48][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_48[5] = layer0[48][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_48[6] = layer0[48][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_48[7] = layer1[48][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_48[8] = layer1[48][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_48[9] = layer1[48][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_48[10] = layer1[48][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_48[11] = layer1[48][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_48[12] = layer1[48][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_48[13] = layer1[48][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_48[14] = layer2[48][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_48[15] = layer2[48][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_48[16] = layer2[48][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_48[17] = layer2[48][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_48[18] = layer2[48][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_48[19] = layer2[48][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_48[20] = layer2[48][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_48[21] = layer3[48][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_48[22] = layer3[48][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_48[23] = layer3[48][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_48[24] = layer3[48][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_48[25] = layer3[48][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_48[26] = layer3[48][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_48[27] = layer3[48][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_48[28] = layer4[48][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_48[29] = layer4[48][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_48[30] = layer4[48][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_48[31] = layer4[48][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_48[32] = layer4[48][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_48[33] = layer4[48][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_48[34] = layer4[48][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_48[35] = layer5[48][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_48[36] = layer5[48][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_48[37] = layer5[48][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_48[38] = layer5[48][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_48[39] = layer5[48][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_48[40] = layer5[48][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_48[41] = layer5[48][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_48[42] = layer6[48][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_48[43] = layer6[48][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_48[44] = layer6[48][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_48[45] = layer6[48][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_48[46] = layer6[48][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_48[47] = layer6[48][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_48[48] = layer6[48][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_48 = kernel_img_mul_48[0] + kernel_img_mul_48[1] + kernel_img_mul_48[2] + 
                kernel_img_mul_48[3] + kernel_img_mul_48[4] + kernel_img_mul_48[5] + 
                kernel_img_mul_48[6] + kernel_img_mul_48[7] + kernel_img_mul_48[8] + 
                kernel_img_mul_48[9] + kernel_img_mul_48[10] + kernel_img_mul_48[11] + 
                kernel_img_mul_48[12] + kernel_img_mul_48[13] + kernel_img_mul_48[14] + 
                kernel_img_mul_48[15] + kernel_img_mul_48[16] + kernel_img_mul_48[17] + 
                kernel_img_mul_48[18] + kernel_img_mul_48[19] + kernel_img_mul_48[20] + 
                kernel_img_mul_48[21] + kernel_img_mul_48[22] + kernel_img_mul_48[23] + 
                kernel_img_mul_48[24] + kernel_img_mul_48[25] + kernel_img_mul_48[26] + 
                kernel_img_mul_48[27] + kernel_img_mul_48[28] + kernel_img_mul_48[29] + 
                kernel_img_mul_48[30] + kernel_img_mul_48[31] + kernel_img_mul_48[32] + 
                kernel_img_mul_48[33] + kernel_img_mul_48[34] + kernel_img_mul_48[35] + 
                kernel_img_mul_48[36] + kernel_img_mul_48[37] + kernel_img_mul_48[38] + 
                kernel_img_mul_48[39] + kernel_img_mul_48[40] + kernel_img_mul_48[41] + 
                kernel_img_mul_48[42] + kernel_img_mul_48[43] + kernel_img_mul_48[44] + 
                kernel_img_mul_48[45] + kernel_img_mul_48[46] + kernel_img_mul_48[47] + 
                kernel_img_mul_48[48];
wire  [39:0]  kernel_img_mul_49[0:48];
assign kernel_img_mul_49[0] = layer0[49][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_49[1] = layer0[49][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_49[2] = layer0[49][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_49[3] = layer0[49][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_49[4] = layer0[49][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_49[5] = layer0[49][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_49[6] = layer0[49][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_49[7] = layer1[49][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_49[8] = layer1[49][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_49[9] = layer1[49][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_49[10] = layer1[49][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_49[11] = layer1[49][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_49[12] = layer1[49][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_49[13] = layer1[49][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_49[14] = layer2[49][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_49[15] = layer2[49][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_49[16] = layer2[49][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_49[17] = layer2[49][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_49[18] = layer2[49][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_49[19] = layer2[49][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_49[20] = layer2[49][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_49[21] = layer3[49][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_49[22] = layer3[49][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_49[23] = layer3[49][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_49[24] = layer3[49][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_49[25] = layer3[49][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_49[26] = layer3[49][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_49[27] = layer3[49][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_49[28] = layer4[49][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_49[29] = layer4[49][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_49[30] = layer4[49][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_49[31] = layer4[49][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_49[32] = layer4[49][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_49[33] = layer4[49][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_49[34] = layer4[49][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_49[35] = layer5[49][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_49[36] = layer5[49][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_49[37] = layer5[49][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_49[38] = layer5[49][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_49[39] = layer5[49][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_49[40] = layer5[49][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_49[41] = layer5[49][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_49[42] = layer6[49][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_49[43] = layer6[49][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_49[44] = layer6[49][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_49[45] = layer6[49][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_49[46] = layer6[49][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_49[47] = layer6[49][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_49[48] = layer6[49][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_49 = kernel_img_mul_49[0] + kernel_img_mul_49[1] + kernel_img_mul_49[2] + 
                kernel_img_mul_49[3] + kernel_img_mul_49[4] + kernel_img_mul_49[5] + 
                kernel_img_mul_49[6] + kernel_img_mul_49[7] + kernel_img_mul_49[8] + 
                kernel_img_mul_49[9] + kernel_img_mul_49[10] + kernel_img_mul_49[11] + 
                kernel_img_mul_49[12] + kernel_img_mul_49[13] + kernel_img_mul_49[14] + 
                kernel_img_mul_49[15] + kernel_img_mul_49[16] + kernel_img_mul_49[17] + 
                kernel_img_mul_49[18] + kernel_img_mul_49[19] + kernel_img_mul_49[20] + 
                kernel_img_mul_49[21] + kernel_img_mul_49[22] + kernel_img_mul_49[23] + 
                kernel_img_mul_49[24] + kernel_img_mul_49[25] + kernel_img_mul_49[26] + 
                kernel_img_mul_49[27] + kernel_img_mul_49[28] + kernel_img_mul_49[29] + 
                kernel_img_mul_49[30] + kernel_img_mul_49[31] + kernel_img_mul_49[32] + 
                kernel_img_mul_49[33] + kernel_img_mul_49[34] + kernel_img_mul_49[35] + 
                kernel_img_mul_49[36] + kernel_img_mul_49[37] + kernel_img_mul_49[38] + 
                kernel_img_mul_49[39] + kernel_img_mul_49[40] + kernel_img_mul_49[41] + 
                kernel_img_mul_49[42] + kernel_img_mul_49[43] + kernel_img_mul_49[44] + 
                kernel_img_mul_49[45] + kernel_img_mul_49[46] + kernel_img_mul_49[47] + 
                kernel_img_mul_49[48];
wire  [39:0]  kernel_img_mul_50[0:48];
assign kernel_img_mul_50[0] = layer0[50][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_50[1] = layer0[50][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_50[2] = layer0[50][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_50[3] = layer0[50][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_50[4] = layer0[50][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_50[5] = layer0[50][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_50[6] = layer0[50][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_50[7] = layer1[50][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_50[8] = layer1[50][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_50[9] = layer1[50][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_50[10] = layer1[50][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_50[11] = layer1[50][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_50[12] = layer1[50][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_50[13] = layer1[50][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_50[14] = layer2[50][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_50[15] = layer2[50][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_50[16] = layer2[50][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_50[17] = layer2[50][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_50[18] = layer2[50][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_50[19] = layer2[50][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_50[20] = layer2[50][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_50[21] = layer3[50][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_50[22] = layer3[50][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_50[23] = layer3[50][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_50[24] = layer3[50][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_50[25] = layer3[50][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_50[26] = layer3[50][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_50[27] = layer3[50][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_50[28] = layer4[50][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_50[29] = layer4[50][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_50[30] = layer4[50][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_50[31] = layer4[50][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_50[32] = layer4[50][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_50[33] = layer4[50][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_50[34] = layer4[50][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_50[35] = layer5[50][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_50[36] = layer5[50][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_50[37] = layer5[50][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_50[38] = layer5[50][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_50[39] = layer5[50][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_50[40] = layer5[50][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_50[41] = layer5[50][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_50[42] = layer6[50][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_50[43] = layer6[50][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_50[44] = layer6[50][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_50[45] = layer6[50][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_50[46] = layer6[50][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_50[47] = layer6[50][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_50[48] = layer6[50][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_50 = kernel_img_mul_50[0] + kernel_img_mul_50[1] + kernel_img_mul_50[2] + 
                kernel_img_mul_50[3] + kernel_img_mul_50[4] + kernel_img_mul_50[5] + 
                kernel_img_mul_50[6] + kernel_img_mul_50[7] + kernel_img_mul_50[8] + 
                kernel_img_mul_50[9] + kernel_img_mul_50[10] + kernel_img_mul_50[11] + 
                kernel_img_mul_50[12] + kernel_img_mul_50[13] + kernel_img_mul_50[14] + 
                kernel_img_mul_50[15] + kernel_img_mul_50[16] + kernel_img_mul_50[17] + 
                kernel_img_mul_50[18] + kernel_img_mul_50[19] + kernel_img_mul_50[20] + 
                kernel_img_mul_50[21] + kernel_img_mul_50[22] + kernel_img_mul_50[23] + 
                kernel_img_mul_50[24] + kernel_img_mul_50[25] + kernel_img_mul_50[26] + 
                kernel_img_mul_50[27] + kernel_img_mul_50[28] + kernel_img_mul_50[29] + 
                kernel_img_mul_50[30] + kernel_img_mul_50[31] + kernel_img_mul_50[32] + 
                kernel_img_mul_50[33] + kernel_img_mul_50[34] + kernel_img_mul_50[35] + 
                kernel_img_mul_50[36] + kernel_img_mul_50[37] + kernel_img_mul_50[38] + 
                kernel_img_mul_50[39] + kernel_img_mul_50[40] + kernel_img_mul_50[41] + 
                kernel_img_mul_50[42] + kernel_img_mul_50[43] + kernel_img_mul_50[44] + 
                kernel_img_mul_50[45] + kernel_img_mul_50[46] + kernel_img_mul_50[47] + 
                kernel_img_mul_50[48];
wire  [39:0]  kernel_img_mul_51[0:48];
assign kernel_img_mul_51[0] = layer0[51][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_51[1] = layer0[51][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_51[2] = layer0[51][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_51[3] = layer0[51][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_51[4] = layer0[51][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_51[5] = layer0[51][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_51[6] = layer0[51][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_51[7] = layer1[51][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_51[8] = layer1[51][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_51[9] = layer1[51][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_51[10] = layer1[51][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_51[11] = layer1[51][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_51[12] = layer1[51][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_51[13] = layer1[51][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_51[14] = layer2[51][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_51[15] = layer2[51][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_51[16] = layer2[51][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_51[17] = layer2[51][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_51[18] = layer2[51][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_51[19] = layer2[51][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_51[20] = layer2[51][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_51[21] = layer3[51][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_51[22] = layer3[51][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_51[23] = layer3[51][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_51[24] = layer3[51][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_51[25] = layer3[51][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_51[26] = layer3[51][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_51[27] = layer3[51][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_51[28] = layer4[51][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_51[29] = layer4[51][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_51[30] = layer4[51][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_51[31] = layer4[51][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_51[32] = layer4[51][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_51[33] = layer4[51][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_51[34] = layer4[51][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_51[35] = layer5[51][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_51[36] = layer5[51][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_51[37] = layer5[51][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_51[38] = layer5[51][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_51[39] = layer5[51][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_51[40] = layer5[51][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_51[41] = layer5[51][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_51[42] = layer6[51][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_51[43] = layer6[51][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_51[44] = layer6[51][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_51[45] = layer6[51][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_51[46] = layer6[51][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_51[47] = layer6[51][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_51[48] = layer6[51][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_51 = kernel_img_mul_51[0] + kernel_img_mul_51[1] + kernel_img_mul_51[2] + 
                kernel_img_mul_51[3] + kernel_img_mul_51[4] + kernel_img_mul_51[5] + 
                kernel_img_mul_51[6] + kernel_img_mul_51[7] + kernel_img_mul_51[8] + 
                kernel_img_mul_51[9] + kernel_img_mul_51[10] + kernel_img_mul_51[11] + 
                kernel_img_mul_51[12] + kernel_img_mul_51[13] + kernel_img_mul_51[14] + 
                kernel_img_mul_51[15] + kernel_img_mul_51[16] + kernel_img_mul_51[17] + 
                kernel_img_mul_51[18] + kernel_img_mul_51[19] + kernel_img_mul_51[20] + 
                kernel_img_mul_51[21] + kernel_img_mul_51[22] + kernel_img_mul_51[23] + 
                kernel_img_mul_51[24] + kernel_img_mul_51[25] + kernel_img_mul_51[26] + 
                kernel_img_mul_51[27] + kernel_img_mul_51[28] + kernel_img_mul_51[29] + 
                kernel_img_mul_51[30] + kernel_img_mul_51[31] + kernel_img_mul_51[32] + 
                kernel_img_mul_51[33] + kernel_img_mul_51[34] + kernel_img_mul_51[35] + 
                kernel_img_mul_51[36] + kernel_img_mul_51[37] + kernel_img_mul_51[38] + 
                kernel_img_mul_51[39] + kernel_img_mul_51[40] + kernel_img_mul_51[41] + 
                kernel_img_mul_51[42] + kernel_img_mul_51[43] + kernel_img_mul_51[44] + 
                kernel_img_mul_51[45] + kernel_img_mul_51[46] + kernel_img_mul_51[47] + 
                kernel_img_mul_51[48];
wire  [39:0]  kernel_img_mul_52[0:48];
assign kernel_img_mul_52[0] = layer0[52][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_52[1] = layer0[52][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_52[2] = layer0[52][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_52[3] = layer0[52][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_52[4] = layer0[52][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_52[5] = layer0[52][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_52[6] = layer0[52][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_52[7] = layer1[52][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_52[8] = layer1[52][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_52[9] = layer1[52][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_52[10] = layer1[52][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_52[11] = layer1[52][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_52[12] = layer1[52][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_52[13] = layer1[52][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_52[14] = layer2[52][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_52[15] = layer2[52][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_52[16] = layer2[52][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_52[17] = layer2[52][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_52[18] = layer2[52][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_52[19] = layer2[52][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_52[20] = layer2[52][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_52[21] = layer3[52][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_52[22] = layer3[52][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_52[23] = layer3[52][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_52[24] = layer3[52][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_52[25] = layer3[52][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_52[26] = layer3[52][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_52[27] = layer3[52][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_52[28] = layer4[52][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_52[29] = layer4[52][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_52[30] = layer4[52][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_52[31] = layer4[52][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_52[32] = layer4[52][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_52[33] = layer4[52][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_52[34] = layer4[52][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_52[35] = layer5[52][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_52[36] = layer5[52][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_52[37] = layer5[52][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_52[38] = layer5[52][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_52[39] = layer5[52][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_52[40] = layer5[52][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_52[41] = layer5[52][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_52[42] = layer6[52][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_52[43] = layer6[52][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_52[44] = layer6[52][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_52[45] = layer6[52][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_52[46] = layer6[52][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_52[47] = layer6[52][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_52[48] = layer6[52][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_52 = kernel_img_mul_52[0] + kernel_img_mul_52[1] + kernel_img_mul_52[2] + 
                kernel_img_mul_52[3] + kernel_img_mul_52[4] + kernel_img_mul_52[5] + 
                kernel_img_mul_52[6] + kernel_img_mul_52[7] + kernel_img_mul_52[8] + 
                kernel_img_mul_52[9] + kernel_img_mul_52[10] + kernel_img_mul_52[11] + 
                kernel_img_mul_52[12] + kernel_img_mul_52[13] + kernel_img_mul_52[14] + 
                kernel_img_mul_52[15] + kernel_img_mul_52[16] + kernel_img_mul_52[17] + 
                kernel_img_mul_52[18] + kernel_img_mul_52[19] + kernel_img_mul_52[20] + 
                kernel_img_mul_52[21] + kernel_img_mul_52[22] + kernel_img_mul_52[23] + 
                kernel_img_mul_52[24] + kernel_img_mul_52[25] + kernel_img_mul_52[26] + 
                kernel_img_mul_52[27] + kernel_img_mul_52[28] + kernel_img_mul_52[29] + 
                kernel_img_mul_52[30] + kernel_img_mul_52[31] + kernel_img_mul_52[32] + 
                kernel_img_mul_52[33] + kernel_img_mul_52[34] + kernel_img_mul_52[35] + 
                kernel_img_mul_52[36] + kernel_img_mul_52[37] + kernel_img_mul_52[38] + 
                kernel_img_mul_52[39] + kernel_img_mul_52[40] + kernel_img_mul_52[41] + 
                kernel_img_mul_52[42] + kernel_img_mul_52[43] + kernel_img_mul_52[44] + 
                kernel_img_mul_52[45] + kernel_img_mul_52[46] + kernel_img_mul_52[47] + 
                kernel_img_mul_52[48];
wire  [39:0]  kernel_img_mul_53[0:48];
assign kernel_img_mul_53[0] = layer0[53][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_53[1] = layer0[53][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_53[2] = layer0[53][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_53[3] = layer0[53][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_53[4] = layer0[53][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_53[5] = layer0[53][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_53[6] = layer0[53][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_53[7] = layer1[53][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_53[8] = layer1[53][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_53[9] = layer1[53][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_53[10] = layer1[53][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_53[11] = layer1[53][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_53[12] = layer1[53][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_53[13] = layer1[53][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_53[14] = layer2[53][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_53[15] = layer2[53][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_53[16] = layer2[53][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_53[17] = layer2[53][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_53[18] = layer2[53][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_53[19] = layer2[53][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_53[20] = layer2[53][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_53[21] = layer3[53][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_53[22] = layer3[53][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_53[23] = layer3[53][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_53[24] = layer3[53][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_53[25] = layer3[53][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_53[26] = layer3[53][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_53[27] = layer3[53][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_53[28] = layer4[53][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_53[29] = layer4[53][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_53[30] = layer4[53][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_53[31] = layer4[53][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_53[32] = layer4[53][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_53[33] = layer4[53][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_53[34] = layer4[53][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_53[35] = layer5[53][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_53[36] = layer5[53][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_53[37] = layer5[53][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_53[38] = layer5[53][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_53[39] = layer5[53][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_53[40] = layer5[53][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_53[41] = layer5[53][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_53[42] = layer6[53][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_53[43] = layer6[53][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_53[44] = layer6[53][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_53[45] = layer6[53][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_53[46] = layer6[53][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_53[47] = layer6[53][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_53[48] = layer6[53][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_53 = kernel_img_mul_53[0] + kernel_img_mul_53[1] + kernel_img_mul_53[2] + 
                kernel_img_mul_53[3] + kernel_img_mul_53[4] + kernel_img_mul_53[5] + 
                kernel_img_mul_53[6] + kernel_img_mul_53[7] + kernel_img_mul_53[8] + 
                kernel_img_mul_53[9] + kernel_img_mul_53[10] + kernel_img_mul_53[11] + 
                kernel_img_mul_53[12] + kernel_img_mul_53[13] + kernel_img_mul_53[14] + 
                kernel_img_mul_53[15] + kernel_img_mul_53[16] + kernel_img_mul_53[17] + 
                kernel_img_mul_53[18] + kernel_img_mul_53[19] + kernel_img_mul_53[20] + 
                kernel_img_mul_53[21] + kernel_img_mul_53[22] + kernel_img_mul_53[23] + 
                kernel_img_mul_53[24] + kernel_img_mul_53[25] + kernel_img_mul_53[26] + 
                kernel_img_mul_53[27] + kernel_img_mul_53[28] + kernel_img_mul_53[29] + 
                kernel_img_mul_53[30] + kernel_img_mul_53[31] + kernel_img_mul_53[32] + 
                kernel_img_mul_53[33] + kernel_img_mul_53[34] + kernel_img_mul_53[35] + 
                kernel_img_mul_53[36] + kernel_img_mul_53[37] + kernel_img_mul_53[38] + 
                kernel_img_mul_53[39] + kernel_img_mul_53[40] + kernel_img_mul_53[41] + 
                kernel_img_mul_53[42] + kernel_img_mul_53[43] + kernel_img_mul_53[44] + 
                kernel_img_mul_53[45] + kernel_img_mul_53[46] + kernel_img_mul_53[47] + 
                kernel_img_mul_53[48];
wire  [39:0]  kernel_img_mul_54[0:48];
assign kernel_img_mul_54[0] = layer0[54][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_54[1] = layer0[54][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_54[2] = layer0[54][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_54[3] = layer0[54][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_54[4] = layer0[54][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_54[5] = layer0[54][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_54[6] = layer0[54][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_54[7] = layer1[54][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_54[8] = layer1[54][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_54[9] = layer1[54][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_54[10] = layer1[54][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_54[11] = layer1[54][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_54[12] = layer1[54][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_54[13] = layer1[54][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_54[14] = layer2[54][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_54[15] = layer2[54][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_54[16] = layer2[54][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_54[17] = layer2[54][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_54[18] = layer2[54][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_54[19] = layer2[54][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_54[20] = layer2[54][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_54[21] = layer3[54][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_54[22] = layer3[54][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_54[23] = layer3[54][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_54[24] = layer3[54][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_54[25] = layer3[54][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_54[26] = layer3[54][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_54[27] = layer3[54][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_54[28] = layer4[54][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_54[29] = layer4[54][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_54[30] = layer4[54][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_54[31] = layer4[54][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_54[32] = layer4[54][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_54[33] = layer4[54][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_54[34] = layer4[54][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_54[35] = layer5[54][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_54[36] = layer5[54][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_54[37] = layer5[54][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_54[38] = layer5[54][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_54[39] = layer5[54][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_54[40] = layer5[54][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_54[41] = layer5[54][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_54[42] = layer6[54][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_54[43] = layer6[54][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_54[44] = layer6[54][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_54[45] = layer6[54][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_54[46] = layer6[54][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_54[47] = layer6[54][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_54[48] = layer6[54][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_54 = kernel_img_mul_54[0] + kernel_img_mul_54[1] + kernel_img_mul_54[2] + 
                kernel_img_mul_54[3] + kernel_img_mul_54[4] + kernel_img_mul_54[5] + 
                kernel_img_mul_54[6] + kernel_img_mul_54[7] + kernel_img_mul_54[8] + 
                kernel_img_mul_54[9] + kernel_img_mul_54[10] + kernel_img_mul_54[11] + 
                kernel_img_mul_54[12] + kernel_img_mul_54[13] + kernel_img_mul_54[14] + 
                kernel_img_mul_54[15] + kernel_img_mul_54[16] + kernel_img_mul_54[17] + 
                kernel_img_mul_54[18] + kernel_img_mul_54[19] + kernel_img_mul_54[20] + 
                kernel_img_mul_54[21] + kernel_img_mul_54[22] + kernel_img_mul_54[23] + 
                kernel_img_mul_54[24] + kernel_img_mul_54[25] + kernel_img_mul_54[26] + 
                kernel_img_mul_54[27] + kernel_img_mul_54[28] + kernel_img_mul_54[29] + 
                kernel_img_mul_54[30] + kernel_img_mul_54[31] + kernel_img_mul_54[32] + 
                kernel_img_mul_54[33] + kernel_img_mul_54[34] + kernel_img_mul_54[35] + 
                kernel_img_mul_54[36] + kernel_img_mul_54[37] + kernel_img_mul_54[38] + 
                kernel_img_mul_54[39] + kernel_img_mul_54[40] + kernel_img_mul_54[41] + 
                kernel_img_mul_54[42] + kernel_img_mul_54[43] + kernel_img_mul_54[44] + 
                kernel_img_mul_54[45] + kernel_img_mul_54[46] + kernel_img_mul_54[47] + 
                kernel_img_mul_54[48];
wire  [39:0]  kernel_img_mul_55[0:48];
assign kernel_img_mul_55[0] = layer0[55][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_55[1] = layer0[55][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_55[2] = layer0[55][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_55[3] = layer0[55][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_55[4] = layer0[55][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_55[5] = layer0[55][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_55[6] = layer0[55][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_55[7] = layer1[55][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_55[8] = layer1[55][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_55[9] = layer1[55][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_55[10] = layer1[55][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_55[11] = layer1[55][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_55[12] = layer1[55][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_55[13] = layer1[55][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_55[14] = layer2[55][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_55[15] = layer2[55][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_55[16] = layer2[55][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_55[17] = layer2[55][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_55[18] = layer2[55][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_55[19] = layer2[55][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_55[20] = layer2[55][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_55[21] = layer3[55][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_55[22] = layer3[55][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_55[23] = layer3[55][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_55[24] = layer3[55][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_55[25] = layer3[55][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_55[26] = layer3[55][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_55[27] = layer3[55][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_55[28] = layer4[55][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_55[29] = layer4[55][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_55[30] = layer4[55][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_55[31] = layer4[55][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_55[32] = layer4[55][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_55[33] = layer4[55][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_55[34] = layer4[55][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_55[35] = layer5[55][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_55[36] = layer5[55][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_55[37] = layer5[55][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_55[38] = layer5[55][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_55[39] = layer5[55][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_55[40] = layer5[55][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_55[41] = layer5[55][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_55[42] = layer6[55][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_55[43] = layer6[55][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_55[44] = layer6[55][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_55[45] = layer6[55][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_55[46] = layer6[55][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_55[47] = layer6[55][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_55[48] = layer6[55][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_55 = kernel_img_mul_55[0] + kernel_img_mul_55[1] + kernel_img_mul_55[2] + 
                kernel_img_mul_55[3] + kernel_img_mul_55[4] + kernel_img_mul_55[5] + 
                kernel_img_mul_55[6] + kernel_img_mul_55[7] + kernel_img_mul_55[8] + 
                kernel_img_mul_55[9] + kernel_img_mul_55[10] + kernel_img_mul_55[11] + 
                kernel_img_mul_55[12] + kernel_img_mul_55[13] + kernel_img_mul_55[14] + 
                kernel_img_mul_55[15] + kernel_img_mul_55[16] + kernel_img_mul_55[17] + 
                kernel_img_mul_55[18] + kernel_img_mul_55[19] + kernel_img_mul_55[20] + 
                kernel_img_mul_55[21] + kernel_img_mul_55[22] + kernel_img_mul_55[23] + 
                kernel_img_mul_55[24] + kernel_img_mul_55[25] + kernel_img_mul_55[26] + 
                kernel_img_mul_55[27] + kernel_img_mul_55[28] + kernel_img_mul_55[29] + 
                kernel_img_mul_55[30] + kernel_img_mul_55[31] + kernel_img_mul_55[32] + 
                kernel_img_mul_55[33] + kernel_img_mul_55[34] + kernel_img_mul_55[35] + 
                kernel_img_mul_55[36] + kernel_img_mul_55[37] + kernel_img_mul_55[38] + 
                kernel_img_mul_55[39] + kernel_img_mul_55[40] + kernel_img_mul_55[41] + 
                kernel_img_mul_55[42] + kernel_img_mul_55[43] + kernel_img_mul_55[44] + 
                kernel_img_mul_55[45] + kernel_img_mul_55[46] + kernel_img_mul_55[47] + 
                kernel_img_mul_55[48];
wire  [39:0]  kernel_img_mul_56[0:48];
assign kernel_img_mul_56[0] = layer0[56][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_56[1] = layer0[56][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_56[2] = layer0[56][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_56[3] = layer0[56][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_56[4] = layer0[56][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_56[5] = layer0[56][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_56[6] = layer0[56][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_56[7] = layer1[56][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_56[8] = layer1[56][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_56[9] = layer1[56][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_56[10] = layer1[56][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_56[11] = layer1[56][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_56[12] = layer1[56][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_56[13] = layer1[56][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_56[14] = layer2[56][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_56[15] = layer2[56][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_56[16] = layer2[56][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_56[17] = layer2[56][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_56[18] = layer2[56][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_56[19] = layer2[56][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_56[20] = layer2[56][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_56[21] = layer3[56][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_56[22] = layer3[56][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_56[23] = layer3[56][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_56[24] = layer3[56][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_56[25] = layer3[56][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_56[26] = layer3[56][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_56[27] = layer3[56][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_56[28] = layer4[56][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_56[29] = layer4[56][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_56[30] = layer4[56][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_56[31] = layer4[56][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_56[32] = layer4[56][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_56[33] = layer4[56][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_56[34] = layer4[56][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_56[35] = layer5[56][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_56[36] = layer5[56][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_56[37] = layer5[56][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_56[38] = layer5[56][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_56[39] = layer5[56][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_56[40] = layer5[56][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_56[41] = layer5[56][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_56[42] = layer6[56][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_56[43] = layer6[56][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_56[44] = layer6[56][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_56[45] = layer6[56][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_56[46] = layer6[56][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_56[47] = layer6[56][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_56[48] = layer6[56][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_56 = kernel_img_mul_56[0] + kernel_img_mul_56[1] + kernel_img_mul_56[2] + 
                kernel_img_mul_56[3] + kernel_img_mul_56[4] + kernel_img_mul_56[5] + 
                kernel_img_mul_56[6] + kernel_img_mul_56[7] + kernel_img_mul_56[8] + 
                kernel_img_mul_56[9] + kernel_img_mul_56[10] + kernel_img_mul_56[11] + 
                kernel_img_mul_56[12] + kernel_img_mul_56[13] + kernel_img_mul_56[14] + 
                kernel_img_mul_56[15] + kernel_img_mul_56[16] + kernel_img_mul_56[17] + 
                kernel_img_mul_56[18] + kernel_img_mul_56[19] + kernel_img_mul_56[20] + 
                kernel_img_mul_56[21] + kernel_img_mul_56[22] + kernel_img_mul_56[23] + 
                kernel_img_mul_56[24] + kernel_img_mul_56[25] + kernel_img_mul_56[26] + 
                kernel_img_mul_56[27] + kernel_img_mul_56[28] + kernel_img_mul_56[29] + 
                kernel_img_mul_56[30] + kernel_img_mul_56[31] + kernel_img_mul_56[32] + 
                kernel_img_mul_56[33] + kernel_img_mul_56[34] + kernel_img_mul_56[35] + 
                kernel_img_mul_56[36] + kernel_img_mul_56[37] + kernel_img_mul_56[38] + 
                kernel_img_mul_56[39] + kernel_img_mul_56[40] + kernel_img_mul_56[41] + 
                kernel_img_mul_56[42] + kernel_img_mul_56[43] + kernel_img_mul_56[44] + 
                kernel_img_mul_56[45] + kernel_img_mul_56[46] + kernel_img_mul_56[47] + 
                kernel_img_mul_56[48];
wire  [39:0]  kernel_img_mul_57[0:48];
assign kernel_img_mul_57[0] = layer0[57][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_57[1] = layer0[57][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_57[2] = layer0[57][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_57[3] = layer0[57][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_57[4] = layer0[57][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_57[5] = layer0[57][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_57[6] = layer0[57][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_57[7] = layer1[57][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_57[8] = layer1[57][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_57[9] = layer1[57][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_57[10] = layer1[57][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_57[11] = layer1[57][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_57[12] = layer1[57][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_57[13] = layer1[57][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_57[14] = layer2[57][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_57[15] = layer2[57][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_57[16] = layer2[57][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_57[17] = layer2[57][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_57[18] = layer2[57][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_57[19] = layer2[57][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_57[20] = layer2[57][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_57[21] = layer3[57][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_57[22] = layer3[57][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_57[23] = layer3[57][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_57[24] = layer3[57][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_57[25] = layer3[57][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_57[26] = layer3[57][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_57[27] = layer3[57][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_57[28] = layer4[57][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_57[29] = layer4[57][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_57[30] = layer4[57][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_57[31] = layer4[57][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_57[32] = layer4[57][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_57[33] = layer4[57][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_57[34] = layer4[57][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_57[35] = layer5[57][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_57[36] = layer5[57][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_57[37] = layer5[57][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_57[38] = layer5[57][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_57[39] = layer5[57][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_57[40] = layer5[57][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_57[41] = layer5[57][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_57[42] = layer6[57][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_57[43] = layer6[57][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_57[44] = layer6[57][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_57[45] = layer6[57][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_57[46] = layer6[57][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_57[47] = layer6[57][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_57[48] = layer6[57][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_57 = kernel_img_mul_57[0] + kernel_img_mul_57[1] + kernel_img_mul_57[2] + 
                kernel_img_mul_57[3] + kernel_img_mul_57[4] + kernel_img_mul_57[5] + 
                kernel_img_mul_57[6] + kernel_img_mul_57[7] + kernel_img_mul_57[8] + 
                kernel_img_mul_57[9] + kernel_img_mul_57[10] + kernel_img_mul_57[11] + 
                kernel_img_mul_57[12] + kernel_img_mul_57[13] + kernel_img_mul_57[14] + 
                kernel_img_mul_57[15] + kernel_img_mul_57[16] + kernel_img_mul_57[17] + 
                kernel_img_mul_57[18] + kernel_img_mul_57[19] + kernel_img_mul_57[20] + 
                kernel_img_mul_57[21] + kernel_img_mul_57[22] + kernel_img_mul_57[23] + 
                kernel_img_mul_57[24] + kernel_img_mul_57[25] + kernel_img_mul_57[26] + 
                kernel_img_mul_57[27] + kernel_img_mul_57[28] + kernel_img_mul_57[29] + 
                kernel_img_mul_57[30] + kernel_img_mul_57[31] + kernel_img_mul_57[32] + 
                kernel_img_mul_57[33] + kernel_img_mul_57[34] + kernel_img_mul_57[35] + 
                kernel_img_mul_57[36] + kernel_img_mul_57[37] + kernel_img_mul_57[38] + 
                kernel_img_mul_57[39] + kernel_img_mul_57[40] + kernel_img_mul_57[41] + 
                kernel_img_mul_57[42] + kernel_img_mul_57[43] + kernel_img_mul_57[44] + 
                kernel_img_mul_57[45] + kernel_img_mul_57[46] + kernel_img_mul_57[47] + 
                kernel_img_mul_57[48];
wire  [39:0]  kernel_img_mul_58[0:48];
assign kernel_img_mul_58[0] = layer0[58][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_58[1] = layer0[58][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_58[2] = layer0[58][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_58[3] = layer0[58][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_58[4] = layer0[58][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_58[5] = layer0[58][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_58[6] = layer0[58][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_58[7] = layer1[58][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_58[8] = layer1[58][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_58[9] = layer1[58][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_58[10] = layer1[58][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_58[11] = layer1[58][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_58[12] = layer1[58][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_58[13] = layer1[58][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_58[14] = layer2[58][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_58[15] = layer2[58][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_58[16] = layer2[58][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_58[17] = layer2[58][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_58[18] = layer2[58][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_58[19] = layer2[58][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_58[20] = layer2[58][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_58[21] = layer3[58][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_58[22] = layer3[58][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_58[23] = layer3[58][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_58[24] = layer3[58][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_58[25] = layer3[58][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_58[26] = layer3[58][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_58[27] = layer3[58][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_58[28] = layer4[58][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_58[29] = layer4[58][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_58[30] = layer4[58][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_58[31] = layer4[58][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_58[32] = layer4[58][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_58[33] = layer4[58][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_58[34] = layer4[58][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_58[35] = layer5[58][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_58[36] = layer5[58][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_58[37] = layer5[58][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_58[38] = layer5[58][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_58[39] = layer5[58][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_58[40] = layer5[58][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_58[41] = layer5[58][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_58[42] = layer6[58][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_58[43] = layer6[58][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_58[44] = layer6[58][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_58[45] = layer6[58][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_58[46] = layer6[58][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_58[47] = layer6[58][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_58[48] = layer6[58][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_58 = kernel_img_mul_58[0] + kernel_img_mul_58[1] + kernel_img_mul_58[2] + 
                kernel_img_mul_58[3] + kernel_img_mul_58[4] + kernel_img_mul_58[5] + 
                kernel_img_mul_58[6] + kernel_img_mul_58[7] + kernel_img_mul_58[8] + 
                kernel_img_mul_58[9] + kernel_img_mul_58[10] + kernel_img_mul_58[11] + 
                kernel_img_mul_58[12] + kernel_img_mul_58[13] + kernel_img_mul_58[14] + 
                kernel_img_mul_58[15] + kernel_img_mul_58[16] + kernel_img_mul_58[17] + 
                kernel_img_mul_58[18] + kernel_img_mul_58[19] + kernel_img_mul_58[20] + 
                kernel_img_mul_58[21] + kernel_img_mul_58[22] + kernel_img_mul_58[23] + 
                kernel_img_mul_58[24] + kernel_img_mul_58[25] + kernel_img_mul_58[26] + 
                kernel_img_mul_58[27] + kernel_img_mul_58[28] + kernel_img_mul_58[29] + 
                kernel_img_mul_58[30] + kernel_img_mul_58[31] + kernel_img_mul_58[32] + 
                kernel_img_mul_58[33] + kernel_img_mul_58[34] + kernel_img_mul_58[35] + 
                kernel_img_mul_58[36] + kernel_img_mul_58[37] + kernel_img_mul_58[38] + 
                kernel_img_mul_58[39] + kernel_img_mul_58[40] + kernel_img_mul_58[41] + 
                kernel_img_mul_58[42] + kernel_img_mul_58[43] + kernel_img_mul_58[44] + 
                kernel_img_mul_58[45] + kernel_img_mul_58[46] + kernel_img_mul_58[47] + 
                kernel_img_mul_58[48];
wire  [39:0]  kernel_img_mul_59[0:48];
assign kernel_img_mul_59[0] = layer0[59][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_59[1] = layer0[59][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_59[2] = layer0[59][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_59[3] = layer0[59][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_59[4] = layer0[59][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_59[5] = layer0[59][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_59[6] = layer0[59][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_59[7] = layer1[59][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_59[8] = layer1[59][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_59[9] = layer1[59][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_59[10] = layer1[59][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_59[11] = layer1[59][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_59[12] = layer1[59][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_59[13] = layer1[59][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_59[14] = layer2[59][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_59[15] = layer2[59][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_59[16] = layer2[59][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_59[17] = layer2[59][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_59[18] = layer2[59][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_59[19] = layer2[59][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_59[20] = layer2[59][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_59[21] = layer3[59][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_59[22] = layer3[59][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_59[23] = layer3[59][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_59[24] = layer3[59][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_59[25] = layer3[59][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_59[26] = layer3[59][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_59[27] = layer3[59][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_59[28] = layer4[59][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_59[29] = layer4[59][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_59[30] = layer4[59][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_59[31] = layer4[59][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_59[32] = layer4[59][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_59[33] = layer4[59][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_59[34] = layer4[59][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_59[35] = layer5[59][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_59[36] = layer5[59][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_59[37] = layer5[59][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_59[38] = layer5[59][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_59[39] = layer5[59][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_59[40] = layer5[59][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_59[41] = layer5[59][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_59[42] = layer6[59][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_59[43] = layer6[59][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_59[44] = layer6[59][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_59[45] = layer6[59][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_59[46] = layer6[59][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_59[47] = layer6[59][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_59[48] = layer6[59][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_59 = kernel_img_mul_59[0] + kernel_img_mul_59[1] + kernel_img_mul_59[2] + 
                kernel_img_mul_59[3] + kernel_img_mul_59[4] + kernel_img_mul_59[5] + 
                kernel_img_mul_59[6] + kernel_img_mul_59[7] + kernel_img_mul_59[8] + 
                kernel_img_mul_59[9] + kernel_img_mul_59[10] + kernel_img_mul_59[11] + 
                kernel_img_mul_59[12] + kernel_img_mul_59[13] + kernel_img_mul_59[14] + 
                kernel_img_mul_59[15] + kernel_img_mul_59[16] + kernel_img_mul_59[17] + 
                kernel_img_mul_59[18] + kernel_img_mul_59[19] + kernel_img_mul_59[20] + 
                kernel_img_mul_59[21] + kernel_img_mul_59[22] + kernel_img_mul_59[23] + 
                kernel_img_mul_59[24] + kernel_img_mul_59[25] + kernel_img_mul_59[26] + 
                kernel_img_mul_59[27] + kernel_img_mul_59[28] + kernel_img_mul_59[29] + 
                kernel_img_mul_59[30] + kernel_img_mul_59[31] + kernel_img_mul_59[32] + 
                kernel_img_mul_59[33] + kernel_img_mul_59[34] + kernel_img_mul_59[35] + 
                kernel_img_mul_59[36] + kernel_img_mul_59[37] + kernel_img_mul_59[38] + 
                kernel_img_mul_59[39] + kernel_img_mul_59[40] + kernel_img_mul_59[41] + 
                kernel_img_mul_59[42] + kernel_img_mul_59[43] + kernel_img_mul_59[44] + 
                kernel_img_mul_59[45] + kernel_img_mul_59[46] + kernel_img_mul_59[47] + 
                kernel_img_mul_59[48];
wire  [39:0]  kernel_img_mul_60[0:48];
assign kernel_img_mul_60[0] = layer0[60][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_60[1] = layer0[60][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_60[2] = layer0[60][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_60[3] = layer0[60][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_60[4] = layer0[60][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_60[5] = layer0[60][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_60[6] = layer0[60][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_60[7] = layer1[60][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_60[8] = layer1[60][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_60[9] = layer1[60][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_60[10] = layer1[60][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_60[11] = layer1[60][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_60[12] = layer1[60][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_60[13] = layer1[60][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_60[14] = layer2[60][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_60[15] = layer2[60][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_60[16] = layer2[60][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_60[17] = layer2[60][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_60[18] = layer2[60][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_60[19] = layer2[60][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_60[20] = layer2[60][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_60[21] = layer3[60][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_60[22] = layer3[60][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_60[23] = layer3[60][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_60[24] = layer3[60][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_60[25] = layer3[60][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_60[26] = layer3[60][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_60[27] = layer3[60][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_60[28] = layer4[60][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_60[29] = layer4[60][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_60[30] = layer4[60][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_60[31] = layer4[60][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_60[32] = layer4[60][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_60[33] = layer4[60][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_60[34] = layer4[60][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_60[35] = layer5[60][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_60[36] = layer5[60][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_60[37] = layer5[60][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_60[38] = layer5[60][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_60[39] = layer5[60][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_60[40] = layer5[60][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_60[41] = layer5[60][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_60[42] = layer6[60][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_60[43] = layer6[60][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_60[44] = layer6[60][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_60[45] = layer6[60][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_60[46] = layer6[60][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_60[47] = layer6[60][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_60[48] = layer6[60][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_60 = kernel_img_mul_60[0] + kernel_img_mul_60[1] + kernel_img_mul_60[2] + 
                kernel_img_mul_60[3] + kernel_img_mul_60[4] + kernel_img_mul_60[5] + 
                kernel_img_mul_60[6] + kernel_img_mul_60[7] + kernel_img_mul_60[8] + 
                kernel_img_mul_60[9] + kernel_img_mul_60[10] + kernel_img_mul_60[11] + 
                kernel_img_mul_60[12] + kernel_img_mul_60[13] + kernel_img_mul_60[14] + 
                kernel_img_mul_60[15] + kernel_img_mul_60[16] + kernel_img_mul_60[17] + 
                kernel_img_mul_60[18] + kernel_img_mul_60[19] + kernel_img_mul_60[20] + 
                kernel_img_mul_60[21] + kernel_img_mul_60[22] + kernel_img_mul_60[23] + 
                kernel_img_mul_60[24] + kernel_img_mul_60[25] + kernel_img_mul_60[26] + 
                kernel_img_mul_60[27] + kernel_img_mul_60[28] + kernel_img_mul_60[29] + 
                kernel_img_mul_60[30] + kernel_img_mul_60[31] + kernel_img_mul_60[32] + 
                kernel_img_mul_60[33] + kernel_img_mul_60[34] + kernel_img_mul_60[35] + 
                kernel_img_mul_60[36] + kernel_img_mul_60[37] + kernel_img_mul_60[38] + 
                kernel_img_mul_60[39] + kernel_img_mul_60[40] + kernel_img_mul_60[41] + 
                kernel_img_mul_60[42] + kernel_img_mul_60[43] + kernel_img_mul_60[44] + 
                kernel_img_mul_60[45] + kernel_img_mul_60[46] + kernel_img_mul_60[47] + 
                kernel_img_mul_60[48];
wire  [39:0]  kernel_img_mul_61[0:48];
assign kernel_img_mul_61[0] = layer0[61][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_61[1] = layer0[61][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_61[2] = layer0[61][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_61[3] = layer0[61][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_61[4] = layer0[61][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_61[5] = layer0[61][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_61[6] = layer0[61][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_61[7] = layer1[61][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_61[8] = layer1[61][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_61[9] = layer1[61][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_61[10] = layer1[61][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_61[11] = layer1[61][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_61[12] = layer1[61][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_61[13] = layer1[61][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_61[14] = layer2[61][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_61[15] = layer2[61][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_61[16] = layer2[61][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_61[17] = layer2[61][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_61[18] = layer2[61][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_61[19] = layer2[61][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_61[20] = layer2[61][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_61[21] = layer3[61][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_61[22] = layer3[61][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_61[23] = layer3[61][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_61[24] = layer3[61][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_61[25] = layer3[61][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_61[26] = layer3[61][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_61[27] = layer3[61][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_61[28] = layer4[61][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_61[29] = layer4[61][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_61[30] = layer4[61][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_61[31] = layer4[61][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_61[32] = layer4[61][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_61[33] = layer4[61][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_61[34] = layer4[61][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_61[35] = layer5[61][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_61[36] = layer5[61][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_61[37] = layer5[61][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_61[38] = layer5[61][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_61[39] = layer5[61][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_61[40] = layer5[61][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_61[41] = layer5[61][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_61[42] = layer6[61][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_61[43] = layer6[61][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_61[44] = layer6[61][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_61[45] = layer6[61][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_61[46] = layer6[61][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_61[47] = layer6[61][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_61[48] = layer6[61][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_61 = kernel_img_mul_61[0] + kernel_img_mul_61[1] + kernel_img_mul_61[2] + 
                kernel_img_mul_61[3] + kernel_img_mul_61[4] + kernel_img_mul_61[5] + 
                kernel_img_mul_61[6] + kernel_img_mul_61[7] + kernel_img_mul_61[8] + 
                kernel_img_mul_61[9] + kernel_img_mul_61[10] + kernel_img_mul_61[11] + 
                kernel_img_mul_61[12] + kernel_img_mul_61[13] + kernel_img_mul_61[14] + 
                kernel_img_mul_61[15] + kernel_img_mul_61[16] + kernel_img_mul_61[17] + 
                kernel_img_mul_61[18] + kernel_img_mul_61[19] + kernel_img_mul_61[20] + 
                kernel_img_mul_61[21] + kernel_img_mul_61[22] + kernel_img_mul_61[23] + 
                kernel_img_mul_61[24] + kernel_img_mul_61[25] + kernel_img_mul_61[26] + 
                kernel_img_mul_61[27] + kernel_img_mul_61[28] + kernel_img_mul_61[29] + 
                kernel_img_mul_61[30] + kernel_img_mul_61[31] + kernel_img_mul_61[32] + 
                kernel_img_mul_61[33] + kernel_img_mul_61[34] + kernel_img_mul_61[35] + 
                kernel_img_mul_61[36] + kernel_img_mul_61[37] + kernel_img_mul_61[38] + 
                kernel_img_mul_61[39] + kernel_img_mul_61[40] + kernel_img_mul_61[41] + 
                kernel_img_mul_61[42] + kernel_img_mul_61[43] + kernel_img_mul_61[44] + 
                kernel_img_mul_61[45] + kernel_img_mul_61[46] + kernel_img_mul_61[47] + 
                kernel_img_mul_61[48];
wire  [39:0]  kernel_img_mul_62[0:48];
assign kernel_img_mul_62[0] = layer0[62][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_62[1] = layer0[62][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_62[2] = layer0[62][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_62[3] = layer0[62][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_62[4] = layer0[62][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_62[5] = layer0[62][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_62[6] = layer0[62][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_62[7] = layer1[62][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_62[8] = layer1[62][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_62[9] = layer1[62][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_62[10] = layer1[62][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_62[11] = layer1[62][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_62[12] = layer1[62][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_62[13] = layer1[62][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_62[14] = layer2[62][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_62[15] = layer2[62][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_62[16] = layer2[62][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_62[17] = layer2[62][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_62[18] = layer2[62][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_62[19] = layer2[62][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_62[20] = layer2[62][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_62[21] = layer3[62][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_62[22] = layer3[62][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_62[23] = layer3[62][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_62[24] = layer3[62][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_62[25] = layer3[62][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_62[26] = layer3[62][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_62[27] = layer3[62][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_62[28] = layer4[62][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_62[29] = layer4[62][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_62[30] = layer4[62][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_62[31] = layer4[62][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_62[32] = layer4[62][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_62[33] = layer4[62][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_62[34] = layer4[62][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_62[35] = layer5[62][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_62[36] = layer5[62][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_62[37] = layer5[62][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_62[38] = layer5[62][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_62[39] = layer5[62][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_62[40] = layer5[62][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_62[41] = layer5[62][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_62[42] = layer6[62][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_62[43] = layer6[62][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_62[44] = layer6[62][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_62[45] = layer6[62][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_62[46] = layer6[62][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_62[47] = layer6[62][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_62[48] = layer6[62][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_62 = kernel_img_mul_62[0] + kernel_img_mul_62[1] + kernel_img_mul_62[2] + 
                kernel_img_mul_62[3] + kernel_img_mul_62[4] + kernel_img_mul_62[5] + 
                kernel_img_mul_62[6] + kernel_img_mul_62[7] + kernel_img_mul_62[8] + 
                kernel_img_mul_62[9] + kernel_img_mul_62[10] + kernel_img_mul_62[11] + 
                kernel_img_mul_62[12] + kernel_img_mul_62[13] + kernel_img_mul_62[14] + 
                kernel_img_mul_62[15] + kernel_img_mul_62[16] + kernel_img_mul_62[17] + 
                kernel_img_mul_62[18] + kernel_img_mul_62[19] + kernel_img_mul_62[20] + 
                kernel_img_mul_62[21] + kernel_img_mul_62[22] + kernel_img_mul_62[23] + 
                kernel_img_mul_62[24] + kernel_img_mul_62[25] + kernel_img_mul_62[26] + 
                kernel_img_mul_62[27] + kernel_img_mul_62[28] + kernel_img_mul_62[29] + 
                kernel_img_mul_62[30] + kernel_img_mul_62[31] + kernel_img_mul_62[32] + 
                kernel_img_mul_62[33] + kernel_img_mul_62[34] + kernel_img_mul_62[35] + 
                kernel_img_mul_62[36] + kernel_img_mul_62[37] + kernel_img_mul_62[38] + 
                kernel_img_mul_62[39] + kernel_img_mul_62[40] + kernel_img_mul_62[41] + 
                kernel_img_mul_62[42] + kernel_img_mul_62[43] + kernel_img_mul_62[44] + 
                kernel_img_mul_62[45] + kernel_img_mul_62[46] + kernel_img_mul_62[47] + 
                kernel_img_mul_62[48];
wire  [39:0]  kernel_img_mul_63[0:48];
assign kernel_img_mul_63[0] = layer0[63][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_63[1] = layer0[63][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_63[2] = layer0[63][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_63[3] = layer0[63][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_63[4] = layer0[63][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_63[5] = layer0[63][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_63[6] = layer0[63][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_63[7] = layer1[63][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_63[8] = layer1[63][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_63[9] = layer1[63][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_63[10] = layer1[63][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_63[11] = layer1[63][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_63[12] = layer1[63][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_63[13] = layer1[63][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_63[14] = layer2[63][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_63[15] = layer2[63][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_63[16] = layer2[63][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_63[17] = layer2[63][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_63[18] = layer2[63][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_63[19] = layer2[63][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_63[20] = layer2[63][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_63[21] = layer3[63][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_63[22] = layer3[63][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_63[23] = layer3[63][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_63[24] = layer3[63][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_63[25] = layer3[63][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_63[26] = layer3[63][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_63[27] = layer3[63][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_63[28] = layer4[63][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_63[29] = layer4[63][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_63[30] = layer4[63][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_63[31] = layer4[63][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_63[32] = layer4[63][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_63[33] = layer4[63][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_63[34] = layer4[63][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_63[35] = layer5[63][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_63[36] = layer5[63][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_63[37] = layer5[63][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_63[38] = layer5[63][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_63[39] = layer5[63][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_63[40] = layer5[63][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_63[41] = layer5[63][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_63[42] = layer6[63][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_63[43] = layer6[63][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_63[44] = layer6[63][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_63[45] = layer6[63][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_63[46] = layer6[63][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_63[47] = layer6[63][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_63[48] = layer6[63][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_63 = kernel_img_mul_63[0] + kernel_img_mul_63[1] + kernel_img_mul_63[2] + 
                kernel_img_mul_63[3] + kernel_img_mul_63[4] + kernel_img_mul_63[5] + 
                kernel_img_mul_63[6] + kernel_img_mul_63[7] + kernel_img_mul_63[8] + 
                kernel_img_mul_63[9] + kernel_img_mul_63[10] + kernel_img_mul_63[11] + 
                kernel_img_mul_63[12] + kernel_img_mul_63[13] + kernel_img_mul_63[14] + 
                kernel_img_mul_63[15] + kernel_img_mul_63[16] + kernel_img_mul_63[17] + 
                kernel_img_mul_63[18] + kernel_img_mul_63[19] + kernel_img_mul_63[20] + 
                kernel_img_mul_63[21] + kernel_img_mul_63[22] + kernel_img_mul_63[23] + 
                kernel_img_mul_63[24] + kernel_img_mul_63[25] + kernel_img_mul_63[26] + 
                kernel_img_mul_63[27] + kernel_img_mul_63[28] + kernel_img_mul_63[29] + 
                kernel_img_mul_63[30] + kernel_img_mul_63[31] + kernel_img_mul_63[32] + 
                kernel_img_mul_63[33] + kernel_img_mul_63[34] + kernel_img_mul_63[35] + 
                kernel_img_mul_63[36] + kernel_img_mul_63[37] + kernel_img_mul_63[38] + 
                kernel_img_mul_63[39] + kernel_img_mul_63[40] + kernel_img_mul_63[41] + 
                kernel_img_mul_63[42] + kernel_img_mul_63[43] + kernel_img_mul_63[44] + 
                kernel_img_mul_63[45] + kernel_img_mul_63[46] + kernel_img_mul_63[47] + 
                kernel_img_mul_63[48];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[7:0] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[7:0] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[7:0] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[15:8] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[15:8] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[15:8] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[23:16] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[23:16] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[23:16] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[31:24] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[31:24] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[31:24] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[39:32] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[39:32] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[39:32] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[47:40] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[47:40] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[47:40] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[55:48] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[55:48] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[55:48] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[63:56] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[63:56] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[63:56] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[71:64] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[71:64] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[71:64] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[79:72] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[79:72] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[79:72] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[87:80] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[87:80] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[87:80] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[95:88] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[95:88] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[95:88] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[103:96] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[103:96] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[103:96] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[111:104] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[111:104] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[111:104] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[119:112] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[119:112] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[119:112] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[127:120] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[127:120] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[127:120] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[135:128] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[135:128] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[135:128] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[143:136] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[143:136] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[143:136] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[151:144] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[151:144] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[151:144] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[159:152] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[159:152] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[159:152] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[167:160] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[167:160] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[167:160] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[175:168] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[175:168] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[175:168] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[183:176] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[183:176] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[183:176] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[191:184] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[191:184] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[191:184] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[199:192] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[199:192] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[199:192] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[207:200] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[207:200] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[207:200] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[215:208] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[215:208] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[215:208] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[223:216] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[223:216] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[223:216] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[231:224] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[231:224] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[231:224] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[239:232] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[239:232] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[239:232] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[247:240] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[247:240] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[247:240] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[255:248] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[255:248] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[255:248] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[263:256] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[263:256] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[263:256] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[271:264] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[271:264] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[271:264] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[279:272] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[279:272] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[279:272] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[287:280] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[287:280] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[287:280] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[295:288] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[295:288] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[295:288] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[303:296] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[303:296] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[303:296] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[311:304] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[311:304] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[311:304] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[319:312] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[319:312] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[319:312] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[327:320] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[327:320] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[327:320] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[335:328] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[335:328] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[335:328] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[343:336] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[343:336] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[343:336] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[351:344] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[351:344] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[351:344] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[359:352] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[359:352] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[359:352] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[367:360] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[367:360] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[367:360] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[375:368] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[375:368] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[375:368] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[383:376] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[383:376] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[383:376] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[391:384] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[391:384] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[391:384] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[399:392] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[399:392] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[399:392] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[407:400] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[407:400] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[407:400] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[415:408] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[415:408] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[415:408] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[423:416] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[423:416] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[423:416] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[431:424] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[431:424] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[431:424] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[439:432] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[439:432] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[439:432] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[447:440] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[447:440] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[447:440] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[455:448] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[455:448] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[455:448] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[463:456] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[463:456] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[463:456] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[471:464] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[471:464] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[471:464] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[479:472] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[479:472] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[479:472] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[487:480] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[487:480] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[487:480] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[495:488] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[495:488] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[495:488] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[503:496] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[503:496] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[503:496] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[511:504] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[511:504] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[511:504] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[519:512] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[519:512] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[519:512] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[527:520] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[527:520] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[527:520] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[535:528] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[535:528] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[535:528] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[543:536] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[543:536] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[543:536] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[551:544] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[551:544] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[551:544] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[559:552] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[559:552] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[559:552] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[567:560] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[567:560] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[567:560] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[575:568] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[575:568] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[575:568] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[583:576] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[583:576] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[583:576] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[591:584] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[591:584] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[591:584] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[599:592] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[599:592] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[599:592] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[607:600] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[607:600] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[607:600] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[615:608] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[615:608] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[615:608] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[623:616] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[623:616] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[623:616] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[631:624] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[631:624] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[631:624] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[639:632] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[639:632] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[639:632] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[647:640] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[647:640] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[647:640] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[655:648] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[655:648] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[655:648] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[663:656] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[663:656] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[663:656] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[671:664] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[671:664] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[671:664] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[679:672] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[679:672] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[679:672] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[687:680] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[687:680] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[687:680] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[695:688] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[695:688] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[695:688] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[703:696] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[703:696] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[703:696] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[711:704] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[711:704] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[711:704] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[719:712] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[719:712] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[719:712] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[727:720] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[727:720] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[727:720] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[735:728] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[735:728] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[735:728] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[743:736] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[743:736] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[743:736] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[751:744] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[751:744] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[751:744] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[759:752] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[759:752] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[759:752] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[767:760] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[767:760] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[767:760] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[775:768] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[775:768] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[775:768] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[783:776] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[783:776] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[783:776] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[791:784] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[791:784] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[791:784] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[799:792] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[799:792] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[799:792] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[807:800] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[807:800] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[807:800] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[815:808] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[815:808] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[815:808] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[823:816] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[823:816] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[823:816] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[831:824] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[831:824] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[831:824] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[839:832] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[839:832] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[839:832] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[847:840] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[847:840] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[847:840] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[855:848] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[855:848] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[855:848] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[863:856] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[863:856] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[863:856] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[871:864] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[871:864] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[871:864] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[879:872] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[879:872] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[879:872] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[887:880] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[887:880] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[887:880] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[895:888] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[895:888] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[895:888] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[903:896] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[903:896] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[903:896] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[911:904] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[911:904] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[911:904] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[919:912] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[919:912] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[919:912] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[927:920] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[927:920] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[927:920] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[935:928] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[935:928] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[935:928] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[943:936] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[943:936] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[943:936] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[951:944] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[951:944] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[951:944] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[959:952] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[959:952] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[959:952] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[967:960] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[967:960] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[967:960] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[975:968] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[975:968] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[975:968] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[983:976] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[983:976] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[983:976] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[991:984] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[991:984] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[991:984] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[999:992] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[999:992] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[999:992] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1007:1000] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[1007:1000] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1007:1000] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1015:1008] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[1015:1008] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1015:1008] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1023:1016] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[1023:1016] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1023:1016] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1031:1024] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1031:1024] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1031:1024] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1039:1032] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1039:1032] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1039:1032] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1047:1040] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1047:1040] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1047:1040] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1055:1048] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1055:1048] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1055:1048] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1063:1056] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1063:1056] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1063:1056] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1071:1064] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1071:1064] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1071:1064] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1079:1072] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1079:1072] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1079:1072] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1087:1080] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1087:1080] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1087:1080] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1095:1088] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1095:1088] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1095:1088] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1103:1096] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1103:1096] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1103:1096] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1111:1104] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1111:1104] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1111:1104] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1119:1112] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1119:1112] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1119:1112] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1127:1120] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1127:1120] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1127:1120] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1135:1128] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1135:1128] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1135:1128] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1143:1136] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1143:1136] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1143:1136] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1151:1144] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1151:1144] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1151:1144] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1159:1152] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1159:1152] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1159:1152] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1167:1160] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1167:1160] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1167:1160] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1175:1168] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1175:1168] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1175:1168] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1183:1176] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1183:1176] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1183:1176] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1191:1184] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1191:1184] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1191:1184] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1199:1192] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1199:1192] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1199:1192] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1207:1200] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1207:1200] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1207:1200] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1215:1208] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1215:1208] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1215:1208] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1223:1216] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1223:1216] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1223:1216] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1231:1224] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1231:1224] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1231:1224] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1239:1232] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1239:1232] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1239:1232] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1247:1240] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1247:1240] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1247:1240] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1255:1248] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1255:1248] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1255:1248] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1263:1256] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1263:1256] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1263:1256] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1271:1264] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1271:1264] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1271:1264] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1279:1272] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1279:1272] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1279:1272] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1287:1280] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1287:1280] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1287:1280] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1295:1288] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1295:1288] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1295:1288] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1303:1296] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1303:1296] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1303:1296] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1311:1304] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1311:1304] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1311:1304] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1319:1312] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1319:1312] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1319:1312] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1327:1320] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1327:1320] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1327:1320] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1335:1328] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1335:1328] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1335:1328] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1343:1336] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1343:1336] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1343:1336] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1351:1344] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1351:1344] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1351:1344] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1359:1352] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1359:1352] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1359:1352] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1367:1360] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1367:1360] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1367:1360] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1375:1368] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1375:1368] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1375:1368] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1383:1376] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1383:1376] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1383:1376] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1391:1384] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1391:1384] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1391:1384] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1399:1392] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1399:1392] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1399:1392] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1407:1400] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1407:1400] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1407:1400] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1415:1408] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1415:1408] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1415:1408] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1423:1416] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1423:1416] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1423:1416] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1431:1424] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1431:1424] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1431:1424] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1439:1432] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1439:1432] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1439:1432] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1447:1440] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1447:1440] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1447:1440] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1455:1448] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1455:1448] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1455:1448] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1463:1456] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1463:1456] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1463:1456] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1471:1464] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1471:1464] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1471:1464] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1479:1472] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1479:1472] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1479:1472] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1487:1480] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1487:1480] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1487:1480] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1495:1488] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1495:1488] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1495:1488] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1503:1496] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1503:1496] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1503:1496] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1511:1504] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1511:1504] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1511:1504] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1519:1512] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1519:1512] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1519:1512] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1527:1520] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1527:1520] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1527:1520] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1535:1528] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1535:1528] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1535:1528] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1543:1536] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1543:1536] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1543:1536] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1551:1544] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1551:1544] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1551:1544] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1559:1552] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1559:1552] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1559:1552] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1567:1560] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1567:1560] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1567:1560] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1575:1568] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1575:1568] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1575:1568] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1583:1576] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1583:1576] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1583:1576] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1591:1584] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1591:1584] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1591:1584] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1599:1592] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1599:1592] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1599:1592] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1607:1600] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1607:1600] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1607:1600] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1615:1608] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1615:1608] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1615:1608] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1623:1616] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1623:1616] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1623:1616] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1631:1624] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1631:1624] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1631:1624] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1639:1632] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1639:1632] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1639:1632] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1647:1640] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1647:1640] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1647:1640] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1655:1648] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1655:1648] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1655:1648] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1663:1656] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1663:1656] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1663:1656] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1671:1664] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1671:1664] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1671:1664] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1679:1672] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1679:1672] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1679:1672] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1687:1680] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1687:1680] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1687:1680] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1695:1688] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1695:1688] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1695:1688] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1703:1696] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1703:1696] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1703:1696] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1711:1704] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1711:1704] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1711:1704] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1719:1712] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1719:1712] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1719:1712] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1727:1720] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1727:1720] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1727:1720] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1735:1728] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1735:1728] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1735:1728] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1743:1736] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1743:1736] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1743:1736] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1751:1744] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1751:1744] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1751:1744] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1759:1752] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1759:1752] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1759:1752] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1767:1760] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1767:1760] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1767:1760] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1775:1768] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1775:1768] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1775:1768] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1783:1776] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1783:1776] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1783:1776] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1791:1784] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1791:1784] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1791:1784] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1799:1792] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1799:1792] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1799:1792] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1807:1800] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1807:1800] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1807:1800] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1815:1808] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1815:1808] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1815:1808] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1823:1816] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1823:1816] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1823:1816] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1831:1824] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1831:1824] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1831:1824] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1839:1832] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1839:1832] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1839:1832] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1847:1840] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1847:1840] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1847:1840] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1855:1848] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1855:1848] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1855:1848] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1863:1856] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1863:1856] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1863:1856] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1871:1864] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1871:1864] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1871:1864] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1879:1872] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1879:1872] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1879:1872] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1887:1880] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1887:1880] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1887:1880] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1895:1888] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1895:1888] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1895:1888] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1903:1896] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1903:1896] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1903:1896] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1911:1904] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1911:1904] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1911:1904] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1919:1912] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1919:1912] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1919:1912] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1927:1920] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1927:1920] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1927:1920] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1935:1928] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1935:1928] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1935:1928] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1943:1936] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1943:1936] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1943:1936] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1951:1944] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1951:1944] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1951:1944] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1959:1952] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1959:1952] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1959:1952] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1967:1960] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1967:1960] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1967:1960] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1975:1968] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1975:1968] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1975:1968] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1983:1976] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1983:1976] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1983:1976] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1991:1984] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1991:1984] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1991:1984] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1999:1992] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1999:1992] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1999:1992] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2007:2000] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[2007:2000] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2007:2000] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2015:2008] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[2015:2008] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2015:2008] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2023:2016] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[2023:2016] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2023:2016] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2031:2024] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[2031:2024] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2031:2024] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2039:2032] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[2039:2032] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2039:2032] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2047:2040] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[2047:2040] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2047:2040] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2055:2048] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2055:2048] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2055:2048] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2063:2056] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2063:2056] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2063:2056] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2071:2064] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2071:2064] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2071:2064] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2079:2072] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2079:2072] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2079:2072] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2087:2080] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2087:2080] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2087:2080] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2095:2088] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2095:2088] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2095:2088] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2103:2096] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2103:2096] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2103:2096] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2111:2104] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2111:2104] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2111:2104] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2119:2112] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2119:2112] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2119:2112] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2127:2120] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2127:2120] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2127:2120] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2135:2128] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2135:2128] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2135:2128] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2143:2136] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2143:2136] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2143:2136] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2151:2144] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2151:2144] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2151:2144] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2159:2152] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2159:2152] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2159:2152] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2167:2160] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2167:2160] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2167:2160] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2175:2168] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2175:2168] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2175:2168] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2183:2176] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2183:2176] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2183:2176] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2191:2184] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2191:2184] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2191:2184] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2199:2192] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2199:2192] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2199:2192] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2207:2200] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2207:2200] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2207:2200] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2215:2208] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2215:2208] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2215:2208] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2223:2216] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2223:2216] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2223:2216] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2231:2224] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2231:2224] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2231:2224] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2239:2232] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2239:2232] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2239:2232] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2247:2240] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2247:2240] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2247:2240] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2255:2248] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2255:2248] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2255:2248] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2263:2256] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2263:2256] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2263:2256] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2271:2264] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2271:2264] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2271:2264] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2279:2272] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2279:2272] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2279:2272] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2287:2280] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2287:2280] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2287:2280] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2295:2288] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2295:2288] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2295:2288] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2303:2296] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2303:2296] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2303:2296] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2311:2304] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2311:2304] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2311:2304] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2319:2312] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2319:2312] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2319:2312] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2327:2320] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2327:2320] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2327:2320] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2335:2328] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2335:2328] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2335:2328] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2343:2336] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2343:2336] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2343:2336] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2351:2344] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2351:2344] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2351:2344] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2359:2352] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2359:2352] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2359:2352] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2367:2360] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2367:2360] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2367:2360] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2375:2368] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2375:2368] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2375:2368] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2383:2376] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2383:2376] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2383:2376] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2391:2384] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2391:2384] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2391:2384] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2399:2392] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2399:2392] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2399:2392] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2407:2400] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2407:2400] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2407:2400] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2415:2408] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2415:2408] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2415:2408] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2423:2416] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2423:2416] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2423:2416] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2431:2424] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2431:2424] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2431:2424] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2439:2432] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2439:2432] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2439:2432] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2447:2440] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2447:2440] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2447:2440] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2455:2448] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2455:2448] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2455:2448] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2463:2456] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2463:2456] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2463:2456] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2471:2464] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2471:2464] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2471:2464] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2479:2472] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2479:2472] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2479:2472] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2487:2480] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2487:2480] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2487:2480] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2495:2488] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2495:2488] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2495:2488] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2503:2496] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2503:2496] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2503:2496] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2511:2504] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2511:2504] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2511:2504] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2519:2512] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2519:2512] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2519:2512] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2527:2520] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2527:2520] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2527:2520] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2535:2528] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2535:2528] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2535:2528] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2543:2536] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2543:2536] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2543:2536] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2551:2544] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2551:2544] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2551:2544] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2559:2552] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2559:2552] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2559:2552] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2567:2560] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2567:2560] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2567:2560] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2575:2568] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2575:2568] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2575:2568] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2583:2576] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2583:2576] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2583:2576] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2591:2584] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2591:2584] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2591:2584] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2599:2592] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2599:2592] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2599:2592] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2607:2600] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2607:2600] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2607:2600] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2615:2608] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2615:2608] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2615:2608] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2623:2616] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2623:2616] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2623:2616] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2631:2624] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2631:2624] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2631:2624] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2639:2632] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2639:2632] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2639:2632] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2647:2640] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2647:2640] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2647:2640] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2655:2648] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2655:2648] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2655:2648] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2663:2656] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2663:2656] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2663:2656] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2671:2664] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2671:2664] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2671:2664] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2679:2672] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2679:2672] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2679:2672] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2687:2680] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2687:2680] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2687:2680] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2695:2688] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2695:2688] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2695:2688] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2703:2696] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2703:2696] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2703:2696] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2711:2704] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2711:2704] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2711:2704] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2719:2712] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2719:2712] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2719:2712] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2727:2720] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2727:2720] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2727:2720] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2735:2728] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2735:2728] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2735:2728] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2743:2736] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2743:2736] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2743:2736] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2751:2744] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2751:2744] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2751:2744] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2759:2752] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2759:2752] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2759:2752] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2767:2760] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2767:2760] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2767:2760] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2775:2768] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2775:2768] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2775:2768] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2783:2776] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2783:2776] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2783:2776] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2791:2784] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2791:2784] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2791:2784] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2799:2792] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2799:2792] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2799:2792] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2807:2800] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2807:2800] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2807:2800] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2815:2808] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2815:2808] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2815:2808] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2823:2816] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2823:2816] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2823:2816] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2831:2824] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2831:2824] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2831:2824] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2839:2832] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2839:2832] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2839:2832] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2847:2840] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2847:2840] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2847:2840] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2855:2848] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2855:2848] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2855:2848] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2863:2856] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2863:2856] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2863:2856] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2871:2864] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2871:2864] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2871:2864] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2879:2872] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2879:2872] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2879:2872] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2887:2880] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2887:2880] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2887:2880] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2895:2888] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2895:2888] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2895:2888] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2903:2896] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2903:2896] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2903:2896] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2911:2904] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2911:2904] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2911:2904] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2919:2912] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2919:2912] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2919:2912] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2927:2920] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2927:2920] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2927:2920] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2935:2928] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2935:2928] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2935:2928] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2943:2936] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2943:2936] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2943:2936] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2951:2944] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2951:2944] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2951:2944] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2959:2952] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2959:2952] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2959:2952] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2967:2960] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2967:2960] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2967:2960] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2975:2968] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2975:2968] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2975:2968] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2983:2976] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2983:2976] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2983:2976] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2991:2984] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2991:2984] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2991:2984] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2999:2992] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2999:2992] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2999:2992] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3007:3000] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3007:3000] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3007:3000] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3015:3008] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3015:3008] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3015:3008] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3023:3016] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3023:3016] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3023:3016] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3031:3024] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3031:3024] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3031:3024] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3039:3032] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3039:3032] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3039:3032] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3047:3040] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3047:3040] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3047:3040] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3055:3048] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3055:3048] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3055:3048] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3063:3056] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3063:3056] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3063:3056] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3071:3064] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3071:3064] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3071:3064] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3079:3072] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3079:3072] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3079:3072] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3087:3080] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3087:3080] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3087:3080] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3095:3088] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3095:3088] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3095:3088] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3103:3096] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3103:3096] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3103:3096] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3111:3104] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3111:3104] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3111:3104] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3119:3112] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3119:3112] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3119:3112] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3127:3120] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3127:3120] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3127:3120] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3135:3128] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3135:3128] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3135:3128] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3143:3136] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3143:3136] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3143:3136] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3151:3144] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3151:3144] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3151:3144] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3159:3152] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3159:3152] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3159:3152] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3167:3160] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3167:3160] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3167:3160] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3175:3168] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3175:3168] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3175:3168] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3183:3176] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3183:3176] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3183:3176] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3191:3184] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3191:3184] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3191:3184] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3199:3192] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3199:3192] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3199:3192] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3207:3200] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3207:3200] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3207:3200] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3215:3208] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3215:3208] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3215:3208] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3223:3216] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3223:3216] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3223:3216] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3231:3224] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3231:3224] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3231:3224] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3239:3232] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3239:3232] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3239:3232] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3247:3240] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3247:3240] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3247:3240] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3255:3248] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3255:3248] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3255:3248] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3263:3256] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3263:3256] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3263:3256] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3271:3264] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3271:3264] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3271:3264] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3279:3272] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3279:3272] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3279:3272] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3287:3280] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3287:3280] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3287:3280] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3295:3288] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3295:3288] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3295:3288] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3303:3296] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3303:3296] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3303:3296] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3311:3304] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3311:3304] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3311:3304] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3319:3312] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3319:3312] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3319:3312] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3327:3320] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3327:3320] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3327:3320] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3335:3328] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3335:3328] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3335:3328] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3343:3336] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3343:3336] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3343:3336] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3351:3344] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3351:3344] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3351:3344] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3359:3352] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3359:3352] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3359:3352] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3367:3360] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3367:3360] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3367:3360] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3375:3368] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3375:3368] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3375:3368] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3383:3376] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3383:3376] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3383:3376] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3391:3384] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3391:3384] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3391:3384] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3399:3392] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3399:3392] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3399:3392] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3407:3400] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3407:3400] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3407:3400] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3415:3408] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3415:3408] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3415:3408] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3423:3416] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3423:3416] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3423:3416] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3431:3424] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3431:3424] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3431:3424] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3439:3432] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3439:3432] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3439:3432] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3447:3440] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3447:3440] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3447:3440] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3455:3448] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3455:3448] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3455:3448] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3463:3456] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3463:3456] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3463:3456] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3471:3464] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3471:3464] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3471:3464] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3479:3472] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3479:3472] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3479:3472] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3487:3480] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3487:3480] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3487:3480] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3495:3488] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3495:3488] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3495:3488] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3503:3496] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3503:3496] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3503:3496] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3511:3504] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3511:3504] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3511:3504] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3519:3512] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3519:3512] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3519:3512] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3527:3520] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3527:3520] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3527:3520] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3535:3528] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3535:3528] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3535:3528] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3543:3536] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3543:3536] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3543:3536] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3551:3544] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3551:3544] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3551:3544] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3559:3552] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3559:3552] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3559:3552] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3567:3560] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3567:3560] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3567:3560] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3575:3568] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3575:3568] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3575:3568] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3583:3576] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3583:3576] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3583:3576] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3591:3584] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3591:3584] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3591:3584] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3599:3592] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3599:3592] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3599:3592] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3607:3600] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3607:3600] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3607:3600] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3615:3608] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3615:3608] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3615:3608] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3623:3616] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3623:3616] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3623:3616] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3631:3624] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3631:3624] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3631:3624] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3639:3632] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3639:3632] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3639:3632] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3647:3640] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3647:3640] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3647:3640] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3655:3648] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3655:3648] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3655:3648] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3663:3656] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3663:3656] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3663:3656] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3671:3664] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3671:3664] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3671:3664] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3679:3672] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3679:3672] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3679:3672] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3687:3680] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3687:3680] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3687:3680] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3695:3688] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3695:3688] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3695:3688] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3703:3696] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3703:3696] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3703:3696] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3711:3704] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3711:3704] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3711:3704] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3719:3712] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3719:3712] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3719:3712] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3727:3720] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3727:3720] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3727:3720] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3735:3728] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3735:3728] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3735:3728] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3743:3736] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3743:3736] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3743:3736] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3751:3744] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3751:3744] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3751:3744] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3759:3752] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3759:3752] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3759:3752] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3767:3760] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3767:3760] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3767:3760] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3775:3768] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3775:3768] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3775:3768] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3783:3776] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3783:3776] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3783:3776] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3791:3784] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3791:3784] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3791:3784] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3799:3792] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3799:3792] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3799:3792] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3807:3800] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3807:3800] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3807:3800] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3815:3808] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3815:3808] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3815:3808] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3823:3816] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3823:3816] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3823:3816] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3831:3824] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3831:3824] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3831:3824] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3839:3832] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3839:3832] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3839:3832] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3847:3840] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3847:3840] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3847:3840] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3855:3848] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3855:3848] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3855:3848] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3863:3856] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3863:3856] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3863:3856] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3871:3864] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3871:3864] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3871:3864] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3879:3872] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3879:3872] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3879:3872] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3887:3880] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3887:3880] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3887:3880] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3895:3888] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3895:3888] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3895:3888] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3903:3896] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3903:3896] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3903:3896] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3911:3904] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3911:3904] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3911:3904] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3919:3912] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3919:3912] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3919:3912] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3927:3920] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3927:3920] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3927:3920] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3935:3928] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3935:3928] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3935:3928] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3943:3936] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3943:3936] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3943:3936] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3951:3944] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3951:3944] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3951:3944] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3959:3952] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3959:3952] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3959:3952] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3967:3960] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3967:3960] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3967:3960] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3975:3968] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3975:3968] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3975:3968] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3983:3976] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3983:3976] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3983:3976] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3991:3984] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3991:3984] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3991:3984] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3999:3992] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3999:3992] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3999:3992] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4007:4000] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4007:4000] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4007:4000] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4015:4008] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4015:4008] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4015:4008] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4023:4016] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4023:4016] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4023:4016] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4031:4024] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4031:4024] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4031:4024] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4039:4032] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4039:4032] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4039:4032] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4047:4040] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4047:4040] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4047:4040] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4055:4048] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4055:4048] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4055:4048] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4063:4056] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4063:4056] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4063:4056] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4071:4064] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4071:4064] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4071:4064] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4079:4072] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4079:4072] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4079:4072] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4087:4080] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4087:4080] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4087:4080] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4095:4088] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4095:4088] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4095:4088] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4103:4096] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4103:4096] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4103:4096] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4111:4104] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4111:4104] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4111:4104] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4119:4112] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4119:4112] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4119:4112] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4127:4120] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4127:4120] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4127:4120] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4135:4128] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4135:4128] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4135:4128] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4143:4136] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4143:4136] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4143:4136] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4151:4144] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4151:4144] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4151:4144] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4159:4152] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4159:4152] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4159:4152] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4167:4160] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4167:4160] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4167:4160] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4175:4168] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4175:4168] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4175:4168] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4183:4176] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4183:4176] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4183:4176] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4191:4184] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4191:4184] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4191:4184] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4199:4192] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4199:4192] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4199:4192] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4207:4200] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4207:4200] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4207:4200] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4215:4208] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4215:4208] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4215:4208] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4223:4216] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4223:4216] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4223:4216] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4231:4224] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4231:4224] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4231:4224] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4239:4232] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4239:4232] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4239:4232] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4247:4240] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4247:4240] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4247:4240] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4255:4248] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4255:4248] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4255:4248] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4263:4256] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4263:4256] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4263:4256] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4271:4264] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4271:4264] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4271:4264] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4279:4272] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4279:4272] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4279:4272] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4287:4280] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4287:4280] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4287:4280] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4295:4288] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4295:4288] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4295:4288] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4303:4296] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4303:4296] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4303:4296] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4311:4304] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4311:4304] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4311:4304] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4319:4312] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4319:4312] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4319:4312] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4327:4320] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4327:4320] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4327:4320] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4335:4328] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4335:4328] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4335:4328] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4343:4336] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4343:4336] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4343:4336] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4351:4344] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4351:4344] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4351:4344] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4359:4352] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4359:4352] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4359:4352] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4367:4360] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4367:4360] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4367:4360] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4375:4368] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4375:4368] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4375:4368] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4383:4376] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4383:4376] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4383:4376] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4391:4384] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4391:4384] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4391:4384] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4399:4392] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4399:4392] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4399:4392] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4407:4400] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4407:4400] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4407:4400] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4415:4408] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4415:4408] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4415:4408] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4423:4416] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4423:4416] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4423:4416] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4431:4424] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4431:4424] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4431:4424] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4439:4432] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4439:4432] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4439:4432] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4447:4440] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4447:4440] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4447:4440] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4455:4448] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4455:4448] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4455:4448] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4463:4456] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4463:4456] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4463:4456] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4471:4464] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4471:4464] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4471:4464] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4479:4472] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4479:4472] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4479:4472] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4487:4480] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4487:4480] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4487:4480] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4495:4488] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4495:4488] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4495:4488] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4503:4496] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4503:4496] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4503:4496] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4511:4504] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4511:4504] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4511:4504] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4519:4512] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4519:4512] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4519:4512] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4527:4520] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4527:4520] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4527:4520] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4535:4528] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4535:4528] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4535:4528] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4543:4536] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4543:4536] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4543:4536] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4551:4544] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4551:4544] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4551:4544] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4559:4552] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4559:4552] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4559:4552] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4567:4560] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4567:4560] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4567:4560] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4575:4568] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4575:4568] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4575:4568] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4583:4576] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4583:4576] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4583:4576] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4591:4584] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4591:4584] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4591:4584] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4599:4592] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4599:4592] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4599:4592] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4607:4600] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4607:4600] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4607:4600] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4615:4608] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4615:4608] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4615:4608] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4623:4616] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4623:4616] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4623:4616] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4631:4624] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4631:4624] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4631:4624] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4639:4632] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4639:4632] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4639:4632] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4647:4640] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4647:4640] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4647:4640] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4655:4648] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4655:4648] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4655:4648] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4663:4656] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4663:4656] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4663:4656] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4671:4664] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4671:4664] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4671:4664] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4679:4672] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4679:4672] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4679:4672] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4687:4680] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4687:4680] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4687:4680] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4695:4688] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4695:4688] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4695:4688] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4703:4696] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4703:4696] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4703:4696] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4711:4704] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4711:4704] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4711:4704] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4719:4712] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4719:4712] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4719:4712] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4727:4720] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4727:4720] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4727:4720] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4735:4728] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4735:4728] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4735:4728] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4743:4736] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4743:4736] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4743:4736] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4751:4744] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4751:4744] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4751:4744] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4759:4752] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4759:4752] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4759:4752] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4767:4760] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4767:4760] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4767:4760] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4775:4768] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4775:4768] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4775:4768] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4783:4776] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4783:4776] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4783:4776] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4791:4784] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4791:4784] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4791:4784] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4799:4792] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4799:4792] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4799:4792] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4807:4800] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4807:4800] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4807:4800] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4815:4808] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4815:4808] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4815:4808] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4823:4816] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4823:4816] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4823:4816] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4831:4824] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4831:4824] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4831:4824] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4839:4832] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4839:4832] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4839:4832] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4847:4840] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4847:4840] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4847:4840] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4855:4848] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4855:4848] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4855:4848] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4863:4856] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4863:4856] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4863:4856] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4871:4864] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4871:4864] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4871:4864] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4879:4872] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4879:4872] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4879:4872] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4887:4880] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4887:4880] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4887:4880] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4895:4888] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4895:4888] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4895:4888] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4903:4896] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4903:4896] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4903:4896] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4911:4904] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4911:4904] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4911:4904] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4919:4912] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4919:4912] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4919:4912] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4927:4920] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4927:4920] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4927:4920] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4935:4928] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4935:4928] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4935:4928] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4943:4936] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4943:4936] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4943:4936] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4951:4944] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4951:4944] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4951:4944] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4959:4952] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4959:4952] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4959:4952] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4967:4960] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4967:4960] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4967:4960] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4975:4968] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4975:4968] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4975:4968] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4983:4976] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4983:4976] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4983:4976] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4991:4984] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4991:4984] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4991:4984] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4999:4992] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4999:4992] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4999:4992] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5007:5000] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5007:5000] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5007:5000] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5015:5008] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5015:5008] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5015:5008] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5023:5016] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5023:5016] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5023:5016] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5031:5024] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5031:5024] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5031:5024] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5039:5032] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5039:5032] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5039:5032] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5047:5040] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5047:5040] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5047:5040] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5055:5048] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5055:5048] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5055:5048] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5063:5056] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5063:5056] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5063:5056] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5071:5064] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5071:5064] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5071:5064] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5079:5072] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5079:5072] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5079:5072] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5087:5080] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5087:5080] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5087:5080] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5095:5088] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5095:5088] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5095:5088] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5103:5096] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5103:5096] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5103:5096] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5111:5104] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5111:5104] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5111:5104] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5119:5112] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5119:5112] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5119:5112] <= 'd0;
end


endmodule