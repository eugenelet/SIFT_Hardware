`timescale 1ns/10ps
module Line_Buffer_10(
  clk,
  rst_n,
  buffer_mode,
  buffer_we,
  fill_zero,
  in_data0,
  in_data1,
  in_data2,
  in_data3,
  in_data4,
  buffer_data_0,
  buffer_data_1,
  buffer_data_2,
  buffer_data_3,
  buffer_data_4,
  buffer_data_5,
  buffer_data_6,
  buffer_data_7,
  buffer_data_8,
  buffer_data_9,
  buffer_col
);
/*SYSTEM*/
input                 clk,
                      rst_n;

/*From SRAM*/
input       [5119:0]  in_data0;
input       [5119:0]  in_data1;
input       [5119:0]  in_data2;
input       [5119:0]  in_data3;
input       [5119:0]  in_data4;

/*Current Column 640/16*/
input[5:0]  buffer_col;

/*From Working Module*/
input                 buffer_mode; /*0: 10 regs as a group   1: 5 groups, 2 each*/
input                 buffer_we;
input                 fill_zero; /*Used in Gaussian blur & Match*/

/*BUFFER OUT*/
output reg  [175:0]   buffer_data_0, // (16 + 6)*8
                      buffer_data_1,
                      buffer_data_2,
                      buffer_data_3,
                      buffer_data_4,
                      buffer_data_5,
                      buffer_data_6,
                      buffer_data_7,
                      buffer_data_8,
                      buffer_data_9;

reg[175:0]  mux_data0,
            mux_data1,
            mux_data2,
            mux_data3,
            mux_data4;

always @(*) begin
  case(buffer_col)
    'd0: begin
      mux_data0[7:0] = 'd0;
      mux_data0[15:8] = 'd0;
      mux_data0[23:16] = 'd0;
      mux_data0[31:24] = in_data0[7:0];
      mux_data0[39:32] = in_data0[15:8];
      mux_data0[47:40] = in_data0[23:16];
      mux_data0[55:48] = in_data0[31:24];
      mux_data0[63:56] = in_data0[39:32];
      mux_data0[71:64] = in_data0[47:40];
      mux_data0[79:72] = in_data0[55:48];
      mux_data0[87:80] = in_data0[63:56];
      mux_data0[95:88] = in_data0[71:64];
      mux_data0[103:96] = in_data0[79:72];
      mux_data0[111:104] = in_data0[87:80];
      mux_data0[119:112] = in_data0[95:88];
      mux_data0[127:120] = in_data0[103:96];
      mux_data0[135:128] = in_data0[111:104];
      mux_data0[143:136] = in_data0[119:112];
      mux_data0[151:144] = in_data0[127:120];
      mux_data0[159:152] = in_data0[135:128];
      mux_data0[167:160] = in_data0[143:136];
      mux_data0[175:168] = in_data0[151:144];
      mux_data1[7:0] = 'd0;
      mux_data1[15:8] = 'd0;
      mux_data1[23:16] = 'd0;
      mux_data1[31:24] = in_data1[7:0];
      mux_data1[39:32] = in_data1[15:8];
      mux_data1[47:40] = in_data1[23:16];
      mux_data1[55:48] = in_data1[31:24];
      mux_data1[63:56] = in_data1[39:32];
      mux_data1[71:64] = in_data1[47:40];
      mux_data1[79:72] = in_data1[55:48];
      mux_data1[87:80] = in_data1[63:56];
      mux_data1[95:88] = in_data1[71:64];
      mux_data1[103:96] = in_data1[79:72];
      mux_data1[111:104] = in_data1[87:80];
      mux_data1[119:112] = in_data1[95:88];
      mux_data1[127:120] = in_data1[103:96];
      mux_data1[135:128] = in_data1[111:104];
      mux_data1[143:136] = in_data1[119:112];
      mux_data1[151:144] = in_data1[127:120];
      mux_data1[159:152] = in_data1[135:128];
      mux_data1[167:160] = in_data1[143:136];
      mux_data1[175:168] = in_data1[151:144];
      mux_data2[7:0] = 'd0;
      mux_data2[15:8] = 'd0;
      mux_data2[23:16] = 'd0;
      mux_data2[31:24] = in_data2[7:0];
      mux_data2[39:32] = in_data2[15:8];
      mux_data2[47:40] = in_data2[23:16];
      mux_data2[55:48] = in_data2[31:24];
      mux_data2[63:56] = in_data2[39:32];
      mux_data2[71:64] = in_data2[47:40];
      mux_data2[79:72] = in_data2[55:48];
      mux_data2[87:80] = in_data2[63:56];
      mux_data2[95:88] = in_data2[71:64];
      mux_data2[103:96] = in_data2[79:72];
      mux_data2[111:104] = in_data2[87:80];
      mux_data2[119:112] = in_data2[95:88];
      mux_data2[127:120] = in_data2[103:96];
      mux_data2[135:128] = in_data2[111:104];
      mux_data2[143:136] = in_data2[119:112];
      mux_data2[151:144] = in_data2[127:120];
      mux_data2[159:152] = in_data2[135:128];
      mux_data2[167:160] = in_data2[143:136];
      mux_data2[175:168] = in_data2[151:144];
      mux_data3[7:0] = 'd0;
      mux_data3[15:8] = 'd0;
      mux_data3[23:16] = 'd0;
      mux_data3[31:24] = in_data3[7:0];
      mux_data3[39:32] = in_data3[15:8];
      mux_data3[47:40] = in_data3[23:16];
      mux_data3[55:48] = in_data3[31:24];
      mux_data3[63:56] = in_data3[39:32];
      mux_data3[71:64] = in_data3[47:40];
      mux_data3[79:72] = in_data3[55:48];
      mux_data3[87:80] = in_data3[63:56];
      mux_data3[95:88] = in_data3[71:64];
      mux_data3[103:96] = in_data3[79:72];
      mux_data3[111:104] = in_data3[87:80];
      mux_data3[119:112] = in_data3[95:88];
      mux_data3[127:120] = in_data3[103:96];
      mux_data3[135:128] = in_data3[111:104];
      mux_data3[143:136] = in_data3[119:112];
      mux_data3[151:144] = in_data3[127:120];
      mux_data3[159:152] = in_data3[135:128];
      mux_data3[167:160] = in_data3[143:136];
      mux_data3[175:168] = in_data3[151:144];
      mux_data4[7:0] = 'd0;
      mux_data4[15:8] = 'd0;
      mux_data4[23:16] = 'd0;
      mux_data4[31:24] = in_data4[7:0];
      mux_data4[39:32] = in_data4[15:8];
      mux_data4[47:40] = in_data4[23:16];
      mux_data4[55:48] = in_data4[31:24];
      mux_data4[63:56] = in_data4[39:32];
      mux_data4[71:64] = in_data4[47:40];
      mux_data4[79:72] = in_data4[55:48];
      mux_data4[87:80] = in_data4[63:56];
      mux_data4[95:88] = in_data4[71:64];
      mux_data4[103:96] = in_data4[79:72];
      mux_data4[111:104] = in_data4[87:80];
      mux_data4[119:112] = in_data4[95:88];
      mux_data4[127:120] = in_data4[103:96];
      mux_data4[135:128] = in_data4[111:104];
      mux_data4[143:136] = in_data4[119:112];
      mux_data4[151:144] = in_data4[127:120];
      mux_data4[159:152] = in_data4[135:128];
      mux_data4[167:160] = in_data4[143:136];
      mux_data4[175:168] = in_data4[151:144];
    end
    'd1: begin
      mux_data0[7:0] = in_data0[111:104];
      mux_data0[15:8] = in_data0[119:112];
      mux_data0[23:16] = in_data0[127:120];
      mux_data0[31:24] = in_data0[135:128];
      mux_data0[39:32] = in_data0[143:136];
      mux_data0[47:40] = in_data0[151:144];
      mux_data0[55:48] = in_data0[159:152];
      mux_data0[63:56] = in_data0[167:160];
      mux_data0[71:64] = in_data0[175:168];
      mux_data0[79:72] = in_data0[183:176];
      mux_data0[87:80] = in_data0[191:184];
      mux_data0[95:88] = in_data0[199:192];
      mux_data0[103:96] = in_data0[207:200];
      mux_data0[111:104] = in_data0[215:208];
      mux_data0[119:112] = in_data0[223:216];
      mux_data0[127:120] = in_data0[231:224];
      mux_data0[135:128] = in_data0[239:232];
      mux_data0[143:136] = in_data0[247:240];
      mux_data0[151:144] = in_data0[255:248];
      mux_data0[159:152] = in_data0[263:256];
      mux_data0[167:160] = in_data0[271:264];
      mux_data0[175:168] = in_data0[279:272];
      mux_data1[7:0] = in_data1[111:104];
      mux_data1[15:8] = in_data1[119:112];
      mux_data1[23:16] = in_data1[127:120];
      mux_data1[31:24] = in_data1[135:128];
      mux_data1[39:32] = in_data1[143:136];
      mux_data1[47:40] = in_data1[151:144];
      mux_data1[55:48] = in_data1[159:152];
      mux_data1[63:56] = in_data1[167:160];
      mux_data1[71:64] = in_data1[175:168];
      mux_data1[79:72] = in_data1[183:176];
      mux_data1[87:80] = in_data1[191:184];
      mux_data1[95:88] = in_data1[199:192];
      mux_data1[103:96] = in_data1[207:200];
      mux_data1[111:104] = in_data1[215:208];
      mux_data1[119:112] = in_data1[223:216];
      mux_data1[127:120] = in_data1[231:224];
      mux_data1[135:128] = in_data1[239:232];
      mux_data1[143:136] = in_data1[247:240];
      mux_data1[151:144] = in_data1[255:248];
      mux_data1[159:152] = in_data1[263:256];
      mux_data1[167:160] = in_data1[271:264];
      mux_data1[175:168] = in_data1[279:272];
      mux_data2[7:0] = in_data2[111:104];
      mux_data2[15:8] = in_data2[119:112];
      mux_data2[23:16] = in_data2[127:120];
      mux_data2[31:24] = in_data2[135:128];
      mux_data2[39:32] = in_data2[143:136];
      mux_data2[47:40] = in_data2[151:144];
      mux_data2[55:48] = in_data2[159:152];
      mux_data2[63:56] = in_data2[167:160];
      mux_data2[71:64] = in_data2[175:168];
      mux_data2[79:72] = in_data2[183:176];
      mux_data2[87:80] = in_data2[191:184];
      mux_data2[95:88] = in_data2[199:192];
      mux_data2[103:96] = in_data2[207:200];
      mux_data2[111:104] = in_data2[215:208];
      mux_data2[119:112] = in_data2[223:216];
      mux_data2[127:120] = in_data2[231:224];
      mux_data2[135:128] = in_data2[239:232];
      mux_data2[143:136] = in_data2[247:240];
      mux_data2[151:144] = in_data2[255:248];
      mux_data2[159:152] = in_data2[263:256];
      mux_data2[167:160] = in_data2[271:264];
      mux_data2[175:168] = in_data2[279:272];
      mux_data3[7:0] = in_data3[111:104];
      mux_data3[15:8] = in_data3[119:112];
      mux_data3[23:16] = in_data3[127:120];
      mux_data3[31:24] = in_data3[135:128];
      mux_data3[39:32] = in_data3[143:136];
      mux_data3[47:40] = in_data3[151:144];
      mux_data3[55:48] = in_data3[159:152];
      mux_data3[63:56] = in_data3[167:160];
      mux_data3[71:64] = in_data3[175:168];
      mux_data3[79:72] = in_data3[183:176];
      mux_data3[87:80] = in_data3[191:184];
      mux_data3[95:88] = in_data3[199:192];
      mux_data3[103:96] = in_data3[207:200];
      mux_data3[111:104] = in_data3[215:208];
      mux_data3[119:112] = in_data3[223:216];
      mux_data3[127:120] = in_data3[231:224];
      mux_data3[135:128] = in_data3[239:232];
      mux_data3[143:136] = in_data3[247:240];
      mux_data3[151:144] = in_data3[255:248];
      mux_data3[159:152] = in_data3[263:256];
      mux_data3[167:160] = in_data3[271:264];
      mux_data3[175:168] = in_data3[279:272];
      mux_data4[7:0] = in_data4[111:104];
      mux_data4[15:8] = in_data4[119:112];
      mux_data4[23:16] = in_data4[127:120];
      mux_data4[31:24] = in_data4[135:128];
      mux_data4[39:32] = in_data4[143:136];
      mux_data4[47:40] = in_data4[151:144];
      mux_data4[55:48] = in_data4[159:152];
      mux_data4[63:56] = in_data4[167:160];
      mux_data4[71:64] = in_data4[175:168];
      mux_data4[79:72] = in_data4[183:176];
      mux_data4[87:80] = in_data4[191:184];
      mux_data4[95:88] = in_data4[199:192];
      mux_data4[103:96] = in_data4[207:200];
      mux_data4[111:104] = in_data4[215:208];
      mux_data4[119:112] = in_data4[223:216];
      mux_data4[127:120] = in_data4[231:224];
      mux_data4[135:128] = in_data4[239:232];
      mux_data4[143:136] = in_data4[247:240];
      mux_data4[151:144] = in_data4[255:248];
      mux_data4[159:152] = in_data4[263:256];
      mux_data4[167:160] = in_data4[271:264];
      mux_data4[175:168] = in_data4[279:272];
    end
    'd2: begin
      mux_data0[7:0] = in_data0[239:232];
      mux_data0[15:8] = in_data0[247:240];
      mux_data0[23:16] = in_data0[255:248];
      mux_data0[31:24] = in_data0[263:256];
      mux_data0[39:32] = in_data0[271:264];
      mux_data0[47:40] = in_data0[279:272];
      mux_data0[55:48] = in_data0[287:280];
      mux_data0[63:56] = in_data0[295:288];
      mux_data0[71:64] = in_data0[303:296];
      mux_data0[79:72] = in_data0[311:304];
      mux_data0[87:80] = in_data0[319:312];
      mux_data0[95:88] = in_data0[327:320];
      mux_data0[103:96] = in_data0[335:328];
      mux_data0[111:104] = in_data0[343:336];
      mux_data0[119:112] = in_data0[351:344];
      mux_data0[127:120] = in_data0[359:352];
      mux_data0[135:128] = in_data0[367:360];
      mux_data0[143:136] = in_data0[375:368];
      mux_data0[151:144] = in_data0[383:376];
      mux_data0[159:152] = in_data0[391:384];
      mux_data0[167:160] = in_data0[399:392];
      mux_data0[175:168] = in_data0[407:400];
      mux_data1[7:0] = in_data1[239:232];
      mux_data1[15:8] = in_data1[247:240];
      mux_data1[23:16] = in_data1[255:248];
      mux_data1[31:24] = in_data1[263:256];
      mux_data1[39:32] = in_data1[271:264];
      mux_data1[47:40] = in_data1[279:272];
      mux_data1[55:48] = in_data1[287:280];
      mux_data1[63:56] = in_data1[295:288];
      mux_data1[71:64] = in_data1[303:296];
      mux_data1[79:72] = in_data1[311:304];
      mux_data1[87:80] = in_data1[319:312];
      mux_data1[95:88] = in_data1[327:320];
      mux_data1[103:96] = in_data1[335:328];
      mux_data1[111:104] = in_data1[343:336];
      mux_data1[119:112] = in_data1[351:344];
      mux_data1[127:120] = in_data1[359:352];
      mux_data1[135:128] = in_data1[367:360];
      mux_data1[143:136] = in_data1[375:368];
      mux_data1[151:144] = in_data1[383:376];
      mux_data1[159:152] = in_data1[391:384];
      mux_data1[167:160] = in_data1[399:392];
      mux_data1[175:168] = in_data1[407:400];
      mux_data2[7:0] = in_data2[239:232];
      mux_data2[15:8] = in_data2[247:240];
      mux_data2[23:16] = in_data2[255:248];
      mux_data2[31:24] = in_data2[263:256];
      mux_data2[39:32] = in_data2[271:264];
      mux_data2[47:40] = in_data2[279:272];
      mux_data2[55:48] = in_data2[287:280];
      mux_data2[63:56] = in_data2[295:288];
      mux_data2[71:64] = in_data2[303:296];
      mux_data2[79:72] = in_data2[311:304];
      mux_data2[87:80] = in_data2[319:312];
      mux_data2[95:88] = in_data2[327:320];
      mux_data2[103:96] = in_data2[335:328];
      mux_data2[111:104] = in_data2[343:336];
      mux_data2[119:112] = in_data2[351:344];
      mux_data2[127:120] = in_data2[359:352];
      mux_data2[135:128] = in_data2[367:360];
      mux_data2[143:136] = in_data2[375:368];
      mux_data2[151:144] = in_data2[383:376];
      mux_data2[159:152] = in_data2[391:384];
      mux_data2[167:160] = in_data2[399:392];
      mux_data2[175:168] = in_data2[407:400];
      mux_data3[7:0] = in_data3[239:232];
      mux_data3[15:8] = in_data3[247:240];
      mux_data3[23:16] = in_data3[255:248];
      mux_data3[31:24] = in_data3[263:256];
      mux_data3[39:32] = in_data3[271:264];
      mux_data3[47:40] = in_data3[279:272];
      mux_data3[55:48] = in_data3[287:280];
      mux_data3[63:56] = in_data3[295:288];
      mux_data3[71:64] = in_data3[303:296];
      mux_data3[79:72] = in_data3[311:304];
      mux_data3[87:80] = in_data3[319:312];
      mux_data3[95:88] = in_data3[327:320];
      mux_data3[103:96] = in_data3[335:328];
      mux_data3[111:104] = in_data3[343:336];
      mux_data3[119:112] = in_data3[351:344];
      mux_data3[127:120] = in_data3[359:352];
      mux_data3[135:128] = in_data3[367:360];
      mux_data3[143:136] = in_data3[375:368];
      mux_data3[151:144] = in_data3[383:376];
      mux_data3[159:152] = in_data3[391:384];
      mux_data3[167:160] = in_data3[399:392];
      mux_data3[175:168] = in_data3[407:400];
      mux_data4[7:0] = in_data4[239:232];
      mux_data4[15:8] = in_data4[247:240];
      mux_data4[23:16] = in_data4[255:248];
      mux_data4[31:24] = in_data4[263:256];
      mux_data4[39:32] = in_data4[271:264];
      mux_data4[47:40] = in_data4[279:272];
      mux_data4[55:48] = in_data4[287:280];
      mux_data4[63:56] = in_data4[295:288];
      mux_data4[71:64] = in_data4[303:296];
      mux_data4[79:72] = in_data4[311:304];
      mux_data4[87:80] = in_data4[319:312];
      mux_data4[95:88] = in_data4[327:320];
      mux_data4[103:96] = in_data4[335:328];
      mux_data4[111:104] = in_data4[343:336];
      mux_data4[119:112] = in_data4[351:344];
      mux_data4[127:120] = in_data4[359:352];
      mux_data4[135:128] = in_data4[367:360];
      mux_data4[143:136] = in_data4[375:368];
      mux_data4[151:144] = in_data4[383:376];
      mux_data4[159:152] = in_data4[391:384];
      mux_data4[167:160] = in_data4[399:392];
      mux_data4[175:168] = in_data4[407:400];
    end
    'd3: begin
      mux_data0[7:0] = in_data0[367:360];
      mux_data0[15:8] = in_data0[375:368];
      mux_data0[23:16] = in_data0[383:376];
      mux_data0[31:24] = in_data0[391:384];
      mux_data0[39:32] = in_data0[399:392];
      mux_data0[47:40] = in_data0[407:400];
      mux_data0[55:48] = in_data0[415:408];
      mux_data0[63:56] = in_data0[423:416];
      mux_data0[71:64] = in_data0[431:424];
      mux_data0[79:72] = in_data0[439:432];
      mux_data0[87:80] = in_data0[447:440];
      mux_data0[95:88] = in_data0[455:448];
      mux_data0[103:96] = in_data0[463:456];
      mux_data0[111:104] = in_data0[471:464];
      mux_data0[119:112] = in_data0[479:472];
      mux_data0[127:120] = in_data0[487:480];
      mux_data0[135:128] = in_data0[495:488];
      mux_data0[143:136] = in_data0[503:496];
      mux_data0[151:144] = in_data0[511:504];
      mux_data0[159:152] = in_data0[519:512];
      mux_data0[167:160] = in_data0[527:520];
      mux_data0[175:168] = in_data0[535:528];
      mux_data1[7:0] = in_data1[367:360];
      mux_data1[15:8] = in_data1[375:368];
      mux_data1[23:16] = in_data1[383:376];
      mux_data1[31:24] = in_data1[391:384];
      mux_data1[39:32] = in_data1[399:392];
      mux_data1[47:40] = in_data1[407:400];
      mux_data1[55:48] = in_data1[415:408];
      mux_data1[63:56] = in_data1[423:416];
      mux_data1[71:64] = in_data1[431:424];
      mux_data1[79:72] = in_data1[439:432];
      mux_data1[87:80] = in_data1[447:440];
      mux_data1[95:88] = in_data1[455:448];
      mux_data1[103:96] = in_data1[463:456];
      mux_data1[111:104] = in_data1[471:464];
      mux_data1[119:112] = in_data1[479:472];
      mux_data1[127:120] = in_data1[487:480];
      mux_data1[135:128] = in_data1[495:488];
      mux_data1[143:136] = in_data1[503:496];
      mux_data1[151:144] = in_data1[511:504];
      mux_data1[159:152] = in_data1[519:512];
      mux_data1[167:160] = in_data1[527:520];
      mux_data1[175:168] = in_data1[535:528];
      mux_data2[7:0] = in_data2[367:360];
      mux_data2[15:8] = in_data2[375:368];
      mux_data2[23:16] = in_data2[383:376];
      mux_data2[31:24] = in_data2[391:384];
      mux_data2[39:32] = in_data2[399:392];
      mux_data2[47:40] = in_data2[407:400];
      mux_data2[55:48] = in_data2[415:408];
      mux_data2[63:56] = in_data2[423:416];
      mux_data2[71:64] = in_data2[431:424];
      mux_data2[79:72] = in_data2[439:432];
      mux_data2[87:80] = in_data2[447:440];
      mux_data2[95:88] = in_data2[455:448];
      mux_data2[103:96] = in_data2[463:456];
      mux_data2[111:104] = in_data2[471:464];
      mux_data2[119:112] = in_data2[479:472];
      mux_data2[127:120] = in_data2[487:480];
      mux_data2[135:128] = in_data2[495:488];
      mux_data2[143:136] = in_data2[503:496];
      mux_data2[151:144] = in_data2[511:504];
      mux_data2[159:152] = in_data2[519:512];
      mux_data2[167:160] = in_data2[527:520];
      mux_data2[175:168] = in_data2[535:528];
      mux_data3[7:0] = in_data3[367:360];
      mux_data3[15:8] = in_data3[375:368];
      mux_data3[23:16] = in_data3[383:376];
      mux_data3[31:24] = in_data3[391:384];
      mux_data3[39:32] = in_data3[399:392];
      mux_data3[47:40] = in_data3[407:400];
      mux_data3[55:48] = in_data3[415:408];
      mux_data3[63:56] = in_data3[423:416];
      mux_data3[71:64] = in_data3[431:424];
      mux_data3[79:72] = in_data3[439:432];
      mux_data3[87:80] = in_data3[447:440];
      mux_data3[95:88] = in_data3[455:448];
      mux_data3[103:96] = in_data3[463:456];
      mux_data3[111:104] = in_data3[471:464];
      mux_data3[119:112] = in_data3[479:472];
      mux_data3[127:120] = in_data3[487:480];
      mux_data3[135:128] = in_data3[495:488];
      mux_data3[143:136] = in_data3[503:496];
      mux_data3[151:144] = in_data3[511:504];
      mux_data3[159:152] = in_data3[519:512];
      mux_data3[167:160] = in_data3[527:520];
      mux_data3[175:168] = in_data3[535:528];
      mux_data4[7:0] = in_data4[367:360];
      mux_data4[15:8] = in_data4[375:368];
      mux_data4[23:16] = in_data4[383:376];
      mux_data4[31:24] = in_data4[391:384];
      mux_data4[39:32] = in_data4[399:392];
      mux_data4[47:40] = in_data4[407:400];
      mux_data4[55:48] = in_data4[415:408];
      mux_data4[63:56] = in_data4[423:416];
      mux_data4[71:64] = in_data4[431:424];
      mux_data4[79:72] = in_data4[439:432];
      mux_data4[87:80] = in_data4[447:440];
      mux_data4[95:88] = in_data4[455:448];
      mux_data4[103:96] = in_data4[463:456];
      mux_data4[111:104] = in_data4[471:464];
      mux_data4[119:112] = in_data4[479:472];
      mux_data4[127:120] = in_data4[487:480];
      mux_data4[135:128] = in_data4[495:488];
      mux_data4[143:136] = in_data4[503:496];
      mux_data4[151:144] = in_data4[511:504];
      mux_data4[159:152] = in_data4[519:512];
      mux_data4[167:160] = in_data4[527:520];
      mux_data4[175:168] = in_data4[535:528];
    end
    'd4: begin
      mux_data0[7:0] = in_data0[495:488];
      mux_data0[15:8] = in_data0[503:496];
      mux_data0[23:16] = in_data0[511:504];
      mux_data0[31:24] = in_data0[519:512];
      mux_data0[39:32] = in_data0[527:520];
      mux_data0[47:40] = in_data0[535:528];
      mux_data0[55:48] = in_data0[543:536];
      mux_data0[63:56] = in_data0[551:544];
      mux_data0[71:64] = in_data0[559:552];
      mux_data0[79:72] = in_data0[567:560];
      mux_data0[87:80] = in_data0[575:568];
      mux_data0[95:88] = in_data0[583:576];
      mux_data0[103:96] = in_data0[591:584];
      mux_data0[111:104] = in_data0[599:592];
      mux_data0[119:112] = in_data0[607:600];
      mux_data0[127:120] = in_data0[615:608];
      mux_data0[135:128] = in_data0[623:616];
      mux_data0[143:136] = in_data0[631:624];
      mux_data0[151:144] = in_data0[639:632];
      mux_data0[159:152] = in_data0[647:640];
      mux_data0[167:160] = in_data0[655:648];
      mux_data0[175:168] = in_data0[663:656];
      mux_data1[7:0] = in_data1[495:488];
      mux_data1[15:8] = in_data1[503:496];
      mux_data1[23:16] = in_data1[511:504];
      mux_data1[31:24] = in_data1[519:512];
      mux_data1[39:32] = in_data1[527:520];
      mux_data1[47:40] = in_data1[535:528];
      mux_data1[55:48] = in_data1[543:536];
      mux_data1[63:56] = in_data1[551:544];
      mux_data1[71:64] = in_data1[559:552];
      mux_data1[79:72] = in_data1[567:560];
      mux_data1[87:80] = in_data1[575:568];
      mux_data1[95:88] = in_data1[583:576];
      mux_data1[103:96] = in_data1[591:584];
      mux_data1[111:104] = in_data1[599:592];
      mux_data1[119:112] = in_data1[607:600];
      mux_data1[127:120] = in_data1[615:608];
      mux_data1[135:128] = in_data1[623:616];
      mux_data1[143:136] = in_data1[631:624];
      mux_data1[151:144] = in_data1[639:632];
      mux_data1[159:152] = in_data1[647:640];
      mux_data1[167:160] = in_data1[655:648];
      mux_data1[175:168] = in_data1[663:656];
      mux_data2[7:0] = in_data2[495:488];
      mux_data2[15:8] = in_data2[503:496];
      mux_data2[23:16] = in_data2[511:504];
      mux_data2[31:24] = in_data2[519:512];
      mux_data2[39:32] = in_data2[527:520];
      mux_data2[47:40] = in_data2[535:528];
      mux_data2[55:48] = in_data2[543:536];
      mux_data2[63:56] = in_data2[551:544];
      mux_data2[71:64] = in_data2[559:552];
      mux_data2[79:72] = in_data2[567:560];
      mux_data2[87:80] = in_data2[575:568];
      mux_data2[95:88] = in_data2[583:576];
      mux_data2[103:96] = in_data2[591:584];
      mux_data2[111:104] = in_data2[599:592];
      mux_data2[119:112] = in_data2[607:600];
      mux_data2[127:120] = in_data2[615:608];
      mux_data2[135:128] = in_data2[623:616];
      mux_data2[143:136] = in_data2[631:624];
      mux_data2[151:144] = in_data2[639:632];
      mux_data2[159:152] = in_data2[647:640];
      mux_data2[167:160] = in_data2[655:648];
      mux_data2[175:168] = in_data2[663:656];
      mux_data3[7:0] = in_data3[495:488];
      mux_data3[15:8] = in_data3[503:496];
      mux_data3[23:16] = in_data3[511:504];
      mux_data3[31:24] = in_data3[519:512];
      mux_data3[39:32] = in_data3[527:520];
      mux_data3[47:40] = in_data3[535:528];
      mux_data3[55:48] = in_data3[543:536];
      mux_data3[63:56] = in_data3[551:544];
      mux_data3[71:64] = in_data3[559:552];
      mux_data3[79:72] = in_data3[567:560];
      mux_data3[87:80] = in_data3[575:568];
      mux_data3[95:88] = in_data3[583:576];
      mux_data3[103:96] = in_data3[591:584];
      mux_data3[111:104] = in_data3[599:592];
      mux_data3[119:112] = in_data3[607:600];
      mux_data3[127:120] = in_data3[615:608];
      mux_data3[135:128] = in_data3[623:616];
      mux_data3[143:136] = in_data3[631:624];
      mux_data3[151:144] = in_data3[639:632];
      mux_data3[159:152] = in_data3[647:640];
      mux_data3[167:160] = in_data3[655:648];
      mux_data3[175:168] = in_data3[663:656];
      mux_data4[7:0] = in_data4[495:488];
      mux_data4[15:8] = in_data4[503:496];
      mux_data4[23:16] = in_data4[511:504];
      mux_data4[31:24] = in_data4[519:512];
      mux_data4[39:32] = in_data4[527:520];
      mux_data4[47:40] = in_data4[535:528];
      mux_data4[55:48] = in_data4[543:536];
      mux_data4[63:56] = in_data4[551:544];
      mux_data4[71:64] = in_data4[559:552];
      mux_data4[79:72] = in_data4[567:560];
      mux_data4[87:80] = in_data4[575:568];
      mux_data4[95:88] = in_data4[583:576];
      mux_data4[103:96] = in_data4[591:584];
      mux_data4[111:104] = in_data4[599:592];
      mux_data4[119:112] = in_data4[607:600];
      mux_data4[127:120] = in_data4[615:608];
      mux_data4[135:128] = in_data4[623:616];
      mux_data4[143:136] = in_data4[631:624];
      mux_data4[151:144] = in_data4[639:632];
      mux_data4[159:152] = in_data4[647:640];
      mux_data4[167:160] = in_data4[655:648];
      mux_data4[175:168] = in_data4[663:656];
    end
    'd5: begin
      mux_data0[7:0] = in_data0[623:616];
      mux_data0[15:8] = in_data0[631:624];
      mux_data0[23:16] = in_data0[639:632];
      mux_data0[31:24] = in_data0[647:640];
      mux_data0[39:32] = in_data0[655:648];
      mux_data0[47:40] = in_data0[663:656];
      mux_data0[55:48] = in_data0[671:664];
      mux_data0[63:56] = in_data0[679:672];
      mux_data0[71:64] = in_data0[687:680];
      mux_data0[79:72] = in_data0[695:688];
      mux_data0[87:80] = in_data0[703:696];
      mux_data0[95:88] = in_data0[711:704];
      mux_data0[103:96] = in_data0[719:712];
      mux_data0[111:104] = in_data0[727:720];
      mux_data0[119:112] = in_data0[735:728];
      mux_data0[127:120] = in_data0[743:736];
      mux_data0[135:128] = in_data0[751:744];
      mux_data0[143:136] = in_data0[759:752];
      mux_data0[151:144] = in_data0[767:760];
      mux_data0[159:152] = in_data0[775:768];
      mux_data0[167:160] = in_data0[783:776];
      mux_data0[175:168] = in_data0[791:784];
      mux_data1[7:0] = in_data1[623:616];
      mux_data1[15:8] = in_data1[631:624];
      mux_data1[23:16] = in_data1[639:632];
      mux_data1[31:24] = in_data1[647:640];
      mux_data1[39:32] = in_data1[655:648];
      mux_data1[47:40] = in_data1[663:656];
      mux_data1[55:48] = in_data1[671:664];
      mux_data1[63:56] = in_data1[679:672];
      mux_data1[71:64] = in_data1[687:680];
      mux_data1[79:72] = in_data1[695:688];
      mux_data1[87:80] = in_data1[703:696];
      mux_data1[95:88] = in_data1[711:704];
      mux_data1[103:96] = in_data1[719:712];
      mux_data1[111:104] = in_data1[727:720];
      mux_data1[119:112] = in_data1[735:728];
      mux_data1[127:120] = in_data1[743:736];
      mux_data1[135:128] = in_data1[751:744];
      mux_data1[143:136] = in_data1[759:752];
      mux_data1[151:144] = in_data1[767:760];
      mux_data1[159:152] = in_data1[775:768];
      mux_data1[167:160] = in_data1[783:776];
      mux_data1[175:168] = in_data1[791:784];
      mux_data2[7:0] = in_data2[623:616];
      mux_data2[15:8] = in_data2[631:624];
      mux_data2[23:16] = in_data2[639:632];
      mux_data2[31:24] = in_data2[647:640];
      mux_data2[39:32] = in_data2[655:648];
      mux_data2[47:40] = in_data2[663:656];
      mux_data2[55:48] = in_data2[671:664];
      mux_data2[63:56] = in_data2[679:672];
      mux_data2[71:64] = in_data2[687:680];
      mux_data2[79:72] = in_data2[695:688];
      mux_data2[87:80] = in_data2[703:696];
      mux_data2[95:88] = in_data2[711:704];
      mux_data2[103:96] = in_data2[719:712];
      mux_data2[111:104] = in_data2[727:720];
      mux_data2[119:112] = in_data2[735:728];
      mux_data2[127:120] = in_data2[743:736];
      mux_data2[135:128] = in_data2[751:744];
      mux_data2[143:136] = in_data2[759:752];
      mux_data2[151:144] = in_data2[767:760];
      mux_data2[159:152] = in_data2[775:768];
      mux_data2[167:160] = in_data2[783:776];
      mux_data2[175:168] = in_data2[791:784];
      mux_data3[7:0] = in_data3[623:616];
      mux_data3[15:8] = in_data3[631:624];
      mux_data3[23:16] = in_data3[639:632];
      mux_data3[31:24] = in_data3[647:640];
      mux_data3[39:32] = in_data3[655:648];
      mux_data3[47:40] = in_data3[663:656];
      mux_data3[55:48] = in_data3[671:664];
      mux_data3[63:56] = in_data3[679:672];
      mux_data3[71:64] = in_data3[687:680];
      mux_data3[79:72] = in_data3[695:688];
      mux_data3[87:80] = in_data3[703:696];
      mux_data3[95:88] = in_data3[711:704];
      mux_data3[103:96] = in_data3[719:712];
      mux_data3[111:104] = in_data3[727:720];
      mux_data3[119:112] = in_data3[735:728];
      mux_data3[127:120] = in_data3[743:736];
      mux_data3[135:128] = in_data3[751:744];
      mux_data3[143:136] = in_data3[759:752];
      mux_data3[151:144] = in_data3[767:760];
      mux_data3[159:152] = in_data3[775:768];
      mux_data3[167:160] = in_data3[783:776];
      mux_data3[175:168] = in_data3[791:784];
      mux_data4[7:0] = in_data4[623:616];
      mux_data4[15:8] = in_data4[631:624];
      mux_data4[23:16] = in_data4[639:632];
      mux_data4[31:24] = in_data4[647:640];
      mux_data4[39:32] = in_data4[655:648];
      mux_data4[47:40] = in_data4[663:656];
      mux_data4[55:48] = in_data4[671:664];
      mux_data4[63:56] = in_data4[679:672];
      mux_data4[71:64] = in_data4[687:680];
      mux_data4[79:72] = in_data4[695:688];
      mux_data4[87:80] = in_data4[703:696];
      mux_data4[95:88] = in_data4[711:704];
      mux_data4[103:96] = in_data4[719:712];
      mux_data4[111:104] = in_data4[727:720];
      mux_data4[119:112] = in_data4[735:728];
      mux_data4[127:120] = in_data4[743:736];
      mux_data4[135:128] = in_data4[751:744];
      mux_data4[143:136] = in_data4[759:752];
      mux_data4[151:144] = in_data4[767:760];
      mux_data4[159:152] = in_data4[775:768];
      mux_data4[167:160] = in_data4[783:776];
      mux_data4[175:168] = in_data4[791:784];
    end
    'd6: begin
      mux_data0[7:0] = in_data0[751:744];
      mux_data0[15:8] = in_data0[759:752];
      mux_data0[23:16] = in_data0[767:760];
      mux_data0[31:24] = in_data0[775:768];
      mux_data0[39:32] = in_data0[783:776];
      mux_data0[47:40] = in_data0[791:784];
      mux_data0[55:48] = in_data0[799:792];
      mux_data0[63:56] = in_data0[807:800];
      mux_data0[71:64] = in_data0[815:808];
      mux_data0[79:72] = in_data0[823:816];
      mux_data0[87:80] = in_data0[831:824];
      mux_data0[95:88] = in_data0[839:832];
      mux_data0[103:96] = in_data0[847:840];
      mux_data0[111:104] = in_data0[855:848];
      mux_data0[119:112] = in_data0[863:856];
      mux_data0[127:120] = in_data0[871:864];
      mux_data0[135:128] = in_data0[879:872];
      mux_data0[143:136] = in_data0[887:880];
      mux_data0[151:144] = in_data0[895:888];
      mux_data0[159:152] = in_data0[903:896];
      mux_data0[167:160] = in_data0[911:904];
      mux_data0[175:168] = in_data0[919:912];
      mux_data1[7:0] = in_data1[751:744];
      mux_data1[15:8] = in_data1[759:752];
      mux_data1[23:16] = in_data1[767:760];
      mux_data1[31:24] = in_data1[775:768];
      mux_data1[39:32] = in_data1[783:776];
      mux_data1[47:40] = in_data1[791:784];
      mux_data1[55:48] = in_data1[799:792];
      mux_data1[63:56] = in_data1[807:800];
      mux_data1[71:64] = in_data1[815:808];
      mux_data1[79:72] = in_data1[823:816];
      mux_data1[87:80] = in_data1[831:824];
      mux_data1[95:88] = in_data1[839:832];
      mux_data1[103:96] = in_data1[847:840];
      mux_data1[111:104] = in_data1[855:848];
      mux_data1[119:112] = in_data1[863:856];
      mux_data1[127:120] = in_data1[871:864];
      mux_data1[135:128] = in_data1[879:872];
      mux_data1[143:136] = in_data1[887:880];
      mux_data1[151:144] = in_data1[895:888];
      mux_data1[159:152] = in_data1[903:896];
      mux_data1[167:160] = in_data1[911:904];
      mux_data1[175:168] = in_data1[919:912];
      mux_data2[7:0] = in_data2[751:744];
      mux_data2[15:8] = in_data2[759:752];
      mux_data2[23:16] = in_data2[767:760];
      mux_data2[31:24] = in_data2[775:768];
      mux_data2[39:32] = in_data2[783:776];
      mux_data2[47:40] = in_data2[791:784];
      mux_data2[55:48] = in_data2[799:792];
      mux_data2[63:56] = in_data2[807:800];
      mux_data2[71:64] = in_data2[815:808];
      mux_data2[79:72] = in_data2[823:816];
      mux_data2[87:80] = in_data2[831:824];
      mux_data2[95:88] = in_data2[839:832];
      mux_data2[103:96] = in_data2[847:840];
      mux_data2[111:104] = in_data2[855:848];
      mux_data2[119:112] = in_data2[863:856];
      mux_data2[127:120] = in_data2[871:864];
      mux_data2[135:128] = in_data2[879:872];
      mux_data2[143:136] = in_data2[887:880];
      mux_data2[151:144] = in_data2[895:888];
      mux_data2[159:152] = in_data2[903:896];
      mux_data2[167:160] = in_data2[911:904];
      mux_data2[175:168] = in_data2[919:912];
      mux_data3[7:0] = in_data3[751:744];
      mux_data3[15:8] = in_data3[759:752];
      mux_data3[23:16] = in_data3[767:760];
      mux_data3[31:24] = in_data3[775:768];
      mux_data3[39:32] = in_data3[783:776];
      mux_data3[47:40] = in_data3[791:784];
      mux_data3[55:48] = in_data3[799:792];
      mux_data3[63:56] = in_data3[807:800];
      mux_data3[71:64] = in_data3[815:808];
      mux_data3[79:72] = in_data3[823:816];
      mux_data3[87:80] = in_data3[831:824];
      mux_data3[95:88] = in_data3[839:832];
      mux_data3[103:96] = in_data3[847:840];
      mux_data3[111:104] = in_data3[855:848];
      mux_data3[119:112] = in_data3[863:856];
      mux_data3[127:120] = in_data3[871:864];
      mux_data3[135:128] = in_data3[879:872];
      mux_data3[143:136] = in_data3[887:880];
      mux_data3[151:144] = in_data3[895:888];
      mux_data3[159:152] = in_data3[903:896];
      mux_data3[167:160] = in_data3[911:904];
      mux_data3[175:168] = in_data3[919:912];
      mux_data4[7:0] = in_data4[751:744];
      mux_data4[15:8] = in_data4[759:752];
      mux_data4[23:16] = in_data4[767:760];
      mux_data4[31:24] = in_data4[775:768];
      mux_data4[39:32] = in_data4[783:776];
      mux_data4[47:40] = in_data4[791:784];
      mux_data4[55:48] = in_data4[799:792];
      mux_data4[63:56] = in_data4[807:800];
      mux_data4[71:64] = in_data4[815:808];
      mux_data4[79:72] = in_data4[823:816];
      mux_data4[87:80] = in_data4[831:824];
      mux_data4[95:88] = in_data4[839:832];
      mux_data4[103:96] = in_data4[847:840];
      mux_data4[111:104] = in_data4[855:848];
      mux_data4[119:112] = in_data4[863:856];
      mux_data4[127:120] = in_data4[871:864];
      mux_data4[135:128] = in_data4[879:872];
      mux_data4[143:136] = in_data4[887:880];
      mux_data4[151:144] = in_data4[895:888];
      mux_data4[159:152] = in_data4[903:896];
      mux_data4[167:160] = in_data4[911:904];
      mux_data4[175:168] = in_data4[919:912];
    end
    'd7: begin
      mux_data0[7:0] = in_data0[879:872];
      mux_data0[15:8] = in_data0[887:880];
      mux_data0[23:16] = in_data0[895:888];
      mux_data0[31:24] = in_data0[903:896];
      mux_data0[39:32] = in_data0[911:904];
      mux_data0[47:40] = in_data0[919:912];
      mux_data0[55:48] = in_data0[927:920];
      mux_data0[63:56] = in_data0[935:928];
      mux_data0[71:64] = in_data0[943:936];
      mux_data0[79:72] = in_data0[951:944];
      mux_data0[87:80] = in_data0[959:952];
      mux_data0[95:88] = in_data0[967:960];
      mux_data0[103:96] = in_data0[975:968];
      mux_data0[111:104] = in_data0[983:976];
      mux_data0[119:112] = in_data0[991:984];
      mux_data0[127:120] = in_data0[999:992];
      mux_data0[135:128] = in_data0[1007:1000];
      mux_data0[143:136] = in_data0[1015:1008];
      mux_data0[151:144] = in_data0[1023:1016];
      mux_data0[159:152] = in_data0[1031:1024];
      mux_data0[167:160] = in_data0[1039:1032];
      mux_data0[175:168] = in_data0[1047:1040];
      mux_data1[7:0] = in_data1[879:872];
      mux_data1[15:8] = in_data1[887:880];
      mux_data1[23:16] = in_data1[895:888];
      mux_data1[31:24] = in_data1[903:896];
      mux_data1[39:32] = in_data1[911:904];
      mux_data1[47:40] = in_data1[919:912];
      mux_data1[55:48] = in_data1[927:920];
      mux_data1[63:56] = in_data1[935:928];
      mux_data1[71:64] = in_data1[943:936];
      mux_data1[79:72] = in_data1[951:944];
      mux_data1[87:80] = in_data1[959:952];
      mux_data1[95:88] = in_data1[967:960];
      mux_data1[103:96] = in_data1[975:968];
      mux_data1[111:104] = in_data1[983:976];
      mux_data1[119:112] = in_data1[991:984];
      mux_data1[127:120] = in_data1[999:992];
      mux_data1[135:128] = in_data1[1007:1000];
      mux_data1[143:136] = in_data1[1015:1008];
      mux_data1[151:144] = in_data1[1023:1016];
      mux_data1[159:152] = in_data1[1031:1024];
      mux_data1[167:160] = in_data1[1039:1032];
      mux_data1[175:168] = in_data1[1047:1040];
      mux_data2[7:0] = in_data2[879:872];
      mux_data2[15:8] = in_data2[887:880];
      mux_data2[23:16] = in_data2[895:888];
      mux_data2[31:24] = in_data2[903:896];
      mux_data2[39:32] = in_data2[911:904];
      mux_data2[47:40] = in_data2[919:912];
      mux_data2[55:48] = in_data2[927:920];
      mux_data2[63:56] = in_data2[935:928];
      mux_data2[71:64] = in_data2[943:936];
      mux_data2[79:72] = in_data2[951:944];
      mux_data2[87:80] = in_data2[959:952];
      mux_data2[95:88] = in_data2[967:960];
      mux_data2[103:96] = in_data2[975:968];
      mux_data2[111:104] = in_data2[983:976];
      mux_data2[119:112] = in_data2[991:984];
      mux_data2[127:120] = in_data2[999:992];
      mux_data2[135:128] = in_data2[1007:1000];
      mux_data2[143:136] = in_data2[1015:1008];
      mux_data2[151:144] = in_data2[1023:1016];
      mux_data2[159:152] = in_data2[1031:1024];
      mux_data2[167:160] = in_data2[1039:1032];
      mux_data2[175:168] = in_data2[1047:1040];
      mux_data3[7:0] = in_data3[879:872];
      mux_data3[15:8] = in_data3[887:880];
      mux_data3[23:16] = in_data3[895:888];
      mux_data3[31:24] = in_data3[903:896];
      mux_data3[39:32] = in_data3[911:904];
      mux_data3[47:40] = in_data3[919:912];
      mux_data3[55:48] = in_data3[927:920];
      mux_data3[63:56] = in_data3[935:928];
      mux_data3[71:64] = in_data3[943:936];
      mux_data3[79:72] = in_data3[951:944];
      mux_data3[87:80] = in_data3[959:952];
      mux_data3[95:88] = in_data3[967:960];
      mux_data3[103:96] = in_data3[975:968];
      mux_data3[111:104] = in_data3[983:976];
      mux_data3[119:112] = in_data3[991:984];
      mux_data3[127:120] = in_data3[999:992];
      mux_data3[135:128] = in_data3[1007:1000];
      mux_data3[143:136] = in_data3[1015:1008];
      mux_data3[151:144] = in_data3[1023:1016];
      mux_data3[159:152] = in_data3[1031:1024];
      mux_data3[167:160] = in_data3[1039:1032];
      mux_data3[175:168] = in_data3[1047:1040];
      mux_data4[7:0] = in_data4[879:872];
      mux_data4[15:8] = in_data4[887:880];
      mux_data4[23:16] = in_data4[895:888];
      mux_data4[31:24] = in_data4[903:896];
      mux_data4[39:32] = in_data4[911:904];
      mux_data4[47:40] = in_data4[919:912];
      mux_data4[55:48] = in_data4[927:920];
      mux_data4[63:56] = in_data4[935:928];
      mux_data4[71:64] = in_data4[943:936];
      mux_data4[79:72] = in_data4[951:944];
      mux_data4[87:80] = in_data4[959:952];
      mux_data4[95:88] = in_data4[967:960];
      mux_data4[103:96] = in_data4[975:968];
      mux_data4[111:104] = in_data4[983:976];
      mux_data4[119:112] = in_data4[991:984];
      mux_data4[127:120] = in_data4[999:992];
      mux_data4[135:128] = in_data4[1007:1000];
      mux_data4[143:136] = in_data4[1015:1008];
      mux_data4[151:144] = in_data4[1023:1016];
      mux_data4[159:152] = in_data4[1031:1024];
      mux_data4[167:160] = in_data4[1039:1032];
      mux_data4[175:168] = in_data4[1047:1040];
    end
    'd8: begin
      mux_data0[7:0] = in_data0[1007:1000];
      mux_data0[15:8] = in_data0[1015:1008];
      mux_data0[23:16] = in_data0[1023:1016];
      mux_data0[31:24] = in_data0[1031:1024];
      mux_data0[39:32] = in_data0[1039:1032];
      mux_data0[47:40] = in_data0[1047:1040];
      mux_data0[55:48] = in_data0[1055:1048];
      mux_data0[63:56] = in_data0[1063:1056];
      mux_data0[71:64] = in_data0[1071:1064];
      mux_data0[79:72] = in_data0[1079:1072];
      mux_data0[87:80] = in_data0[1087:1080];
      mux_data0[95:88] = in_data0[1095:1088];
      mux_data0[103:96] = in_data0[1103:1096];
      mux_data0[111:104] = in_data0[1111:1104];
      mux_data0[119:112] = in_data0[1119:1112];
      mux_data0[127:120] = in_data0[1127:1120];
      mux_data0[135:128] = in_data0[1135:1128];
      mux_data0[143:136] = in_data0[1143:1136];
      mux_data0[151:144] = in_data0[1151:1144];
      mux_data0[159:152] = in_data0[1159:1152];
      mux_data0[167:160] = in_data0[1167:1160];
      mux_data0[175:168] = in_data0[1175:1168];
      mux_data1[7:0] = in_data1[1007:1000];
      mux_data1[15:8] = in_data1[1015:1008];
      mux_data1[23:16] = in_data1[1023:1016];
      mux_data1[31:24] = in_data1[1031:1024];
      mux_data1[39:32] = in_data1[1039:1032];
      mux_data1[47:40] = in_data1[1047:1040];
      mux_data1[55:48] = in_data1[1055:1048];
      mux_data1[63:56] = in_data1[1063:1056];
      mux_data1[71:64] = in_data1[1071:1064];
      mux_data1[79:72] = in_data1[1079:1072];
      mux_data1[87:80] = in_data1[1087:1080];
      mux_data1[95:88] = in_data1[1095:1088];
      mux_data1[103:96] = in_data1[1103:1096];
      mux_data1[111:104] = in_data1[1111:1104];
      mux_data1[119:112] = in_data1[1119:1112];
      mux_data1[127:120] = in_data1[1127:1120];
      mux_data1[135:128] = in_data1[1135:1128];
      mux_data1[143:136] = in_data1[1143:1136];
      mux_data1[151:144] = in_data1[1151:1144];
      mux_data1[159:152] = in_data1[1159:1152];
      mux_data1[167:160] = in_data1[1167:1160];
      mux_data1[175:168] = in_data1[1175:1168];
      mux_data2[7:0] = in_data2[1007:1000];
      mux_data2[15:8] = in_data2[1015:1008];
      mux_data2[23:16] = in_data2[1023:1016];
      mux_data2[31:24] = in_data2[1031:1024];
      mux_data2[39:32] = in_data2[1039:1032];
      mux_data2[47:40] = in_data2[1047:1040];
      mux_data2[55:48] = in_data2[1055:1048];
      mux_data2[63:56] = in_data2[1063:1056];
      mux_data2[71:64] = in_data2[1071:1064];
      mux_data2[79:72] = in_data2[1079:1072];
      mux_data2[87:80] = in_data2[1087:1080];
      mux_data2[95:88] = in_data2[1095:1088];
      mux_data2[103:96] = in_data2[1103:1096];
      mux_data2[111:104] = in_data2[1111:1104];
      mux_data2[119:112] = in_data2[1119:1112];
      mux_data2[127:120] = in_data2[1127:1120];
      mux_data2[135:128] = in_data2[1135:1128];
      mux_data2[143:136] = in_data2[1143:1136];
      mux_data2[151:144] = in_data2[1151:1144];
      mux_data2[159:152] = in_data2[1159:1152];
      mux_data2[167:160] = in_data2[1167:1160];
      mux_data2[175:168] = in_data2[1175:1168];
      mux_data3[7:0] = in_data3[1007:1000];
      mux_data3[15:8] = in_data3[1015:1008];
      mux_data3[23:16] = in_data3[1023:1016];
      mux_data3[31:24] = in_data3[1031:1024];
      mux_data3[39:32] = in_data3[1039:1032];
      mux_data3[47:40] = in_data3[1047:1040];
      mux_data3[55:48] = in_data3[1055:1048];
      mux_data3[63:56] = in_data3[1063:1056];
      mux_data3[71:64] = in_data3[1071:1064];
      mux_data3[79:72] = in_data3[1079:1072];
      mux_data3[87:80] = in_data3[1087:1080];
      mux_data3[95:88] = in_data3[1095:1088];
      mux_data3[103:96] = in_data3[1103:1096];
      mux_data3[111:104] = in_data3[1111:1104];
      mux_data3[119:112] = in_data3[1119:1112];
      mux_data3[127:120] = in_data3[1127:1120];
      mux_data3[135:128] = in_data3[1135:1128];
      mux_data3[143:136] = in_data3[1143:1136];
      mux_data3[151:144] = in_data3[1151:1144];
      mux_data3[159:152] = in_data3[1159:1152];
      mux_data3[167:160] = in_data3[1167:1160];
      mux_data3[175:168] = in_data3[1175:1168];
      mux_data4[7:0] = in_data4[1007:1000];
      mux_data4[15:8] = in_data4[1015:1008];
      mux_data4[23:16] = in_data4[1023:1016];
      mux_data4[31:24] = in_data4[1031:1024];
      mux_data4[39:32] = in_data4[1039:1032];
      mux_data4[47:40] = in_data4[1047:1040];
      mux_data4[55:48] = in_data4[1055:1048];
      mux_data4[63:56] = in_data4[1063:1056];
      mux_data4[71:64] = in_data4[1071:1064];
      mux_data4[79:72] = in_data4[1079:1072];
      mux_data4[87:80] = in_data4[1087:1080];
      mux_data4[95:88] = in_data4[1095:1088];
      mux_data4[103:96] = in_data4[1103:1096];
      mux_data4[111:104] = in_data4[1111:1104];
      mux_data4[119:112] = in_data4[1119:1112];
      mux_data4[127:120] = in_data4[1127:1120];
      mux_data4[135:128] = in_data4[1135:1128];
      mux_data4[143:136] = in_data4[1143:1136];
      mux_data4[151:144] = in_data4[1151:1144];
      mux_data4[159:152] = in_data4[1159:1152];
      mux_data4[167:160] = in_data4[1167:1160];
      mux_data4[175:168] = in_data4[1175:1168];
    end
    'd9: begin
      mux_data0[7:0] = in_data0[1135:1128];
      mux_data0[15:8] = in_data0[1143:1136];
      mux_data0[23:16] = in_data0[1151:1144];
      mux_data0[31:24] = in_data0[1159:1152];
      mux_data0[39:32] = in_data0[1167:1160];
      mux_data0[47:40] = in_data0[1175:1168];
      mux_data0[55:48] = in_data0[1183:1176];
      mux_data0[63:56] = in_data0[1191:1184];
      mux_data0[71:64] = in_data0[1199:1192];
      mux_data0[79:72] = in_data0[1207:1200];
      mux_data0[87:80] = in_data0[1215:1208];
      mux_data0[95:88] = in_data0[1223:1216];
      mux_data0[103:96] = in_data0[1231:1224];
      mux_data0[111:104] = in_data0[1239:1232];
      mux_data0[119:112] = in_data0[1247:1240];
      mux_data0[127:120] = in_data0[1255:1248];
      mux_data0[135:128] = in_data0[1263:1256];
      mux_data0[143:136] = in_data0[1271:1264];
      mux_data0[151:144] = in_data0[1279:1272];
      mux_data0[159:152] = in_data0[1287:1280];
      mux_data0[167:160] = in_data0[1295:1288];
      mux_data0[175:168] = in_data0[1303:1296];
      mux_data1[7:0] = in_data1[1135:1128];
      mux_data1[15:8] = in_data1[1143:1136];
      mux_data1[23:16] = in_data1[1151:1144];
      mux_data1[31:24] = in_data1[1159:1152];
      mux_data1[39:32] = in_data1[1167:1160];
      mux_data1[47:40] = in_data1[1175:1168];
      mux_data1[55:48] = in_data1[1183:1176];
      mux_data1[63:56] = in_data1[1191:1184];
      mux_data1[71:64] = in_data1[1199:1192];
      mux_data1[79:72] = in_data1[1207:1200];
      mux_data1[87:80] = in_data1[1215:1208];
      mux_data1[95:88] = in_data1[1223:1216];
      mux_data1[103:96] = in_data1[1231:1224];
      mux_data1[111:104] = in_data1[1239:1232];
      mux_data1[119:112] = in_data1[1247:1240];
      mux_data1[127:120] = in_data1[1255:1248];
      mux_data1[135:128] = in_data1[1263:1256];
      mux_data1[143:136] = in_data1[1271:1264];
      mux_data1[151:144] = in_data1[1279:1272];
      mux_data1[159:152] = in_data1[1287:1280];
      mux_data1[167:160] = in_data1[1295:1288];
      mux_data1[175:168] = in_data1[1303:1296];
      mux_data2[7:0] = in_data2[1135:1128];
      mux_data2[15:8] = in_data2[1143:1136];
      mux_data2[23:16] = in_data2[1151:1144];
      mux_data2[31:24] = in_data2[1159:1152];
      mux_data2[39:32] = in_data2[1167:1160];
      mux_data2[47:40] = in_data2[1175:1168];
      mux_data2[55:48] = in_data2[1183:1176];
      mux_data2[63:56] = in_data2[1191:1184];
      mux_data2[71:64] = in_data2[1199:1192];
      mux_data2[79:72] = in_data2[1207:1200];
      mux_data2[87:80] = in_data2[1215:1208];
      mux_data2[95:88] = in_data2[1223:1216];
      mux_data2[103:96] = in_data2[1231:1224];
      mux_data2[111:104] = in_data2[1239:1232];
      mux_data2[119:112] = in_data2[1247:1240];
      mux_data2[127:120] = in_data2[1255:1248];
      mux_data2[135:128] = in_data2[1263:1256];
      mux_data2[143:136] = in_data2[1271:1264];
      mux_data2[151:144] = in_data2[1279:1272];
      mux_data2[159:152] = in_data2[1287:1280];
      mux_data2[167:160] = in_data2[1295:1288];
      mux_data2[175:168] = in_data2[1303:1296];
      mux_data3[7:0] = in_data3[1135:1128];
      mux_data3[15:8] = in_data3[1143:1136];
      mux_data3[23:16] = in_data3[1151:1144];
      mux_data3[31:24] = in_data3[1159:1152];
      mux_data3[39:32] = in_data3[1167:1160];
      mux_data3[47:40] = in_data3[1175:1168];
      mux_data3[55:48] = in_data3[1183:1176];
      mux_data3[63:56] = in_data3[1191:1184];
      mux_data3[71:64] = in_data3[1199:1192];
      mux_data3[79:72] = in_data3[1207:1200];
      mux_data3[87:80] = in_data3[1215:1208];
      mux_data3[95:88] = in_data3[1223:1216];
      mux_data3[103:96] = in_data3[1231:1224];
      mux_data3[111:104] = in_data3[1239:1232];
      mux_data3[119:112] = in_data3[1247:1240];
      mux_data3[127:120] = in_data3[1255:1248];
      mux_data3[135:128] = in_data3[1263:1256];
      mux_data3[143:136] = in_data3[1271:1264];
      mux_data3[151:144] = in_data3[1279:1272];
      mux_data3[159:152] = in_data3[1287:1280];
      mux_data3[167:160] = in_data3[1295:1288];
      mux_data3[175:168] = in_data3[1303:1296];
      mux_data4[7:0] = in_data4[1135:1128];
      mux_data4[15:8] = in_data4[1143:1136];
      mux_data4[23:16] = in_data4[1151:1144];
      mux_data4[31:24] = in_data4[1159:1152];
      mux_data4[39:32] = in_data4[1167:1160];
      mux_data4[47:40] = in_data4[1175:1168];
      mux_data4[55:48] = in_data4[1183:1176];
      mux_data4[63:56] = in_data4[1191:1184];
      mux_data4[71:64] = in_data4[1199:1192];
      mux_data4[79:72] = in_data4[1207:1200];
      mux_data4[87:80] = in_data4[1215:1208];
      mux_data4[95:88] = in_data4[1223:1216];
      mux_data4[103:96] = in_data4[1231:1224];
      mux_data4[111:104] = in_data4[1239:1232];
      mux_data4[119:112] = in_data4[1247:1240];
      mux_data4[127:120] = in_data4[1255:1248];
      mux_data4[135:128] = in_data4[1263:1256];
      mux_data4[143:136] = in_data4[1271:1264];
      mux_data4[151:144] = in_data4[1279:1272];
      mux_data4[159:152] = in_data4[1287:1280];
      mux_data4[167:160] = in_data4[1295:1288];
      mux_data4[175:168] = in_data4[1303:1296];
    end
    'd10: begin
      mux_data0[7:0] = in_data0[1263:1256];
      mux_data0[15:8] = in_data0[1271:1264];
      mux_data0[23:16] = in_data0[1279:1272];
      mux_data0[31:24] = in_data0[1287:1280];
      mux_data0[39:32] = in_data0[1295:1288];
      mux_data0[47:40] = in_data0[1303:1296];
      mux_data0[55:48] = in_data0[1311:1304];
      mux_data0[63:56] = in_data0[1319:1312];
      mux_data0[71:64] = in_data0[1327:1320];
      mux_data0[79:72] = in_data0[1335:1328];
      mux_data0[87:80] = in_data0[1343:1336];
      mux_data0[95:88] = in_data0[1351:1344];
      mux_data0[103:96] = in_data0[1359:1352];
      mux_data0[111:104] = in_data0[1367:1360];
      mux_data0[119:112] = in_data0[1375:1368];
      mux_data0[127:120] = in_data0[1383:1376];
      mux_data0[135:128] = in_data0[1391:1384];
      mux_data0[143:136] = in_data0[1399:1392];
      mux_data0[151:144] = in_data0[1407:1400];
      mux_data0[159:152] = in_data0[1415:1408];
      mux_data0[167:160] = in_data0[1423:1416];
      mux_data0[175:168] = in_data0[1431:1424];
      mux_data1[7:0] = in_data1[1263:1256];
      mux_data1[15:8] = in_data1[1271:1264];
      mux_data1[23:16] = in_data1[1279:1272];
      mux_data1[31:24] = in_data1[1287:1280];
      mux_data1[39:32] = in_data1[1295:1288];
      mux_data1[47:40] = in_data1[1303:1296];
      mux_data1[55:48] = in_data1[1311:1304];
      mux_data1[63:56] = in_data1[1319:1312];
      mux_data1[71:64] = in_data1[1327:1320];
      mux_data1[79:72] = in_data1[1335:1328];
      mux_data1[87:80] = in_data1[1343:1336];
      mux_data1[95:88] = in_data1[1351:1344];
      mux_data1[103:96] = in_data1[1359:1352];
      mux_data1[111:104] = in_data1[1367:1360];
      mux_data1[119:112] = in_data1[1375:1368];
      mux_data1[127:120] = in_data1[1383:1376];
      mux_data1[135:128] = in_data1[1391:1384];
      mux_data1[143:136] = in_data1[1399:1392];
      mux_data1[151:144] = in_data1[1407:1400];
      mux_data1[159:152] = in_data1[1415:1408];
      mux_data1[167:160] = in_data1[1423:1416];
      mux_data1[175:168] = in_data1[1431:1424];
      mux_data2[7:0] = in_data2[1263:1256];
      mux_data2[15:8] = in_data2[1271:1264];
      mux_data2[23:16] = in_data2[1279:1272];
      mux_data2[31:24] = in_data2[1287:1280];
      mux_data2[39:32] = in_data2[1295:1288];
      mux_data2[47:40] = in_data2[1303:1296];
      mux_data2[55:48] = in_data2[1311:1304];
      mux_data2[63:56] = in_data2[1319:1312];
      mux_data2[71:64] = in_data2[1327:1320];
      mux_data2[79:72] = in_data2[1335:1328];
      mux_data2[87:80] = in_data2[1343:1336];
      mux_data2[95:88] = in_data2[1351:1344];
      mux_data2[103:96] = in_data2[1359:1352];
      mux_data2[111:104] = in_data2[1367:1360];
      mux_data2[119:112] = in_data2[1375:1368];
      mux_data2[127:120] = in_data2[1383:1376];
      mux_data2[135:128] = in_data2[1391:1384];
      mux_data2[143:136] = in_data2[1399:1392];
      mux_data2[151:144] = in_data2[1407:1400];
      mux_data2[159:152] = in_data2[1415:1408];
      mux_data2[167:160] = in_data2[1423:1416];
      mux_data2[175:168] = in_data2[1431:1424];
      mux_data3[7:0] = in_data3[1263:1256];
      mux_data3[15:8] = in_data3[1271:1264];
      mux_data3[23:16] = in_data3[1279:1272];
      mux_data3[31:24] = in_data3[1287:1280];
      mux_data3[39:32] = in_data3[1295:1288];
      mux_data3[47:40] = in_data3[1303:1296];
      mux_data3[55:48] = in_data3[1311:1304];
      mux_data3[63:56] = in_data3[1319:1312];
      mux_data3[71:64] = in_data3[1327:1320];
      mux_data3[79:72] = in_data3[1335:1328];
      mux_data3[87:80] = in_data3[1343:1336];
      mux_data3[95:88] = in_data3[1351:1344];
      mux_data3[103:96] = in_data3[1359:1352];
      mux_data3[111:104] = in_data3[1367:1360];
      mux_data3[119:112] = in_data3[1375:1368];
      mux_data3[127:120] = in_data3[1383:1376];
      mux_data3[135:128] = in_data3[1391:1384];
      mux_data3[143:136] = in_data3[1399:1392];
      mux_data3[151:144] = in_data3[1407:1400];
      mux_data3[159:152] = in_data3[1415:1408];
      mux_data3[167:160] = in_data3[1423:1416];
      mux_data3[175:168] = in_data3[1431:1424];
      mux_data4[7:0] = in_data4[1263:1256];
      mux_data4[15:8] = in_data4[1271:1264];
      mux_data4[23:16] = in_data4[1279:1272];
      mux_data4[31:24] = in_data4[1287:1280];
      mux_data4[39:32] = in_data4[1295:1288];
      mux_data4[47:40] = in_data4[1303:1296];
      mux_data4[55:48] = in_data4[1311:1304];
      mux_data4[63:56] = in_data4[1319:1312];
      mux_data4[71:64] = in_data4[1327:1320];
      mux_data4[79:72] = in_data4[1335:1328];
      mux_data4[87:80] = in_data4[1343:1336];
      mux_data4[95:88] = in_data4[1351:1344];
      mux_data4[103:96] = in_data4[1359:1352];
      mux_data4[111:104] = in_data4[1367:1360];
      mux_data4[119:112] = in_data4[1375:1368];
      mux_data4[127:120] = in_data4[1383:1376];
      mux_data4[135:128] = in_data4[1391:1384];
      mux_data4[143:136] = in_data4[1399:1392];
      mux_data4[151:144] = in_data4[1407:1400];
      mux_data4[159:152] = in_data4[1415:1408];
      mux_data4[167:160] = in_data4[1423:1416];
      mux_data4[175:168] = in_data4[1431:1424];
    end
    'd11: begin
      mux_data0[7:0] = in_data0[1391:1384];
      mux_data0[15:8] = in_data0[1399:1392];
      mux_data0[23:16] = in_data0[1407:1400];
      mux_data0[31:24] = in_data0[1415:1408];
      mux_data0[39:32] = in_data0[1423:1416];
      mux_data0[47:40] = in_data0[1431:1424];
      mux_data0[55:48] = in_data0[1439:1432];
      mux_data0[63:56] = in_data0[1447:1440];
      mux_data0[71:64] = in_data0[1455:1448];
      mux_data0[79:72] = in_data0[1463:1456];
      mux_data0[87:80] = in_data0[1471:1464];
      mux_data0[95:88] = in_data0[1479:1472];
      mux_data0[103:96] = in_data0[1487:1480];
      mux_data0[111:104] = in_data0[1495:1488];
      mux_data0[119:112] = in_data0[1503:1496];
      mux_data0[127:120] = in_data0[1511:1504];
      mux_data0[135:128] = in_data0[1519:1512];
      mux_data0[143:136] = in_data0[1527:1520];
      mux_data0[151:144] = in_data0[1535:1528];
      mux_data0[159:152] = in_data0[1543:1536];
      mux_data0[167:160] = in_data0[1551:1544];
      mux_data0[175:168] = in_data0[1559:1552];
      mux_data1[7:0] = in_data1[1391:1384];
      mux_data1[15:8] = in_data1[1399:1392];
      mux_data1[23:16] = in_data1[1407:1400];
      mux_data1[31:24] = in_data1[1415:1408];
      mux_data1[39:32] = in_data1[1423:1416];
      mux_data1[47:40] = in_data1[1431:1424];
      mux_data1[55:48] = in_data1[1439:1432];
      mux_data1[63:56] = in_data1[1447:1440];
      mux_data1[71:64] = in_data1[1455:1448];
      mux_data1[79:72] = in_data1[1463:1456];
      mux_data1[87:80] = in_data1[1471:1464];
      mux_data1[95:88] = in_data1[1479:1472];
      mux_data1[103:96] = in_data1[1487:1480];
      mux_data1[111:104] = in_data1[1495:1488];
      mux_data1[119:112] = in_data1[1503:1496];
      mux_data1[127:120] = in_data1[1511:1504];
      mux_data1[135:128] = in_data1[1519:1512];
      mux_data1[143:136] = in_data1[1527:1520];
      mux_data1[151:144] = in_data1[1535:1528];
      mux_data1[159:152] = in_data1[1543:1536];
      mux_data1[167:160] = in_data1[1551:1544];
      mux_data1[175:168] = in_data1[1559:1552];
      mux_data2[7:0] = in_data2[1391:1384];
      mux_data2[15:8] = in_data2[1399:1392];
      mux_data2[23:16] = in_data2[1407:1400];
      mux_data2[31:24] = in_data2[1415:1408];
      mux_data2[39:32] = in_data2[1423:1416];
      mux_data2[47:40] = in_data2[1431:1424];
      mux_data2[55:48] = in_data2[1439:1432];
      mux_data2[63:56] = in_data2[1447:1440];
      mux_data2[71:64] = in_data2[1455:1448];
      mux_data2[79:72] = in_data2[1463:1456];
      mux_data2[87:80] = in_data2[1471:1464];
      mux_data2[95:88] = in_data2[1479:1472];
      mux_data2[103:96] = in_data2[1487:1480];
      mux_data2[111:104] = in_data2[1495:1488];
      mux_data2[119:112] = in_data2[1503:1496];
      mux_data2[127:120] = in_data2[1511:1504];
      mux_data2[135:128] = in_data2[1519:1512];
      mux_data2[143:136] = in_data2[1527:1520];
      mux_data2[151:144] = in_data2[1535:1528];
      mux_data2[159:152] = in_data2[1543:1536];
      mux_data2[167:160] = in_data2[1551:1544];
      mux_data2[175:168] = in_data2[1559:1552];
      mux_data3[7:0] = in_data3[1391:1384];
      mux_data3[15:8] = in_data3[1399:1392];
      mux_data3[23:16] = in_data3[1407:1400];
      mux_data3[31:24] = in_data3[1415:1408];
      mux_data3[39:32] = in_data3[1423:1416];
      mux_data3[47:40] = in_data3[1431:1424];
      mux_data3[55:48] = in_data3[1439:1432];
      mux_data3[63:56] = in_data3[1447:1440];
      mux_data3[71:64] = in_data3[1455:1448];
      mux_data3[79:72] = in_data3[1463:1456];
      mux_data3[87:80] = in_data3[1471:1464];
      mux_data3[95:88] = in_data3[1479:1472];
      mux_data3[103:96] = in_data3[1487:1480];
      mux_data3[111:104] = in_data3[1495:1488];
      mux_data3[119:112] = in_data3[1503:1496];
      mux_data3[127:120] = in_data3[1511:1504];
      mux_data3[135:128] = in_data3[1519:1512];
      mux_data3[143:136] = in_data3[1527:1520];
      mux_data3[151:144] = in_data3[1535:1528];
      mux_data3[159:152] = in_data3[1543:1536];
      mux_data3[167:160] = in_data3[1551:1544];
      mux_data3[175:168] = in_data3[1559:1552];
      mux_data4[7:0] = in_data4[1391:1384];
      mux_data4[15:8] = in_data4[1399:1392];
      mux_data4[23:16] = in_data4[1407:1400];
      mux_data4[31:24] = in_data4[1415:1408];
      mux_data4[39:32] = in_data4[1423:1416];
      mux_data4[47:40] = in_data4[1431:1424];
      mux_data4[55:48] = in_data4[1439:1432];
      mux_data4[63:56] = in_data4[1447:1440];
      mux_data4[71:64] = in_data4[1455:1448];
      mux_data4[79:72] = in_data4[1463:1456];
      mux_data4[87:80] = in_data4[1471:1464];
      mux_data4[95:88] = in_data4[1479:1472];
      mux_data4[103:96] = in_data4[1487:1480];
      mux_data4[111:104] = in_data4[1495:1488];
      mux_data4[119:112] = in_data4[1503:1496];
      mux_data4[127:120] = in_data4[1511:1504];
      mux_data4[135:128] = in_data4[1519:1512];
      mux_data4[143:136] = in_data4[1527:1520];
      mux_data4[151:144] = in_data4[1535:1528];
      mux_data4[159:152] = in_data4[1543:1536];
      mux_data4[167:160] = in_data4[1551:1544];
      mux_data4[175:168] = in_data4[1559:1552];
    end
    'd12: begin
      mux_data0[7:0] = in_data0[1519:1512];
      mux_data0[15:8] = in_data0[1527:1520];
      mux_data0[23:16] = in_data0[1535:1528];
      mux_data0[31:24] = in_data0[1543:1536];
      mux_data0[39:32] = in_data0[1551:1544];
      mux_data0[47:40] = in_data0[1559:1552];
      mux_data0[55:48] = in_data0[1567:1560];
      mux_data0[63:56] = in_data0[1575:1568];
      mux_data0[71:64] = in_data0[1583:1576];
      mux_data0[79:72] = in_data0[1591:1584];
      mux_data0[87:80] = in_data0[1599:1592];
      mux_data0[95:88] = in_data0[1607:1600];
      mux_data0[103:96] = in_data0[1615:1608];
      mux_data0[111:104] = in_data0[1623:1616];
      mux_data0[119:112] = in_data0[1631:1624];
      mux_data0[127:120] = in_data0[1639:1632];
      mux_data0[135:128] = in_data0[1647:1640];
      mux_data0[143:136] = in_data0[1655:1648];
      mux_data0[151:144] = in_data0[1663:1656];
      mux_data0[159:152] = in_data0[1671:1664];
      mux_data0[167:160] = in_data0[1679:1672];
      mux_data0[175:168] = in_data0[1687:1680];
      mux_data1[7:0] = in_data1[1519:1512];
      mux_data1[15:8] = in_data1[1527:1520];
      mux_data1[23:16] = in_data1[1535:1528];
      mux_data1[31:24] = in_data1[1543:1536];
      mux_data1[39:32] = in_data1[1551:1544];
      mux_data1[47:40] = in_data1[1559:1552];
      mux_data1[55:48] = in_data1[1567:1560];
      mux_data1[63:56] = in_data1[1575:1568];
      mux_data1[71:64] = in_data1[1583:1576];
      mux_data1[79:72] = in_data1[1591:1584];
      mux_data1[87:80] = in_data1[1599:1592];
      mux_data1[95:88] = in_data1[1607:1600];
      mux_data1[103:96] = in_data1[1615:1608];
      mux_data1[111:104] = in_data1[1623:1616];
      mux_data1[119:112] = in_data1[1631:1624];
      mux_data1[127:120] = in_data1[1639:1632];
      mux_data1[135:128] = in_data1[1647:1640];
      mux_data1[143:136] = in_data1[1655:1648];
      mux_data1[151:144] = in_data1[1663:1656];
      mux_data1[159:152] = in_data1[1671:1664];
      mux_data1[167:160] = in_data1[1679:1672];
      mux_data1[175:168] = in_data1[1687:1680];
      mux_data2[7:0] = in_data2[1519:1512];
      mux_data2[15:8] = in_data2[1527:1520];
      mux_data2[23:16] = in_data2[1535:1528];
      mux_data2[31:24] = in_data2[1543:1536];
      mux_data2[39:32] = in_data2[1551:1544];
      mux_data2[47:40] = in_data2[1559:1552];
      mux_data2[55:48] = in_data2[1567:1560];
      mux_data2[63:56] = in_data2[1575:1568];
      mux_data2[71:64] = in_data2[1583:1576];
      mux_data2[79:72] = in_data2[1591:1584];
      mux_data2[87:80] = in_data2[1599:1592];
      mux_data2[95:88] = in_data2[1607:1600];
      mux_data2[103:96] = in_data2[1615:1608];
      mux_data2[111:104] = in_data2[1623:1616];
      mux_data2[119:112] = in_data2[1631:1624];
      mux_data2[127:120] = in_data2[1639:1632];
      mux_data2[135:128] = in_data2[1647:1640];
      mux_data2[143:136] = in_data2[1655:1648];
      mux_data2[151:144] = in_data2[1663:1656];
      mux_data2[159:152] = in_data2[1671:1664];
      mux_data2[167:160] = in_data2[1679:1672];
      mux_data2[175:168] = in_data2[1687:1680];
      mux_data3[7:0] = in_data3[1519:1512];
      mux_data3[15:8] = in_data3[1527:1520];
      mux_data3[23:16] = in_data3[1535:1528];
      mux_data3[31:24] = in_data3[1543:1536];
      mux_data3[39:32] = in_data3[1551:1544];
      mux_data3[47:40] = in_data3[1559:1552];
      mux_data3[55:48] = in_data3[1567:1560];
      mux_data3[63:56] = in_data3[1575:1568];
      mux_data3[71:64] = in_data3[1583:1576];
      mux_data3[79:72] = in_data3[1591:1584];
      mux_data3[87:80] = in_data3[1599:1592];
      mux_data3[95:88] = in_data3[1607:1600];
      mux_data3[103:96] = in_data3[1615:1608];
      mux_data3[111:104] = in_data3[1623:1616];
      mux_data3[119:112] = in_data3[1631:1624];
      mux_data3[127:120] = in_data3[1639:1632];
      mux_data3[135:128] = in_data3[1647:1640];
      mux_data3[143:136] = in_data3[1655:1648];
      mux_data3[151:144] = in_data3[1663:1656];
      mux_data3[159:152] = in_data3[1671:1664];
      mux_data3[167:160] = in_data3[1679:1672];
      mux_data3[175:168] = in_data3[1687:1680];
      mux_data4[7:0] = in_data4[1519:1512];
      mux_data4[15:8] = in_data4[1527:1520];
      mux_data4[23:16] = in_data4[1535:1528];
      mux_data4[31:24] = in_data4[1543:1536];
      mux_data4[39:32] = in_data4[1551:1544];
      mux_data4[47:40] = in_data4[1559:1552];
      mux_data4[55:48] = in_data4[1567:1560];
      mux_data4[63:56] = in_data4[1575:1568];
      mux_data4[71:64] = in_data4[1583:1576];
      mux_data4[79:72] = in_data4[1591:1584];
      mux_data4[87:80] = in_data4[1599:1592];
      mux_data4[95:88] = in_data4[1607:1600];
      mux_data4[103:96] = in_data4[1615:1608];
      mux_data4[111:104] = in_data4[1623:1616];
      mux_data4[119:112] = in_data4[1631:1624];
      mux_data4[127:120] = in_data4[1639:1632];
      mux_data4[135:128] = in_data4[1647:1640];
      mux_data4[143:136] = in_data4[1655:1648];
      mux_data4[151:144] = in_data4[1663:1656];
      mux_data4[159:152] = in_data4[1671:1664];
      mux_data4[167:160] = in_data4[1679:1672];
      mux_data4[175:168] = in_data4[1687:1680];
    end
    'd13: begin
      mux_data0[7:0] = in_data0[1647:1640];
      mux_data0[15:8] = in_data0[1655:1648];
      mux_data0[23:16] = in_data0[1663:1656];
      mux_data0[31:24] = in_data0[1671:1664];
      mux_data0[39:32] = in_data0[1679:1672];
      mux_data0[47:40] = in_data0[1687:1680];
      mux_data0[55:48] = in_data0[1695:1688];
      mux_data0[63:56] = in_data0[1703:1696];
      mux_data0[71:64] = in_data0[1711:1704];
      mux_data0[79:72] = in_data0[1719:1712];
      mux_data0[87:80] = in_data0[1727:1720];
      mux_data0[95:88] = in_data0[1735:1728];
      mux_data0[103:96] = in_data0[1743:1736];
      mux_data0[111:104] = in_data0[1751:1744];
      mux_data0[119:112] = in_data0[1759:1752];
      mux_data0[127:120] = in_data0[1767:1760];
      mux_data0[135:128] = in_data0[1775:1768];
      mux_data0[143:136] = in_data0[1783:1776];
      mux_data0[151:144] = in_data0[1791:1784];
      mux_data0[159:152] = in_data0[1799:1792];
      mux_data0[167:160] = in_data0[1807:1800];
      mux_data0[175:168] = in_data0[1815:1808];
      mux_data1[7:0] = in_data1[1647:1640];
      mux_data1[15:8] = in_data1[1655:1648];
      mux_data1[23:16] = in_data1[1663:1656];
      mux_data1[31:24] = in_data1[1671:1664];
      mux_data1[39:32] = in_data1[1679:1672];
      mux_data1[47:40] = in_data1[1687:1680];
      mux_data1[55:48] = in_data1[1695:1688];
      mux_data1[63:56] = in_data1[1703:1696];
      mux_data1[71:64] = in_data1[1711:1704];
      mux_data1[79:72] = in_data1[1719:1712];
      mux_data1[87:80] = in_data1[1727:1720];
      mux_data1[95:88] = in_data1[1735:1728];
      mux_data1[103:96] = in_data1[1743:1736];
      mux_data1[111:104] = in_data1[1751:1744];
      mux_data1[119:112] = in_data1[1759:1752];
      mux_data1[127:120] = in_data1[1767:1760];
      mux_data1[135:128] = in_data1[1775:1768];
      mux_data1[143:136] = in_data1[1783:1776];
      mux_data1[151:144] = in_data1[1791:1784];
      mux_data1[159:152] = in_data1[1799:1792];
      mux_data1[167:160] = in_data1[1807:1800];
      mux_data1[175:168] = in_data1[1815:1808];
      mux_data2[7:0] = in_data2[1647:1640];
      mux_data2[15:8] = in_data2[1655:1648];
      mux_data2[23:16] = in_data2[1663:1656];
      mux_data2[31:24] = in_data2[1671:1664];
      mux_data2[39:32] = in_data2[1679:1672];
      mux_data2[47:40] = in_data2[1687:1680];
      mux_data2[55:48] = in_data2[1695:1688];
      mux_data2[63:56] = in_data2[1703:1696];
      mux_data2[71:64] = in_data2[1711:1704];
      mux_data2[79:72] = in_data2[1719:1712];
      mux_data2[87:80] = in_data2[1727:1720];
      mux_data2[95:88] = in_data2[1735:1728];
      mux_data2[103:96] = in_data2[1743:1736];
      mux_data2[111:104] = in_data2[1751:1744];
      mux_data2[119:112] = in_data2[1759:1752];
      mux_data2[127:120] = in_data2[1767:1760];
      mux_data2[135:128] = in_data2[1775:1768];
      mux_data2[143:136] = in_data2[1783:1776];
      mux_data2[151:144] = in_data2[1791:1784];
      mux_data2[159:152] = in_data2[1799:1792];
      mux_data2[167:160] = in_data2[1807:1800];
      mux_data2[175:168] = in_data2[1815:1808];
      mux_data3[7:0] = in_data3[1647:1640];
      mux_data3[15:8] = in_data3[1655:1648];
      mux_data3[23:16] = in_data3[1663:1656];
      mux_data3[31:24] = in_data3[1671:1664];
      mux_data3[39:32] = in_data3[1679:1672];
      mux_data3[47:40] = in_data3[1687:1680];
      mux_data3[55:48] = in_data3[1695:1688];
      mux_data3[63:56] = in_data3[1703:1696];
      mux_data3[71:64] = in_data3[1711:1704];
      mux_data3[79:72] = in_data3[1719:1712];
      mux_data3[87:80] = in_data3[1727:1720];
      mux_data3[95:88] = in_data3[1735:1728];
      mux_data3[103:96] = in_data3[1743:1736];
      mux_data3[111:104] = in_data3[1751:1744];
      mux_data3[119:112] = in_data3[1759:1752];
      mux_data3[127:120] = in_data3[1767:1760];
      mux_data3[135:128] = in_data3[1775:1768];
      mux_data3[143:136] = in_data3[1783:1776];
      mux_data3[151:144] = in_data3[1791:1784];
      mux_data3[159:152] = in_data3[1799:1792];
      mux_data3[167:160] = in_data3[1807:1800];
      mux_data3[175:168] = in_data3[1815:1808];
      mux_data4[7:0] = in_data4[1647:1640];
      mux_data4[15:8] = in_data4[1655:1648];
      mux_data4[23:16] = in_data4[1663:1656];
      mux_data4[31:24] = in_data4[1671:1664];
      mux_data4[39:32] = in_data4[1679:1672];
      mux_data4[47:40] = in_data4[1687:1680];
      mux_data4[55:48] = in_data4[1695:1688];
      mux_data4[63:56] = in_data4[1703:1696];
      mux_data4[71:64] = in_data4[1711:1704];
      mux_data4[79:72] = in_data4[1719:1712];
      mux_data4[87:80] = in_data4[1727:1720];
      mux_data4[95:88] = in_data4[1735:1728];
      mux_data4[103:96] = in_data4[1743:1736];
      mux_data4[111:104] = in_data4[1751:1744];
      mux_data4[119:112] = in_data4[1759:1752];
      mux_data4[127:120] = in_data4[1767:1760];
      mux_data4[135:128] = in_data4[1775:1768];
      mux_data4[143:136] = in_data4[1783:1776];
      mux_data4[151:144] = in_data4[1791:1784];
      mux_data4[159:152] = in_data4[1799:1792];
      mux_data4[167:160] = in_data4[1807:1800];
      mux_data4[175:168] = in_data4[1815:1808];
    end
    'd14: begin
      mux_data0[7:0] = in_data0[1775:1768];
      mux_data0[15:8] = in_data0[1783:1776];
      mux_data0[23:16] = in_data0[1791:1784];
      mux_data0[31:24] = in_data0[1799:1792];
      mux_data0[39:32] = in_data0[1807:1800];
      mux_data0[47:40] = in_data0[1815:1808];
      mux_data0[55:48] = in_data0[1823:1816];
      mux_data0[63:56] = in_data0[1831:1824];
      mux_data0[71:64] = in_data0[1839:1832];
      mux_data0[79:72] = in_data0[1847:1840];
      mux_data0[87:80] = in_data0[1855:1848];
      mux_data0[95:88] = in_data0[1863:1856];
      mux_data0[103:96] = in_data0[1871:1864];
      mux_data0[111:104] = in_data0[1879:1872];
      mux_data0[119:112] = in_data0[1887:1880];
      mux_data0[127:120] = in_data0[1895:1888];
      mux_data0[135:128] = in_data0[1903:1896];
      mux_data0[143:136] = in_data0[1911:1904];
      mux_data0[151:144] = in_data0[1919:1912];
      mux_data0[159:152] = in_data0[1927:1920];
      mux_data0[167:160] = in_data0[1935:1928];
      mux_data0[175:168] = in_data0[1943:1936];
      mux_data1[7:0] = in_data1[1775:1768];
      mux_data1[15:8] = in_data1[1783:1776];
      mux_data1[23:16] = in_data1[1791:1784];
      mux_data1[31:24] = in_data1[1799:1792];
      mux_data1[39:32] = in_data1[1807:1800];
      mux_data1[47:40] = in_data1[1815:1808];
      mux_data1[55:48] = in_data1[1823:1816];
      mux_data1[63:56] = in_data1[1831:1824];
      mux_data1[71:64] = in_data1[1839:1832];
      mux_data1[79:72] = in_data1[1847:1840];
      mux_data1[87:80] = in_data1[1855:1848];
      mux_data1[95:88] = in_data1[1863:1856];
      mux_data1[103:96] = in_data1[1871:1864];
      mux_data1[111:104] = in_data1[1879:1872];
      mux_data1[119:112] = in_data1[1887:1880];
      mux_data1[127:120] = in_data1[1895:1888];
      mux_data1[135:128] = in_data1[1903:1896];
      mux_data1[143:136] = in_data1[1911:1904];
      mux_data1[151:144] = in_data1[1919:1912];
      mux_data1[159:152] = in_data1[1927:1920];
      mux_data1[167:160] = in_data1[1935:1928];
      mux_data1[175:168] = in_data1[1943:1936];
      mux_data2[7:0] = in_data2[1775:1768];
      mux_data2[15:8] = in_data2[1783:1776];
      mux_data2[23:16] = in_data2[1791:1784];
      mux_data2[31:24] = in_data2[1799:1792];
      mux_data2[39:32] = in_data2[1807:1800];
      mux_data2[47:40] = in_data2[1815:1808];
      mux_data2[55:48] = in_data2[1823:1816];
      mux_data2[63:56] = in_data2[1831:1824];
      mux_data2[71:64] = in_data2[1839:1832];
      mux_data2[79:72] = in_data2[1847:1840];
      mux_data2[87:80] = in_data2[1855:1848];
      mux_data2[95:88] = in_data2[1863:1856];
      mux_data2[103:96] = in_data2[1871:1864];
      mux_data2[111:104] = in_data2[1879:1872];
      mux_data2[119:112] = in_data2[1887:1880];
      mux_data2[127:120] = in_data2[1895:1888];
      mux_data2[135:128] = in_data2[1903:1896];
      mux_data2[143:136] = in_data2[1911:1904];
      mux_data2[151:144] = in_data2[1919:1912];
      mux_data2[159:152] = in_data2[1927:1920];
      mux_data2[167:160] = in_data2[1935:1928];
      mux_data2[175:168] = in_data2[1943:1936];
      mux_data3[7:0] = in_data3[1775:1768];
      mux_data3[15:8] = in_data3[1783:1776];
      mux_data3[23:16] = in_data3[1791:1784];
      mux_data3[31:24] = in_data3[1799:1792];
      mux_data3[39:32] = in_data3[1807:1800];
      mux_data3[47:40] = in_data3[1815:1808];
      mux_data3[55:48] = in_data3[1823:1816];
      mux_data3[63:56] = in_data3[1831:1824];
      mux_data3[71:64] = in_data3[1839:1832];
      mux_data3[79:72] = in_data3[1847:1840];
      mux_data3[87:80] = in_data3[1855:1848];
      mux_data3[95:88] = in_data3[1863:1856];
      mux_data3[103:96] = in_data3[1871:1864];
      mux_data3[111:104] = in_data3[1879:1872];
      mux_data3[119:112] = in_data3[1887:1880];
      mux_data3[127:120] = in_data3[1895:1888];
      mux_data3[135:128] = in_data3[1903:1896];
      mux_data3[143:136] = in_data3[1911:1904];
      mux_data3[151:144] = in_data3[1919:1912];
      mux_data3[159:152] = in_data3[1927:1920];
      mux_data3[167:160] = in_data3[1935:1928];
      mux_data3[175:168] = in_data3[1943:1936];
      mux_data4[7:0] = in_data4[1775:1768];
      mux_data4[15:8] = in_data4[1783:1776];
      mux_data4[23:16] = in_data4[1791:1784];
      mux_data4[31:24] = in_data4[1799:1792];
      mux_data4[39:32] = in_data4[1807:1800];
      mux_data4[47:40] = in_data4[1815:1808];
      mux_data4[55:48] = in_data4[1823:1816];
      mux_data4[63:56] = in_data4[1831:1824];
      mux_data4[71:64] = in_data4[1839:1832];
      mux_data4[79:72] = in_data4[1847:1840];
      mux_data4[87:80] = in_data4[1855:1848];
      mux_data4[95:88] = in_data4[1863:1856];
      mux_data4[103:96] = in_data4[1871:1864];
      mux_data4[111:104] = in_data4[1879:1872];
      mux_data4[119:112] = in_data4[1887:1880];
      mux_data4[127:120] = in_data4[1895:1888];
      mux_data4[135:128] = in_data4[1903:1896];
      mux_data4[143:136] = in_data4[1911:1904];
      mux_data4[151:144] = in_data4[1919:1912];
      mux_data4[159:152] = in_data4[1927:1920];
      mux_data4[167:160] = in_data4[1935:1928];
      mux_data4[175:168] = in_data4[1943:1936];
    end
    'd15: begin
      mux_data0[7:0] = in_data0[1903:1896];
      mux_data0[15:8] = in_data0[1911:1904];
      mux_data0[23:16] = in_data0[1919:1912];
      mux_data0[31:24] = in_data0[1927:1920];
      mux_data0[39:32] = in_data0[1935:1928];
      mux_data0[47:40] = in_data0[1943:1936];
      mux_data0[55:48] = in_data0[1951:1944];
      mux_data0[63:56] = in_data0[1959:1952];
      mux_data0[71:64] = in_data0[1967:1960];
      mux_data0[79:72] = in_data0[1975:1968];
      mux_data0[87:80] = in_data0[1983:1976];
      mux_data0[95:88] = in_data0[1991:1984];
      mux_data0[103:96] = in_data0[1999:1992];
      mux_data0[111:104] = in_data0[2007:2000];
      mux_data0[119:112] = in_data0[2015:2008];
      mux_data0[127:120] = in_data0[2023:2016];
      mux_data0[135:128] = in_data0[2031:2024];
      mux_data0[143:136] = in_data0[2039:2032];
      mux_data0[151:144] = in_data0[2047:2040];
      mux_data0[159:152] = in_data0[2055:2048];
      mux_data0[167:160] = in_data0[2063:2056];
      mux_data0[175:168] = in_data0[2071:2064];
      mux_data1[7:0] = in_data1[1903:1896];
      mux_data1[15:8] = in_data1[1911:1904];
      mux_data1[23:16] = in_data1[1919:1912];
      mux_data1[31:24] = in_data1[1927:1920];
      mux_data1[39:32] = in_data1[1935:1928];
      mux_data1[47:40] = in_data1[1943:1936];
      mux_data1[55:48] = in_data1[1951:1944];
      mux_data1[63:56] = in_data1[1959:1952];
      mux_data1[71:64] = in_data1[1967:1960];
      mux_data1[79:72] = in_data1[1975:1968];
      mux_data1[87:80] = in_data1[1983:1976];
      mux_data1[95:88] = in_data1[1991:1984];
      mux_data1[103:96] = in_data1[1999:1992];
      mux_data1[111:104] = in_data1[2007:2000];
      mux_data1[119:112] = in_data1[2015:2008];
      mux_data1[127:120] = in_data1[2023:2016];
      mux_data1[135:128] = in_data1[2031:2024];
      mux_data1[143:136] = in_data1[2039:2032];
      mux_data1[151:144] = in_data1[2047:2040];
      mux_data1[159:152] = in_data1[2055:2048];
      mux_data1[167:160] = in_data1[2063:2056];
      mux_data1[175:168] = in_data1[2071:2064];
      mux_data2[7:0] = in_data2[1903:1896];
      mux_data2[15:8] = in_data2[1911:1904];
      mux_data2[23:16] = in_data2[1919:1912];
      mux_data2[31:24] = in_data2[1927:1920];
      mux_data2[39:32] = in_data2[1935:1928];
      mux_data2[47:40] = in_data2[1943:1936];
      mux_data2[55:48] = in_data2[1951:1944];
      mux_data2[63:56] = in_data2[1959:1952];
      mux_data2[71:64] = in_data2[1967:1960];
      mux_data2[79:72] = in_data2[1975:1968];
      mux_data2[87:80] = in_data2[1983:1976];
      mux_data2[95:88] = in_data2[1991:1984];
      mux_data2[103:96] = in_data2[1999:1992];
      mux_data2[111:104] = in_data2[2007:2000];
      mux_data2[119:112] = in_data2[2015:2008];
      mux_data2[127:120] = in_data2[2023:2016];
      mux_data2[135:128] = in_data2[2031:2024];
      mux_data2[143:136] = in_data2[2039:2032];
      mux_data2[151:144] = in_data2[2047:2040];
      mux_data2[159:152] = in_data2[2055:2048];
      mux_data2[167:160] = in_data2[2063:2056];
      mux_data2[175:168] = in_data2[2071:2064];
      mux_data3[7:0] = in_data3[1903:1896];
      mux_data3[15:8] = in_data3[1911:1904];
      mux_data3[23:16] = in_data3[1919:1912];
      mux_data3[31:24] = in_data3[1927:1920];
      mux_data3[39:32] = in_data3[1935:1928];
      mux_data3[47:40] = in_data3[1943:1936];
      mux_data3[55:48] = in_data3[1951:1944];
      mux_data3[63:56] = in_data3[1959:1952];
      mux_data3[71:64] = in_data3[1967:1960];
      mux_data3[79:72] = in_data3[1975:1968];
      mux_data3[87:80] = in_data3[1983:1976];
      mux_data3[95:88] = in_data3[1991:1984];
      mux_data3[103:96] = in_data3[1999:1992];
      mux_data3[111:104] = in_data3[2007:2000];
      mux_data3[119:112] = in_data3[2015:2008];
      mux_data3[127:120] = in_data3[2023:2016];
      mux_data3[135:128] = in_data3[2031:2024];
      mux_data3[143:136] = in_data3[2039:2032];
      mux_data3[151:144] = in_data3[2047:2040];
      mux_data3[159:152] = in_data3[2055:2048];
      mux_data3[167:160] = in_data3[2063:2056];
      mux_data3[175:168] = in_data3[2071:2064];
      mux_data4[7:0] = in_data4[1903:1896];
      mux_data4[15:8] = in_data4[1911:1904];
      mux_data4[23:16] = in_data4[1919:1912];
      mux_data4[31:24] = in_data4[1927:1920];
      mux_data4[39:32] = in_data4[1935:1928];
      mux_data4[47:40] = in_data4[1943:1936];
      mux_data4[55:48] = in_data4[1951:1944];
      mux_data4[63:56] = in_data4[1959:1952];
      mux_data4[71:64] = in_data4[1967:1960];
      mux_data4[79:72] = in_data4[1975:1968];
      mux_data4[87:80] = in_data4[1983:1976];
      mux_data4[95:88] = in_data4[1991:1984];
      mux_data4[103:96] = in_data4[1999:1992];
      mux_data4[111:104] = in_data4[2007:2000];
      mux_data4[119:112] = in_data4[2015:2008];
      mux_data4[127:120] = in_data4[2023:2016];
      mux_data4[135:128] = in_data4[2031:2024];
      mux_data4[143:136] = in_data4[2039:2032];
      mux_data4[151:144] = in_data4[2047:2040];
      mux_data4[159:152] = in_data4[2055:2048];
      mux_data4[167:160] = in_data4[2063:2056];
      mux_data4[175:168] = in_data4[2071:2064];
    end
    'd16: begin
      mux_data0[7:0] = in_data0[2031:2024];
      mux_data0[15:8] = in_data0[2039:2032];
      mux_data0[23:16] = in_data0[2047:2040];
      mux_data0[31:24] = in_data0[2055:2048];
      mux_data0[39:32] = in_data0[2063:2056];
      mux_data0[47:40] = in_data0[2071:2064];
      mux_data0[55:48] = in_data0[2079:2072];
      mux_data0[63:56] = in_data0[2087:2080];
      mux_data0[71:64] = in_data0[2095:2088];
      mux_data0[79:72] = in_data0[2103:2096];
      mux_data0[87:80] = in_data0[2111:2104];
      mux_data0[95:88] = in_data0[2119:2112];
      mux_data0[103:96] = in_data0[2127:2120];
      mux_data0[111:104] = in_data0[2135:2128];
      mux_data0[119:112] = in_data0[2143:2136];
      mux_data0[127:120] = in_data0[2151:2144];
      mux_data0[135:128] = in_data0[2159:2152];
      mux_data0[143:136] = in_data0[2167:2160];
      mux_data0[151:144] = in_data0[2175:2168];
      mux_data0[159:152] = in_data0[2183:2176];
      mux_data0[167:160] = in_data0[2191:2184];
      mux_data0[175:168] = in_data0[2199:2192];
      mux_data1[7:0] = in_data1[2031:2024];
      mux_data1[15:8] = in_data1[2039:2032];
      mux_data1[23:16] = in_data1[2047:2040];
      mux_data1[31:24] = in_data1[2055:2048];
      mux_data1[39:32] = in_data1[2063:2056];
      mux_data1[47:40] = in_data1[2071:2064];
      mux_data1[55:48] = in_data1[2079:2072];
      mux_data1[63:56] = in_data1[2087:2080];
      mux_data1[71:64] = in_data1[2095:2088];
      mux_data1[79:72] = in_data1[2103:2096];
      mux_data1[87:80] = in_data1[2111:2104];
      mux_data1[95:88] = in_data1[2119:2112];
      mux_data1[103:96] = in_data1[2127:2120];
      mux_data1[111:104] = in_data1[2135:2128];
      mux_data1[119:112] = in_data1[2143:2136];
      mux_data1[127:120] = in_data1[2151:2144];
      mux_data1[135:128] = in_data1[2159:2152];
      mux_data1[143:136] = in_data1[2167:2160];
      mux_data1[151:144] = in_data1[2175:2168];
      mux_data1[159:152] = in_data1[2183:2176];
      mux_data1[167:160] = in_data1[2191:2184];
      mux_data1[175:168] = in_data1[2199:2192];
      mux_data2[7:0] = in_data2[2031:2024];
      mux_data2[15:8] = in_data2[2039:2032];
      mux_data2[23:16] = in_data2[2047:2040];
      mux_data2[31:24] = in_data2[2055:2048];
      mux_data2[39:32] = in_data2[2063:2056];
      mux_data2[47:40] = in_data2[2071:2064];
      mux_data2[55:48] = in_data2[2079:2072];
      mux_data2[63:56] = in_data2[2087:2080];
      mux_data2[71:64] = in_data2[2095:2088];
      mux_data2[79:72] = in_data2[2103:2096];
      mux_data2[87:80] = in_data2[2111:2104];
      mux_data2[95:88] = in_data2[2119:2112];
      mux_data2[103:96] = in_data2[2127:2120];
      mux_data2[111:104] = in_data2[2135:2128];
      mux_data2[119:112] = in_data2[2143:2136];
      mux_data2[127:120] = in_data2[2151:2144];
      mux_data2[135:128] = in_data2[2159:2152];
      mux_data2[143:136] = in_data2[2167:2160];
      mux_data2[151:144] = in_data2[2175:2168];
      mux_data2[159:152] = in_data2[2183:2176];
      mux_data2[167:160] = in_data2[2191:2184];
      mux_data2[175:168] = in_data2[2199:2192];
      mux_data3[7:0] = in_data3[2031:2024];
      mux_data3[15:8] = in_data3[2039:2032];
      mux_data3[23:16] = in_data3[2047:2040];
      mux_data3[31:24] = in_data3[2055:2048];
      mux_data3[39:32] = in_data3[2063:2056];
      mux_data3[47:40] = in_data3[2071:2064];
      mux_data3[55:48] = in_data3[2079:2072];
      mux_data3[63:56] = in_data3[2087:2080];
      mux_data3[71:64] = in_data3[2095:2088];
      mux_data3[79:72] = in_data3[2103:2096];
      mux_data3[87:80] = in_data3[2111:2104];
      mux_data3[95:88] = in_data3[2119:2112];
      mux_data3[103:96] = in_data3[2127:2120];
      mux_data3[111:104] = in_data3[2135:2128];
      mux_data3[119:112] = in_data3[2143:2136];
      mux_data3[127:120] = in_data3[2151:2144];
      mux_data3[135:128] = in_data3[2159:2152];
      mux_data3[143:136] = in_data3[2167:2160];
      mux_data3[151:144] = in_data3[2175:2168];
      mux_data3[159:152] = in_data3[2183:2176];
      mux_data3[167:160] = in_data3[2191:2184];
      mux_data3[175:168] = in_data3[2199:2192];
      mux_data4[7:0] = in_data4[2031:2024];
      mux_data4[15:8] = in_data4[2039:2032];
      mux_data4[23:16] = in_data4[2047:2040];
      mux_data4[31:24] = in_data4[2055:2048];
      mux_data4[39:32] = in_data4[2063:2056];
      mux_data4[47:40] = in_data4[2071:2064];
      mux_data4[55:48] = in_data4[2079:2072];
      mux_data4[63:56] = in_data4[2087:2080];
      mux_data4[71:64] = in_data4[2095:2088];
      mux_data4[79:72] = in_data4[2103:2096];
      mux_data4[87:80] = in_data4[2111:2104];
      mux_data4[95:88] = in_data4[2119:2112];
      mux_data4[103:96] = in_data4[2127:2120];
      mux_data4[111:104] = in_data4[2135:2128];
      mux_data4[119:112] = in_data4[2143:2136];
      mux_data4[127:120] = in_data4[2151:2144];
      mux_data4[135:128] = in_data4[2159:2152];
      mux_data4[143:136] = in_data4[2167:2160];
      mux_data4[151:144] = in_data4[2175:2168];
      mux_data4[159:152] = in_data4[2183:2176];
      mux_data4[167:160] = in_data4[2191:2184];
      mux_data4[175:168] = in_data4[2199:2192];
    end
    'd17: begin
      mux_data0[7:0] = in_data0[2159:2152];
      mux_data0[15:8] = in_data0[2167:2160];
      mux_data0[23:16] = in_data0[2175:2168];
      mux_data0[31:24] = in_data0[2183:2176];
      mux_data0[39:32] = in_data0[2191:2184];
      mux_data0[47:40] = in_data0[2199:2192];
      mux_data0[55:48] = in_data0[2207:2200];
      mux_data0[63:56] = in_data0[2215:2208];
      mux_data0[71:64] = in_data0[2223:2216];
      mux_data0[79:72] = in_data0[2231:2224];
      mux_data0[87:80] = in_data0[2239:2232];
      mux_data0[95:88] = in_data0[2247:2240];
      mux_data0[103:96] = in_data0[2255:2248];
      mux_data0[111:104] = in_data0[2263:2256];
      mux_data0[119:112] = in_data0[2271:2264];
      mux_data0[127:120] = in_data0[2279:2272];
      mux_data0[135:128] = in_data0[2287:2280];
      mux_data0[143:136] = in_data0[2295:2288];
      mux_data0[151:144] = in_data0[2303:2296];
      mux_data0[159:152] = in_data0[2311:2304];
      mux_data0[167:160] = in_data0[2319:2312];
      mux_data0[175:168] = in_data0[2327:2320];
      mux_data1[7:0] = in_data1[2159:2152];
      mux_data1[15:8] = in_data1[2167:2160];
      mux_data1[23:16] = in_data1[2175:2168];
      mux_data1[31:24] = in_data1[2183:2176];
      mux_data1[39:32] = in_data1[2191:2184];
      mux_data1[47:40] = in_data1[2199:2192];
      mux_data1[55:48] = in_data1[2207:2200];
      mux_data1[63:56] = in_data1[2215:2208];
      mux_data1[71:64] = in_data1[2223:2216];
      mux_data1[79:72] = in_data1[2231:2224];
      mux_data1[87:80] = in_data1[2239:2232];
      mux_data1[95:88] = in_data1[2247:2240];
      mux_data1[103:96] = in_data1[2255:2248];
      mux_data1[111:104] = in_data1[2263:2256];
      mux_data1[119:112] = in_data1[2271:2264];
      mux_data1[127:120] = in_data1[2279:2272];
      mux_data1[135:128] = in_data1[2287:2280];
      mux_data1[143:136] = in_data1[2295:2288];
      mux_data1[151:144] = in_data1[2303:2296];
      mux_data1[159:152] = in_data1[2311:2304];
      mux_data1[167:160] = in_data1[2319:2312];
      mux_data1[175:168] = in_data1[2327:2320];
      mux_data2[7:0] = in_data2[2159:2152];
      mux_data2[15:8] = in_data2[2167:2160];
      mux_data2[23:16] = in_data2[2175:2168];
      mux_data2[31:24] = in_data2[2183:2176];
      mux_data2[39:32] = in_data2[2191:2184];
      mux_data2[47:40] = in_data2[2199:2192];
      mux_data2[55:48] = in_data2[2207:2200];
      mux_data2[63:56] = in_data2[2215:2208];
      mux_data2[71:64] = in_data2[2223:2216];
      mux_data2[79:72] = in_data2[2231:2224];
      mux_data2[87:80] = in_data2[2239:2232];
      mux_data2[95:88] = in_data2[2247:2240];
      mux_data2[103:96] = in_data2[2255:2248];
      mux_data2[111:104] = in_data2[2263:2256];
      mux_data2[119:112] = in_data2[2271:2264];
      mux_data2[127:120] = in_data2[2279:2272];
      mux_data2[135:128] = in_data2[2287:2280];
      mux_data2[143:136] = in_data2[2295:2288];
      mux_data2[151:144] = in_data2[2303:2296];
      mux_data2[159:152] = in_data2[2311:2304];
      mux_data2[167:160] = in_data2[2319:2312];
      mux_data2[175:168] = in_data2[2327:2320];
      mux_data3[7:0] = in_data3[2159:2152];
      mux_data3[15:8] = in_data3[2167:2160];
      mux_data3[23:16] = in_data3[2175:2168];
      mux_data3[31:24] = in_data3[2183:2176];
      mux_data3[39:32] = in_data3[2191:2184];
      mux_data3[47:40] = in_data3[2199:2192];
      mux_data3[55:48] = in_data3[2207:2200];
      mux_data3[63:56] = in_data3[2215:2208];
      mux_data3[71:64] = in_data3[2223:2216];
      mux_data3[79:72] = in_data3[2231:2224];
      mux_data3[87:80] = in_data3[2239:2232];
      mux_data3[95:88] = in_data3[2247:2240];
      mux_data3[103:96] = in_data3[2255:2248];
      mux_data3[111:104] = in_data3[2263:2256];
      mux_data3[119:112] = in_data3[2271:2264];
      mux_data3[127:120] = in_data3[2279:2272];
      mux_data3[135:128] = in_data3[2287:2280];
      mux_data3[143:136] = in_data3[2295:2288];
      mux_data3[151:144] = in_data3[2303:2296];
      mux_data3[159:152] = in_data3[2311:2304];
      mux_data3[167:160] = in_data3[2319:2312];
      mux_data3[175:168] = in_data3[2327:2320];
      mux_data4[7:0] = in_data4[2159:2152];
      mux_data4[15:8] = in_data4[2167:2160];
      mux_data4[23:16] = in_data4[2175:2168];
      mux_data4[31:24] = in_data4[2183:2176];
      mux_data4[39:32] = in_data4[2191:2184];
      mux_data4[47:40] = in_data4[2199:2192];
      mux_data4[55:48] = in_data4[2207:2200];
      mux_data4[63:56] = in_data4[2215:2208];
      mux_data4[71:64] = in_data4[2223:2216];
      mux_data4[79:72] = in_data4[2231:2224];
      mux_data4[87:80] = in_data4[2239:2232];
      mux_data4[95:88] = in_data4[2247:2240];
      mux_data4[103:96] = in_data4[2255:2248];
      mux_data4[111:104] = in_data4[2263:2256];
      mux_data4[119:112] = in_data4[2271:2264];
      mux_data4[127:120] = in_data4[2279:2272];
      mux_data4[135:128] = in_data4[2287:2280];
      mux_data4[143:136] = in_data4[2295:2288];
      mux_data4[151:144] = in_data4[2303:2296];
      mux_data4[159:152] = in_data4[2311:2304];
      mux_data4[167:160] = in_data4[2319:2312];
      mux_data4[175:168] = in_data4[2327:2320];
    end
    'd18: begin
      mux_data0[7:0] = in_data0[2287:2280];
      mux_data0[15:8] = in_data0[2295:2288];
      mux_data0[23:16] = in_data0[2303:2296];
      mux_data0[31:24] = in_data0[2311:2304];
      mux_data0[39:32] = in_data0[2319:2312];
      mux_data0[47:40] = in_data0[2327:2320];
      mux_data0[55:48] = in_data0[2335:2328];
      mux_data0[63:56] = in_data0[2343:2336];
      mux_data0[71:64] = in_data0[2351:2344];
      mux_data0[79:72] = in_data0[2359:2352];
      mux_data0[87:80] = in_data0[2367:2360];
      mux_data0[95:88] = in_data0[2375:2368];
      mux_data0[103:96] = in_data0[2383:2376];
      mux_data0[111:104] = in_data0[2391:2384];
      mux_data0[119:112] = in_data0[2399:2392];
      mux_data0[127:120] = in_data0[2407:2400];
      mux_data0[135:128] = in_data0[2415:2408];
      mux_data0[143:136] = in_data0[2423:2416];
      mux_data0[151:144] = in_data0[2431:2424];
      mux_data0[159:152] = in_data0[2439:2432];
      mux_data0[167:160] = in_data0[2447:2440];
      mux_data0[175:168] = in_data0[2455:2448];
      mux_data1[7:0] = in_data1[2287:2280];
      mux_data1[15:8] = in_data1[2295:2288];
      mux_data1[23:16] = in_data1[2303:2296];
      mux_data1[31:24] = in_data1[2311:2304];
      mux_data1[39:32] = in_data1[2319:2312];
      mux_data1[47:40] = in_data1[2327:2320];
      mux_data1[55:48] = in_data1[2335:2328];
      mux_data1[63:56] = in_data1[2343:2336];
      mux_data1[71:64] = in_data1[2351:2344];
      mux_data1[79:72] = in_data1[2359:2352];
      mux_data1[87:80] = in_data1[2367:2360];
      mux_data1[95:88] = in_data1[2375:2368];
      mux_data1[103:96] = in_data1[2383:2376];
      mux_data1[111:104] = in_data1[2391:2384];
      mux_data1[119:112] = in_data1[2399:2392];
      mux_data1[127:120] = in_data1[2407:2400];
      mux_data1[135:128] = in_data1[2415:2408];
      mux_data1[143:136] = in_data1[2423:2416];
      mux_data1[151:144] = in_data1[2431:2424];
      mux_data1[159:152] = in_data1[2439:2432];
      mux_data1[167:160] = in_data1[2447:2440];
      mux_data1[175:168] = in_data1[2455:2448];
      mux_data2[7:0] = in_data2[2287:2280];
      mux_data2[15:8] = in_data2[2295:2288];
      mux_data2[23:16] = in_data2[2303:2296];
      mux_data2[31:24] = in_data2[2311:2304];
      mux_data2[39:32] = in_data2[2319:2312];
      mux_data2[47:40] = in_data2[2327:2320];
      mux_data2[55:48] = in_data2[2335:2328];
      mux_data2[63:56] = in_data2[2343:2336];
      mux_data2[71:64] = in_data2[2351:2344];
      mux_data2[79:72] = in_data2[2359:2352];
      mux_data2[87:80] = in_data2[2367:2360];
      mux_data2[95:88] = in_data2[2375:2368];
      mux_data2[103:96] = in_data2[2383:2376];
      mux_data2[111:104] = in_data2[2391:2384];
      mux_data2[119:112] = in_data2[2399:2392];
      mux_data2[127:120] = in_data2[2407:2400];
      mux_data2[135:128] = in_data2[2415:2408];
      mux_data2[143:136] = in_data2[2423:2416];
      mux_data2[151:144] = in_data2[2431:2424];
      mux_data2[159:152] = in_data2[2439:2432];
      mux_data2[167:160] = in_data2[2447:2440];
      mux_data2[175:168] = in_data2[2455:2448];
      mux_data3[7:0] = in_data3[2287:2280];
      mux_data3[15:8] = in_data3[2295:2288];
      mux_data3[23:16] = in_data3[2303:2296];
      mux_data3[31:24] = in_data3[2311:2304];
      mux_data3[39:32] = in_data3[2319:2312];
      mux_data3[47:40] = in_data3[2327:2320];
      mux_data3[55:48] = in_data3[2335:2328];
      mux_data3[63:56] = in_data3[2343:2336];
      mux_data3[71:64] = in_data3[2351:2344];
      mux_data3[79:72] = in_data3[2359:2352];
      mux_data3[87:80] = in_data3[2367:2360];
      mux_data3[95:88] = in_data3[2375:2368];
      mux_data3[103:96] = in_data3[2383:2376];
      mux_data3[111:104] = in_data3[2391:2384];
      mux_data3[119:112] = in_data3[2399:2392];
      mux_data3[127:120] = in_data3[2407:2400];
      mux_data3[135:128] = in_data3[2415:2408];
      mux_data3[143:136] = in_data3[2423:2416];
      mux_data3[151:144] = in_data3[2431:2424];
      mux_data3[159:152] = in_data3[2439:2432];
      mux_data3[167:160] = in_data3[2447:2440];
      mux_data3[175:168] = in_data3[2455:2448];
      mux_data4[7:0] = in_data4[2287:2280];
      mux_data4[15:8] = in_data4[2295:2288];
      mux_data4[23:16] = in_data4[2303:2296];
      mux_data4[31:24] = in_data4[2311:2304];
      mux_data4[39:32] = in_data4[2319:2312];
      mux_data4[47:40] = in_data4[2327:2320];
      mux_data4[55:48] = in_data4[2335:2328];
      mux_data4[63:56] = in_data4[2343:2336];
      mux_data4[71:64] = in_data4[2351:2344];
      mux_data4[79:72] = in_data4[2359:2352];
      mux_data4[87:80] = in_data4[2367:2360];
      mux_data4[95:88] = in_data4[2375:2368];
      mux_data4[103:96] = in_data4[2383:2376];
      mux_data4[111:104] = in_data4[2391:2384];
      mux_data4[119:112] = in_data4[2399:2392];
      mux_data4[127:120] = in_data4[2407:2400];
      mux_data4[135:128] = in_data4[2415:2408];
      mux_data4[143:136] = in_data4[2423:2416];
      mux_data4[151:144] = in_data4[2431:2424];
      mux_data4[159:152] = in_data4[2439:2432];
      mux_data4[167:160] = in_data4[2447:2440];
      mux_data4[175:168] = in_data4[2455:2448];
    end
    'd19: begin
      mux_data0[7:0] = in_data0[2415:2408];
      mux_data0[15:8] = in_data0[2423:2416];
      mux_data0[23:16] = in_data0[2431:2424];
      mux_data0[31:24] = in_data0[2439:2432];
      mux_data0[39:32] = in_data0[2447:2440];
      mux_data0[47:40] = in_data0[2455:2448];
      mux_data0[55:48] = in_data0[2463:2456];
      mux_data0[63:56] = in_data0[2471:2464];
      mux_data0[71:64] = in_data0[2479:2472];
      mux_data0[79:72] = in_data0[2487:2480];
      mux_data0[87:80] = in_data0[2495:2488];
      mux_data0[95:88] = in_data0[2503:2496];
      mux_data0[103:96] = in_data0[2511:2504];
      mux_data0[111:104] = in_data0[2519:2512];
      mux_data0[119:112] = in_data0[2527:2520];
      mux_data0[127:120] = in_data0[2535:2528];
      mux_data0[135:128] = in_data0[2543:2536];
      mux_data0[143:136] = in_data0[2551:2544];
      mux_data0[151:144] = in_data0[2559:2552];
      mux_data0[159:152] = in_data0[2567:2560];
      mux_data0[167:160] = in_data0[2575:2568];
      mux_data0[175:168] = in_data0[2583:2576];
      mux_data1[7:0] = in_data1[2415:2408];
      mux_data1[15:8] = in_data1[2423:2416];
      mux_data1[23:16] = in_data1[2431:2424];
      mux_data1[31:24] = in_data1[2439:2432];
      mux_data1[39:32] = in_data1[2447:2440];
      mux_data1[47:40] = in_data1[2455:2448];
      mux_data1[55:48] = in_data1[2463:2456];
      mux_data1[63:56] = in_data1[2471:2464];
      mux_data1[71:64] = in_data1[2479:2472];
      mux_data1[79:72] = in_data1[2487:2480];
      mux_data1[87:80] = in_data1[2495:2488];
      mux_data1[95:88] = in_data1[2503:2496];
      mux_data1[103:96] = in_data1[2511:2504];
      mux_data1[111:104] = in_data1[2519:2512];
      mux_data1[119:112] = in_data1[2527:2520];
      mux_data1[127:120] = in_data1[2535:2528];
      mux_data1[135:128] = in_data1[2543:2536];
      mux_data1[143:136] = in_data1[2551:2544];
      mux_data1[151:144] = in_data1[2559:2552];
      mux_data1[159:152] = in_data1[2567:2560];
      mux_data1[167:160] = in_data1[2575:2568];
      mux_data1[175:168] = in_data1[2583:2576];
      mux_data2[7:0] = in_data2[2415:2408];
      mux_data2[15:8] = in_data2[2423:2416];
      mux_data2[23:16] = in_data2[2431:2424];
      mux_data2[31:24] = in_data2[2439:2432];
      mux_data2[39:32] = in_data2[2447:2440];
      mux_data2[47:40] = in_data2[2455:2448];
      mux_data2[55:48] = in_data2[2463:2456];
      mux_data2[63:56] = in_data2[2471:2464];
      mux_data2[71:64] = in_data2[2479:2472];
      mux_data2[79:72] = in_data2[2487:2480];
      mux_data2[87:80] = in_data2[2495:2488];
      mux_data2[95:88] = in_data2[2503:2496];
      mux_data2[103:96] = in_data2[2511:2504];
      mux_data2[111:104] = in_data2[2519:2512];
      mux_data2[119:112] = in_data2[2527:2520];
      mux_data2[127:120] = in_data2[2535:2528];
      mux_data2[135:128] = in_data2[2543:2536];
      mux_data2[143:136] = in_data2[2551:2544];
      mux_data2[151:144] = in_data2[2559:2552];
      mux_data2[159:152] = in_data2[2567:2560];
      mux_data2[167:160] = in_data2[2575:2568];
      mux_data2[175:168] = in_data2[2583:2576];
      mux_data3[7:0] = in_data3[2415:2408];
      mux_data3[15:8] = in_data3[2423:2416];
      mux_data3[23:16] = in_data3[2431:2424];
      mux_data3[31:24] = in_data3[2439:2432];
      mux_data3[39:32] = in_data3[2447:2440];
      mux_data3[47:40] = in_data3[2455:2448];
      mux_data3[55:48] = in_data3[2463:2456];
      mux_data3[63:56] = in_data3[2471:2464];
      mux_data3[71:64] = in_data3[2479:2472];
      mux_data3[79:72] = in_data3[2487:2480];
      mux_data3[87:80] = in_data3[2495:2488];
      mux_data3[95:88] = in_data3[2503:2496];
      mux_data3[103:96] = in_data3[2511:2504];
      mux_data3[111:104] = in_data3[2519:2512];
      mux_data3[119:112] = in_data3[2527:2520];
      mux_data3[127:120] = in_data3[2535:2528];
      mux_data3[135:128] = in_data3[2543:2536];
      mux_data3[143:136] = in_data3[2551:2544];
      mux_data3[151:144] = in_data3[2559:2552];
      mux_data3[159:152] = in_data3[2567:2560];
      mux_data3[167:160] = in_data3[2575:2568];
      mux_data3[175:168] = in_data3[2583:2576];
      mux_data4[7:0] = in_data4[2415:2408];
      mux_data4[15:8] = in_data4[2423:2416];
      mux_data4[23:16] = in_data4[2431:2424];
      mux_data4[31:24] = in_data4[2439:2432];
      mux_data4[39:32] = in_data4[2447:2440];
      mux_data4[47:40] = in_data4[2455:2448];
      mux_data4[55:48] = in_data4[2463:2456];
      mux_data4[63:56] = in_data4[2471:2464];
      mux_data4[71:64] = in_data4[2479:2472];
      mux_data4[79:72] = in_data4[2487:2480];
      mux_data4[87:80] = in_data4[2495:2488];
      mux_data4[95:88] = in_data4[2503:2496];
      mux_data4[103:96] = in_data4[2511:2504];
      mux_data4[111:104] = in_data4[2519:2512];
      mux_data4[119:112] = in_data4[2527:2520];
      mux_data4[127:120] = in_data4[2535:2528];
      mux_data4[135:128] = in_data4[2543:2536];
      mux_data4[143:136] = in_data4[2551:2544];
      mux_data4[151:144] = in_data4[2559:2552];
      mux_data4[159:152] = in_data4[2567:2560];
      mux_data4[167:160] = in_data4[2575:2568];
      mux_data4[175:168] = in_data4[2583:2576];
    end
    'd20: begin
      mux_data0[7:0] = in_data0[2543:2536];
      mux_data0[15:8] = in_data0[2551:2544];
      mux_data0[23:16] = in_data0[2559:2552];
      mux_data0[31:24] = in_data0[2567:2560];
      mux_data0[39:32] = in_data0[2575:2568];
      mux_data0[47:40] = in_data0[2583:2576];
      mux_data0[55:48] = in_data0[2591:2584];
      mux_data0[63:56] = in_data0[2599:2592];
      mux_data0[71:64] = in_data0[2607:2600];
      mux_data0[79:72] = in_data0[2615:2608];
      mux_data0[87:80] = in_data0[2623:2616];
      mux_data0[95:88] = in_data0[2631:2624];
      mux_data0[103:96] = in_data0[2639:2632];
      mux_data0[111:104] = in_data0[2647:2640];
      mux_data0[119:112] = in_data0[2655:2648];
      mux_data0[127:120] = in_data0[2663:2656];
      mux_data0[135:128] = in_data0[2671:2664];
      mux_data0[143:136] = in_data0[2679:2672];
      mux_data0[151:144] = in_data0[2687:2680];
      mux_data0[159:152] = in_data0[2695:2688];
      mux_data0[167:160] = in_data0[2703:2696];
      mux_data0[175:168] = in_data0[2711:2704];
      mux_data1[7:0] = in_data1[2543:2536];
      mux_data1[15:8] = in_data1[2551:2544];
      mux_data1[23:16] = in_data1[2559:2552];
      mux_data1[31:24] = in_data1[2567:2560];
      mux_data1[39:32] = in_data1[2575:2568];
      mux_data1[47:40] = in_data1[2583:2576];
      mux_data1[55:48] = in_data1[2591:2584];
      mux_data1[63:56] = in_data1[2599:2592];
      mux_data1[71:64] = in_data1[2607:2600];
      mux_data1[79:72] = in_data1[2615:2608];
      mux_data1[87:80] = in_data1[2623:2616];
      mux_data1[95:88] = in_data1[2631:2624];
      mux_data1[103:96] = in_data1[2639:2632];
      mux_data1[111:104] = in_data1[2647:2640];
      mux_data1[119:112] = in_data1[2655:2648];
      mux_data1[127:120] = in_data1[2663:2656];
      mux_data1[135:128] = in_data1[2671:2664];
      mux_data1[143:136] = in_data1[2679:2672];
      mux_data1[151:144] = in_data1[2687:2680];
      mux_data1[159:152] = in_data1[2695:2688];
      mux_data1[167:160] = in_data1[2703:2696];
      mux_data1[175:168] = in_data1[2711:2704];
      mux_data2[7:0] = in_data2[2543:2536];
      mux_data2[15:8] = in_data2[2551:2544];
      mux_data2[23:16] = in_data2[2559:2552];
      mux_data2[31:24] = in_data2[2567:2560];
      mux_data2[39:32] = in_data2[2575:2568];
      mux_data2[47:40] = in_data2[2583:2576];
      mux_data2[55:48] = in_data2[2591:2584];
      mux_data2[63:56] = in_data2[2599:2592];
      mux_data2[71:64] = in_data2[2607:2600];
      mux_data2[79:72] = in_data2[2615:2608];
      mux_data2[87:80] = in_data2[2623:2616];
      mux_data2[95:88] = in_data2[2631:2624];
      mux_data2[103:96] = in_data2[2639:2632];
      mux_data2[111:104] = in_data2[2647:2640];
      mux_data2[119:112] = in_data2[2655:2648];
      mux_data2[127:120] = in_data2[2663:2656];
      mux_data2[135:128] = in_data2[2671:2664];
      mux_data2[143:136] = in_data2[2679:2672];
      mux_data2[151:144] = in_data2[2687:2680];
      mux_data2[159:152] = in_data2[2695:2688];
      mux_data2[167:160] = in_data2[2703:2696];
      mux_data2[175:168] = in_data2[2711:2704];
      mux_data3[7:0] = in_data3[2543:2536];
      mux_data3[15:8] = in_data3[2551:2544];
      mux_data3[23:16] = in_data3[2559:2552];
      mux_data3[31:24] = in_data3[2567:2560];
      mux_data3[39:32] = in_data3[2575:2568];
      mux_data3[47:40] = in_data3[2583:2576];
      mux_data3[55:48] = in_data3[2591:2584];
      mux_data3[63:56] = in_data3[2599:2592];
      mux_data3[71:64] = in_data3[2607:2600];
      mux_data3[79:72] = in_data3[2615:2608];
      mux_data3[87:80] = in_data3[2623:2616];
      mux_data3[95:88] = in_data3[2631:2624];
      mux_data3[103:96] = in_data3[2639:2632];
      mux_data3[111:104] = in_data3[2647:2640];
      mux_data3[119:112] = in_data3[2655:2648];
      mux_data3[127:120] = in_data3[2663:2656];
      mux_data3[135:128] = in_data3[2671:2664];
      mux_data3[143:136] = in_data3[2679:2672];
      mux_data3[151:144] = in_data3[2687:2680];
      mux_data3[159:152] = in_data3[2695:2688];
      mux_data3[167:160] = in_data3[2703:2696];
      mux_data3[175:168] = in_data3[2711:2704];
      mux_data4[7:0] = in_data4[2543:2536];
      mux_data4[15:8] = in_data4[2551:2544];
      mux_data4[23:16] = in_data4[2559:2552];
      mux_data4[31:24] = in_data4[2567:2560];
      mux_data4[39:32] = in_data4[2575:2568];
      mux_data4[47:40] = in_data4[2583:2576];
      mux_data4[55:48] = in_data4[2591:2584];
      mux_data4[63:56] = in_data4[2599:2592];
      mux_data4[71:64] = in_data4[2607:2600];
      mux_data4[79:72] = in_data4[2615:2608];
      mux_data4[87:80] = in_data4[2623:2616];
      mux_data4[95:88] = in_data4[2631:2624];
      mux_data4[103:96] = in_data4[2639:2632];
      mux_data4[111:104] = in_data4[2647:2640];
      mux_data4[119:112] = in_data4[2655:2648];
      mux_data4[127:120] = in_data4[2663:2656];
      mux_data4[135:128] = in_data4[2671:2664];
      mux_data4[143:136] = in_data4[2679:2672];
      mux_data4[151:144] = in_data4[2687:2680];
      mux_data4[159:152] = in_data4[2695:2688];
      mux_data4[167:160] = in_data4[2703:2696];
      mux_data4[175:168] = in_data4[2711:2704];
    end
    'd21: begin
      mux_data0[7:0] = in_data0[2671:2664];
      mux_data0[15:8] = in_data0[2679:2672];
      mux_data0[23:16] = in_data0[2687:2680];
      mux_data0[31:24] = in_data0[2695:2688];
      mux_data0[39:32] = in_data0[2703:2696];
      mux_data0[47:40] = in_data0[2711:2704];
      mux_data0[55:48] = in_data0[2719:2712];
      mux_data0[63:56] = in_data0[2727:2720];
      mux_data0[71:64] = in_data0[2735:2728];
      mux_data0[79:72] = in_data0[2743:2736];
      mux_data0[87:80] = in_data0[2751:2744];
      mux_data0[95:88] = in_data0[2759:2752];
      mux_data0[103:96] = in_data0[2767:2760];
      mux_data0[111:104] = in_data0[2775:2768];
      mux_data0[119:112] = in_data0[2783:2776];
      mux_data0[127:120] = in_data0[2791:2784];
      mux_data0[135:128] = in_data0[2799:2792];
      mux_data0[143:136] = in_data0[2807:2800];
      mux_data0[151:144] = in_data0[2815:2808];
      mux_data0[159:152] = in_data0[2823:2816];
      mux_data0[167:160] = in_data0[2831:2824];
      mux_data0[175:168] = in_data0[2839:2832];
      mux_data1[7:0] = in_data1[2671:2664];
      mux_data1[15:8] = in_data1[2679:2672];
      mux_data1[23:16] = in_data1[2687:2680];
      mux_data1[31:24] = in_data1[2695:2688];
      mux_data1[39:32] = in_data1[2703:2696];
      mux_data1[47:40] = in_data1[2711:2704];
      mux_data1[55:48] = in_data1[2719:2712];
      mux_data1[63:56] = in_data1[2727:2720];
      mux_data1[71:64] = in_data1[2735:2728];
      mux_data1[79:72] = in_data1[2743:2736];
      mux_data1[87:80] = in_data1[2751:2744];
      mux_data1[95:88] = in_data1[2759:2752];
      mux_data1[103:96] = in_data1[2767:2760];
      mux_data1[111:104] = in_data1[2775:2768];
      mux_data1[119:112] = in_data1[2783:2776];
      mux_data1[127:120] = in_data1[2791:2784];
      mux_data1[135:128] = in_data1[2799:2792];
      mux_data1[143:136] = in_data1[2807:2800];
      mux_data1[151:144] = in_data1[2815:2808];
      mux_data1[159:152] = in_data1[2823:2816];
      mux_data1[167:160] = in_data1[2831:2824];
      mux_data1[175:168] = in_data1[2839:2832];
      mux_data2[7:0] = in_data2[2671:2664];
      mux_data2[15:8] = in_data2[2679:2672];
      mux_data2[23:16] = in_data2[2687:2680];
      mux_data2[31:24] = in_data2[2695:2688];
      mux_data2[39:32] = in_data2[2703:2696];
      mux_data2[47:40] = in_data2[2711:2704];
      mux_data2[55:48] = in_data2[2719:2712];
      mux_data2[63:56] = in_data2[2727:2720];
      mux_data2[71:64] = in_data2[2735:2728];
      mux_data2[79:72] = in_data2[2743:2736];
      mux_data2[87:80] = in_data2[2751:2744];
      mux_data2[95:88] = in_data2[2759:2752];
      mux_data2[103:96] = in_data2[2767:2760];
      mux_data2[111:104] = in_data2[2775:2768];
      mux_data2[119:112] = in_data2[2783:2776];
      mux_data2[127:120] = in_data2[2791:2784];
      mux_data2[135:128] = in_data2[2799:2792];
      mux_data2[143:136] = in_data2[2807:2800];
      mux_data2[151:144] = in_data2[2815:2808];
      mux_data2[159:152] = in_data2[2823:2816];
      mux_data2[167:160] = in_data2[2831:2824];
      mux_data2[175:168] = in_data2[2839:2832];
      mux_data3[7:0] = in_data3[2671:2664];
      mux_data3[15:8] = in_data3[2679:2672];
      mux_data3[23:16] = in_data3[2687:2680];
      mux_data3[31:24] = in_data3[2695:2688];
      mux_data3[39:32] = in_data3[2703:2696];
      mux_data3[47:40] = in_data3[2711:2704];
      mux_data3[55:48] = in_data3[2719:2712];
      mux_data3[63:56] = in_data3[2727:2720];
      mux_data3[71:64] = in_data3[2735:2728];
      mux_data3[79:72] = in_data3[2743:2736];
      mux_data3[87:80] = in_data3[2751:2744];
      mux_data3[95:88] = in_data3[2759:2752];
      mux_data3[103:96] = in_data3[2767:2760];
      mux_data3[111:104] = in_data3[2775:2768];
      mux_data3[119:112] = in_data3[2783:2776];
      mux_data3[127:120] = in_data3[2791:2784];
      mux_data3[135:128] = in_data3[2799:2792];
      mux_data3[143:136] = in_data3[2807:2800];
      mux_data3[151:144] = in_data3[2815:2808];
      mux_data3[159:152] = in_data3[2823:2816];
      mux_data3[167:160] = in_data3[2831:2824];
      mux_data3[175:168] = in_data3[2839:2832];
      mux_data4[7:0] = in_data4[2671:2664];
      mux_data4[15:8] = in_data4[2679:2672];
      mux_data4[23:16] = in_data4[2687:2680];
      mux_data4[31:24] = in_data4[2695:2688];
      mux_data4[39:32] = in_data4[2703:2696];
      mux_data4[47:40] = in_data4[2711:2704];
      mux_data4[55:48] = in_data4[2719:2712];
      mux_data4[63:56] = in_data4[2727:2720];
      mux_data4[71:64] = in_data4[2735:2728];
      mux_data4[79:72] = in_data4[2743:2736];
      mux_data4[87:80] = in_data4[2751:2744];
      mux_data4[95:88] = in_data4[2759:2752];
      mux_data4[103:96] = in_data4[2767:2760];
      mux_data4[111:104] = in_data4[2775:2768];
      mux_data4[119:112] = in_data4[2783:2776];
      mux_data4[127:120] = in_data4[2791:2784];
      mux_data4[135:128] = in_data4[2799:2792];
      mux_data4[143:136] = in_data4[2807:2800];
      mux_data4[151:144] = in_data4[2815:2808];
      mux_data4[159:152] = in_data4[2823:2816];
      mux_data4[167:160] = in_data4[2831:2824];
      mux_data4[175:168] = in_data4[2839:2832];
    end
    'd22: begin
      mux_data0[7:0] = in_data0[2799:2792];
      mux_data0[15:8] = in_data0[2807:2800];
      mux_data0[23:16] = in_data0[2815:2808];
      mux_data0[31:24] = in_data0[2823:2816];
      mux_data0[39:32] = in_data0[2831:2824];
      mux_data0[47:40] = in_data0[2839:2832];
      mux_data0[55:48] = in_data0[2847:2840];
      mux_data0[63:56] = in_data0[2855:2848];
      mux_data0[71:64] = in_data0[2863:2856];
      mux_data0[79:72] = in_data0[2871:2864];
      mux_data0[87:80] = in_data0[2879:2872];
      mux_data0[95:88] = in_data0[2887:2880];
      mux_data0[103:96] = in_data0[2895:2888];
      mux_data0[111:104] = in_data0[2903:2896];
      mux_data0[119:112] = in_data0[2911:2904];
      mux_data0[127:120] = in_data0[2919:2912];
      mux_data0[135:128] = in_data0[2927:2920];
      mux_data0[143:136] = in_data0[2935:2928];
      mux_data0[151:144] = in_data0[2943:2936];
      mux_data0[159:152] = in_data0[2951:2944];
      mux_data0[167:160] = in_data0[2959:2952];
      mux_data0[175:168] = in_data0[2967:2960];
      mux_data1[7:0] = in_data1[2799:2792];
      mux_data1[15:8] = in_data1[2807:2800];
      mux_data1[23:16] = in_data1[2815:2808];
      mux_data1[31:24] = in_data1[2823:2816];
      mux_data1[39:32] = in_data1[2831:2824];
      mux_data1[47:40] = in_data1[2839:2832];
      mux_data1[55:48] = in_data1[2847:2840];
      mux_data1[63:56] = in_data1[2855:2848];
      mux_data1[71:64] = in_data1[2863:2856];
      mux_data1[79:72] = in_data1[2871:2864];
      mux_data1[87:80] = in_data1[2879:2872];
      mux_data1[95:88] = in_data1[2887:2880];
      mux_data1[103:96] = in_data1[2895:2888];
      mux_data1[111:104] = in_data1[2903:2896];
      mux_data1[119:112] = in_data1[2911:2904];
      mux_data1[127:120] = in_data1[2919:2912];
      mux_data1[135:128] = in_data1[2927:2920];
      mux_data1[143:136] = in_data1[2935:2928];
      mux_data1[151:144] = in_data1[2943:2936];
      mux_data1[159:152] = in_data1[2951:2944];
      mux_data1[167:160] = in_data1[2959:2952];
      mux_data1[175:168] = in_data1[2967:2960];
      mux_data2[7:0] = in_data2[2799:2792];
      mux_data2[15:8] = in_data2[2807:2800];
      mux_data2[23:16] = in_data2[2815:2808];
      mux_data2[31:24] = in_data2[2823:2816];
      mux_data2[39:32] = in_data2[2831:2824];
      mux_data2[47:40] = in_data2[2839:2832];
      mux_data2[55:48] = in_data2[2847:2840];
      mux_data2[63:56] = in_data2[2855:2848];
      mux_data2[71:64] = in_data2[2863:2856];
      mux_data2[79:72] = in_data2[2871:2864];
      mux_data2[87:80] = in_data2[2879:2872];
      mux_data2[95:88] = in_data2[2887:2880];
      mux_data2[103:96] = in_data2[2895:2888];
      mux_data2[111:104] = in_data2[2903:2896];
      mux_data2[119:112] = in_data2[2911:2904];
      mux_data2[127:120] = in_data2[2919:2912];
      mux_data2[135:128] = in_data2[2927:2920];
      mux_data2[143:136] = in_data2[2935:2928];
      mux_data2[151:144] = in_data2[2943:2936];
      mux_data2[159:152] = in_data2[2951:2944];
      mux_data2[167:160] = in_data2[2959:2952];
      mux_data2[175:168] = in_data2[2967:2960];
      mux_data3[7:0] = in_data3[2799:2792];
      mux_data3[15:8] = in_data3[2807:2800];
      mux_data3[23:16] = in_data3[2815:2808];
      mux_data3[31:24] = in_data3[2823:2816];
      mux_data3[39:32] = in_data3[2831:2824];
      mux_data3[47:40] = in_data3[2839:2832];
      mux_data3[55:48] = in_data3[2847:2840];
      mux_data3[63:56] = in_data3[2855:2848];
      mux_data3[71:64] = in_data3[2863:2856];
      mux_data3[79:72] = in_data3[2871:2864];
      mux_data3[87:80] = in_data3[2879:2872];
      mux_data3[95:88] = in_data3[2887:2880];
      mux_data3[103:96] = in_data3[2895:2888];
      mux_data3[111:104] = in_data3[2903:2896];
      mux_data3[119:112] = in_data3[2911:2904];
      mux_data3[127:120] = in_data3[2919:2912];
      mux_data3[135:128] = in_data3[2927:2920];
      mux_data3[143:136] = in_data3[2935:2928];
      mux_data3[151:144] = in_data3[2943:2936];
      mux_data3[159:152] = in_data3[2951:2944];
      mux_data3[167:160] = in_data3[2959:2952];
      mux_data3[175:168] = in_data3[2967:2960];
      mux_data4[7:0] = in_data4[2799:2792];
      mux_data4[15:8] = in_data4[2807:2800];
      mux_data4[23:16] = in_data4[2815:2808];
      mux_data4[31:24] = in_data4[2823:2816];
      mux_data4[39:32] = in_data4[2831:2824];
      mux_data4[47:40] = in_data4[2839:2832];
      mux_data4[55:48] = in_data4[2847:2840];
      mux_data4[63:56] = in_data4[2855:2848];
      mux_data4[71:64] = in_data4[2863:2856];
      mux_data4[79:72] = in_data4[2871:2864];
      mux_data4[87:80] = in_data4[2879:2872];
      mux_data4[95:88] = in_data4[2887:2880];
      mux_data4[103:96] = in_data4[2895:2888];
      mux_data4[111:104] = in_data4[2903:2896];
      mux_data4[119:112] = in_data4[2911:2904];
      mux_data4[127:120] = in_data4[2919:2912];
      mux_data4[135:128] = in_data4[2927:2920];
      mux_data4[143:136] = in_data4[2935:2928];
      mux_data4[151:144] = in_data4[2943:2936];
      mux_data4[159:152] = in_data4[2951:2944];
      mux_data4[167:160] = in_data4[2959:2952];
      mux_data4[175:168] = in_data4[2967:2960];
    end
    'd23: begin
      mux_data0[7:0] = in_data0[2927:2920];
      mux_data0[15:8] = in_data0[2935:2928];
      mux_data0[23:16] = in_data0[2943:2936];
      mux_data0[31:24] = in_data0[2951:2944];
      mux_data0[39:32] = in_data0[2959:2952];
      mux_data0[47:40] = in_data0[2967:2960];
      mux_data0[55:48] = in_data0[2975:2968];
      mux_data0[63:56] = in_data0[2983:2976];
      mux_data0[71:64] = in_data0[2991:2984];
      mux_data0[79:72] = in_data0[2999:2992];
      mux_data0[87:80] = in_data0[3007:3000];
      mux_data0[95:88] = in_data0[3015:3008];
      mux_data0[103:96] = in_data0[3023:3016];
      mux_data0[111:104] = in_data0[3031:3024];
      mux_data0[119:112] = in_data0[3039:3032];
      mux_data0[127:120] = in_data0[3047:3040];
      mux_data0[135:128] = in_data0[3055:3048];
      mux_data0[143:136] = in_data0[3063:3056];
      mux_data0[151:144] = in_data0[3071:3064];
      mux_data0[159:152] = in_data0[3079:3072];
      mux_data0[167:160] = in_data0[3087:3080];
      mux_data0[175:168] = in_data0[3095:3088];
      mux_data1[7:0] = in_data1[2927:2920];
      mux_data1[15:8] = in_data1[2935:2928];
      mux_data1[23:16] = in_data1[2943:2936];
      mux_data1[31:24] = in_data1[2951:2944];
      mux_data1[39:32] = in_data1[2959:2952];
      mux_data1[47:40] = in_data1[2967:2960];
      mux_data1[55:48] = in_data1[2975:2968];
      mux_data1[63:56] = in_data1[2983:2976];
      mux_data1[71:64] = in_data1[2991:2984];
      mux_data1[79:72] = in_data1[2999:2992];
      mux_data1[87:80] = in_data1[3007:3000];
      mux_data1[95:88] = in_data1[3015:3008];
      mux_data1[103:96] = in_data1[3023:3016];
      mux_data1[111:104] = in_data1[3031:3024];
      mux_data1[119:112] = in_data1[3039:3032];
      mux_data1[127:120] = in_data1[3047:3040];
      mux_data1[135:128] = in_data1[3055:3048];
      mux_data1[143:136] = in_data1[3063:3056];
      mux_data1[151:144] = in_data1[3071:3064];
      mux_data1[159:152] = in_data1[3079:3072];
      mux_data1[167:160] = in_data1[3087:3080];
      mux_data1[175:168] = in_data1[3095:3088];
      mux_data2[7:0] = in_data2[2927:2920];
      mux_data2[15:8] = in_data2[2935:2928];
      mux_data2[23:16] = in_data2[2943:2936];
      mux_data2[31:24] = in_data2[2951:2944];
      mux_data2[39:32] = in_data2[2959:2952];
      mux_data2[47:40] = in_data2[2967:2960];
      mux_data2[55:48] = in_data2[2975:2968];
      mux_data2[63:56] = in_data2[2983:2976];
      mux_data2[71:64] = in_data2[2991:2984];
      mux_data2[79:72] = in_data2[2999:2992];
      mux_data2[87:80] = in_data2[3007:3000];
      mux_data2[95:88] = in_data2[3015:3008];
      mux_data2[103:96] = in_data2[3023:3016];
      mux_data2[111:104] = in_data2[3031:3024];
      mux_data2[119:112] = in_data2[3039:3032];
      mux_data2[127:120] = in_data2[3047:3040];
      mux_data2[135:128] = in_data2[3055:3048];
      mux_data2[143:136] = in_data2[3063:3056];
      mux_data2[151:144] = in_data2[3071:3064];
      mux_data2[159:152] = in_data2[3079:3072];
      mux_data2[167:160] = in_data2[3087:3080];
      mux_data2[175:168] = in_data2[3095:3088];
      mux_data3[7:0] = in_data3[2927:2920];
      mux_data3[15:8] = in_data3[2935:2928];
      mux_data3[23:16] = in_data3[2943:2936];
      mux_data3[31:24] = in_data3[2951:2944];
      mux_data3[39:32] = in_data3[2959:2952];
      mux_data3[47:40] = in_data3[2967:2960];
      mux_data3[55:48] = in_data3[2975:2968];
      mux_data3[63:56] = in_data3[2983:2976];
      mux_data3[71:64] = in_data3[2991:2984];
      mux_data3[79:72] = in_data3[2999:2992];
      mux_data3[87:80] = in_data3[3007:3000];
      mux_data3[95:88] = in_data3[3015:3008];
      mux_data3[103:96] = in_data3[3023:3016];
      mux_data3[111:104] = in_data3[3031:3024];
      mux_data3[119:112] = in_data3[3039:3032];
      mux_data3[127:120] = in_data3[3047:3040];
      mux_data3[135:128] = in_data3[3055:3048];
      mux_data3[143:136] = in_data3[3063:3056];
      mux_data3[151:144] = in_data3[3071:3064];
      mux_data3[159:152] = in_data3[3079:3072];
      mux_data3[167:160] = in_data3[3087:3080];
      mux_data3[175:168] = in_data3[3095:3088];
      mux_data4[7:0] = in_data4[2927:2920];
      mux_data4[15:8] = in_data4[2935:2928];
      mux_data4[23:16] = in_data4[2943:2936];
      mux_data4[31:24] = in_data4[2951:2944];
      mux_data4[39:32] = in_data4[2959:2952];
      mux_data4[47:40] = in_data4[2967:2960];
      mux_data4[55:48] = in_data4[2975:2968];
      mux_data4[63:56] = in_data4[2983:2976];
      mux_data4[71:64] = in_data4[2991:2984];
      mux_data4[79:72] = in_data4[2999:2992];
      mux_data4[87:80] = in_data4[3007:3000];
      mux_data4[95:88] = in_data4[3015:3008];
      mux_data4[103:96] = in_data4[3023:3016];
      mux_data4[111:104] = in_data4[3031:3024];
      mux_data4[119:112] = in_data4[3039:3032];
      mux_data4[127:120] = in_data4[3047:3040];
      mux_data4[135:128] = in_data4[3055:3048];
      mux_data4[143:136] = in_data4[3063:3056];
      mux_data4[151:144] = in_data4[3071:3064];
      mux_data4[159:152] = in_data4[3079:3072];
      mux_data4[167:160] = in_data4[3087:3080];
      mux_data4[175:168] = in_data4[3095:3088];
    end
    'd24: begin
      mux_data0[7:0] = in_data0[3055:3048];
      mux_data0[15:8] = in_data0[3063:3056];
      mux_data0[23:16] = in_data0[3071:3064];
      mux_data0[31:24] = in_data0[3079:3072];
      mux_data0[39:32] = in_data0[3087:3080];
      mux_data0[47:40] = in_data0[3095:3088];
      mux_data0[55:48] = in_data0[3103:3096];
      mux_data0[63:56] = in_data0[3111:3104];
      mux_data0[71:64] = in_data0[3119:3112];
      mux_data0[79:72] = in_data0[3127:3120];
      mux_data0[87:80] = in_data0[3135:3128];
      mux_data0[95:88] = in_data0[3143:3136];
      mux_data0[103:96] = in_data0[3151:3144];
      mux_data0[111:104] = in_data0[3159:3152];
      mux_data0[119:112] = in_data0[3167:3160];
      mux_data0[127:120] = in_data0[3175:3168];
      mux_data0[135:128] = in_data0[3183:3176];
      mux_data0[143:136] = in_data0[3191:3184];
      mux_data0[151:144] = in_data0[3199:3192];
      mux_data0[159:152] = in_data0[3207:3200];
      mux_data0[167:160] = in_data0[3215:3208];
      mux_data0[175:168] = in_data0[3223:3216];
      mux_data1[7:0] = in_data1[3055:3048];
      mux_data1[15:8] = in_data1[3063:3056];
      mux_data1[23:16] = in_data1[3071:3064];
      mux_data1[31:24] = in_data1[3079:3072];
      mux_data1[39:32] = in_data1[3087:3080];
      mux_data1[47:40] = in_data1[3095:3088];
      mux_data1[55:48] = in_data1[3103:3096];
      mux_data1[63:56] = in_data1[3111:3104];
      mux_data1[71:64] = in_data1[3119:3112];
      mux_data1[79:72] = in_data1[3127:3120];
      mux_data1[87:80] = in_data1[3135:3128];
      mux_data1[95:88] = in_data1[3143:3136];
      mux_data1[103:96] = in_data1[3151:3144];
      mux_data1[111:104] = in_data1[3159:3152];
      mux_data1[119:112] = in_data1[3167:3160];
      mux_data1[127:120] = in_data1[3175:3168];
      mux_data1[135:128] = in_data1[3183:3176];
      mux_data1[143:136] = in_data1[3191:3184];
      mux_data1[151:144] = in_data1[3199:3192];
      mux_data1[159:152] = in_data1[3207:3200];
      mux_data1[167:160] = in_data1[3215:3208];
      mux_data1[175:168] = in_data1[3223:3216];
      mux_data2[7:0] = in_data2[3055:3048];
      mux_data2[15:8] = in_data2[3063:3056];
      mux_data2[23:16] = in_data2[3071:3064];
      mux_data2[31:24] = in_data2[3079:3072];
      mux_data2[39:32] = in_data2[3087:3080];
      mux_data2[47:40] = in_data2[3095:3088];
      mux_data2[55:48] = in_data2[3103:3096];
      mux_data2[63:56] = in_data2[3111:3104];
      mux_data2[71:64] = in_data2[3119:3112];
      mux_data2[79:72] = in_data2[3127:3120];
      mux_data2[87:80] = in_data2[3135:3128];
      mux_data2[95:88] = in_data2[3143:3136];
      mux_data2[103:96] = in_data2[3151:3144];
      mux_data2[111:104] = in_data2[3159:3152];
      mux_data2[119:112] = in_data2[3167:3160];
      mux_data2[127:120] = in_data2[3175:3168];
      mux_data2[135:128] = in_data2[3183:3176];
      mux_data2[143:136] = in_data2[3191:3184];
      mux_data2[151:144] = in_data2[3199:3192];
      mux_data2[159:152] = in_data2[3207:3200];
      mux_data2[167:160] = in_data2[3215:3208];
      mux_data2[175:168] = in_data2[3223:3216];
      mux_data3[7:0] = in_data3[3055:3048];
      mux_data3[15:8] = in_data3[3063:3056];
      mux_data3[23:16] = in_data3[3071:3064];
      mux_data3[31:24] = in_data3[3079:3072];
      mux_data3[39:32] = in_data3[3087:3080];
      mux_data3[47:40] = in_data3[3095:3088];
      mux_data3[55:48] = in_data3[3103:3096];
      mux_data3[63:56] = in_data3[3111:3104];
      mux_data3[71:64] = in_data3[3119:3112];
      mux_data3[79:72] = in_data3[3127:3120];
      mux_data3[87:80] = in_data3[3135:3128];
      mux_data3[95:88] = in_data3[3143:3136];
      mux_data3[103:96] = in_data3[3151:3144];
      mux_data3[111:104] = in_data3[3159:3152];
      mux_data3[119:112] = in_data3[3167:3160];
      mux_data3[127:120] = in_data3[3175:3168];
      mux_data3[135:128] = in_data3[3183:3176];
      mux_data3[143:136] = in_data3[3191:3184];
      mux_data3[151:144] = in_data3[3199:3192];
      mux_data3[159:152] = in_data3[3207:3200];
      mux_data3[167:160] = in_data3[3215:3208];
      mux_data3[175:168] = in_data3[3223:3216];
      mux_data4[7:0] = in_data4[3055:3048];
      mux_data4[15:8] = in_data4[3063:3056];
      mux_data4[23:16] = in_data4[3071:3064];
      mux_data4[31:24] = in_data4[3079:3072];
      mux_data4[39:32] = in_data4[3087:3080];
      mux_data4[47:40] = in_data4[3095:3088];
      mux_data4[55:48] = in_data4[3103:3096];
      mux_data4[63:56] = in_data4[3111:3104];
      mux_data4[71:64] = in_data4[3119:3112];
      mux_data4[79:72] = in_data4[3127:3120];
      mux_data4[87:80] = in_data4[3135:3128];
      mux_data4[95:88] = in_data4[3143:3136];
      mux_data4[103:96] = in_data4[3151:3144];
      mux_data4[111:104] = in_data4[3159:3152];
      mux_data4[119:112] = in_data4[3167:3160];
      mux_data4[127:120] = in_data4[3175:3168];
      mux_data4[135:128] = in_data4[3183:3176];
      mux_data4[143:136] = in_data4[3191:3184];
      mux_data4[151:144] = in_data4[3199:3192];
      mux_data4[159:152] = in_data4[3207:3200];
      mux_data4[167:160] = in_data4[3215:3208];
      mux_data4[175:168] = in_data4[3223:3216];
    end
    'd25: begin
      mux_data0[7:0] = in_data0[3183:3176];
      mux_data0[15:8] = in_data0[3191:3184];
      mux_data0[23:16] = in_data0[3199:3192];
      mux_data0[31:24] = in_data0[3207:3200];
      mux_data0[39:32] = in_data0[3215:3208];
      mux_data0[47:40] = in_data0[3223:3216];
      mux_data0[55:48] = in_data0[3231:3224];
      mux_data0[63:56] = in_data0[3239:3232];
      mux_data0[71:64] = in_data0[3247:3240];
      mux_data0[79:72] = in_data0[3255:3248];
      mux_data0[87:80] = in_data0[3263:3256];
      mux_data0[95:88] = in_data0[3271:3264];
      mux_data0[103:96] = in_data0[3279:3272];
      mux_data0[111:104] = in_data0[3287:3280];
      mux_data0[119:112] = in_data0[3295:3288];
      mux_data0[127:120] = in_data0[3303:3296];
      mux_data0[135:128] = in_data0[3311:3304];
      mux_data0[143:136] = in_data0[3319:3312];
      mux_data0[151:144] = in_data0[3327:3320];
      mux_data0[159:152] = in_data0[3335:3328];
      mux_data0[167:160] = in_data0[3343:3336];
      mux_data0[175:168] = in_data0[3351:3344];
      mux_data1[7:0] = in_data1[3183:3176];
      mux_data1[15:8] = in_data1[3191:3184];
      mux_data1[23:16] = in_data1[3199:3192];
      mux_data1[31:24] = in_data1[3207:3200];
      mux_data1[39:32] = in_data1[3215:3208];
      mux_data1[47:40] = in_data1[3223:3216];
      mux_data1[55:48] = in_data1[3231:3224];
      mux_data1[63:56] = in_data1[3239:3232];
      mux_data1[71:64] = in_data1[3247:3240];
      mux_data1[79:72] = in_data1[3255:3248];
      mux_data1[87:80] = in_data1[3263:3256];
      mux_data1[95:88] = in_data1[3271:3264];
      mux_data1[103:96] = in_data1[3279:3272];
      mux_data1[111:104] = in_data1[3287:3280];
      mux_data1[119:112] = in_data1[3295:3288];
      mux_data1[127:120] = in_data1[3303:3296];
      mux_data1[135:128] = in_data1[3311:3304];
      mux_data1[143:136] = in_data1[3319:3312];
      mux_data1[151:144] = in_data1[3327:3320];
      mux_data1[159:152] = in_data1[3335:3328];
      mux_data1[167:160] = in_data1[3343:3336];
      mux_data1[175:168] = in_data1[3351:3344];
      mux_data2[7:0] = in_data2[3183:3176];
      mux_data2[15:8] = in_data2[3191:3184];
      mux_data2[23:16] = in_data2[3199:3192];
      mux_data2[31:24] = in_data2[3207:3200];
      mux_data2[39:32] = in_data2[3215:3208];
      mux_data2[47:40] = in_data2[3223:3216];
      mux_data2[55:48] = in_data2[3231:3224];
      mux_data2[63:56] = in_data2[3239:3232];
      mux_data2[71:64] = in_data2[3247:3240];
      mux_data2[79:72] = in_data2[3255:3248];
      mux_data2[87:80] = in_data2[3263:3256];
      mux_data2[95:88] = in_data2[3271:3264];
      mux_data2[103:96] = in_data2[3279:3272];
      mux_data2[111:104] = in_data2[3287:3280];
      mux_data2[119:112] = in_data2[3295:3288];
      mux_data2[127:120] = in_data2[3303:3296];
      mux_data2[135:128] = in_data2[3311:3304];
      mux_data2[143:136] = in_data2[3319:3312];
      mux_data2[151:144] = in_data2[3327:3320];
      mux_data2[159:152] = in_data2[3335:3328];
      mux_data2[167:160] = in_data2[3343:3336];
      mux_data2[175:168] = in_data2[3351:3344];
      mux_data3[7:0] = in_data3[3183:3176];
      mux_data3[15:8] = in_data3[3191:3184];
      mux_data3[23:16] = in_data3[3199:3192];
      mux_data3[31:24] = in_data3[3207:3200];
      mux_data3[39:32] = in_data3[3215:3208];
      mux_data3[47:40] = in_data3[3223:3216];
      mux_data3[55:48] = in_data3[3231:3224];
      mux_data3[63:56] = in_data3[3239:3232];
      mux_data3[71:64] = in_data3[3247:3240];
      mux_data3[79:72] = in_data3[3255:3248];
      mux_data3[87:80] = in_data3[3263:3256];
      mux_data3[95:88] = in_data3[3271:3264];
      mux_data3[103:96] = in_data3[3279:3272];
      mux_data3[111:104] = in_data3[3287:3280];
      mux_data3[119:112] = in_data3[3295:3288];
      mux_data3[127:120] = in_data3[3303:3296];
      mux_data3[135:128] = in_data3[3311:3304];
      mux_data3[143:136] = in_data3[3319:3312];
      mux_data3[151:144] = in_data3[3327:3320];
      mux_data3[159:152] = in_data3[3335:3328];
      mux_data3[167:160] = in_data3[3343:3336];
      mux_data3[175:168] = in_data3[3351:3344];
      mux_data4[7:0] = in_data4[3183:3176];
      mux_data4[15:8] = in_data4[3191:3184];
      mux_data4[23:16] = in_data4[3199:3192];
      mux_data4[31:24] = in_data4[3207:3200];
      mux_data4[39:32] = in_data4[3215:3208];
      mux_data4[47:40] = in_data4[3223:3216];
      mux_data4[55:48] = in_data4[3231:3224];
      mux_data4[63:56] = in_data4[3239:3232];
      mux_data4[71:64] = in_data4[3247:3240];
      mux_data4[79:72] = in_data4[3255:3248];
      mux_data4[87:80] = in_data4[3263:3256];
      mux_data4[95:88] = in_data4[3271:3264];
      mux_data4[103:96] = in_data4[3279:3272];
      mux_data4[111:104] = in_data4[3287:3280];
      mux_data4[119:112] = in_data4[3295:3288];
      mux_data4[127:120] = in_data4[3303:3296];
      mux_data4[135:128] = in_data4[3311:3304];
      mux_data4[143:136] = in_data4[3319:3312];
      mux_data4[151:144] = in_data4[3327:3320];
      mux_data4[159:152] = in_data4[3335:3328];
      mux_data4[167:160] = in_data4[3343:3336];
      mux_data4[175:168] = in_data4[3351:3344];
    end
    'd26: begin
      mux_data0[7:0] = in_data0[3311:3304];
      mux_data0[15:8] = in_data0[3319:3312];
      mux_data0[23:16] = in_data0[3327:3320];
      mux_data0[31:24] = in_data0[3335:3328];
      mux_data0[39:32] = in_data0[3343:3336];
      mux_data0[47:40] = in_data0[3351:3344];
      mux_data0[55:48] = in_data0[3359:3352];
      mux_data0[63:56] = in_data0[3367:3360];
      mux_data0[71:64] = in_data0[3375:3368];
      mux_data0[79:72] = in_data0[3383:3376];
      mux_data0[87:80] = in_data0[3391:3384];
      mux_data0[95:88] = in_data0[3399:3392];
      mux_data0[103:96] = in_data0[3407:3400];
      mux_data0[111:104] = in_data0[3415:3408];
      mux_data0[119:112] = in_data0[3423:3416];
      mux_data0[127:120] = in_data0[3431:3424];
      mux_data0[135:128] = in_data0[3439:3432];
      mux_data0[143:136] = in_data0[3447:3440];
      mux_data0[151:144] = in_data0[3455:3448];
      mux_data0[159:152] = in_data0[3463:3456];
      mux_data0[167:160] = in_data0[3471:3464];
      mux_data0[175:168] = in_data0[3479:3472];
      mux_data1[7:0] = in_data1[3311:3304];
      mux_data1[15:8] = in_data1[3319:3312];
      mux_data1[23:16] = in_data1[3327:3320];
      mux_data1[31:24] = in_data1[3335:3328];
      mux_data1[39:32] = in_data1[3343:3336];
      mux_data1[47:40] = in_data1[3351:3344];
      mux_data1[55:48] = in_data1[3359:3352];
      mux_data1[63:56] = in_data1[3367:3360];
      mux_data1[71:64] = in_data1[3375:3368];
      mux_data1[79:72] = in_data1[3383:3376];
      mux_data1[87:80] = in_data1[3391:3384];
      mux_data1[95:88] = in_data1[3399:3392];
      mux_data1[103:96] = in_data1[3407:3400];
      mux_data1[111:104] = in_data1[3415:3408];
      mux_data1[119:112] = in_data1[3423:3416];
      mux_data1[127:120] = in_data1[3431:3424];
      mux_data1[135:128] = in_data1[3439:3432];
      mux_data1[143:136] = in_data1[3447:3440];
      mux_data1[151:144] = in_data1[3455:3448];
      mux_data1[159:152] = in_data1[3463:3456];
      mux_data1[167:160] = in_data1[3471:3464];
      mux_data1[175:168] = in_data1[3479:3472];
      mux_data2[7:0] = in_data2[3311:3304];
      mux_data2[15:8] = in_data2[3319:3312];
      mux_data2[23:16] = in_data2[3327:3320];
      mux_data2[31:24] = in_data2[3335:3328];
      mux_data2[39:32] = in_data2[3343:3336];
      mux_data2[47:40] = in_data2[3351:3344];
      mux_data2[55:48] = in_data2[3359:3352];
      mux_data2[63:56] = in_data2[3367:3360];
      mux_data2[71:64] = in_data2[3375:3368];
      mux_data2[79:72] = in_data2[3383:3376];
      mux_data2[87:80] = in_data2[3391:3384];
      mux_data2[95:88] = in_data2[3399:3392];
      mux_data2[103:96] = in_data2[3407:3400];
      mux_data2[111:104] = in_data2[3415:3408];
      mux_data2[119:112] = in_data2[3423:3416];
      mux_data2[127:120] = in_data2[3431:3424];
      mux_data2[135:128] = in_data2[3439:3432];
      mux_data2[143:136] = in_data2[3447:3440];
      mux_data2[151:144] = in_data2[3455:3448];
      mux_data2[159:152] = in_data2[3463:3456];
      mux_data2[167:160] = in_data2[3471:3464];
      mux_data2[175:168] = in_data2[3479:3472];
      mux_data3[7:0] = in_data3[3311:3304];
      mux_data3[15:8] = in_data3[3319:3312];
      mux_data3[23:16] = in_data3[3327:3320];
      mux_data3[31:24] = in_data3[3335:3328];
      mux_data3[39:32] = in_data3[3343:3336];
      mux_data3[47:40] = in_data3[3351:3344];
      mux_data3[55:48] = in_data3[3359:3352];
      mux_data3[63:56] = in_data3[3367:3360];
      mux_data3[71:64] = in_data3[3375:3368];
      mux_data3[79:72] = in_data3[3383:3376];
      mux_data3[87:80] = in_data3[3391:3384];
      mux_data3[95:88] = in_data3[3399:3392];
      mux_data3[103:96] = in_data3[3407:3400];
      mux_data3[111:104] = in_data3[3415:3408];
      mux_data3[119:112] = in_data3[3423:3416];
      mux_data3[127:120] = in_data3[3431:3424];
      mux_data3[135:128] = in_data3[3439:3432];
      mux_data3[143:136] = in_data3[3447:3440];
      mux_data3[151:144] = in_data3[3455:3448];
      mux_data3[159:152] = in_data3[3463:3456];
      mux_data3[167:160] = in_data3[3471:3464];
      mux_data3[175:168] = in_data3[3479:3472];
      mux_data4[7:0] = in_data4[3311:3304];
      mux_data4[15:8] = in_data4[3319:3312];
      mux_data4[23:16] = in_data4[3327:3320];
      mux_data4[31:24] = in_data4[3335:3328];
      mux_data4[39:32] = in_data4[3343:3336];
      mux_data4[47:40] = in_data4[3351:3344];
      mux_data4[55:48] = in_data4[3359:3352];
      mux_data4[63:56] = in_data4[3367:3360];
      mux_data4[71:64] = in_data4[3375:3368];
      mux_data4[79:72] = in_data4[3383:3376];
      mux_data4[87:80] = in_data4[3391:3384];
      mux_data4[95:88] = in_data4[3399:3392];
      mux_data4[103:96] = in_data4[3407:3400];
      mux_data4[111:104] = in_data4[3415:3408];
      mux_data4[119:112] = in_data4[3423:3416];
      mux_data4[127:120] = in_data4[3431:3424];
      mux_data4[135:128] = in_data4[3439:3432];
      mux_data4[143:136] = in_data4[3447:3440];
      mux_data4[151:144] = in_data4[3455:3448];
      mux_data4[159:152] = in_data4[3463:3456];
      mux_data4[167:160] = in_data4[3471:3464];
      mux_data4[175:168] = in_data4[3479:3472];
    end
    'd27: begin
      mux_data0[7:0] = in_data0[3439:3432];
      mux_data0[15:8] = in_data0[3447:3440];
      mux_data0[23:16] = in_data0[3455:3448];
      mux_data0[31:24] = in_data0[3463:3456];
      mux_data0[39:32] = in_data0[3471:3464];
      mux_data0[47:40] = in_data0[3479:3472];
      mux_data0[55:48] = in_data0[3487:3480];
      mux_data0[63:56] = in_data0[3495:3488];
      mux_data0[71:64] = in_data0[3503:3496];
      mux_data0[79:72] = in_data0[3511:3504];
      mux_data0[87:80] = in_data0[3519:3512];
      mux_data0[95:88] = in_data0[3527:3520];
      mux_data0[103:96] = in_data0[3535:3528];
      mux_data0[111:104] = in_data0[3543:3536];
      mux_data0[119:112] = in_data0[3551:3544];
      mux_data0[127:120] = in_data0[3559:3552];
      mux_data0[135:128] = in_data0[3567:3560];
      mux_data0[143:136] = in_data0[3575:3568];
      mux_data0[151:144] = in_data0[3583:3576];
      mux_data0[159:152] = in_data0[3591:3584];
      mux_data0[167:160] = in_data0[3599:3592];
      mux_data0[175:168] = in_data0[3607:3600];
      mux_data1[7:0] = in_data1[3439:3432];
      mux_data1[15:8] = in_data1[3447:3440];
      mux_data1[23:16] = in_data1[3455:3448];
      mux_data1[31:24] = in_data1[3463:3456];
      mux_data1[39:32] = in_data1[3471:3464];
      mux_data1[47:40] = in_data1[3479:3472];
      mux_data1[55:48] = in_data1[3487:3480];
      mux_data1[63:56] = in_data1[3495:3488];
      mux_data1[71:64] = in_data1[3503:3496];
      mux_data1[79:72] = in_data1[3511:3504];
      mux_data1[87:80] = in_data1[3519:3512];
      mux_data1[95:88] = in_data1[3527:3520];
      mux_data1[103:96] = in_data1[3535:3528];
      mux_data1[111:104] = in_data1[3543:3536];
      mux_data1[119:112] = in_data1[3551:3544];
      mux_data1[127:120] = in_data1[3559:3552];
      mux_data1[135:128] = in_data1[3567:3560];
      mux_data1[143:136] = in_data1[3575:3568];
      mux_data1[151:144] = in_data1[3583:3576];
      mux_data1[159:152] = in_data1[3591:3584];
      mux_data1[167:160] = in_data1[3599:3592];
      mux_data1[175:168] = in_data1[3607:3600];
      mux_data2[7:0] = in_data2[3439:3432];
      mux_data2[15:8] = in_data2[3447:3440];
      mux_data2[23:16] = in_data2[3455:3448];
      mux_data2[31:24] = in_data2[3463:3456];
      mux_data2[39:32] = in_data2[3471:3464];
      mux_data2[47:40] = in_data2[3479:3472];
      mux_data2[55:48] = in_data2[3487:3480];
      mux_data2[63:56] = in_data2[3495:3488];
      mux_data2[71:64] = in_data2[3503:3496];
      mux_data2[79:72] = in_data2[3511:3504];
      mux_data2[87:80] = in_data2[3519:3512];
      mux_data2[95:88] = in_data2[3527:3520];
      mux_data2[103:96] = in_data2[3535:3528];
      mux_data2[111:104] = in_data2[3543:3536];
      mux_data2[119:112] = in_data2[3551:3544];
      mux_data2[127:120] = in_data2[3559:3552];
      mux_data2[135:128] = in_data2[3567:3560];
      mux_data2[143:136] = in_data2[3575:3568];
      mux_data2[151:144] = in_data2[3583:3576];
      mux_data2[159:152] = in_data2[3591:3584];
      mux_data2[167:160] = in_data2[3599:3592];
      mux_data2[175:168] = in_data2[3607:3600];
      mux_data3[7:0] = in_data3[3439:3432];
      mux_data3[15:8] = in_data3[3447:3440];
      mux_data3[23:16] = in_data3[3455:3448];
      mux_data3[31:24] = in_data3[3463:3456];
      mux_data3[39:32] = in_data3[3471:3464];
      mux_data3[47:40] = in_data3[3479:3472];
      mux_data3[55:48] = in_data3[3487:3480];
      mux_data3[63:56] = in_data3[3495:3488];
      mux_data3[71:64] = in_data3[3503:3496];
      mux_data3[79:72] = in_data3[3511:3504];
      mux_data3[87:80] = in_data3[3519:3512];
      mux_data3[95:88] = in_data3[3527:3520];
      mux_data3[103:96] = in_data3[3535:3528];
      mux_data3[111:104] = in_data3[3543:3536];
      mux_data3[119:112] = in_data3[3551:3544];
      mux_data3[127:120] = in_data3[3559:3552];
      mux_data3[135:128] = in_data3[3567:3560];
      mux_data3[143:136] = in_data3[3575:3568];
      mux_data3[151:144] = in_data3[3583:3576];
      mux_data3[159:152] = in_data3[3591:3584];
      mux_data3[167:160] = in_data3[3599:3592];
      mux_data3[175:168] = in_data3[3607:3600];
      mux_data4[7:0] = in_data4[3439:3432];
      mux_data4[15:8] = in_data4[3447:3440];
      mux_data4[23:16] = in_data4[3455:3448];
      mux_data4[31:24] = in_data4[3463:3456];
      mux_data4[39:32] = in_data4[3471:3464];
      mux_data4[47:40] = in_data4[3479:3472];
      mux_data4[55:48] = in_data4[3487:3480];
      mux_data4[63:56] = in_data4[3495:3488];
      mux_data4[71:64] = in_data4[3503:3496];
      mux_data4[79:72] = in_data4[3511:3504];
      mux_data4[87:80] = in_data4[3519:3512];
      mux_data4[95:88] = in_data4[3527:3520];
      mux_data4[103:96] = in_data4[3535:3528];
      mux_data4[111:104] = in_data4[3543:3536];
      mux_data4[119:112] = in_data4[3551:3544];
      mux_data4[127:120] = in_data4[3559:3552];
      mux_data4[135:128] = in_data4[3567:3560];
      mux_data4[143:136] = in_data4[3575:3568];
      mux_data4[151:144] = in_data4[3583:3576];
      mux_data4[159:152] = in_data4[3591:3584];
      mux_data4[167:160] = in_data4[3599:3592];
      mux_data4[175:168] = in_data4[3607:3600];
    end
    'd28: begin
      mux_data0[7:0] = in_data0[3567:3560];
      mux_data0[15:8] = in_data0[3575:3568];
      mux_data0[23:16] = in_data0[3583:3576];
      mux_data0[31:24] = in_data0[3591:3584];
      mux_data0[39:32] = in_data0[3599:3592];
      mux_data0[47:40] = in_data0[3607:3600];
      mux_data0[55:48] = in_data0[3615:3608];
      mux_data0[63:56] = in_data0[3623:3616];
      mux_data0[71:64] = in_data0[3631:3624];
      mux_data0[79:72] = in_data0[3639:3632];
      mux_data0[87:80] = in_data0[3647:3640];
      mux_data0[95:88] = in_data0[3655:3648];
      mux_data0[103:96] = in_data0[3663:3656];
      mux_data0[111:104] = in_data0[3671:3664];
      mux_data0[119:112] = in_data0[3679:3672];
      mux_data0[127:120] = in_data0[3687:3680];
      mux_data0[135:128] = in_data0[3695:3688];
      mux_data0[143:136] = in_data0[3703:3696];
      mux_data0[151:144] = in_data0[3711:3704];
      mux_data0[159:152] = in_data0[3719:3712];
      mux_data0[167:160] = in_data0[3727:3720];
      mux_data0[175:168] = in_data0[3735:3728];
      mux_data1[7:0] = in_data1[3567:3560];
      mux_data1[15:8] = in_data1[3575:3568];
      mux_data1[23:16] = in_data1[3583:3576];
      mux_data1[31:24] = in_data1[3591:3584];
      mux_data1[39:32] = in_data1[3599:3592];
      mux_data1[47:40] = in_data1[3607:3600];
      mux_data1[55:48] = in_data1[3615:3608];
      mux_data1[63:56] = in_data1[3623:3616];
      mux_data1[71:64] = in_data1[3631:3624];
      mux_data1[79:72] = in_data1[3639:3632];
      mux_data1[87:80] = in_data1[3647:3640];
      mux_data1[95:88] = in_data1[3655:3648];
      mux_data1[103:96] = in_data1[3663:3656];
      mux_data1[111:104] = in_data1[3671:3664];
      mux_data1[119:112] = in_data1[3679:3672];
      mux_data1[127:120] = in_data1[3687:3680];
      mux_data1[135:128] = in_data1[3695:3688];
      mux_data1[143:136] = in_data1[3703:3696];
      mux_data1[151:144] = in_data1[3711:3704];
      mux_data1[159:152] = in_data1[3719:3712];
      mux_data1[167:160] = in_data1[3727:3720];
      mux_data1[175:168] = in_data1[3735:3728];
      mux_data2[7:0] = in_data2[3567:3560];
      mux_data2[15:8] = in_data2[3575:3568];
      mux_data2[23:16] = in_data2[3583:3576];
      mux_data2[31:24] = in_data2[3591:3584];
      mux_data2[39:32] = in_data2[3599:3592];
      mux_data2[47:40] = in_data2[3607:3600];
      mux_data2[55:48] = in_data2[3615:3608];
      mux_data2[63:56] = in_data2[3623:3616];
      mux_data2[71:64] = in_data2[3631:3624];
      mux_data2[79:72] = in_data2[3639:3632];
      mux_data2[87:80] = in_data2[3647:3640];
      mux_data2[95:88] = in_data2[3655:3648];
      mux_data2[103:96] = in_data2[3663:3656];
      mux_data2[111:104] = in_data2[3671:3664];
      mux_data2[119:112] = in_data2[3679:3672];
      mux_data2[127:120] = in_data2[3687:3680];
      mux_data2[135:128] = in_data2[3695:3688];
      mux_data2[143:136] = in_data2[3703:3696];
      mux_data2[151:144] = in_data2[3711:3704];
      mux_data2[159:152] = in_data2[3719:3712];
      mux_data2[167:160] = in_data2[3727:3720];
      mux_data2[175:168] = in_data2[3735:3728];
      mux_data3[7:0] = in_data3[3567:3560];
      mux_data3[15:8] = in_data3[3575:3568];
      mux_data3[23:16] = in_data3[3583:3576];
      mux_data3[31:24] = in_data3[3591:3584];
      mux_data3[39:32] = in_data3[3599:3592];
      mux_data3[47:40] = in_data3[3607:3600];
      mux_data3[55:48] = in_data3[3615:3608];
      mux_data3[63:56] = in_data3[3623:3616];
      mux_data3[71:64] = in_data3[3631:3624];
      mux_data3[79:72] = in_data3[3639:3632];
      mux_data3[87:80] = in_data3[3647:3640];
      mux_data3[95:88] = in_data3[3655:3648];
      mux_data3[103:96] = in_data3[3663:3656];
      mux_data3[111:104] = in_data3[3671:3664];
      mux_data3[119:112] = in_data3[3679:3672];
      mux_data3[127:120] = in_data3[3687:3680];
      mux_data3[135:128] = in_data3[3695:3688];
      mux_data3[143:136] = in_data3[3703:3696];
      mux_data3[151:144] = in_data3[3711:3704];
      mux_data3[159:152] = in_data3[3719:3712];
      mux_data3[167:160] = in_data3[3727:3720];
      mux_data3[175:168] = in_data3[3735:3728];
      mux_data4[7:0] = in_data4[3567:3560];
      mux_data4[15:8] = in_data4[3575:3568];
      mux_data4[23:16] = in_data4[3583:3576];
      mux_data4[31:24] = in_data4[3591:3584];
      mux_data4[39:32] = in_data4[3599:3592];
      mux_data4[47:40] = in_data4[3607:3600];
      mux_data4[55:48] = in_data4[3615:3608];
      mux_data4[63:56] = in_data4[3623:3616];
      mux_data4[71:64] = in_data4[3631:3624];
      mux_data4[79:72] = in_data4[3639:3632];
      mux_data4[87:80] = in_data4[3647:3640];
      mux_data4[95:88] = in_data4[3655:3648];
      mux_data4[103:96] = in_data4[3663:3656];
      mux_data4[111:104] = in_data4[3671:3664];
      mux_data4[119:112] = in_data4[3679:3672];
      mux_data4[127:120] = in_data4[3687:3680];
      mux_data4[135:128] = in_data4[3695:3688];
      mux_data4[143:136] = in_data4[3703:3696];
      mux_data4[151:144] = in_data4[3711:3704];
      mux_data4[159:152] = in_data4[3719:3712];
      mux_data4[167:160] = in_data4[3727:3720];
      mux_data4[175:168] = in_data4[3735:3728];
    end
    'd29: begin
      mux_data0[7:0] = in_data0[3695:3688];
      mux_data0[15:8] = in_data0[3703:3696];
      mux_data0[23:16] = in_data0[3711:3704];
      mux_data0[31:24] = in_data0[3719:3712];
      mux_data0[39:32] = in_data0[3727:3720];
      mux_data0[47:40] = in_data0[3735:3728];
      mux_data0[55:48] = in_data0[3743:3736];
      mux_data0[63:56] = in_data0[3751:3744];
      mux_data0[71:64] = in_data0[3759:3752];
      mux_data0[79:72] = in_data0[3767:3760];
      mux_data0[87:80] = in_data0[3775:3768];
      mux_data0[95:88] = in_data0[3783:3776];
      mux_data0[103:96] = in_data0[3791:3784];
      mux_data0[111:104] = in_data0[3799:3792];
      mux_data0[119:112] = in_data0[3807:3800];
      mux_data0[127:120] = in_data0[3815:3808];
      mux_data0[135:128] = in_data0[3823:3816];
      mux_data0[143:136] = in_data0[3831:3824];
      mux_data0[151:144] = in_data0[3839:3832];
      mux_data0[159:152] = in_data0[3847:3840];
      mux_data0[167:160] = in_data0[3855:3848];
      mux_data0[175:168] = in_data0[3863:3856];
      mux_data1[7:0] = in_data1[3695:3688];
      mux_data1[15:8] = in_data1[3703:3696];
      mux_data1[23:16] = in_data1[3711:3704];
      mux_data1[31:24] = in_data1[3719:3712];
      mux_data1[39:32] = in_data1[3727:3720];
      mux_data1[47:40] = in_data1[3735:3728];
      mux_data1[55:48] = in_data1[3743:3736];
      mux_data1[63:56] = in_data1[3751:3744];
      mux_data1[71:64] = in_data1[3759:3752];
      mux_data1[79:72] = in_data1[3767:3760];
      mux_data1[87:80] = in_data1[3775:3768];
      mux_data1[95:88] = in_data1[3783:3776];
      mux_data1[103:96] = in_data1[3791:3784];
      mux_data1[111:104] = in_data1[3799:3792];
      mux_data1[119:112] = in_data1[3807:3800];
      mux_data1[127:120] = in_data1[3815:3808];
      mux_data1[135:128] = in_data1[3823:3816];
      mux_data1[143:136] = in_data1[3831:3824];
      mux_data1[151:144] = in_data1[3839:3832];
      mux_data1[159:152] = in_data1[3847:3840];
      mux_data1[167:160] = in_data1[3855:3848];
      mux_data1[175:168] = in_data1[3863:3856];
      mux_data2[7:0] = in_data2[3695:3688];
      mux_data2[15:8] = in_data2[3703:3696];
      mux_data2[23:16] = in_data2[3711:3704];
      mux_data2[31:24] = in_data2[3719:3712];
      mux_data2[39:32] = in_data2[3727:3720];
      mux_data2[47:40] = in_data2[3735:3728];
      mux_data2[55:48] = in_data2[3743:3736];
      mux_data2[63:56] = in_data2[3751:3744];
      mux_data2[71:64] = in_data2[3759:3752];
      mux_data2[79:72] = in_data2[3767:3760];
      mux_data2[87:80] = in_data2[3775:3768];
      mux_data2[95:88] = in_data2[3783:3776];
      mux_data2[103:96] = in_data2[3791:3784];
      mux_data2[111:104] = in_data2[3799:3792];
      mux_data2[119:112] = in_data2[3807:3800];
      mux_data2[127:120] = in_data2[3815:3808];
      mux_data2[135:128] = in_data2[3823:3816];
      mux_data2[143:136] = in_data2[3831:3824];
      mux_data2[151:144] = in_data2[3839:3832];
      mux_data2[159:152] = in_data2[3847:3840];
      mux_data2[167:160] = in_data2[3855:3848];
      mux_data2[175:168] = in_data2[3863:3856];
      mux_data3[7:0] = in_data3[3695:3688];
      mux_data3[15:8] = in_data3[3703:3696];
      mux_data3[23:16] = in_data3[3711:3704];
      mux_data3[31:24] = in_data3[3719:3712];
      mux_data3[39:32] = in_data3[3727:3720];
      mux_data3[47:40] = in_data3[3735:3728];
      mux_data3[55:48] = in_data3[3743:3736];
      mux_data3[63:56] = in_data3[3751:3744];
      mux_data3[71:64] = in_data3[3759:3752];
      mux_data3[79:72] = in_data3[3767:3760];
      mux_data3[87:80] = in_data3[3775:3768];
      mux_data3[95:88] = in_data3[3783:3776];
      mux_data3[103:96] = in_data3[3791:3784];
      mux_data3[111:104] = in_data3[3799:3792];
      mux_data3[119:112] = in_data3[3807:3800];
      mux_data3[127:120] = in_data3[3815:3808];
      mux_data3[135:128] = in_data3[3823:3816];
      mux_data3[143:136] = in_data3[3831:3824];
      mux_data3[151:144] = in_data3[3839:3832];
      mux_data3[159:152] = in_data3[3847:3840];
      mux_data3[167:160] = in_data3[3855:3848];
      mux_data3[175:168] = in_data3[3863:3856];
      mux_data4[7:0] = in_data4[3695:3688];
      mux_data4[15:8] = in_data4[3703:3696];
      mux_data4[23:16] = in_data4[3711:3704];
      mux_data4[31:24] = in_data4[3719:3712];
      mux_data4[39:32] = in_data4[3727:3720];
      mux_data4[47:40] = in_data4[3735:3728];
      mux_data4[55:48] = in_data4[3743:3736];
      mux_data4[63:56] = in_data4[3751:3744];
      mux_data4[71:64] = in_data4[3759:3752];
      mux_data4[79:72] = in_data4[3767:3760];
      mux_data4[87:80] = in_data4[3775:3768];
      mux_data4[95:88] = in_data4[3783:3776];
      mux_data4[103:96] = in_data4[3791:3784];
      mux_data4[111:104] = in_data4[3799:3792];
      mux_data4[119:112] = in_data4[3807:3800];
      mux_data4[127:120] = in_data4[3815:3808];
      mux_data4[135:128] = in_data4[3823:3816];
      mux_data4[143:136] = in_data4[3831:3824];
      mux_data4[151:144] = in_data4[3839:3832];
      mux_data4[159:152] = in_data4[3847:3840];
      mux_data4[167:160] = in_data4[3855:3848];
      mux_data4[175:168] = in_data4[3863:3856];
    end
    'd30: begin
      mux_data0[7:0] = in_data0[3823:3816];
      mux_data0[15:8] = in_data0[3831:3824];
      mux_data0[23:16] = in_data0[3839:3832];
      mux_data0[31:24] = in_data0[3847:3840];
      mux_data0[39:32] = in_data0[3855:3848];
      mux_data0[47:40] = in_data0[3863:3856];
      mux_data0[55:48] = in_data0[3871:3864];
      mux_data0[63:56] = in_data0[3879:3872];
      mux_data0[71:64] = in_data0[3887:3880];
      mux_data0[79:72] = in_data0[3895:3888];
      mux_data0[87:80] = in_data0[3903:3896];
      mux_data0[95:88] = in_data0[3911:3904];
      mux_data0[103:96] = in_data0[3919:3912];
      mux_data0[111:104] = in_data0[3927:3920];
      mux_data0[119:112] = in_data0[3935:3928];
      mux_data0[127:120] = in_data0[3943:3936];
      mux_data0[135:128] = in_data0[3951:3944];
      mux_data0[143:136] = in_data0[3959:3952];
      mux_data0[151:144] = in_data0[3967:3960];
      mux_data0[159:152] = in_data0[3975:3968];
      mux_data0[167:160] = in_data0[3983:3976];
      mux_data0[175:168] = in_data0[3991:3984];
      mux_data1[7:0] = in_data1[3823:3816];
      mux_data1[15:8] = in_data1[3831:3824];
      mux_data1[23:16] = in_data1[3839:3832];
      mux_data1[31:24] = in_data1[3847:3840];
      mux_data1[39:32] = in_data1[3855:3848];
      mux_data1[47:40] = in_data1[3863:3856];
      mux_data1[55:48] = in_data1[3871:3864];
      mux_data1[63:56] = in_data1[3879:3872];
      mux_data1[71:64] = in_data1[3887:3880];
      mux_data1[79:72] = in_data1[3895:3888];
      mux_data1[87:80] = in_data1[3903:3896];
      mux_data1[95:88] = in_data1[3911:3904];
      mux_data1[103:96] = in_data1[3919:3912];
      mux_data1[111:104] = in_data1[3927:3920];
      mux_data1[119:112] = in_data1[3935:3928];
      mux_data1[127:120] = in_data1[3943:3936];
      mux_data1[135:128] = in_data1[3951:3944];
      mux_data1[143:136] = in_data1[3959:3952];
      mux_data1[151:144] = in_data1[3967:3960];
      mux_data1[159:152] = in_data1[3975:3968];
      mux_data1[167:160] = in_data1[3983:3976];
      mux_data1[175:168] = in_data1[3991:3984];
      mux_data2[7:0] = in_data2[3823:3816];
      mux_data2[15:8] = in_data2[3831:3824];
      mux_data2[23:16] = in_data2[3839:3832];
      mux_data2[31:24] = in_data2[3847:3840];
      mux_data2[39:32] = in_data2[3855:3848];
      mux_data2[47:40] = in_data2[3863:3856];
      mux_data2[55:48] = in_data2[3871:3864];
      mux_data2[63:56] = in_data2[3879:3872];
      mux_data2[71:64] = in_data2[3887:3880];
      mux_data2[79:72] = in_data2[3895:3888];
      mux_data2[87:80] = in_data2[3903:3896];
      mux_data2[95:88] = in_data2[3911:3904];
      mux_data2[103:96] = in_data2[3919:3912];
      mux_data2[111:104] = in_data2[3927:3920];
      mux_data2[119:112] = in_data2[3935:3928];
      mux_data2[127:120] = in_data2[3943:3936];
      mux_data2[135:128] = in_data2[3951:3944];
      mux_data2[143:136] = in_data2[3959:3952];
      mux_data2[151:144] = in_data2[3967:3960];
      mux_data2[159:152] = in_data2[3975:3968];
      mux_data2[167:160] = in_data2[3983:3976];
      mux_data2[175:168] = in_data2[3991:3984];
      mux_data3[7:0] = in_data3[3823:3816];
      mux_data3[15:8] = in_data3[3831:3824];
      mux_data3[23:16] = in_data3[3839:3832];
      mux_data3[31:24] = in_data3[3847:3840];
      mux_data3[39:32] = in_data3[3855:3848];
      mux_data3[47:40] = in_data3[3863:3856];
      mux_data3[55:48] = in_data3[3871:3864];
      mux_data3[63:56] = in_data3[3879:3872];
      mux_data3[71:64] = in_data3[3887:3880];
      mux_data3[79:72] = in_data3[3895:3888];
      mux_data3[87:80] = in_data3[3903:3896];
      mux_data3[95:88] = in_data3[3911:3904];
      mux_data3[103:96] = in_data3[3919:3912];
      mux_data3[111:104] = in_data3[3927:3920];
      mux_data3[119:112] = in_data3[3935:3928];
      mux_data3[127:120] = in_data3[3943:3936];
      mux_data3[135:128] = in_data3[3951:3944];
      mux_data3[143:136] = in_data3[3959:3952];
      mux_data3[151:144] = in_data3[3967:3960];
      mux_data3[159:152] = in_data3[3975:3968];
      mux_data3[167:160] = in_data3[3983:3976];
      mux_data3[175:168] = in_data3[3991:3984];
      mux_data4[7:0] = in_data4[3823:3816];
      mux_data4[15:8] = in_data4[3831:3824];
      mux_data4[23:16] = in_data4[3839:3832];
      mux_data4[31:24] = in_data4[3847:3840];
      mux_data4[39:32] = in_data4[3855:3848];
      mux_data4[47:40] = in_data4[3863:3856];
      mux_data4[55:48] = in_data4[3871:3864];
      mux_data4[63:56] = in_data4[3879:3872];
      mux_data4[71:64] = in_data4[3887:3880];
      mux_data4[79:72] = in_data4[3895:3888];
      mux_data4[87:80] = in_data4[3903:3896];
      mux_data4[95:88] = in_data4[3911:3904];
      mux_data4[103:96] = in_data4[3919:3912];
      mux_data4[111:104] = in_data4[3927:3920];
      mux_data4[119:112] = in_data4[3935:3928];
      mux_data4[127:120] = in_data4[3943:3936];
      mux_data4[135:128] = in_data4[3951:3944];
      mux_data4[143:136] = in_data4[3959:3952];
      mux_data4[151:144] = in_data4[3967:3960];
      mux_data4[159:152] = in_data4[3975:3968];
      mux_data4[167:160] = in_data4[3983:3976];
      mux_data4[175:168] = in_data4[3991:3984];
    end
    'd31: begin
      mux_data0[7:0] = in_data0[3951:3944];
      mux_data0[15:8] = in_data0[3959:3952];
      mux_data0[23:16] = in_data0[3967:3960];
      mux_data0[31:24] = in_data0[3975:3968];
      mux_data0[39:32] = in_data0[3983:3976];
      mux_data0[47:40] = in_data0[3991:3984];
      mux_data0[55:48] = in_data0[3999:3992];
      mux_data0[63:56] = in_data0[4007:4000];
      mux_data0[71:64] = in_data0[4015:4008];
      mux_data0[79:72] = in_data0[4023:4016];
      mux_data0[87:80] = in_data0[4031:4024];
      mux_data0[95:88] = in_data0[4039:4032];
      mux_data0[103:96] = in_data0[4047:4040];
      mux_data0[111:104] = in_data0[4055:4048];
      mux_data0[119:112] = in_data0[4063:4056];
      mux_data0[127:120] = in_data0[4071:4064];
      mux_data0[135:128] = in_data0[4079:4072];
      mux_data0[143:136] = in_data0[4087:4080];
      mux_data0[151:144] = in_data0[4095:4088];
      mux_data0[159:152] = in_data0[4103:4096];
      mux_data0[167:160] = in_data0[4111:4104];
      mux_data0[175:168] = in_data0[4119:4112];
      mux_data1[7:0] = in_data1[3951:3944];
      mux_data1[15:8] = in_data1[3959:3952];
      mux_data1[23:16] = in_data1[3967:3960];
      mux_data1[31:24] = in_data1[3975:3968];
      mux_data1[39:32] = in_data1[3983:3976];
      mux_data1[47:40] = in_data1[3991:3984];
      mux_data1[55:48] = in_data1[3999:3992];
      mux_data1[63:56] = in_data1[4007:4000];
      mux_data1[71:64] = in_data1[4015:4008];
      mux_data1[79:72] = in_data1[4023:4016];
      mux_data1[87:80] = in_data1[4031:4024];
      mux_data1[95:88] = in_data1[4039:4032];
      mux_data1[103:96] = in_data1[4047:4040];
      mux_data1[111:104] = in_data1[4055:4048];
      mux_data1[119:112] = in_data1[4063:4056];
      mux_data1[127:120] = in_data1[4071:4064];
      mux_data1[135:128] = in_data1[4079:4072];
      mux_data1[143:136] = in_data1[4087:4080];
      mux_data1[151:144] = in_data1[4095:4088];
      mux_data1[159:152] = in_data1[4103:4096];
      mux_data1[167:160] = in_data1[4111:4104];
      mux_data1[175:168] = in_data1[4119:4112];
      mux_data2[7:0] = in_data2[3951:3944];
      mux_data2[15:8] = in_data2[3959:3952];
      mux_data2[23:16] = in_data2[3967:3960];
      mux_data2[31:24] = in_data2[3975:3968];
      mux_data2[39:32] = in_data2[3983:3976];
      mux_data2[47:40] = in_data2[3991:3984];
      mux_data2[55:48] = in_data2[3999:3992];
      mux_data2[63:56] = in_data2[4007:4000];
      mux_data2[71:64] = in_data2[4015:4008];
      mux_data2[79:72] = in_data2[4023:4016];
      mux_data2[87:80] = in_data2[4031:4024];
      mux_data2[95:88] = in_data2[4039:4032];
      mux_data2[103:96] = in_data2[4047:4040];
      mux_data2[111:104] = in_data2[4055:4048];
      mux_data2[119:112] = in_data2[4063:4056];
      mux_data2[127:120] = in_data2[4071:4064];
      mux_data2[135:128] = in_data2[4079:4072];
      mux_data2[143:136] = in_data2[4087:4080];
      mux_data2[151:144] = in_data2[4095:4088];
      mux_data2[159:152] = in_data2[4103:4096];
      mux_data2[167:160] = in_data2[4111:4104];
      mux_data2[175:168] = in_data2[4119:4112];
      mux_data3[7:0] = in_data3[3951:3944];
      mux_data3[15:8] = in_data3[3959:3952];
      mux_data3[23:16] = in_data3[3967:3960];
      mux_data3[31:24] = in_data3[3975:3968];
      mux_data3[39:32] = in_data3[3983:3976];
      mux_data3[47:40] = in_data3[3991:3984];
      mux_data3[55:48] = in_data3[3999:3992];
      mux_data3[63:56] = in_data3[4007:4000];
      mux_data3[71:64] = in_data3[4015:4008];
      mux_data3[79:72] = in_data3[4023:4016];
      mux_data3[87:80] = in_data3[4031:4024];
      mux_data3[95:88] = in_data3[4039:4032];
      mux_data3[103:96] = in_data3[4047:4040];
      mux_data3[111:104] = in_data3[4055:4048];
      mux_data3[119:112] = in_data3[4063:4056];
      mux_data3[127:120] = in_data3[4071:4064];
      mux_data3[135:128] = in_data3[4079:4072];
      mux_data3[143:136] = in_data3[4087:4080];
      mux_data3[151:144] = in_data3[4095:4088];
      mux_data3[159:152] = in_data3[4103:4096];
      mux_data3[167:160] = in_data3[4111:4104];
      mux_data3[175:168] = in_data3[4119:4112];
      mux_data4[7:0] = in_data4[3951:3944];
      mux_data4[15:8] = in_data4[3959:3952];
      mux_data4[23:16] = in_data4[3967:3960];
      mux_data4[31:24] = in_data4[3975:3968];
      mux_data4[39:32] = in_data4[3983:3976];
      mux_data4[47:40] = in_data4[3991:3984];
      mux_data4[55:48] = in_data4[3999:3992];
      mux_data4[63:56] = in_data4[4007:4000];
      mux_data4[71:64] = in_data4[4015:4008];
      mux_data4[79:72] = in_data4[4023:4016];
      mux_data4[87:80] = in_data4[4031:4024];
      mux_data4[95:88] = in_data4[4039:4032];
      mux_data4[103:96] = in_data4[4047:4040];
      mux_data4[111:104] = in_data4[4055:4048];
      mux_data4[119:112] = in_data4[4063:4056];
      mux_data4[127:120] = in_data4[4071:4064];
      mux_data4[135:128] = in_data4[4079:4072];
      mux_data4[143:136] = in_data4[4087:4080];
      mux_data4[151:144] = in_data4[4095:4088];
      mux_data4[159:152] = in_data4[4103:4096];
      mux_data4[167:160] = in_data4[4111:4104];
      mux_data4[175:168] = in_data4[4119:4112];
    end
    'd32: begin
      mux_data0[7:0] = in_data0[4079:4072];
      mux_data0[15:8] = in_data0[4087:4080];
      mux_data0[23:16] = in_data0[4095:4088];
      mux_data0[31:24] = in_data0[4103:4096];
      mux_data0[39:32] = in_data0[4111:4104];
      mux_data0[47:40] = in_data0[4119:4112];
      mux_data0[55:48] = in_data0[4127:4120];
      mux_data0[63:56] = in_data0[4135:4128];
      mux_data0[71:64] = in_data0[4143:4136];
      mux_data0[79:72] = in_data0[4151:4144];
      mux_data0[87:80] = in_data0[4159:4152];
      mux_data0[95:88] = in_data0[4167:4160];
      mux_data0[103:96] = in_data0[4175:4168];
      mux_data0[111:104] = in_data0[4183:4176];
      mux_data0[119:112] = in_data0[4191:4184];
      mux_data0[127:120] = in_data0[4199:4192];
      mux_data0[135:128] = in_data0[4207:4200];
      mux_data0[143:136] = in_data0[4215:4208];
      mux_data0[151:144] = in_data0[4223:4216];
      mux_data0[159:152] = in_data0[4231:4224];
      mux_data0[167:160] = in_data0[4239:4232];
      mux_data0[175:168] = in_data0[4247:4240];
      mux_data1[7:0] = in_data1[4079:4072];
      mux_data1[15:8] = in_data1[4087:4080];
      mux_data1[23:16] = in_data1[4095:4088];
      mux_data1[31:24] = in_data1[4103:4096];
      mux_data1[39:32] = in_data1[4111:4104];
      mux_data1[47:40] = in_data1[4119:4112];
      mux_data1[55:48] = in_data1[4127:4120];
      mux_data1[63:56] = in_data1[4135:4128];
      mux_data1[71:64] = in_data1[4143:4136];
      mux_data1[79:72] = in_data1[4151:4144];
      mux_data1[87:80] = in_data1[4159:4152];
      mux_data1[95:88] = in_data1[4167:4160];
      mux_data1[103:96] = in_data1[4175:4168];
      mux_data1[111:104] = in_data1[4183:4176];
      mux_data1[119:112] = in_data1[4191:4184];
      mux_data1[127:120] = in_data1[4199:4192];
      mux_data1[135:128] = in_data1[4207:4200];
      mux_data1[143:136] = in_data1[4215:4208];
      mux_data1[151:144] = in_data1[4223:4216];
      mux_data1[159:152] = in_data1[4231:4224];
      mux_data1[167:160] = in_data1[4239:4232];
      mux_data1[175:168] = in_data1[4247:4240];
      mux_data2[7:0] = in_data2[4079:4072];
      mux_data2[15:8] = in_data2[4087:4080];
      mux_data2[23:16] = in_data2[4095:4088];
      mux_data2[31:24] = in_data2[4103:4096];
      mux_data2[39:32] = in_data2[4111:4104];
      mux_data2[47:40] = in_data2[4119:4112];
      mux_data2[55:48] = in_data2[4127:4120];
      mux_data2[63:56] = in_data2[4135:4128];
      mux_data2[71:64] = in_data2[4143:4136];
      mux_data2[79:72] = in_data2[4151:4144];
      mux_data2[87:80] = in_data2[4159:4152];
      mux_data2[95:88] = in_data2[4167:4160];
      mux_data2[103:96] = in_data2[4175:4168];
      mux_data2[111:104] = in_data2[4183:4176];
      mux_data2[119:112] = in_data2[4191:4184];
      mux_data2[127:120] = in_data2[4199:4192];
      mux_data2[135:128] = in_data2[4207:4200];
      mux_data2[143:136] = in_data2[4215:4208];
      mux_data2[151:144] = in_data2[4223:4216];
      mux_data2[159:152] = in_data2[4231:4224];
      mux_data2[167:160] = in_data2[4239:4232];
      mux_data2[175:168] = in_data2[4247:4240];
      mux_data3[7:0] = in_data3[4079:4072];
      mux_data3[15:8] = in_data3[4087:4080];
      mux_data3[23:16] = in_data3[4095:4088];
      mux_data3[31:24] = in_data3[4103:4096];
      mux_data3[39:32] = in_data3[4111:4104];
      mux_data3[47:40] = in_data3[4119:4112];
      mux_data3[55:48] = in_data3[4127:4120];
      mux_data3[63:56] = in_data3[4135:4128];
      mux_data3[71:64] = in_data3[4143:4136];
      mux_data3[79:72] = in_data3[4151:4144];
      mux_data3[87:80] = in_data3[4159:4152];
      mux_data3[95:88] = in_data3[4167:4160];
      mux_data3[103:96] = in_data3[4175:4168];
      mux_data3[111:104] = in_data3[4183:4176];
      mux_data3[119:112] = in_data3[4191:4184];
      mux_data3[127:120] = in_data3[4199:4192];
      mux_data3[135:128] = in_data3[4207:4200];
      mux_data3[143:136] = in_data3[4215:4208];
      mux_data3[151:144] = in_data3[4223:4216];
      mux_data3[159:152] = in_data3[4231:4224];
      mux_data3[167:160] = in_data3[4239:4232];
      mux_data3[175:168] = in_data3[4247:4240];
      mux_data4[7:0] = in_data4[4079:4072];
      mux_data4[15:8] = in_data4[4087:4080];
      mux_data4[23:16] = in_data4[4095:4088];
      mux_data4[31:24] = in_data4[4103:4096];
      mux_data4[39:32] = in_data4[4111:4104];
      mux_data4[47:40] = in_data4[4119:4112];
      mux_data4[55:48] = in_data4[4127:4120];
      mux_data4[63:56] = in_data4[4135:4128];
      mux_data4[71:64] = in_data4[4143:4136];
      mux_data4[79:72] = in_data4[4151:4144];
      mux_data4[87:80] = in_data4[4159:4152];
      mux_data4[95:88] = in_data4[4167:4160];
      mux_data4[103:96] = in_data4[4175:4168];
      mux_data4[111:104] = in_data4[4183:4176];
      mux_data4[119:112] = in_data4[4191:4184];
      mux_data4[127:120] = in_data4[4199:4192];
      mux_data4[135:128] = in_data4[4207:4200];
      mux_data4[143:136] = in_data4[4215:4208];
      mux_data4[151:144] = in_data4[4223:4216];
      mux_data4[159:152] = in_data4[4231:4224];
      mux_data4[167:160] = in_data4[4239:4232];
      mux_data4[175:168] = in_data4[4247:4240];
    end
    'd33: begin
      mux_data0[7:0] = in_data0[4207:4200];
      mux_data0[15:8] = in_data0[4215:4208];
      mux_data0[23:16] = in_data0[4223:4216];
      mux_data0[31:24] = in_data0[4231:4224];
      mux_data0[39:32] = in_data0[4239:4232];
      mux_data0[47:40] = in_data0[4247:4240];
      mux_data0[55:48] = in_data0[4255:4248];
      mux_data0[63:56] = in_data0[4263:4256];
      mux_data0[71:64] = in_data0[4271:4264];
      mux_data0[79:72] = in_data0[4279:4272];
      mux_data0[87:80] = in_data0[4287:4280];
      mux_data0[95:88] = in_data0[4295:4288];
      mux_data0[103:96] = in_data0[4303:4296];
      mux_data0[111:104] = in_data0[4311:4304];
      mux_data0[119:112] = in_data0[4319:4312];
      mux_data0[127:120] = in_data0[4327:4320];
      mux_data0[135:128] = in_data0[4335:4328];
      mux_data0[143:136] = in_data0[4343:4336];
      mux_data0[151:144] = in_data0[4351:4344];
      mux_data0[159:152] = in_data0[4359:4352];
      mux_data0[167:160] = in_data0[4367:4360];
      mux_data0[175:168] = in_data0[4375:4368];
      mux_data1[7:0] = in_data1[4207:4200];
      mux_data1[15:8] = in_data1[4215:4208];
      mux_data1[23:16] = in_data1[4223:4216];
      mux_data1[31:24] = in_data1[4231:4224];
      mux_data1[39:32] = in_data1[4239:4232];
      mux_data1[47:40] = in_data1[4247:4240];
      mux_data1[55:48] = in_data1[4255:4248];
      mux_data1[63:56] = in_data1[4263:4256];
      mux_data1[71:64] = in_data1[4271:4264];
      mux_data1[79:72] = in_data1[4279:4272];
      mux_data1[87:80] = in_data1[4287:4280];
      mux_data1[95:88] = in_data1[4295:4288];
      mux_data1[103:96] = in_data1[4303:4296];
      mux_data1[111:104] = in_data1[4311:4304];
      mux_data1[119:112] = in_data1[4319:4312];
      mux_data1[127:120] = in_data1[4327:4320];
      mux_data1[135:128] = in_data1[4335:4328];
      mux_data1[143:136] = in_data1[4343:4336];
      mux_data1[151:144] = in_data1[4351:4344];
      mux_data1[159:152] = in_data1[4359:4352];
      mux_data1[167:160] = in_data1[4367:4360];
      mux_data1[175:168] = in_data1[4375:4368];
      mux_data2[7:0] = in_data2[4207:4200];
      mux_data2[15:8] = in_data2[4215:4208];
      mux_data2[23:16] = in_data2[4223:4216];
      mux_data2[31:24] = in_data2[4231:4224];
      mux_data2[39:32] = in_data2[4239:4232];
      mux_data2[47:40] = in_data2[4247:4240];
      mux_data2[55:48] = in_data2[4255:4248];
      mux_data2[63:56] = in_data2[4263:4256];
      mux_data2[71:64] = in_data2[4271:4264];
      mux_data2[79:72] = in_data2[4279:4272];
      mux_data2[87:80] = in_data2[4287:4280];
      mux_data2[95:88] = in_data2[4295:4288];
      mux_data2[103:96] = in_data2[4303:4296];
      mux_data2[111:104] = in_data2[4311:4304];
      mux_data2[119:112] = in_data2[4319:4312];
      mux_data2[127:120] = in_data2[4327:4320];
      mux_data2[135:128] = in_data2[4335:4328];
      mux_data2[143:136] = in_data2[4343:4336];
      mux_data2[151:144] = in_data2[4351:4344];
      mux_data2[159:152] = in_data2[4359:4352];
      mux_data2[167:160] = in_data2[4367:4360];
      mux_data2[175:168] = in_data2[4375:4368];
      mux_data3[7:0] = in_data3[4207:4200];
      mux_data3[15:8] = in_data3[4215:4208];
      mux_data3[23:16] = in_data3[4223:4216];
      mux_data3[31:24] = in_data3[4231:4224];
      mux_data3[39:32] = in_data3[4239:4232];
      mux_data3[47:40] = in_data3[4247:4240];
      mux_data3[55:48] = in_data3[4255:4248];
      mux_data3[63:56] = in_data3[4263:4256];
      mux_data3[71:64] = in_data3[4271:4264];
      mux_data3[79:72] = in_data3[4279:4272];
      mux_data3[87:80] = in_data3[4287:4280];
      mux_data3[95:88] = in_data3[4295:4288];
      mux_data3[103:96] = in_data3[4303:4296];
      mux_data3[111:104] = in_data3[4311:4304];
      mux_data3[119:112] = in_data3[4319:4312];
      mux_data3[127:120] = in_data3[4327:4320];
      mux_data3[135:128] = in_data3[4335:4328];
      mux_data3[143:136] = in_data3[4343:4336];
      mux_data3[151:144] = in_data3[4351:4344];
      mux_data3[159:152] = in_data3[4359:4352];
      mux_data3[167:160] = in_data3[4367:4360];
      mux_data3[175:168] = in_data3[4375:4368];
      mux_data4[7:0] = in_data4[4207:4200];
      mux_data4[15:8] = in_data4[4215:4208];
      mux_data4[23:16] = in_data4[4223:4216];
      mux_data4[31:24] = in_data4[4231:4224];
      mux_data4[39:32] = in_data4[4239:4232];
      mux_data4[47:40] = in_data4[4247:4240];
      mux_data4[55:48] = in_data4[4255:4248];
      mux_data4[63:56] = in_data4[4263:4256];
      mux_data4[71:64] = in_data4[4271:4264];
      mux_data4[79:72] = in_data4[4279:4272];
      mux_data4[87:80] = in_data4[4287:4280];
      mux_data4[95:88] = in_data4[4295:4288];
      mux_data4[103:96] = in_data4[4303:4296];
      mux_data4[111:104] = in_data4[4311:4304];
      mux_data4[119:112] = in_data4[4319:4312];
      mux_data4[127:120] = in_data4[4327:4320];
      mux_data4[135:128] = in_data4[4335:4328];
      mux_data4[143:136] = in_data4[4343:4336];
      mux_data4[151:144] = in_data4[4351:4344];
      mux_data4[159:152] = in_data4[4359:4352];
      mux_data4[167:160] = in_data4[4367:4360];
      mux_data4[175:168] = in_data4[4375:4368];
    end
    'd34: begin
      mux_data0[7:0] = in_data0[4335:4328];
      mux_data0[15:8] = in_data0[4343:4336];
      mux_data0[23:16] = in_data0[4351:4344];
      mux_data0[31:24] = in_data0[4359:4352];
      mux_data0[39:32] = in_data0[4367:4360];
      mux_data0[47:40] = in_data0[4375:4368];
      mux_data0[55:48] = in_data0[4383:4376];
      mux_data0[63:56] = in_data0[4391:4384];
      mux_data0[71:64] = in_data0[4399:4392];
      mux_data0[79:72] = in_data0[4407:4400];
      mux_data0[87:80] = in_data0[4415:4408];
      mux_data0[95:88] = in_data0[4423:4416];
      mux_data0[103:96] = in_data0[4431:4424];
      mux_data0[111:104] = in_data0[4439:4432];
      mux_data0[119:112] = in_data0[4447:4440];
      mux_data0[127:120] = in_data0[4455:4448];
      mux_data0[135:128] = in_data0[4463:4456];
      mux_data0[143:136] = in_data0[4471:4464];
      mux_data0[151:144] = in_data0[4479:4472];
      mux_data0[159:152] = in_data0[4487:4480];
      mux_data0[167:160] = in_data0[4495:4488];
      mux_data0[175:168] = in_data0[4503:4496];
      mux_data1[7:0] = in_data1[4335:4328];
      mux_data1[15:8] = in_data1[4343:4336];
      mux_data1[23:16] = in_data1[4351:4344];
      mux_data1[31:24] = in_data1[4359:4352];
      mux_data1[39:32] = in_data1[4367:4360];
      mux_data1[47:40] = in_data1[4375:4368];
      mux_data1[55:48] = in_data1[4383:4376];
      mux_data1[63:56] = in_data1[4391:4384];
      mux_data1[71:64] = in_data1[4399:4392];
      mux_data1[79:72] = in_data1[4407:4400];
      mux_data1[87:80] = in_data1[4415:4408];
      mux_data1[95:88] = in_data1[4423:4416];
      mux_data1[103:96] = in_data1[4431:4424];
      mux_data1[111:104] = in_data1[4439:4432];
      mux_data1[119:112] = in_data1[4447:4440];
      mux_data1[127:120] = in_data1[4455:4448];
      mux_data1[135:128] = in_data1[4463:4456];
      mux_data1[143:136] = in_data1[4471:4464];
      mux_data1[151:144] = in_data1[4479:4472];
      mux_data1[159:152] = in_data1[4487:4480];
      mux_data1[167:160] = in_data1[4495:4488];
      mux_data1[175:168] = in_data1[4503:4496];
      mux_data2[7:0] = in_data2[4335:4328];
      mux_data2[15:8] = in_data2[4343:4336];
      mux_data2[23:16] = in_data2[4351:4344];
      mux_data2[31:24] = in_data2[4359:4352];
      mux_data2[39:32] = in_data2[4367:4360];
      mux_data2[47:40] = in_data2[4375:4368];
      mux_data2[55:48] = in_data2[4383:4376];
      mux_data2[63:56] = in_data2[4391:4384];
      mux_data2[71:64] = in_data2[4399:4392];
      mux_data2[79:72] = in_data2[4407:4400];
      mux_data2[87:80] = in_data2[4415:4408];
      mux_data2[95:88] = in_data2[4423:4416];
      mux_data2[103:96] = in_data2[4431:4424];
      mux_data2[111:104] = in_data2[4439:4432];
      mux_data2[119:112] = in_data2[4447:4440];
      mux_data2[127:120] = in_data2[4455:4448];
      mux_data2[135:128] = in_data2[4463:4456];
      mux_data2[143:136] = in_data2[4471:4464];
      mux_data2[151:144] = in_data2[4479:4472];
      mux_data2[159:152] = in_data2[4487:4480];
      mux_data2[167:160] = in_data2[4495:4488];
      mux_data2[175:168] = in_data2[4503:4496];
      mux_data3[7:0] = in_data3[4335:4328];
      mux_data3[15:8] = in_data3[4343:4336];
      mux_data3[23:16] = in_data3[4351:4344];
      mux_data3[31:24] = in_data3[4359:4352];
      mux_data3[39:32] = in_data3[4367:4360];
      mux_data3[47:40] = in_data3[4375:4368];
      mux_data3[55:48] = in_data3[4383:4376];
      mux_data3[63:56] = in_data3[4391:4384];
      mux_data3[71:64] = in_data3[4399:4392];
      mux_data3[79:72] = in_data3[4407:4400];
      mux_data3[87:80] = in_data3[4415:4408];
      mux_data3[95:88] = in_data3[4423:4416];
      mux_data3[103:96] = in_data3[4431:4424];
      mux_data3[111:104] = in_data3[4439:4432];
      mux_data3[119:112] = in_data3[4447:4440];
      mux_data3[127:120] = in_data3[4455:4448];
      mux_data3[135:128] = in_data3[4463:4456];
      mux_data3[143:136] = in_data3[4471:4464];
      mux_data3[151:144] = in_data3[4479:4472];
      mux_data3[159:152] = in_data3[4487:4480];
      mux_data3[167:160] = in_data3[4495:4488];
      mux_data3[175:168] = in_data3[4503:4496];
      mux_data4[7:0] = in_data4[4335:4328];
      mux_data4[15:8] = in_data4[4343:4336];
      mux_data4[23:16] = in_data4[4351:4344];
      mux_data4[31:24] = in_data4[4359:4352];
      mux_data4[39:32] = in_data4[4367:4360];
      mux_data4[47:40] = in_data4[4375:4368];
      mux_data4[55:48] = in_data4[4383:4376];
      mux_data4[63:56] = in_data4[4391:4384];
      mux_data4[71:64] = in_data4[4399:4392];
      mux_data4[79:72] = in_data4[4407:4400];
      mux_data4[87:80] = in_data4[4415:4408];
      mux_data4[95:88] = in_data4[4423:4416];
      mux_data4[103:96] = in_data4[4431:4424];
      mux_data4[111:104] = in_data4[4439:4432];
      mux_data4[119:112] = in_data4[4447:4440];
      mux_data4[127:120] = in_data4[4455:4448];
      mux_data4[135:128] = in_data4[4463:4456];
      mux_data4[143:136] = in_data4[4471:4464];
      mux_data4[151:144] = in_data4[4479:4472];
      mux_data4[159:152] = in_data4[4487:4480];
      mux_data4[167:160] = in_data4[4495:4488];
      mux_data4[175:168] = in_data4[4503:4496];
    end
    'd35: begin
      mux_data0[7:0] = in_data0[4463:4456];
      mux_data0[15:8] = in_data0[4471:4464];
      mux_data0[23:16] = in_data0[4479:4472];
      mux_data0[31:24] = in_data0[4487:4480];
      mux_data0[39:32] = in_data0[4495:4488];
      mux_data0[47:40] = in_data0[4503:4496];
      mux_data0[55:48] = in_data0[4511:4504];
      mux_data0[63:56] = in_data0[4519:4512];
      mux_data0[71:64] = in_data0[4527:4520];
      mux_data0[79:72] = in_data0[4535:4528];
      mux_data0[87:80] = in_data0[4543:4536];
      mux_data0[95:88] = in_data0[4551:4544];
      mux_data0[103:96] = in_data0[4559:4552];
      mux_data0[111:104] = in_data0[4567:4560];
      mux_data0[119:112] = in_data0[4575:4568];
      mux_data0[127:120] = in_data0[4583:4576];
      mux_data0[135:128] = in_data0[4591:4584];
      mux_data0[143:136] = in_data0[4599:4592];
      mux_data0[151:144] = in_data0[4607:4600];
      mux_data0[159:152] = in_data0[4615:4608];
      mux_data0[167:160] = in_data0[4623:4616];
      mux_data0[175:168] = in_data0[4631:4624];
      mux_data1[7:0] = in_data1[4463:4456];
      mux_data1[15:8] = in_data1[4471:4464];
      mux_data1[23:16] = in_data1[4479:4472];
      mux_data1[31:24] = in_data1[4487:4480];
      mux_data1[39:32] = in_data1[4495:4488];
      mux_data1[47:40] = in_data1[4503:4496];
      mux_data1[55:48] = in_data1[4511:4504];
      mux_data1[63:56] = in_data1[4519:4512];
      mux_data1[71:64] = in_data1[4527:4520];
      mux_data1[79:72] = in_data1[4535:4528];
      mux_data1[87:80] = in_data1[4543:4536];
      mux_data1[95:88] = in_data1[4551:4544];
      mux_data1[103:96] = in_data1[4559:4552];
      mux_data1[111:104] = in_data1[4567:4560];
      mux_data1[119:112] = in_data1[4575:4568];
      mux_data1[127:120] = in_data1[4583:4576];
      mux_data1[135:128] = in_data1[4591:4584];
      mux_data1[143:136] = in_data1[4599:4592];
      mux_data1[151:144] = in_data1[4607:4600];
      mux_data1[159:152] = in_data1[4615:4608];
      mux_data1[167:160] = in_data1[4623:4616];
      mux_data1[175:168] = in_data1[4631:4624];
      mux_data2[7:0] = in_data2[4463:4456];
      mux_data2[15:8] = in_data2[4471:4464];
      mux_data2[23:16] = in_data2[4479:4472];
      mux_data2[31:24] = in_data2[4487:4480];
      mux_data2[39:32] = in_data2[4495:4488];
      mux_data2[47:40] = in_data2[4503:4496];
      mux_data2[55:48] = in_data2[4511:4504];
      mux_data2[63:56] = in_data2[4519:4512];
      mux_data2[71:64] = in_data2[4527:4520];
      mux_data2[79:72] = in_data2[4535:4528];
      mux_data2[87:80] = in_data2[4543:4536];
      mux_data2[95:88] = in_data2[4551:4544];
      mux_data2[103:96] = in_data2[4559:4552];
      mux_data2[111:104] = in_data2[4567:4560];
      mux_data2[119:112] = in_data2[4575:4568];
      mux_data2[127:120] = in_data2[4583:4576];
      mux_data2[135:128] = in_data2[4591:4584];
      mux_data2[143:136] = in_data2[4599:4592];
      mux_data2[151:144] = in_data2[4607:4600];
      mux_data2[159:152] = in_data2[4615:4608];
      mux_data2[167:160] = in_data2[4623:4616];
      mux_data2[175:168] = in_data2[4631:4624];
      mux_data3[7:0] = in_data3[4463:4456];
      mux_data3[15:8] = in_data3[4471:4464];
      mux_data3[23:16] = in_data3[4479:4472];
      mux_data3[31:24] = in_data3[4487:4480];
      mux_data3[39:32] = in_data3[4495:4488];
      mux_data3[47:40] = in_data3[4503:4496];
      mux_data3[55:48] = in_data3[4511:4504];
      mux_data3[63:56] = in_data3[4519:4512];
      mux_data3[71:64] = in_data3[4527:4520];
      mux_data3[79:72] = in_data3[4535:4528];
      mux_data3[87:80] = in_data3[4543:4536];
      mux_data3[95:88] = in_data3[4551:4544];
      mux_data3[103:96] = in_data3[4559:4552];
      mux_data3[111:104] = in_data3[4567:4560];
      mux_data3[119:112] = in_data3[4575:4568];
      mux_data3[127:120] = in_data3[4583:4576];
      mux_data3[135:128] = in_data3[4591:4584];
      mux_data3[143:136] = in_data3[4599:4592];
      mux_data3[151:144] = in_data3[4607:4600];
      mux_data3[159:152] = in_data3[4615:4608];
      mux_data3[167:160] = in_data3[4623:4616];
      mux_data3[175:168] = in_data3[4631:4624];
      mux_data4[7:0] = in_data4[4463:4456];
      mux_data4[15:8] = in_data4[4471:4464];
      mux_data4[23:16] = in_data4[4479:4472];
      mux_data4[31:24] = in_data4[4487:4480];
      mux_data4[39:32] = in_data4[4495:4488];
      mux_data4[47:40] = in_data4[4503:4496];
      mux_data4[55:48] = in_data4[4511:4504];
      mux_data4[63:56] = in_data4[4519:4512];
      mux_data4[71:64] = in_data4[4527:4520];
      mux_data4[79:72] = in_data4[4535:4528];
      mux_data4[87:80] = in_data4[4543:4536];
      mux_data4[95:88] = in_data4[4551:4544];
      mux_data4[103:96] = in_data4[4559:4552];
      mux_data4[111:104] = in_data4[4567:4560];
      mux_data4[119:112] = in_data4[4575:4568];
      mux_data4[127:120] = in_data4[4583:4576];
      mux_data4[135:128] = in_data4[4591:4584];
      mux_data4[143:136] = in_data4[4599:4592];
      mux_data4[151:144] = in_data4[4607:4600];
      mux_data4[159:152] = in_data4[4615:4608];
      mux_data4[167:160] = in_data4[4623:4616];
      mux_data4[175:168] = in_data4[4631:4624];
    end
    'd36: begin
      mux_data0[7:0] = in_data0[4591:4584];
      mux_data0[15:8] = in_data0[4599:4592];
      mux_data0[23:16] = in_data0[4607:4600];
      mux_data0[31:24] = in_data0[4615:4608];
      mux_data0[39:32] = in_data0[4623:4616];
      mux_data0[47:40] = in_data0[4631:4624];
      mux_data0[55:48] = in_data0[4639:4632];
      mux_data0[63:56] = in_data0[4647:4640];
      mux_data0[71:64] = in_data0[4655:4648];
      mux_data0[79:72] = in_data0[4663:4656];
      mux_data0[87:80] = in_data0[4671:4664];
      mux_data0[95:88] = in_data0[4679:4672];
      mux_data0[103:96] = in_data0[4687:4680];
      mux_data0[111:104] = in_data0[4695:4688];
      mux_data0[119:112] = in_data0[4703:4696];
      mux_data0[127:120] = in_data0[4711:4704];
      mux_data0[135:128] = in_data0[4719:4712];
      mux_data0[143:136] = in_data0[4727:4720];
      mux_data0[151:144] = in_data0[4735:4728];
      mux_data0[159:152] = in_data0[4743:4736];
      mux_data0[167:160] = in_data0[4751:4744];
      mux_data0[175:168] = in_data0[4759:4752];
      mux_data1[7:0] = in_data1[4591:4584];
      mux_data1[15:8] = in_data1[4599:4592];
      mux_data1[23:16] = in_data1[4607:4600];
      mux_data1[31:24] = in_data1[4615:4608];
      mux_data1[39:32] = in_data1[4623:4616];
      mux_data1[47:40] = in_data1[4631:4624];
      mux_data1[55:48] = in_data1[4639:4632];
      mux_data1[63:56] = in_data1[4647:4640];
      mux_data1[71:64] = in_data1[4655:4648];
      mux_data1[79:72] = in_data1[4663:4656];
      mux_data1[87:80] = in_data1[4671:4664];
      mux_data1[95:88] = in_data1[4679:4672];
      mux_data1[103:96] = in_data1[4687:4680];
      mux_data1[111:104] = in_data1[4695:4688];
      mux_data1[119:112] = in_data1[4703:4696];
      mux_data1[127:120] = in_data1[4711:4704];
      mux_data1[135:128] = in_data1[4719:4712];
      mux_data1[143:136] = in_data1[4727:4720];
      mux_data1[151:144] = in_data1[4735:4728];
      mux_data1[159:152] = in_data1[4743:4736];
      mux_data1[167:160] = in_data1[4751:4744];
      mux_data1[175:168] = in_data1[4759:4752];
      mux_data2[7:0] = in_data2[4591:4584];
      mux_data2[15:8] = in_data2[4599:4592];
      mux_data2[23:16] = in_data2[4607:4600];
      mux_data2[31:24] = in_data2[4615:4608];
      mux_data2[39:32] = in_data2[4623:4616];
      mux_data2[47:40] = in_data2[4631:4624];
      mux_data2[55:48] = in_data2[4639:4632];
      mux_data2[63:56] = in_data2[4647:4640];
      mux_data2[71:64] = in_data2[4655:4648];
      mux_data2[79:72] = in_data2[4663:4656];
      mux_data2[87:80] = in_data2[4671:4664];
      mux_data2[95:88] = in_data2[4679:4672];
      mux_data2[103:96] = in_data2[4687:4680];
      mux_data2[111:104] = in_data2[4695:4688];
      mux_data2[119:112] = in_data2[4703:4696];
      mux_data2[127:120] = in_data2[4711:4704];
      mux_data2[135:128] = in_data2[4719:4712];
      mux_data2[143:136] = in_data2[4727:4720];
      mux_data2[151:144] = in_data2[4735:4728];
      mux_data2[159:152] = in_data2[4743:4736];
      mux_data2[167:160] = in_data2[4751:4744];
      mux_data2[175:168] = in_data2[4759:4752];
      mux_data3[7:0] = in_data3[4591:4584];
      mux_data3[15:8] = in_data3[4599:4592];
      mux_data3[23:16] = in_data3[4607:4600];
      mux_data3[31:24] = in_data3[4615:4608];
      mux_data3[39:32] = in_data3[4623:4616];
      mux_data3[47:40] = in_data3[4631:4624];
      mux_data3[55:48] = in_data3[4639:4632];
      mux_data3[63:56] = in_data3[4647:4640];
      mux_data3[71:64] = in_data3[4655:4648];
      mux_data3[79:72] = in_data3[4663:4656];
      mux_data3[87:80] = in_data3[4671:4664];
      mux_data3[95:88] = in_data3[4679:4672];
      mux_data3[103:96] = in_data3[4687:4680];
      mux_data3[111:104] = in_data3[4695:4688];
      mux_data3[119:112] = in_data3[4703:4696];
      mux_data3[127:120] = in_data3[4711:4704];
      mux_data3[135:128] = in_data3[4719:4712];
      mux_data3[143:136] = in_data3[4727:4720];
      mux_data3[151:144] = in_data3[4735:4728];
      mux_data3[159:152] = in_data3[4743:4736];
      mux_data3[167:160] = in_data3[4751:4744];
      mux_data3[175:168] = in_data3[4759:4752];
      mux_data4[7:0] = in_data4[4591:4584];
      mux_data4[15:8] = in_data4[4599:4592];
      mux_data4[23:16] = in_data4[4607:4600];
      mux_data4[31:24] = in_data4[4615:4608];
      mux_data4[39:32] = in_data4[4623:4616];
      mux_data4[47:40] = in_data4[4631:4624];
      mux_data4[55:48] = in_data4[4639:4632];
      mux_data4[63:56] = in_data4[4647:4640];
      mux_data4[71:64] = in_data4[4655:4648];
      mux_data4[79:72] = in_data4[4663:4656];
      mux_data4[87:80] = in_data4[4671:4664];
      mux_data4[95:88] = in_data4[4679:4672];
      mux_data4[103:96] = in_data4[4687:4680];
      mux_data4[111:104] = in_data4[4695:4688];
      mux_data4[119:112] = in_data4[4703:4696];
      mux_data4[127:120] = in_data4[4711:4704];
      mux_data4[135:128] = in_data4[4719:4712];
      mux_data4[143:136] = in_data4[4727:4720];
      mux_data4[151:144] = in_data4[4735:4728];
      mux_data4[159:152] = in_data4[4743:4736];
      mux_data4[167:160] = in_data4[4751:4744];
      mux_data4[175:168] = in_data4[4759:4752];
    end
    'd37: begin
      mux_data0[7:0] = in_data0[4719:4712];
      mux_data0[15:8] = in_data0[4727:4720];
      mux_data0[23:16] = in_data0[4735:4728];
      mux_data0[31:24] = in_data0[4743:4736];
      mux_data0[39:32] = in_data0[4751:4744];
      mux_data0[47:40] = in_data0[4759:4752];
      mux_data0[55:48] = in_data0[4767:4760];
      mux_data0[63:56] = in_data0[4775:4768];
      mux_data0[71:64] = in_data0[4783:4776];
      mux_data0[79:72] = in_data0[4791:4784];
      mux_data0[87:80] = in_data0[4799:4792];
      mux_data0[95:88] = in_data0[4807:4800];
      mux_data0[103:96] = in_data0[4815:4808];
      mux_data0[111:104] = in_data0[4823:4816];
      mux_data0[119:112] = in_data0[4831:4824];
      mux_data0[127:120] = in_data0[4839:4832];
      mux_data0[135:128] = in_data0[4847:4840];
      mux_data0[143:136] = in_data0[4855:4848];
      mux_data0[151:144] = in_data0[4863:4856];
      mux_data0[159:152] = in_data0[4871:4864];
      mux_data0[167:160] = in_data0[4879:4872];
      mux_data0[175:168] = in_data0[4887:4880];
      mux_data1[7:0] = in_data1[4719:4712];
      mux_data1[15:8] = in_data1[4727:4720];
      mux_data1[23:16] = in_data1[4735:4728];
      mux_data1[31:24] = in_data1[4743:4736];
      mux_data1[39:32] = in_data1[4751:4744];
      mux_data1[47:40] = in_data1[4759:4752];
      mux_data1[55:48] = in_data1[4767:4760];
      mux_data1[63:56] = in_data1[4775:4768];
      mux_data1[71:64] = in_data1[4783:4776];
      mux_data1[79:72] = in_data1[4791:4784];
      mux_data1[87:80] = in_data1[4799:4792];
      mux_data1[95:88] = in_data1[4807:4800];
      mux_data1[103:96] = in_data1[4815:4808];
      mux_data1[111:104] = in_data1[4823:4816];
      mux_data1[119:112] = in_data1[4831:4824];
      mux_data1[127:120] = in_data1[4839:4832];
      mux_data1[135:128] = in_data1[4847:4840];
      mux_data1[143:136] = in_data1[4855:4848];
      mux_data1[151:144] = in_data1[4863:4856];
      mux_data1[159:152] = in_data1[4871:4864];
      mux_data1[167:160] = in_data1[4879:4872];
      mux_data1[175:168] = in_data1[4887:4880];
      mux_data2[7:0] = in_data2[4719:4712];
      mux_data2[15:8] = in_data2[4727:4720];
      mux_data2[23:16] = in_data2[4735:4728];
      mux_data2[31:24] = in_data2[4743:4736];
      mux_data2[39:32] = in_data2[4751:4744];
      mux_data2[47:40] = in_data2[4759:4752];
      mux_data2[55:48] = in_data2[4767:4760];
      mux_data2[63:56] = in_data2[4775:4768];
      mux_data2[71:64] = in_data2[4783:4776];
      mux_data2[79:72] = in_data2[4791:4784];
      mux_data2[87:80] = in_data2[4799:4792];
      mux_data2[95:88] = in_data2[4807:4800];
      mux_data2[103:96] = in_data2[4815:4808];
      mux_data2[111:104] = in_data2[4823:4816];
      mux_data2[119:112] = in_data2[4831:4824];
      mux_data2[127:120] = in_data2[4839:4832];
      mux_data2[135:128] = in_data2[4847:4840];
      mux_data2[143:136] = in_data2[4855:4848];
      mux_data2[151:144] = in_data2[4863:4856];
      mux_data2[159:152] = in_data2[4871:4864];
      mux_data2[167:160] = in_data2[4879:4872];
      mux_data2[175:168] = in_data2[4887:4880];
      mux_data3[7:0] = in_data3[4719:4712];
      mux_data3[15:8] = in_data3[4727:4720];
      mux_data3[23:16] = in_data3[4735:4728];
      mux_data3[31:24] = in_data3[4743:4736];
      mux_data3[39:32] = in_data3[4751:4744];
      mux_data3[47:40] = in_data3[4759:4752];
      mux_data3[55:48] = in_data3[4767:4760];
      mux_data3[63:56] = in_data3[4775:4768];
      mux_data3[71:64] = in_data3[4783:4776];
      mux_data3[79:72] = in_data3[4791:4784];
      mux_data3[87:80] = in_data3[4799:4792];
      mux_data3[95:88] = in_data3[4807:4800];
      mux_data3[103:96] = in_data3[4815:4808];
      mux_data3[111:104] = in_data3[4823:4816];
      mux_data3[119:112] = in_data3[4831:4824];
      mux_data3[127:120] = in_data3[4839:4832];
      mux_data3[135:128] = in_data3[4847:4840];
      mux_data3[143:136] = in_data3[4855:4848];
      mux_data3[151:144] = in_data3[4863:4856];
      mux_data3[159:152] = in_data3[4871:4864];
      mux_data3[167:160] = in_data3[4879:4872];
      mux_data3[175:168] = in_data3[4887:4880];
      mux_data4[7:0] = in_data4[4719:4712];
      mux_data4[15:8] = in_data4[4727:4720];
      mux_data4[23:16] = in_data4[4735:4728];
      mux_data4[31:24] = in_data4[4743:4736];
      mux_data4[39:32] = in_data4[4751:4744];
      mux_data4[47:40] = in_data4[4759:4752];
      mux_data4[55:48] = in_data4[4767:4760];
      mux_data4[63:56] = in_data4[4775:4768];
      mux_data4[71:64] = in_data4[4783:4776];
      mux_data4[79:72] = in_data4[4791:4784];
      mux_data4[87:80] = in_data4[4799:4792];
      mux_data4[95:88] = in_data4[4807:4800];
      mux_data4[103:96] = in_data4[4815:4808];
      mux_data4[111:104] = in_data4[4823:4816];
      mux_data4[119:112] = in_data4[4831:4824];
      mux_data4[127:120] = in_data4[4839:4832];
      mux_data4[135:128] = in_data4[4847:4840];
      mux_data4[143:136] = in_data4[4855:4848];
      mux_data4[151:144] = in_data4[4863:4856];
      mux_data4[159:152] = in_data4[4871:4864];
      mux_data4[167:160] = in_data4[4879:4872];
      mux_data4[175:168] = in_data4[4887:4880];
    end
    'd38: begin
      mux_data0[7:0] = in_data0[4847:4840];
      mux_data0[15:8] = in_data0[4855:4848];
      mux_data0[23:16] = in_data0[4863:4856];
      mux_data0[31:24] = in_data0[4871:4864];
      mux_data0[39:32] = in_data0[4879:4872];
      mux_data0[47:40] = in_data0[4887:4880];
      mux_data0[55:48] = in_data0[4895:4888];
      mux_data0[63:56] = in_data0[4903:4896];
      mux_data0[71:64] = in_data0[4911:4904];
      mux_data0[79:72] = in_data0[4919:4912];
      mux_data0[87:80] = in_data0[4927:4920];
      mux_data0[95:88] = in_data0[4935:4928];
      mux_data0[103:96] = in_data0[4943:4936];
      mux_data0[111:104] = in_data0[4951:4944];
      mux_data0[119:112] = in_data0[4959:4952];
      mux_data0[127:120] = in_data0[4967:4960];
      mux_data0[135:128] = in_data0[4975:4968];
      mux_data0[143:136] = in_data0[4983:4976];
      mux_data0[151:144] = in_data0[4991:4984];
      mux_data0[159:152] = in_data0[4999:4992];
      mux_data0[167:160] = in_data0[5007:5000];
      mux_data0[175:168] = in_data0[5015:5008];
      mux_data1[7:0] = in_data1[4847:4840];
      mux_data1[15:8] = in_data1[4855:4848];
      mux_data1[23:16] = in_data1[4863:4856];
      mux_data1[31:24] = in_data1[4871:4864];
      mux_data1[39:32] = in_data1[4879:4872];
      mux_data1[47:40] = in_data1[4887:4880];
      mux_data1[55:48] = in_data1[4895:4888];
      mux_data1[63:56] = in_data1[4903:4896];
      mux_data1[71:64] = in_data1[4911:4904];
      mux_data1[79:72] = in_data1[4919:4912];
      mux_data1[87:80] = in_data1[4927:4920];
      mux_data1[95:88] = in_data1[4935:4928];
      mux_data1[103:96] = in_data1[4943:4936];
      mux_data1[111:104] = in_data1[4951:4944];
      mux_data1[119:112] = in_data1[4959:4952];
      mux_data1[127:120] = in_data1[4967:4960];
      mux_data1[135:128] = in_data1[4975:4968];
      mux_data1[143:136] = in_data1[4983:4976];
      mux_data1[151:144] = in_data1[4991:4984];
      mux_data1[159:152] = in_data1[4999:4992];
      mux_data1[167:160] = in_data1[5007:5000];
      mux_data1[175:168] = in_data1[5015:5008];
      mux_data2[7:0] = in_data2[4847:4840];
      mux_data2[15:8] = in_data2[4855:4848];
      mux_data2[23:16] = in_data2[4863:4856];
      mux_data2[31:24] = in_data2[4871:4864];
      mux_data2[39:32] = in_data2[4879:4872];
      mux_data2[47:40] = in_data2[4887:4880];
      mux_data2[55:48] = in_data2[4895:4888];
      mux_data2[63:56] = in_data2[4903:4896];
      mux_data2[71:64] = in_data2[4911:4904];
      mux_data2[79:72] = in_data2[4919:4912];
      mux_data2[87:80] = in_data2[4927:4920];
      mux_data2[95:88] = in_data2[4935:4928];
      mux_data2[103:96] = in_data2[4943:4936];
      mux_data2[111:104] = in_data2[4951:4944];
      mux_data2[119:112] = in_data2[4959:4952];
      mux_data2[127:120] = in_data2[4967:4960];
      mux_data2[135:128] = in_data2[4975:4968];
      mux_data2[143:136] = in_data2[4983:4976];
      mux_data2[151:144] = in_data2[4991:4984];
      mux_data2[159:152] = in_data2[4999:4992];
      mux_data2[167:160] = in_data2[5007:5000];
      mux_data2[175:168] = in_data2[5015:5008];
      mux_data3[7:0] = in_data3[4847:4840];
      mux_data3[15:8] = in_data3[4855:4848];
      mux_data3[23:16] = in_data3[4863:4856];
      mux_data3[31:24] = in_data3[4871:4864];
      mux_data3[39:32] = in_data3[4879:4872];
      mux_data3[47:40] = in_data3[4887:4880];
      mux_data3[55:48] = in_data3[4895:4888];
      mux_data3[63:56] = in_data3[4903:4896];
      mux_data3[71:64] = in_data3[4911:4904];
      mux_data3[79:72] = in_data3[4919:4912];
      mux_data3[87:80] = in_data3[4927:4920];
      mux_data3[95:88] = in_data3[4935:4928];
      mux_data3[103:96] = in_data3[4943:4936];
      mux_data3[111:104] = in_data3[4951:4944];
      mux_data3[119:112] = in_data3[4959:4952];
      mux_data3[127:120] = in_data3[4967:4960];
      mux_data3[135:128] = in_data3[4975:4968];
      mux_data3[143:136] = in_data3[4983:4976];
      mux_data3[151:144] = in_data3[4991:4984];
      mux_data3[159:152] = in_data3[4999:4992];
      mux_data3[167:160] = in_data3[5007:5000];
      mux_data3[175:168] = in_data3[5015:5008];
      mux_data4[7:0] = in_data4[4847:4840];
      mux_data4[15:8] = in_data4[4855:4848];
      mux_data4[23:16] = in_data4[4863:4856];
      mux_data4[31:24] = in_data4[4871:4864];
      mux_data4[39:32] = in_data4[4879:4872];
      mux_data4[47:40] = in_data4[4887:4880];
      mux_data4[55:48] = in_data4[4895:4888];
      mux_data4[63:56] = in_data4[4903:4896];
      mux_data4[71:64] = in_data4[4911:4904];
      mux_data4[79:72] = in_data4[4919:4912];
      mux_data4[87:80] = in_data4[4927:4920];
      mux_data4[95:88] = in_data4[4935:4928];
      mux_data4[103:96] = in_data4[4943:4936];
      mux_data4[111:104] = in_data4[4951:4944];
      mux_data4[119:112] = in_data4[4959:4952];
      mux_data4[127:120] = in_data4[4967:4960];
      mux_data4[135:128] = in_data4[4975:4968];
      mux_data4[143:136] = in_data4[4983:4976];
      mux_data4[151:144] = in_data4[4991:4984];
      mux_data4[159:152] = in_data4[4999:4992];
      mux_data4[167:160] = in_data4[5007:5000];
      mux_data4[175:168] = in_data4[5015:5008];
    end
    'd39: begin
      mux_data0[7:0] = in_data0[4975:4968];
      mux_data0[15:8] = in_data0[4983:4976];
      mux_data0[23:16] = in_data0[4991:4984];
      mux_data0[31:24] = in_data0[4999:4992];
      mux_data0[39:32] = in_data0[5007:5000];
      mux_data0[47:40] = in_data0[5015:5008];
      mux_data0[55:48] = in_data0[5023:5016];
      mux_data0[63:56] = in_data0[5031:5024];
      mux_data0[71:64] = in_data0[5039:5032];
      mux_data0[79:72] = in_data0[5047:5040];
      mux_data0[87:80] = in_data0[5055:5048];
      mux_data0[95:88] = in_data0[5063:5056];
      mux_data0[103:96] = in_data0[5071:5064];
      mux_data0[111:104] = in_data0[5079:5072];
      mux_data0[119:112] = in_data0[5087:5080];
      mux_data0[127:120] = in_data0[5095:5088];
      mux_data0[135:128] = in_data0[5103:5096];
      mux_data0[143:136] = in_data0[5111:5104];
      mux_data0[151:144] = in_data0[5119:5112];
      mux_data0[159:152] = 'd0;
      mux_data0[167:160] = 'd0;
      mux_data0[175:168] = 'd0;
      mux_data1[7:0] = in_data1[4975:4968];
      mux_data1[15:8] = in_data1[4983:4976];
      mux_data1[23:16] = in_data1[4991:4984];
      mux_data1[31:24] = in_data1[4999:4992];
      mux_data1[39:32] = in_data1[5007:5000];
      mux_data1[47:40] = in_data1[5015:5008];
      mux_data1[55:48] = in_data1[5023:5016];
      mux_data1[63:56] = in_data1[5031:5024];
      mux_data1[71:64] = in_data1[5039:5032];
      mux_data1[79:72] = in_data1[5047:5040];
      mux_data1[87:80] = in_data1[5055:5048];
      mux_data1[95:88] = in_data1[5063:5056];
      mux_data1[103:96] = in_data1[5071:5064];
      mux_data1[111:104] = in_data1[5079:5072];
      mux_data1[119:112] = in_data1[5087:5080];
      mux_data1[127:120] = in_data1[5095:5088];
      mux_data1[135:128] = in_data1[5103:5096];
      mux_data1[143:136] = in_data1[5111:5104];
      mux_data1[151:144] = in_data1[5119:5112];
      mux_data1[159:152] = 'd0;
      mux_data1[167:160] = 'd0;
      mux_data1[175:168] = 'd0;
      mux_data2[7:0] = in_data2[4975:4968];
      mux_data2[15:8] = in_data2[4983:4976];
      mux_data2[23:16] = in_data2[4991:4984];
      mux_data2[31:24] = in_data2[4999:4992];
      mux_data2[39:32] = in_data2[5007:5000];
      mux_data2[47:40] = in_data2[5015:5008];
      mux_data2[55:48] = in_data2[5023:5016];
      mux_data2[63:56] = in_data2[5031:5024];
      mux_data2[71:64] = in_data2[5039:5032];
      mux_data2[79:72] = in_data2[5047:5040];
      mux_data2[87:80] = in_data2[5055:5048];
      mux_data2[95:88] = in_data2[5063:5056];
      mux_data2[103:96] = in_data2[5071:5064];
      mux_data2[111:104] = in_data2[5079:5072];
      mux_data2[119:112] = in_data2[5087:5080];
      mux_data2[127:120] = in_data2[5095:5088];
      mux_data2[135:128] = in_data2[5103:5096];
      mux_data2[143:136] = in_data2[5111:5104];
      mux_data2[151:144] = in_data2[5119:5112];
      mux_data2[159:152] = 'd0;
      mux_data2[167:160] = 'd0;
      mux_data2[175:168] = 'd0;
      mux_data3[7:0] = in_data3[4975:4968];
      mux_data3[15:8] = in_data3[4983:4976];
      mux_data3[23:16] = in_data3[4991:4984];
      mux_data3[31:24] = in_data3[4999:4992];
      mux_data3[39:32] = in_data3[5007:5000];
      mux_data3[47:40] = in_data3[5015:5008];
      mux_data3[55:48] = in_data3[5023:5016];
      mux_data3[63:56] = in_data3[5031:5024];
      mux_data3[71:64] = in_data3[5039:5032];
      mux_data3[79:72] = in_data3[5047:5040];
      mux_data3[87:80] = in_data3[5055:5048];
      mux_data3[95:88] = in_data3[5063:5056];
      mux_data3[103:96] = in_data3[5071:5064];
      mux_data3[111:104] = in_data3[5079:5072];
      mux_data3[119:112] = in_data3[5087:5080];
      mux_data3[127:120] = in_data3[5095:5088];
      mux_data3[135:128] = in_data3[5103:5096];
      mux_data3[143:136] = in_data3[5111:5104];
      mux_data3[151:144] = in_data3[5119:5112];
      mux_data3[159:152] = 'd0;
      mux_data3[167:160] = 'd0;
      mux_data3[175:168] = 'd0;
      mux_data4[7:0] = in_data4[4975:4968];
      mux_data4[15:8] = in_data4[4983:4976];
      mux_data4[23:16] = in_data4[4991:4984];
      mux_data4[31:24] = in_data4[4999:4992];
      mux_data4[39:32] = in_data4[5007:5000];
      mux_data4[47:40] = in_data4[5015:5008];
      mux_data4[55:48] = in_data4[5023:5016];
      mux_data4[63:56] = in_data4[5031:5024];
      mux_data4[71:64] = in_data4[5039:5032];
      mux_data4[79:72] = in_data4[5047:5040];
      mux_data4[87:80] = in_data4[5055:5048];
      mux_data4[95:88] = in_data4[5063:5056];
      mux_data4[103:96] = in_data4[5071:5064];
      mux_data4[111:104] = in_data4[5079:5072];
      mux_data4[119:112] = in_data4[5087:5080];
      mux_data4[127:120] = in_data4[5095:5088];
      mux_data4[135:128] = in_data4[5103:5096];
      mux_data4[143:136] = in_data4[5111:5104];
      mux_data4[151:144] = in_data4[5119:5112];
      mux_data4[159:152] = 'd0;
      mux_data4[167:160] = 'd0;
      mux_data4[175:168] = 'd0;
    end
    default: begin
      mux_data0[7:0] = 'd0;
      mux_data0[15:8] = 'd0;
      mux_data0[23:16] = 'd0;
      mux_data0[31:24] = 'd0;
      mux_data0[39:32] = 'd0;
      mux_data0[47:40] = 'd0;
      mux_data0[55:48] = 'd0;
      mux_data0[63:56] = 'd0;
      mux_data0[71:64] = 'd0;
      mux_data0[79:72] = 'd0;
      mux_data0[87:80] = 'd0;
      mux_data0[95:88] = 'd0;
      mux_data0[103:96] = 'd0;
      mux_data0[111:104] = 'd0;
      mux_data0[119:112] = 'd0;
      mux_data0[127:120] = 'd0;
      mux_data0[135:128] = 'd0;
      mux_data0[143:136] = 'd0;
      mux_data0[151:144] = 'd0;
      mux_data0[159:152] = 'd0;
      mux_data0[167:160] = 'd0;
      mux_data0[175:168] = 'd0;
      mux_data1[7:0] = 'd0;
      mux_data1[15:8] = 'd0;
      mux_data1[23:16] = 'd0;
      mux_data1[31:24] = 'd0;
      mux_data1[39:32] = 'd0;
      mux_data1[47:40] = 'd0;
      mux_data1[55:48] = 'd0;
      mux_data1[63:56] = 'd0;
      mux_data1[71:64] = 'd0;
      mux_data1[79:72] = 'd0;
      mux_data1[87:80] = 'd0;
      mux_data1[95:88] = 'd0;
      mux_data1[103:96] = 'd0;
      mux_data1[111:104] = 'd0;
      mux_data1[119:112] = 'd0;
      mux_data1[127:120] = 'd0;
      mux_data1[135:128] = 'd0;
      mux_data1[143:136] = 'd0;
      mux_data1[151:144] = 'd0;
      mux_data1[159:152] = 'd0;
      mux_data1[167:160] = 'd0;
      mux_data1[175:168] = 'd0;
      mux_data2[7:0] = 'd0;
      mux_data2[15:8] = 'd0;
      mux_data2[23:16] = 'd0;
      mux_data2[31:24] = 'd0;
      mux_data2[39:32] = 'd0;
      mux_data2[47:40] = 'd0;
      mux_data2[55:48] = 'd0;
      mux_data2[63:56] = 'd0;
      mux_data2[71:64] = 'd0;
      mux_data2[79:72] = 'd0;
      mux_data2[87:80] = 'd0;
      mux_data2[95:88] = 'd0;
      mux_data2[103:96] = 'd0;
      mux_data2[111:104] = 'd0;
      mux_data2[119:112] = 'd0;
      mux_data2[127:120] = 'd0;
      mux_data2[135:128] = 'd0;
      mux_data2[143:136] = 'd0;
      mux_data2[151:144] = 'd0;
      mux_data2[159:152] = 'd0;
      mux_data2[167:160] = 'd0;
      mux_data2[175:168] = 'd0;
      mux_data3[7:0] = 'd0;
      mux_data3[15:8] = 'd0;
      mux_data3[23:16] = 'd0;
      mux_data3[31:24] = 'd0;
      mux_data3[39:32] = 'd0;
      mux_data3[47:40] = 'd0;
      mux_data3[55:48] = 'd0;
      mux_data3[63:56] = 'd0;
      mux_data3[71:64] = 'd0;
      mux_data3[79:72] = 'd0;
      mux_data3[87:80] = 'd0;
      mux_data3[95:88] = 'd0;
      mux_data3[103:96] = 'd0;
      mux_data3[111:104] = 'd0;
      mux_data3[119:112] = 'd0;
      mux_data3[127:120] = 'd0;
      mux_data3[135:128] = 'd0;
      mux_data3[143:136] = 'd0;
      mux_data3[151:144] = 'd0;
      mux_data3[159:152] = 'd0;
      mux_data3[167:160] = 'd0;
      mux_data3[175:168] = 'd0;
      mux_data4[7:0] = 'd0;
      mux_data4[15:8] = 'd0;
      mux_data4[23:16] = 'd0;
      mux_data4[31:24] = 'd0;
      mux_data4[39:32] = 'd0;
      mux_data4[47:40] = 'd0;
      mux_data4[55:48] = 'd0;
      mux_data4[63:56] = 'd0;
      mux_data4[71:64] = 'd0;
      mux_data4[79:72] = 'd0;
      mux_data4[87:80] = 'd0;
      mux_data4[95:88] = 'd0;
      mux_data4[103:96] = 'd0;
      mux_data4[111:104] = 'd0;
      mux_data4[119:112] = 'd0;
      mux_data4[127:120] = 'd0;
      mux_data4[135:128] = 'd0;
      mux_data4[143:136] = 'd0;
      mux_data4[151:144] = 'd0;
      mux_data4[159:152] = 'd0;
      mux_data4[167:160] = 'd0;
      mux_data4[175:168] = 'd0;
    end
  endcase
end



always @(posedge clk) begin
  if (!rst_n) 
    buffer_data_0 <= 'd0;
  else if (!buffer_mode && fill_zero)
    buffer_data_0 <= 'd0;
  else if (!buffer_mode && buffer_we)
    buffer_data_0 <= mux_data0;
  else if (buffer_mode && buffer_we)
    buffer_data_0 <= mux_data0;
end

always @(posedge clk) begin
  if (!rst_n) 
    buffer_data_1 <= 'd0; 
  else if (buffer_we)
    buffer_data_1 <= buffer_data_0;
end

always @(posedge clk) begin
  if (!rst_n) 
    buffer_data_2 <= 'd0;    
  else if (!buffer_mode && buffer_we)
    buffer_data_2 <= buffer_data_1;
  else if (buffer_mode && buffer_we)
    buffer_data_2 <= mux_data1;
end

always @(posedge clk) begin
  if (!rst_n) 
    buffer_data_3 <= 'd0;    
  else if (buffer_we)
    buffer_data_3 <= buffer_data_2;
end

always @(posedge clk) begin
  if (!rst_n) 
    buffer_data_4 <= 'd0;    
  else if (!buffer_mode && buffer_we)
    buffer_data_4 <= buffer_data_3;
  else if (buffer_mode && buffer_we)
    buffer_data_4 <= mux_data2;
end

always @(posedge clk) begin
  if (!rst_n) 
    buffer_data_5 <= 'd0;    
  else if (buffer_we)
    buffer_data_5 <= buffer_data_4;
end


always @(posedge clk) begin
  if (!rst_n) 
    buffer_data_6 <= 'd0;    
  else if (!buffer_mode && buffer_we)
    buffer_data_6 <= buffer_data_5;
  else if (buffer_mode && buffer_we)
    buffer_data_6 <= mux_data3;
end

always @(posedge clk) begin
  if (!rst_n) 
    buffer_data_7 <= 'd0;    
  else if (buffer_we)
    buffer_data_7 <= buffer_data_6;
end

always @(posedge clk) begin
  if (!rst_n) 
    buffer_data_8 <= 'd0;    
  else if (!buffer_mode && buffer_we)
    buffer_data_8 <= buffer_data_7;
  else if (buffer_mode && buffer_we)
    buffer_data_8 <= mux_data4;
end

always @(posedge clk) begin
  if (!rst_n) 
    buffer_data_9 <= 'd0;    
  else if (buffer_we)
    buffer_data_9 <= buffer_data_8;
end


endmodule 