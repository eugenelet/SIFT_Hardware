module Gaussian_Blur_3x3(
  clk,
  rst_n,
  buffer_data_0,
  buffer_data_1,
  buffer_data_2,
  current_col,
  blur_out,
  start,
  done
);

input                 clk;
input                 rst_n;
input                 start;
output                done;
input         [5:0]   current_col;
input       [175:0]   buffer_data_0;
input       [175:0]   buffer_data_1;
input       [175:0]   buffer_data_2;
output reg  [127:0]   blur_out; // wire

parameter  ST_MUX         = 0,
           ST_MUL         = 1,
           ST_ADD         = 2,
           ST_UPDATE      = 3;
reg     [2:0] current_state,
              next_state;
assign done = (current_state==ST_UPDATE) ? 1 : 0;

wire       [23:0]  G_Kernel_3x3_0;
wire       [23:0]  G_Kernel_3x3_1;
assign  G_Kernel_3x3_0[7:0]   = 8'h17; //BC5428; //18'b00_0101_1110_1111_0001;//'d092717;
assign  G_Kernel_3x3_0[15:8]  = 8'h1E; //7ABFF3; //18'b00_0111_1001_1110_1010;//'d119061;
assign  G_Kernel_3x3_0[23:16] = 8'h17; //BC5428; //18'b00_0101_1110_1111_0001;//'d092717;
assign  G_Kernel_3x3_1[7:0]   = 8'h1E; //7ABFF3; //18'b00_0111_1001_1110_1010;//'d119061;
assign  G_Kernel_3x3_1[15:8]  = 8'h27; //23AF8E; //18'b00_1001_1100_1000_1110;//'d152888;
assign  G_Kernel_3x3_1[23:16] = 8'h1E; //7ABFF3; //18'b00_0111_1001_1110_1011;//'d119061;

reg    [23:0]    layer0[0:15]; //wire
reg    [23:0]    layer1[0:15]; //wire
reg    [23:0]    layer2[0:15]; //wire
always @(posedge clk) begin
  if(!rst_n) begin
    layer0[0] <= 'd0;
    layer0[1] <= 'd0;
    layer0[2] <= 'd0;
    layer0[3] <= 'd0;
    layer0[4] <= 'd0;
    layer0[5] <= 'd0;
    layer0[6] <= 'd0;
    layer0[7] <= 'd0;
    layer0[8] <= 'd0;
    layer0[9] <= 'd0;
    layer0[10] <= 'd0;
    layer0[11] <= 'd0;
    layer0[12] <= 'd0;
    layer0[13] <= 'd0;
    layer0[14] <= 'd0;
    layer0[15] <= 'd0;
    layer1[0] <= 'd0;
    layer1[1] <= 'd0;
    layer1[2] <= 'd0;
    layer1[3] <= 'd0;
    layer1[4] <= 'd0;
    layer1[5] <= 'd0;
    layer1[6] <= 'd0;
    layer1[7] <= 'd0;
    layer1[8] <= 'd0;
    layer1[9] <= 'd0;
    layer1[10] <= 'd0;
    layer1[11] <= 'd0;
    layer1[12] <= 'd0;
    layer1[13] <= 'd0;
    layer1[14] <= 'd0;
    layer1[15] <= 'd0;
    layer2[0] <= 'd0;
    layer2[1] <= 'd0;
    layer2[2] <= 'd0;
    layer2[3] <= 'd0;
    layer2[4] <= 'd0;
    layer2[5] <= 'd0;
    layer2[6] <= 'd0;
    layer2[7] <= 'd0;
    layer2[8] <= 'd0;
    layer2[9] <= 'd0;
    layer2[10] <= 'd0;
    layer2[11] <= 'd0;
    layer2[12] <= 'd0;
    layer2[13] <= 'd0;
    layer2[14] <= 'd0;
    layer2[15] <= 'd0;
  end
  else if(current_state==ST_MUX) begin
    case(current_col)
      'd0: begin
        layer0[0][7:0] <= 0;
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= 0;
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= 0;
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd1: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd2: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd3: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd4: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd5: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd6: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd7: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd8: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd9: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd10: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd11: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd12: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd13: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd14: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd15: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd16: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd17: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd18: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd19: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd20: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd21: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd22: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd23: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd24: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd25: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd26: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd27: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd28: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd29: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd30: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd31: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd32: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd33: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd34: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd35: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd36: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd37: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd38: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= buffer_data_2[159:152];
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= buffer_data_1[159:152];
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= buffer_data_0[159:152];
    end
      'd39: begin
        layer0[0][7:0] <= buffer_data_2[23:16];
        layer0[0][15:8] <= buffer_data_2[31:24];
        layer0[0][23:16] <= buffer_data_2[39:32];
        layer1[0][7:0] <= buffer_data_1[23:16];
        layer1[0][15:8] <= buffer_data_1[31:24];
        layer1[0][23:16] <= buffer_data_1[39:32];
        layer2[0][7:0] <= buffer_data_0[23:16];
        layer2[0][15:8] <= buffer_data_0[31:24];
        layer2[0][23:16] <= buffer_data_0[39:32];
        layer0[1][7:0] <= buffer_data_2[31:24];
        layer0[1][15:8] <= buffer_data_2[39:32];
        layer0[1][23:16] <= buffer_data_2[47:40];
        layer1[1][7:0] <= buffer_data_1[31:24];
        layer1[1][15:8] <= buffer_data_1[39:32];
        layer1[1][23:16] <= buffer_data_1[47:40];
        layer2[1][7:0] <= buffer_data_0[31:24];
        layer2[1][15:8] <= buffer_data_0[39:32];
        layer2[1][23:16] <= buffer_data_0[47:40];
        layer0[2][7:0] <= buffer_data_2[39:32];
        layer0[2][15:8] <= buffer_data_2[47:40];
        layer0[2][23:16] <= buffer_data_2[55:48];
        layer1[2][7:0] <= buffer_data_1[39:32];
        layer1[2][15:8] <= buffer_data_1[47:40];
        layer1[2][23:16] <= buffer_data_1[55:48];
        layer2[2][7:0] <= buffer_data_0[39:32];
        layer2[2][15:8] <= buffer_data_0[47:40];
        layer2[2][23:16] <= buffer_data_0[55:48];
        layer0[3][7:0] <= buffer_data_2[47:40];
        layer0[3][15:8] <= buffer_data_2[55:48];
        layer0[3][23:16] <= buffer_data_2[63:56];
        layer1[3][7:0] <= buffer_data_1[47:40];
        layer1[3][15:8] <= buffer_data_1[55:48];
        layer1[3][23:16] <= buffer_data_1[63:56];
        layer2[3][7:0] <= buffer_data_0[47:40];
        layer2[3][15:8] <= buffer_data_0[55:48];
        layer2[3][23:16] <= buffer_data_0[63:56];
        layer0[4][7:0] <= buffer_data_2[55:48];
        layer0[4][15:8] <= buffer_data_2[63:56];
        layer0[4][23:16] <= buffer_data_2[71:64];
        layer1[4][7:0] <= buffer_data_1[55:48];
        layer1[4][15:8] <= buffer_data_1[63:56];
        layer1[4][23:16] <= buffer_data_1[71:64];
        layer2[4][7:0] <= buffer_data_0[55:48];
        layer2[4][15:8] <= buffer_data_0[63:56];
        layer2[4][23:16] <= buffer_data_0[71:64];
        layer0[5][7:0] <= buffer_data_2[63:56];
        layer0[5][15:8] <= buffer_data_2[71:64];
        layer0[5][23:16] <= buffer_data_2[79:72];
        layer1[5][7:0] <= buffer_data_1[63:56];
        layer1[5][15:8] <= buffer_data_1[71:64];
        layer1[5][23:16] <= buffer_data_1[79:72];
        layer2[5][7:0] <= buffer_data_0[63:56];
        layer2[5][15:8] <= buffer_data_0[71:64];
        layer2[5][23:16] <= buffer_data_0[79:72];
        layer0[6][7:0] <= buffer_data_2[71:64];
        layer0[6][15:8] <= buffer_data_2[79:72];
        layer0[6][23:16] <= buffer_data_2[87:80];
        layer1[6][7:0] <= buffer_data_1[71:64];
        layer1[6][15:8] <= buffer_data_1[79:72];
        layer1[6][23:16] <= buffer_data_1[87:80];
        layer2[6][7:0] <= buffer_data_0[71:64];
        layer2[6][15:8] <= buffer_data_0[79:72];
        layer2[6][23:16] <= buffer_data_0[87:80];
        layer0[7][7:0] <= buffer_data_2[79:72];
        layer0[7][15:8] <= buffer_data_2[87:80];
        layer0[7][23:16] <= buffer_data_2[95:88];
        layer1[7][7:0] <= buffer_data_1[79:72];
        layer1[7][15:8] <= buffer_data_1[87:80];
        layer1[7][23:16] <= buffer_data_1[95:88];
        layer2[7][7:0] <= buffer_data_0[79:72];
        layer2[7][15:8] <= buffer_data_0[87:80];
        layer2[7][23:16] <= buffer_data_0[95:88];
        layer0[8][7:0] <= buffer_data_2[87:80];
        layer0[8][15:8] <= buffer_data_2[95:88];
        layer0[8][23:16] <= buffer_data_2[103:96];
        layer1[8][7:0] <= buffer_data_1[87:80];
        layer1[8][15:8] <= buffer_data_1[95:88];
        layer1[8][23:16] <= buffer_data_1[103:96];
        layer2[8][7:0] <= buffer_data_0[87:80];
        layer2[8][15:8] <= buffer_data_0[95:88];
        layer2[8][23:16] <= buffer_data_0[103:96];
        layer0[9][7:0] <= buffer_data_2[95:88];
        layer0[9][15:8] <= buffer_data_2[103:96];
        layer0[9][23:16] <= buffer_data_2[111:104];
        layer1[9][7:0] <= buffer_data_1[95:88];
        layer1[9][15:8] <= buffer_data_1[103:96];
        layer1[9][23:16] <= buffer_data_1[111:104];
        layer2[9][7:0] <= buffer_data_0[95:88];
        layer2[9][15:8] <= buffer_data_0[103:96];
        layer2[9][23:16] <= buffer_data_0[111:104];
        layer0[10][7:0] <= buffer_data_2[103:96];
        layer0[10][15:8] <= buffer_data_2[111:104];
        layer0[10][23:16] <= buffer_data_2[119:112];
        layer1[10][7:0] <= buffer_data_1[103:96];
        layer1[10][15:8] <= buffer_data_1[111:104];
        layer1[10][23:16] <= buffer_data_1[119:112];
        layer2[10][7:0] <= buffer_data_0[103:96];
        layer2[10][15:8] <= buffer_data_0[111:104];
        layer2[10][23:16] <= buffer_data_0[119:112];
        layer0[11][7:0] <= buffer_data_2[111:104];
        layer0[11][15:8] <= buffer_data_2[119:112];
        layer0[11][23:16] <= buffer_data_2[127:120];
        layer1[11][7:0] <= buffer_data_1[111:104];
        layer1[11][15:8] <= buffer_data_1[119:112];
        layer1[11][23:16] <= buffer_data_1[127:120];
        layer2[11][7:0] <= buffer_data_0[111:104];
        layer2[11][15:8] <= buffer_data_0[119:112];
        layer2[11][23:16] <= buffer_data_0[127:120];
        layer0[12][7:0] <= buffer_data_2[119:112];
        layer0[12][15:8] <= buffer_data_2[127:120];
        layer0[12][23:16] <= buffer_data_2[135:128];
        layer1[12][7:0] <= buffer_data_1[119:112];
        layer1[12][15:8] <= buffer_data_1[127:120];
        layer1[12][23:16] <= buffer_data_1[135:128];
        layer2[12][7:0] <= buffer_data_0[119:112];
        layer2[12][15:8] <= buffer_data_0[127:120];
        layer2[12][23:16] <= buffer_data_0[135:128];
        layer0[13][7:0] <= buffer_data_2[127:120];
        layer0[13][15:8] <= buffer_data_2[135:128];
        layer0[13][23:16] <= buffer_data_2[143:136];
        layer1[13][7:0] <= buffer_data_1[127:120];
        layer1[13][15:8] <= buffer_data_1[135:128];
        layer1[13][23:16] <= buffer_data_1[143:136];
        layer2[13][7:0] <= buffer_data_0[127:120];
        layer2[13][15:8] <= buffer_data_0[135:128];
        layer2[13][23:16] <= buffer_data_0[143:136];
        layer0[14][7:0] <= buffer_data_2[135:128];
        layer0[14][15:8] <= buffer_data_2[143:136];
        layer0[14][23:16] <= buffer_data_2[151:144];
        layer1[14][7:0] <= buffer_data_1[135:128];
        layer1[14][15:8] <= buffer_data_1[143:136];
        layer1[14][23:16] <= buffer_data_1[151:144];
        layer2[14][7:0] <= buffer_data_0[135:128];
        layer2[14][15:8] <= buffer_data_0[143:136];
        layer2[14][23:16] <= buffer_data_0[151:144];
        layer0[15][7:0] <= buffer_data_2[143:136];
        layer0[15][15:8] <= buffer_data_2[151:144];
        layer0[15][23:16] <= 0;
        layer1[15][7:0] <= buffer_data_1[143:136];
        layer1[15][15:8] <= buffer_data_1[151:144];
        layer1[15][23:16] <= 0;
        layer2[15][7:0] <= buffer_data_0[143:136];
        layer2[15][15:8] <= buffer_data_0[151:144];
        layer2[15][23:16] <= 0;
    end
      default: begin
        layer0[0][7:0] <= 'd0;
        layer0[0][15:8] <= 'd0;
        layer0[0][23:16] <= 'd0;
        layer1[0][7:0] <= 'd0;
        layer1[0][15:8] <= 'd0;
        layer1[0][23:16] <= 'd0;
        layer2[0][7:0] <= 'd0;
        layer2[0][15:8] <= 'd0;
        layer2[0][23:16] <= 'd0;
        layer0[1][7:0] <= 'd0;
        layer0[1][15:8] <= 'd0;
        layer0[1][23:16] <= 'd0;
        layer1[1][7:0] <= 'd0;
        layer1[1][15:8] <= 'd0;
        layer1[1][23:16] <= 'd0;
        layer2[1][7:0] <= 'd0;
        layer2[1][15:8] <= 'd0;
        layer2[1][23:16] <= 'd0;
        layer0[2][7:0] <= 'd0;
        layer0[2][15:8] <= 'd0;
        layer0[2][23:16] <= 'd0;
        layer1[2][7:0] <= 'd0;
        layer1[2][15:8] <= 'd0;
        layer1[2][23:16] <= 'd0;
        layer2[2][7:0] <= 'd0;
        layer2[2][15:8] <= 'd0;
        layer2[2][23:16] <= 'd0;
        layer0[3][7:0] <= 'd0;
        layer0[3][15:8] <= 'd0;
        layer0[3][23:16] <= 'd0;
        layer1[3][7:0] <= 'd0;
        layer1[3][15:8] <= 'd0;
        layer1[3][23:16] <= 'd0;
        layer2[3][7:0] <= 'd0;
        layer2[3][15:8] <= 'd0;
        layer2[3][23:16] <= 'd0;
        layer0[4][7:0] <= 'd0;
        layer0[4][15:8] <= 'd0;
        layer0[4][23:16] <= 'd0;
        layer1[4][7:0] <= 'd0;
        layer1[4][15:8] <= 'd0;
        layer1[4][23:16] <= 'd0;
        layer2[4][7:0] <= 'd0;
        layer2[4][15:8] <= 'd0;
        layer2[4][23:16] <= 'd0;
        layer0[5][7:0] <= 'd0;
        layer0[5][15:8] <= 'd0;
        layer0[5][23:16] <= 'd0;
        layer1[5][7:0] <= 'd0;
        layer1[5][15:8] <= 'd0;
        layer1[5][23:16] <= 'd0;
        layer2[5][7:0] <= 'd0;
        layer2[5][15:8] <= 'd0;
        layer2[5][23:16] <= 'd0;
        layer0[6][7:0] <= 'd0;
        layer0[6][15:8] <= 'd0;
        layer0[6][23:16] <= 'd0;
        layer1[6][7:0] <= 'd0;
        layer1[6][15:8] <= 'd0;
        layer1[6][23:16] <= 'd0;
        layer2[6][7:0] <= 'd0;
        layer2[6][15:8] <= 'd0;
        layer2[6][23:16] <= 'd0;
        layer0[7][7:0] <= 'd0;
        layer0[7][15:8] <= 'd0;
        layer0[7][23:16] <= 'd0;
        layer1[7][7:0] <= 'd0;
        layer1[7][15:8] <= 'd0;
        layer1[7][23:16] <= 'd0;
        layer2[7][7:0] <= 'd0;
        layer2[7][15:8] <= 'd0;
        layer2[7][23:16] <= 'd0;
        layer0[8][7:0] <= 'd0;
        layer0[8][15:8] <= 'd0;
        layer0[8][23:16] <= 'd0;
        layer1[8][7:0] <= 'd0;
        layer1[8][15:8] <= 'd0;
        layer1[8][23:16] <= 'd0;
        layer2[8][7:0] <= 'd0;
        layer2[8][15:8] <= 'd0;
        layer2[8][23:16] <= 'd0;
        layer0[9][7:0] <= 'd0;
        layer0[9][15:8] <= 'd0;
        layer0[9][23:16] <= 'd0;
        layer1[9][7:0] <= 'd0;
        layer1[9][15:8] <= 'd0;
        layer1[9][23:16] <= 'd0;
        layer2[9][7:0] <= 'd0;
        layer2[9][15:8] <= 'd0;
        layer2[9][23:16] <= 'd0;
        layer0[10][7:0] <= 'd0;
        layer0[10][15:8] <= 'd0;
        layer0[10][23:16] <= 'd0;
        layer1[10][7:0] <= 'd0;
        layer1[10][15:8] <= 'd0;
        layer1[10][23:16] <= 'd0;
        layer2[10][7:0] <= 'd0;
        layer2[10][15:8] <= 'd0;
        layer2[10][23:16] <= 'd0;
        layer0[11][7:0] <= 'd0;
        layer0[11][15:8] <= 'd0;
        layer0[11][23:16] <= 'd0;
        layer1[11][7:0] <= 'd0;
        layer1[11][15:8] <= 'd0;
        layer1[11][23:16] <= 'd0;
        layer2[11][7:0] <= 'd0;
        layer2[11][15:8] <= 'd0;
        layer2[11][23:16] <= 'd0;
        layer0[12][7:0] <= 'd0;
        layer0[12][15:8] <= 'd0;
        layer0[12][23:16] <= 'd0;
        layer1[12][7:0] <= 'd0;
        layer1[12][15:8] <= 'd0;
        layer1[12][23:16] <= 'd0;
        layer2[12][7:0] <= 'd0;
        layer2[12][15:8] <= 'd0;
        layer2[12][23:16] <= 'd0;
        layer0[13][7:0] <= 'd0;
        layer0[13][15:8] <= 'd0;
        layer0[13][23:16] <= 'd0;
        layer1[13][7:0] <= 'd0;
        layer1[13][15:8] <= 'd0;
        layer1[13][23:16] <= 'd0;
        layer2[13][7:0] <= 'd0;
        layer2[13][15:8] <= 'd0;
        layer2[13][23:16] <= 'd0;
        layer0[14][7:0] <= 'd0;
        layer0[14][15:8] <= 'd0;
        layer0[14][23:16] <= 'd0;
        layer1[14][7:0] <= 'd0;
        layer1[14][15:8] <= 'd0;
        layer1[14][23:16] <= 'd0;
        layer2[14][7:0] <= 'd0;
        layer2[14][15:8] <= 'd0;
        layer2[14][23:16] <= 'd0;
        layer0[15][7:0] <= 'd0;
        layer0[15][15:8] <= 'd0;
        layer0[15][23:16] <= 'd0;
        layer1[15][7:0] <= 'd0;
        layer1[15][15:8] <= 'd0;
        layer1[15][23:16] <= 'd0;
        layer2[15][7:0] <= 'd0;
        layer2[15][15:8] <= 'd0;
        layer2[15][23:16] <= 'd0;
      end
    endcase
  end
end

reg  [15:0]  kernel_img_mul_0[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_0[0] <= 'd0;
    kernel_img_mul_0[1] <= 'd0;
    kernel_img_mul_0[2] <= 'd0;
    kernel_img_mul_0[3] <= 'd0;
    kernel_img_mul_0[4] <= 'd0;
    kernel_img_mul_0[5] <= 'd0;
    kernel_img_mul_0[6] <= 'd0;
    kernel_img_mul_0[7] <= 'd0;
    kernel_img_mul_0[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_0[0] <= { {8{1'b0}},layer0[0][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_0[1] <= { {8{1'b0}},layer0[0][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_0[2] <= { {8{1'b0}},layer0[0][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_0[3] <= { {8{1'b0}},layer1[0][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_0[4] <= { {8{1'b0}},layer1[0][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_0[5] <= { {8{1'b0}},layer1[0][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_0[6] <= { {8{1'b0}},layer2[0][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_0[7] <= { {8{1'b0}},layer2[0][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_0[8] <= { {8{1'b0}},layer2[0][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_0;
reg  [15:0]  kernel_img_sum_2_0;
reg  [15:0]  kernel_img_sum_3_0;
reg  [15:0]  kernel_img_sum_4_0;
reg  [15:0]  kernel_img_sum_5_0;
reg  [15:0]  kernel_img_sum_6_0;
reg  [15:0]  kernel_img_sum_7_0;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_0 <= kernel_img_mul_0[0] + kernel_img_mul_0[1] + kernel_img_mul_0[2] + kernel_img_mul_0[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_0 <= kernel_img_mul_0[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_0 <= kernel_img_mul_0[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_0 <= kernel_img_mul_0[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_0 <= kernel_img_mul_0[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_0 <= kernel_img_mul_0[8];
  end
end
always@(*) begin
  kernel_img_sum_7_0 = kernel_img_sum_1_0 + kernel_img_sum_2_0 + kernel_img_sum_3_0 + kernel_img_sum_4_0 + kernel_img_sum_5_0 + kernel_img_sum_6_0;
end
reg  [15:0]  kernel_img_mul_1[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_1[0] <= 'd0;
    kernel_img_mul_1[1] <= 'd0;
    kernel_img_mul_1[2] <= 'd0;
    kernel_img_mul_1[3] <= 'd0;
    kernel_img_mul_1[4] <= 'd0;
    kernel_img_mul_1[5] <= 'd0;
    kernel_img_mul_1[6] <= 'd0;
    kernel_img_mul_1[7] <= 'd0;
    kernel_img_mul_1[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_1[0] <= { {8{1'b0}},layer0[1][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_1[1] <= { {8{1'b0}},layer0[1][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_1[2] <= { {8{1'b0}},layer0[1][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_1[3] <= { {8{1'b0}},layer1[1][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_1[4] <= { {8{1'b0}},layer1[1][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_1[5] <= { {8{1'b0}},layer1[1][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_1[6] <= { {8{1'b0}},layer2[1][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_1[7] <= { {8{1'b0}},layer2[1][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_1[8] <= { {8{1'b0}},layer2[1][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_1;
reg  [15:0]  kernel_img_sum_2_1;
reg  [15:0]  kernel_img_sum_3_1;
reg  [15:0]  kernel_img_sum_4_1;
reg  [15:0]  kernel_img_sum_5_1;
reg  [15:0]  kernel_img_sum_6_1;
reg  [15:0]  kernel_img_sum_7_1;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_1 <= kernel_img_mul_1[0] + kernel_img_mul_1[1] + kernel_img_mul_1[2] + kernel_img_mul_1[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_1 <= kernel_img_mul_1[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_1 <= kernel_img_mul_1[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_1 <= kernel_img_mul_1[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_1 <= kernel_img_mul_1[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_1 <= kernel_img_mul_1[8];
  end
end
always@(*) begin
  kernel_img_sum_7_1 = kernel_img_sum_1_1 + kernel_img_sum_2_1 + kernel_img_sum_3_1 + kernel_img_sum_4_1 + kernel_img_sum_5_1 + kernel_img_sum_6_1;
end
reg  [15:0]  kernel_img_mul_2[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_2[0] <= 'd0;
    kernel_img_mul_2[1] <= 'd0;
    kernel_img_mul_2[2] <= 'd0;
    kernel_img_mul_2[3] <= 'd0;
    kernel_img_mul_2[4] <= 'd0;
    kernel_img_mul_2[5] <= 'd0;
    kernel_img_mul_2[6] <= 'd0;
    kernel_img_mul_2[7] <= 'd0;
    kernel_img_mul_2[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_2[0] <= { {8{1'b0}},layer0[2][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_2[1] <= { {8{1'b0}},layer0[2][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_2[2] <= { {8{1'b0}},layer0[2][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_2[3] <= { {8{1'b0}},layer1[2][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_2[4] <= { {8{1'b0}},layer1[2][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_2[5] <= { {8{1'b0}},layer1[2][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_2[6] <= { {8{1'b0}},layer2[2][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_2[7] <= { {8{1'b0}},layer2[2][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_2[8] <= { {8{1'b0}},layer2[2][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_2;
reg  [15:0]  kernel_img_sum_2_2;
reg  [15:0]  kernel_img_sum_3_2;
reg  [15:0]  kernel_img_sum_4_2;
reg  [15:0]  kernel_img_sum_5_2;
reg  [15:0]  kernel_img_sum_6_2;
reg  [15:0]  kernel_img_sum_7_2;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_2 <= kernel_img_mul_2[0] + kernel_img_mul_2[1] + kernel_img_mul_2[2] + kernel_img_mul_2[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_2 <= kernel_img_mul_2[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_2 <= kernel_img_mul_2[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_2 <= kernel_img_mul_2[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_2 <= kernel_img_mul_2[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_2 <= kernel_img_mul_2[8];
  end
end
always@(*) begin
  kernel_img_sum_7_2 = kernel_img_sum_1_2 + kernel_img_sum_2_2 + kernel_img_sum_3_2 + kernel_img_sum_4_2 + kernel_img_sum_5_2 + kernel_img_sum_6_2;
end
reg  [15:0]  kernel_img_mul_3[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_3[0] <= 'd0;
    kernel_img_mul_3[1] <= 'd0;
    kernel_img_mul_3[2] <= 'd0;
    kernel_img_mul_3[3] <= 'd0;
    kernel_img_mul_3[4] <= 'd0;
    kernel_img_mul_3[5] <= 'd0;
    kernel_img_mul_3[6] <= 'd0;
    kernel_img_mul_3[7] <= 'd0;
    kernel_img_mul_3[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_3[0] <= { {8{1'b0}},layer0[3][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_3[1] <= { {8{1'b0}},layer0[3][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_3[2] <= { {8{1'b0}},layer0[3][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_3[3] <= { {8{1'b0}},layer1[3][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_3[4] <= { {8{1'b0}},layer1[3][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_3[5] <= { {8{1'b0}},layer1[3][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_3[6] <= { {8{1'b0}},layer2[3][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_3[7] <= { {8{1'b0}},layer2[3][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_3[8] <= { {8{1'b0}},layer2[3][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_3;
reg  [15:0]  kernel_img_sum_2_3;
reg  [15:0]  kernel_img_sum_3_3;
reg  [15:0]  kernel_img_sum_4_3;
reg  [15:0]  kernel_img_sum_5_3;
reg  [15:0]  kernel_img_sum_6_3;
reg  [15:0]  kernel_img_sum_7_3;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_3 <= kernel_img_mul_3[0] + kernel_img_mul_3[1] + kernel_img_mul_3[2] + kernel_img_mul_3[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_3 <= kernel_img_mul_3[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_3 <= kernel_img_mul_3[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_3 <= kernel_img_mul_3[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_3 <= kernel_img_mul_3[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_3 <= kernel_img_mul_3[8];
  end
end
always@(*) begin
  kernel_img_sum_7_3 = kernel_img_sum_1_3 + kernel_img_sum_2_3 + kernel_img_sum_3_3 + kernel_img_sum_4_3 + kernel_img_sum_5_3 + kernel_img_sum_6_3;
end
reg  [15:0]  kernel_img_mul_4[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_4[0] <= 'd0;
    kernel_img_mul_4[1] <= 'd0;
    kernel_img_mul_4[2] <= 'd0;
    kernel_img_mul_4[3] <= 'd0;
    kernel_img_mul_4[4] <= 'd0;
    kernel_img_mul_4[5] <= 'd0;
    kernel_img_mul_4[6] <= 'd0;
    kernel_img_mul_4[7] <= 'd0;
    kernel_img_mul_4[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_4[0] <= { {8{1'b0}},layer0[4][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_4[1] <= { {8{1'b0}},layer0[4][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_4[2] <= { {8{1'b0}},layer0[4][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_4[3] <= { {8{1'b0}},layer1[4][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_4[4] <= { {8{1'b0}},layer1[4][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_4[5] <= { {8{1'b0}},layer1[4][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_4[6] <= { {8{1'b0}},layer2[4][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_4[7] <= { {8{1'b0}},layer2[4][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_4[8] <= { {8{1'b0}},layer2[4][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_4;
reg  [15:0]  kernel_img_sum_2_4;
reg  [15:0]  kernel_img_sum_3_4;
reg  [15:0]  kernel_img_sum_4_4;
reg  [15:0]  kernel_img_sum_5_4;
reg  [15:0]  kernel_img_sum_6_4;
reg  [15:0]  kernel_img_sum_7_4;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_4 <= kernel_img_mul_4[0] + kernel_img_mul_4[1] + kernel_img_mul_4[2] + kernel_img_mul_4[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_4 <= kernel_img_mul_4[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_4 <= kernel_img_mul_4[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_4 <= kernel_img_mul_4[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_4 <= kernel_img_mul_4[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_4 <= kernel_img_mul_4[8];
  end
end
always@(*) begin
  kernel_img_sum_7_4 = kernel_img_sum_1_4 + kernel_img_sum_2_4 + kernel_img_sum_3_4 + kernel_img_sum_4_4 + kernel_img_sum_5_4 + kernel_img_sum_6_4;
end
reg  [15:0]  kernel_img_mul_5[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_5[0] <= 'd0;
    kernel_img_mul_5[1] <= 'd0;
    kernel_img_mul_5[2] <= 'd0;
    kernel_img_mul_5[3] <= 'd0;
    kernel_img_mul_5[4] <= 'd0;
    kernel_img_mul_5[5] <= 'd0;
    kernel_img_mul_5[6] <= 'd0;
    kernel_img_mul_5[7] <= 'd0;
    kernel_img_mul_5[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_5[0] <= { {8{1'b0}},layer0[5][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_5[1] <= { {8{1'b0}},layer0[5][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_5[2] <= { {8{1'b0}},layer0[5][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_5[3] <= { {8{1'b0}},layer1[5][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_5[4] <= { {8{1'b0}},layer1[5][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_5[5] <= { {8{1'b0}},layer1[5][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_5[6] <= { {8{1'b0}},layer2[5][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_5[7] <= { {8{1'b0}},layer2[5][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_5[8] <= { {8{1'b0}},layer2[5][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_5;
reg  [15:0]  kernel_img_sum_2_5;
reg  [15:0]  kernel_img_sum_3_5;
reg  [15:0]  kernel_img_sum_4_5;
reg  [15:0]  kernel_img_sum_5_5;
reg  [15:0]  kernel_img_sum_6_5;
reg  [15:0]  kernel_img_sum_7_5;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_5 <= kernel_img_mul_5[0] + kernel_img_mul_5[1] + kernel_img_mul_5[2] + kernel_img_mul_5[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_5 <= kernel_img_mul_5[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_5 <= kernel_img_mul_5[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_5 <= kernel_img_mul_5[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_5 <= kernel_img_mul_5[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_5 <= kernel_img_mul_5[8];
  end
end
always@(*) begin
  kernel_img_sum_7_5 = kernel_img_sum_1_5 + kernel_img_sum_2_5 + kernel_img_sum_3_5 + kernel_img_sum_4_5 + kernel_img_sum_5_5 + kernel_img_sum_6_5;
end
reg  [15:0]  kernel_img_mul_6[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_6[0] <= 'd0;
    kernel_img_mul_6[1] <= 'd0;
    kernel_img_mul_6[2] <= 'd0;
    kernel_img_mul_6[3] <= 'd0;
    kernel_img_mul_6[4] <= 'd0;
    kernel_img_mul_6[5] <= 'd0;
    kernel_img_mul_6[6] <= 'd0;
    kernel_img_mul_6[7] <= 'd0;
    kernel_img_mul_6[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_6[0] <= { {8{1'b0}},layer0[6][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_6[1] <= { {8{1'b0}},layer0[6][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_6[2] <= { {8{1'b0}},layer0[6][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_6[3] <= { {8{1'b0}},layer1[6][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_6[4] <= { {8{1'b0}},layer1[6][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_6[5] <= { {8{1'b0}},layer1[6][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_6[6] <= { {8{1'b0}},layer2[6][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_6[7] <= { {8{1'b0}},layer2[6][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_6[8] <= { {8{1'b0}},layer2[6][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_6;
reg  [15:0]  kernel_img_sum_2_6;
reg  [15:0]  kernel_img_sum_3_6;
reg  [15:0]  kernel_img_sum_4_6;
reg  [15:0]  kernel_img_sum_5_6;
reg  [15:0]  kernel_img_sum_6_6;
reg  [15:0]  kernel_img_sum_7_6;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_6 <= kernel_img_mul_6[0] + kernel_img_mul_6[1] + kernel_img_mul_6[2] + kernel_img_mul_6[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_6 <= kernel_img_mul_6[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_6 <= kernel_img_mul_6[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_6 <= kernel_img_mul_6[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_6 <= kernel_img_mul_6[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_6 <= kernel_img_mul_6[8];
  end
end
always@(*) begin
  kernel_img_sum_7_6 = kernel_img_sum_1_6 + kernel_img_sum_2_6 + kernel_img_sum_3_6 + kernel_img_sum_4_6 + kernel_img_sum_5_6 + kernel_img_sum_6_6;
end
reg  [15:0]  kernel_img_mul_7[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_7[0] <= 'd0;
    kernel_img_mul_7[1] <= 'd0;
    kernel_img_mul_7[2] <= 'd0;
    kernel_img_mul_7[3] <= 'd0;
    kernel_img_mul_7[4] <= 'd0;
    kernel_img_mul_7[5] <= 'd0;
    kernel_img_mul_7[6] <= 'd0;
    kernel_img_mul_7[7] <= 'd0;
    kernel_img_mul_7[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_7[0] <= { {8{1'b0}},layer0[7][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_7[1] <= { {8{1'b0}},layer0[7][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_7[2] <= { {8{1'b0}},layer0[7][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_7[3] <= { {8{1'b0}},layer1[7][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_7[4] <= { {8{1'b0}},layer1[7][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_7[5] <= { {8{1'b0}},layer1[7][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_7[6] <= { {8{1'b0}},layer2[7][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_7[7] <= { {8{1'b0}},layer2[7][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_7[8] <= { {8{1'b0}},layer2[7][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_7;
reg  [15:0]  kernel_img_sum_2_7;
reg  [15:0]  kernel_img_sum_3_7;
reg  [15:0]  kernel_img_sum_4_7;
reg  [15:0]  kernel_img_sum_5_7;
reg  [15:0]  kernel_img_sum_6_7;
reg  [15:0]  kernel_img_sum_7_7;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_7 <= kernel_img_mul_7[0] + kernel_img_mul_7[1] + kernel_img_mul_7[2] + kernel_img_mul_7[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_7 <= kernel_img_mul_7[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_7 <= kernel_img_mul_7[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_7 <= kernel_img_mul_7[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_7 <= kernel_img_mul_7[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_7 <= kernel_img_mul_7[8];
  end
end
always@(*) begin
  kernel_img_sum_7_7 = kernel_img_sum_1_7 + kernel_img_sum_2_7 + kernel_img_sum_3_7 + kernel_img_sum_4_7 + kernel_img_sum_5_7 + kernel_img_sum_6_7;
end
reg  [15:0]  kernel_img_mul_8[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_8[0] <= 'd0;
    kernel_img_mul_8[1] <= 'd0;
    kernel_img_mul_8[2] <= 'd0;
    kernel_img_mul_8[3] <= 'd0;
    kernel_img_mul_8[4] <= 'd0;
    kernel_img_mul_8[5] <= 'd0;
    kernel_img_mul_8[6] <= 'd0;
    kernel_img_mul_8[7] <= 'd0;
    kernel_img_mul_8[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_8[0] <= { {8{1'b0}},layer0[8][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_8[1] <= { {8{1'b0}},layer0[8][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_8[2] <= { {8{1'b0}},layer0[8][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_8[3] <= { {8{1'b0}},layer1[8][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_8[4] <= { {8{1'b0}},layer1[8][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_8[5] <= { {8{1'b0}},layer1[8][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_8[6] <= { {8{1'b0}},layer2[8][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_8[7] <= { {8{1'b0}},layer2[8][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_8[8] <= { {8{1'b0}},layer2[8][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_8;
reg  [15:0]  kernel_img_sum_2_8;
reg  [15:0]  kernel_img_sum_3_8;
reg  [15:0]  kernel_img_sum_4_8;
reg  [15:0]  kernel_img_sum_5_8;
reg  [15:0]  kernel_img_sum_6_8;
reg  [15:0]  kernel_img_sum_7_8;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_8 <= kernel_img_mul_8[0] + kernel_img_mul_8[1] + kernel_img_mul_8[2] + kernel_img_mul_8[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_8 <= kernel_img_mul_8[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_8 <= kernel_img_mul_8[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_8 <= kernel_img_mul_8[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_8 <= kernel_img_mul_8[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_8 <= kernel_img_mul_8[8];
  end
end
always@(*) begin
  kernel_img_sum_7_8 = kernel_img_sum_1_8 + kernel_img_sum_2_8 + kernel_img_sum_3_8 + kernel_img_sum_4_8 + kernel_img_sum_5_8 + kernel_img_sum_6_8;
end
reg  [15:0]  kernel_img_mul_9[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_9[0] <= 'd0;
    kernel_img_mul_9[1] <= 'd0;
    kernel_img_mul_9[2] <= 'd0;
    kernel_img_mul_9[3] <= 'd0;
    kernel_img_mul_9[4] <= 'd0;
    kernel_img_mul_9[5] <= 'd0;
    kernel_img_mul_9[6] <= 'd0;
    kernel_img_mul_9[7] <= 'd0;
    kernel_img_mul_9[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_9[0] <= { {8{1'b0}},layer0[9][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_9[1] <= { {8{1'b0}},layer0[9][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_9[2] <= { {8{1'b0}},layer0[9][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_9[3] <= { {8{1'b0}},layer1[9][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_9[4] <= { {8{1'b0}},layer1[9][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_9[5] <= { {8{1'b0}},layer1[9][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_9[6] <= { {8{1'b0}},layer2[9][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_9[7] <= { {8{1'b0}},layer2[9][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_9[8] <= { {8{1'b0}},layer2[9][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_9;
reg  [15:0]  kernel_img_sum_2_9;
reg  [15:0]  kernel_img_sum_3_9;
reg  [15:0]  kernel_img_sum_4_9;
reg  [15:0]  kernel_img_sum_5_9;
reg  [15:0]  kernel_img_sum_6_9;
reg  [15:0]  kernel_img_sum_7_9;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_9 <= kernel_img_mul_9[0] + kernel_img_mul_9[1] + kernel_img_mul_9[2] + kernel_img_mul_9[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_9 <= kernel_img_mul_9[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_9 <= kernel_img_mul_9[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_9 <= kernel_img_mul_9[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_9 <= kernel_img_mul_9[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_9 <= kernel_img_mul_9[8];
  end
end
always@(*) begin
  kernel_img_sum_7_9 = kernel_img_sum_1_9 + kernel_img_sum_2_9 + kernel_img_sum_3_9 + kernel_img_sum_4_9 + kernel_img_sum_5_9 + kernel_img_sum_6_9;
end
reg  [15:0]  kernel_img_mul_10[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_10[0] <= 'd0;
    kernel_img_mul_10[1] <= 'd0;
    kernel_img_mul_10[2] <= 'd0;
    kernel_img_mul_10[3] <= 'd0;
    kernel_img_mul_10[4] <= 'd0;
    kernel_img_mul_10[5] <= 'd0;
    kernel_img_mul_10[6] <= 'd0;
    kernel_img_mul_10[7] <= 'd0;
    kernel_img_mul_10[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_10[0] <= { {8{1'b0}},layer0[10][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_10[1] <= { {8{1'b0}},layer0[10][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_10[2] <= { {8{1'b0}},layer0[10][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_10[3] <= { {8{1'b0}},layer1[10][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_10[4] <= { {8{1'b0}},layer1[10][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_10[5] <= { {8{1'b0}},layer1[10][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_10[6] <= { {8{1'b0}},layer2[10][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_10[7] <= { {8{1'b0}},layer2[10][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_10[8] <= { {8{1'b0}},layer2[10][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_10;
reg  [15:0]  kernel_img_sum_2_10;
reg  [15:0]  kernel_img_sum_3_10;
reg  [15:0]  kernel_img_sum_4_10;
reg  [15:0]  kernel_img_sum_5_10;
reg  [15:0]  kernel_img_sum_6_10;
reg  [15:0]  kernel_img_sum_7_10;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_10 <= kernel_img_mul_10[0] + kernel_img_mul_10[1] + kernel_img_mul_10[2] + kernel_img_mul_10[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_10 <= kernel_img_mul_10[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_10 <= kernel_img_mul_10[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_10 <= kernel_img_mul_10[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_10 <= kernel_img_mul_10[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_10 <= kernel_img_mul_10[8];
  end
end
always@(*) begin
  kernel_img_sum_7_10 = kernel_img_sum_1_10 + kernel_img_sum_2_10 + kernel_img_sum_3_10 + kernel_img_sum_4_10 + kernel_img_sum_5_10 + kernel_img_sum_6_10;
end
reg  [15:0]  kernel_img_mul_11[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_11[0] <= 'd0;
    kernel_img_mul_11[1] <= 'd0;
    kernel_img_mul_11[2] <= 'd0;
    kernel_img_mul_11[3] <= 'd0;
    kernel_img_mul_11[4] <= 'd0;
    kernel_img_mul_11[5] <= 'd0;
    kernel_img_mul_11[6] <= 'd0;
    kernel_img_mul_11[7] <= 'd0;
    kernel_img_mul_11[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_11[0] <= { {8{1'b0}},layer0[11][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_11[1] <= { {8{1'b0}},layer0[11][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_11[2] <= { {8{1'b0}},layer0[11][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_11[3] <= { {8{1'b0}},layer1[11][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_11[4] <= { {8{1'b0}},layer1[11][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_11[5] <= { {8{1'b0}},layer1[11][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_11[6] <= { {8{1'b0}},layer2[11][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_11[7] <= { {8{1'b0}},layer2[11][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_11[8] <= { {8{1'b0}},layer2[11][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_11;
reg  [15:0]  kernel_img_sum_2_11;
reg  [15:0]  kernel_img_sum_3_11;
reg  [15:0]  kernel_img_sum_4_11;
reg  [15:0]  kernel_img_sum_5_11;
reg  [15:0]  kernel_img_sum_6_11;
reg  [15:0]  kernel_img_sum_7_11;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_11 <= kernel_img_mul_11[0] + kernel_img_mul_11[1] + kernel_img_mul_11[2] + kernel_img_mul_11[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_11 <= kernel_img_mul_11[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_11 <= kernel_img_mul_11[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_11 <= kernel_img_mul_11[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_11 <= kernel_img_mul_11[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_11 <= kernel_img_mul_11[8];
  end
end
always@(*) begin
  kernel_img_sum_7_11 = kernel_img_sum_1_11 + kernel_img_sum_2_11 + kernel_img_sum_3_11 + kernel_img_sum_4_11 + kernel_img_sum_5_11 + kernel_img_sum_6_11;
end
reg  [15:0]  kernel_img_mul_12[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_12[0] <= 'd0;
    kernel_img_mul_12[1] <= 'd0;
    kernel_img_mul_12[2] <= 'd0;
    kernel_img_mul_12[3] <= 'd0;
    kernel_img_mul_12[4] <= 'd0;
    kernel_img_mul_12[5] <= 'd0;
    kernel_img_mul_12[6] <= 'd0;
    kernel_img_mul_12[7] <= 'd0;
    kernel_img_mul_12[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_12[0] <= { {8{1'b0}},layer0[12][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_12[1] <= { {8{1'b0}},layer0[12][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_12[2] <= { {8{1'b0}},layer0[12][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_12[3] <= { {8{1'b0}},layer1[12][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_12[4] <= { {8{1'b0}},layer1[12][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_12[5] <= { {8{1'b0}},layer1[12][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_12[6] <= { {8{1'b0}},layer2[12][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_12[7] <= { {8{1'b0}},layer2[12][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_12[8] <= { {8{1'b0}},layer2[12][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_12;
reg  [15:0]  kernel_img_sum_2_12;
reg  [15:0]  kernel_img_sum_3_12;
reg  [15:0]  kernel_img_sum_4_12;
reg  [15:0]  kernel_img_sum_5_12;
reg  [15:0]  kernel_img_sum_6_12;
reg  [15:0]  kernel_img_sum_7_12;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_12 <= kernel_img_mul_12[0] + kernel_img_mul_12[1] + kernel_img_mul_12[2] + kernel_img_mul_12[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_12 <= kernel_img_mul_12[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_12 <= kernel_img_mul_12[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_12 <= kernel_img_mul_12[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_12 <= kernel_img_mul_12[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_12 <= kernel_img_mul_12[8];
  end
end
always@(*) begin
  kernel_img_sum_7_12 = kernel_img_sum_1_12 + kernel_img_sum_2_12 + kernel_img_sum_3_12 + kernel_img_sum_4_12 + kernel_img_sum_5_12 + kernel_img_sum_6_12;
end
reg  [15:0]  kernel_img_mul_13[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_13[0] <= 'd0;
    kernel_img_mul_13[1] <= 'd0;
    kernel_img_mul_13[2] <= 'd0;
    kernel_img_mul_13[3] <= 'd0;
    kernel_img_mul_13[4] <= 'd0;
    kernel_img_mul_13[5] <= 'd0;
    kernel_img_mul_13[6] <= 'd0;
    kernel_img_mul_13[7] <= 'd0;
    kernel_img_mul_13[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_13[0] <= { {8{1'b0}},layer0[13][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_13[1] <= { {8{1'b0}},layer0[13][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_13[2] <= { {8{1'b0}},layer0[13][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_13[3] <= { {8{1'b0}},layer1[13][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_13[4] <= { {8{1'b0}},layer1[13][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_13[5] <= { {8{1'b0}},layer1[13][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_13[6] <= { {8{1'b0}},layer2[13][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_13[7] <= { {8{1'b0}},layer2[13][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_13[8] <= { {8{1'b0}},layer2[13][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_13;
reg  [15:0]  kernel_img_sum_2_13;
reg  [15:0]  kernel_img_sum_3_13;
reg  [15:0]  kernel_img_sum_4_13;
reg  [15:0]  kernel_img_sum_5_13;
reg  [15:0]  kernel_img_sum_6_13;
reg  [15:0]  kernel_img_sum_7_13;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_13 <= kernel_img_mul_13[0] + kernel_img_mul_13[1] + kernel_img_mul_13[2] + kernel_img_mul_13[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_13 <= kernel_img_mul_13[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_13 <= kernel_img_mul_13[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_13 <= kernel_img_mul_13[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_13 <= kernel_img_mul_13[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_13 <= kernel_img_mul_13[8];
  end
end
always@(*) begin
  kernel_img_sum_7_13 = kernel_img_sum_1_13 + kernel_img_sum_2_13 + kernel_img_sum_3_13 + kernel_img_sum_4_13 + kernel_img_sum_5_13 + kernel_img_sum_6_13;
end
reg  [15:0]  kernel_img_mul_14[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_14[0] <= 'd0;
    kernel_img_mul_14[1] <= 'd0;
    kernel_img_mul_14[2] <= 'd0;
    kernel_img_mul_14[3] <= 'd0;
    kernel_img_mul_14[4] <= 'd0;
    kernel_img_mul_14[5] <= 'd0;
    kernel_img_mul_14[6] <= 'd0;
    kernel_img_mul_14[7] <= 'd0;
    kernel_img_mul_14[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_14[0] <= { {8{1'b0}},layer0[14][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_14[1] <= { {8{1'b0}},layer0[14][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_14[2] <= { {8{1'b0}},layer0[14][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_14[3] <= { {8{1'b0}},layer1[14][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_14[4] <= { {8{1'b0}},layer1[14][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_14[5] <= { {8{1'b0}},layer1[14][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_14[6] <= { {8{1'b0}},layer2[14][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_14[7] <= { {8{1'b0}},layer2[14][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_14[8] <= { {8{1'b0}},layer2[14][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_14;
reg  [15:0]  kernel_img_sum_2_14;
reg  [15:0]  kernel_img_sum_3_14;
reg  [15:0]  kernel_img_sum_4_14;
reg  [15:0]  kernel_img_sum_5_14;
reg  [15:0]  kernel_img_sum_6_14;
reg  [15:0]  kernel_img_sum_7_14;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_14 <= kernel_img_mul_14[0] + kernel_img_mul_14[1] + kernel_img_mul_14[2] + kernel_img_mul_14[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_14 <= kernel_img_mul_14[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_14 <= kernel_img_mul_14[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_14 <= kernel_img_mul_14[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_14 <= kernel_img_mul_14[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_14 <= kernel_img_mul_14[8];
  end
end
always@(*) begin
  kernel_img_sum_7_14 = kernel_img_sum_1_14 + kernel_img_sum_2_14 + kernel_img_sum_3_14 + kernel_img_sum_4_14 + kernel_img_sum_5_14 + kernel_img_sum_6_14;
end
reg  [15:0]  kernel_img_mul_15[0:8];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_15[0] <= 'd0;
    kernel_img_mul_15[1] <= 'd0;
    kernel_img_mul_15[2] <= 'd0;
    kernel_img_mul_15[3] <= 'd0;
    kernel_img_mul_15[4] <= 'd0;
    kernel_img_mul_15[5] <= 'd0;
    kernel_img_mul_15[6] <= 'd0;
    kernel_img_mul_15[7] <= 'd0;
    kernel_img_mul_15[8] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_15[0] <= { {8{1'b0}},layer0[15][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_15[1] <= { {8{1'b0}},layer0[15][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_15[2] <= { {8{1'b0}},layer0[15][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
    kernel_img_mul_15[3] <= { {8{1'b0}},layer1[15][7:0]} * { {8{1'b0}}, G_Kernel_3x3_1[7:0]};
    kernel_img_mul_15[4] <= { {8{1'b0}},layer1[15][15:8]} * { {8{1'b0}}, G_Kernel_3x3_1[15:8]};
    kernel_img_mul_15[5] <= { {8{1'b0}},layer1[15][23:16]} * { {8{1'b0}}, G_Kernel_3x3_1[23:16]};
    kernel_img_mul_15[6] <= { {8{1'b0}},layer2[15][7:0]} * { {8{1'b0}}, G_Kernel_3x3_0[7:0]};
    kernel_img_mul_15[7] <= { {8{1'b0}},layer2[15][15:8]} * { {8{1'b0}}, G_Kernel_3x3_0[15:8]};
    kernel_img_mul_15[8] <= { {8{1'b0}},layer2[15][23:16]} * { {8{1'b0}}, G_Kernel_3x3_0[23:16]};
  end
end
reg  [15:0]  kernel_img_sum_1_15;
reg  [15:0]  kernel_img_sum_2_15;
reg  [15:0]  kernel_img_sum_3_15;
reg  [15:0]  kernel_img_sum_4_15;
reg  [15:0]  kernel_img_sum_5_15;
reg  [15:0]  kernel_img_sum_6_15;
reg  [15:0]  kernel_img_sum_7_15;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_15 <= kernel_img_mul_15[0] + kernel_img_mul_15[1] + kernel_img_mul_15[2] + kernel_img_mul_15[3];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_15 <= kernel_img_mul_15[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_15 <= kernel_img_mul_15[5];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_15 <= kernel_img_mul_15[6];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_15 <= kernel_img_mul_15[7];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_15 <= kernel_img_mul_15[8];
  end
end
always@(*) begin
  kernel_img_sum_7_15 = kernel_img_sum_1_15 + kernel_img_sum_2_15 + kernel_img_sum_3_15 + kernel_img_sum_4_15 + kernel_img_sum_5_15 + kernel_img_sum_6_15;
end
always @(posedge clk) begin
  if(!rst_n) begin
    blur_out[7:0] <= 'd0;
    blur_out[15:8] <= 'd0;
    blur_out[23:16] <= 'd0;
    blur_out[31:24] <= 'd0;
    blur_out[39:32] <= 'd0;
    blur_out[47:40] <= 'd0;
    blur_out[55:48] <= 'd0;
    blur_out[63:56] <= 'd0;
    blur_out[71:64] <= 'd0;
    blur_out[79:72] <= 'd0;
    blur_out[87:80] <= 'd0;
    blur_out[95:88] <= 'd0;
    blur_out[103:96] <= 'd0;
    blur_out[111:104] <= 'd0;
    blur_out[119:112] <= 'd0;
    blur_out[127:120] <= 'd0;
  end
  else if(current_state==ST_UPDATE) begin
    blur_out[7:0] <= kernel_img_sum_7_0[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[15:8] <= kernel_img_sum_7_1[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[23:16] <= kernel_img_sum_7_2[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[31:24] <= kernel_img_sum_7_3[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[39:32] <= kernel_img_sum_7_4[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[47:40] <= kernel_img_sum_7_5[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[55:48] <= kernel_img_sum_7_6[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[63:56] <= kernel_img_sum_7_7[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[71:64] <= kernel_img_sum_7_8[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[79:72] <= kernel_img_sum_7_9[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[87:80] <= kernel_img_sum_7_10[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[95:88] <= kernel_img_sum_7_11[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[103:96] <= kernel_img_sum_7_12[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[111:104] <= kernel_img_sum_7_13[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[119:112] <= kernel_img_sum_7_14[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[127:120] <= kernel_img_sum_7_15[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
  end
end

/*
 *  FSM
 *
 */
always @(posedge clk) begin
  if (!rst_n) begin
    current_state <= ST_MUX;    
  end
  else begin
    current_state <= next_state;
  end
end
always @(*) begin
  case(current_state)
    ST_MUX: begin
      if(start)
        next_state = ST_MUL;
      else
        next_state = ST_MUX;
    end
    ST_MUL: begin
      if(current_state==ST_MUL)
        next_state = ST_ADD;
      else 
        next_state = ST_MUL;
    end
    ST_ADD: begin
      if(current_state==ST_ADD)
        next_state = ST_UPDATE;
      else 
        next_state = ST_ADD;
    end
    ST_UPDATE: begin
      if(current_state==ST_UPDATE)
        next_state = ST_MUL;
      else 
        next_state = ST_UPDATE;
    end
    default:
      next_state = ST_MUL;
  endcase
end

endmodule